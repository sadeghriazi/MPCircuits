
module knn_comb_BMR_W16_K2_N128 ( p_input, o );
  input [2063:0] p_input;
  output [31:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][15] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
         n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
         n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
         n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
         n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
         n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
         n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
         n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
         n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
         n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
         n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
         n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459,
         n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
         n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
         n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483,
         n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
         n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
         n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507,
         n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
         n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
         n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
         n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
         n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
         n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555,
         n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
         n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
         n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579,
         n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
         n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
         n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603,
         n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
         n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
         n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
         n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635,
         n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643,
         n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651,
         n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
         n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
         n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675,
         n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683,
         n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691,
         n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699,
         n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707,
         n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715,
         n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723,
         n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
         n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
         n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747,
         n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755,
         n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763,
         n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771,
         n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
         n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787,
         n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795,
         n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
         n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
         n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819,
         n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827,
         n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835,
         n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843,
         n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851,
         n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859,
         n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867,
         n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
         n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
         n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891,
         n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899,
         n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
         n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915,
         n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923,
         n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931,
         n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939,
         n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947,
         n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955,
         n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963,
         n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971,
         n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979,
         n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987,
         n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995,
         n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003,
         n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011,
         n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019,
         n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027,
         n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035,
         n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043,
         n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
         n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059,
         n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067,
         n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075,
         n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083,
         n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091,
         n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099,
         n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107,
         n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115,
         n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
         n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131,
         n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139,
         n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147,
         n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155,
         n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163,
         n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171,
         n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179,
         n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187,
         n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
         n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203,
         n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211,
         n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219,
         n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227,
         n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235,
         n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243,
         n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251,
         n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259,
         n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267,
         n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275,
         n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283,
         n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291,
         n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299,
         n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307,
         n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315,
         n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323,
         n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331,
         n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339,
         n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347,
         n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355,
         n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363,
         n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371,
         n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379,
         n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387,
         n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395,
         n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403,
         n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411,
         n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419,
         n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427,
         n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435,
         n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443,
         n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451,
         n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459,
         n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467,
         n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475,
         n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483,
         n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491,
         n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499,
         n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507,
         n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515,
         n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523,
         n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531,
         n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539,
         n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547,
         n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555,
         n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563,
         n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571,
         n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579,
         n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587,
         n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595,
         n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603,
         n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611,
         n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619,
         n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627,
         n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635,
         n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643,
         n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651,
         n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659,
         n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667,
         n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675,
         n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683,
         n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691,
         n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699,
         n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707,
         n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715,
         n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723,
         n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731,
         n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739,
         n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747,
         n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755,
         n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763,
         n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771,
         n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779,
         n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787,
         n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795,
         n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803,
         n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811,
         n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819,
         n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827,
         n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835,
         n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843,
         n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851,
         n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859,
         n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867,
         n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875,
         n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883,
         n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891,
         n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899,
         n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907,
         n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915,
         n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923,
         n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931,
         n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939,
         n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947,
         n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955,
         n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963,
         n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971,
         n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979,
         n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987,
         n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995,
         n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003,
         n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011,
         n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019,
         n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027,
         n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035,
         n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043,
         n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051,
         n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059,
         n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067,
         n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075,
         n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083,
         n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091,
         n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099,
         n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107,
         n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115,
         n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123,
         n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131,
         n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139,
         n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147,
         n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155,
         n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163,
         n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171,
         n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179,
         n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187,
         n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195,
         n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203,
         n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211,
         n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219,
         n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227,
         n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235,
         n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243,
         n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251,
         n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259,
         n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267,
         n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275,
         n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283,
         n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291,
         n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299,
         n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307,
         n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315,
         n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323,
         n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331,
         n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339,
         n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347,
         n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355,
         n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363,
         n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371,
         n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379,
         n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387,
         n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395,
         n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403,
         n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411,
         n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419,
         n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427,
         n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435,
         n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443,
         n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451,
         n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459,
         n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467,
         n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475,
         n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483,
         n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491,
         n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499,
         n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507,
         n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515,
         n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523,
         n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531,
         n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539,
         n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547,
         n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555,
         n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563,
         n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571,
         n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579,
         n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587,
         n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595,
         n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603,
         n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611,
         n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619,
         n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627,
         n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635,
         n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643,
         n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651,
         n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659,
         n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667,
         n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675,
         n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683,
         n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691,
         n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699,
         n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707,
         n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715,
         n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723,
         n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731,
         n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739,
         n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747,
         n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755,
         n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763,
         n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771,
         n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779,
         n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787,
         n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795,
         n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803,
         n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811,
         n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819,
         n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827,
         n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835,
         n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843,
         n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851,
         n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859,
         n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867,
         n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875,
         n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883,
         n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891,
         n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899,
         n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907,
         n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915,
         n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923,
         n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931,
         n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939,
         n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
         n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955,
         n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963,
         n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971,
         n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979,
         n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987,
         n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995,
         n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003,
         n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011,
         n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019,
         n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027,
         n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035,
         n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043,
         n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051,
         n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059,
         n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067,
         n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075,
         n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083,
         n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091,
         n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099,
         n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107,
         n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115,
         n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123,
         n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131,
         n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139,
         n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147,
         n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155,
         n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163,
         n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171,
         n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179,
         n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187,
         n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195,
         n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203,
         n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211,
         n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219,
         n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227,
         n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235,
         n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243,
         n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251,
         n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259,
         n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267,
         n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275,
         n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283,
         n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291,
         n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299,
         n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307,
         n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315,
         n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323,
         n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331,
         n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339,
         n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347,
         n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355,
         n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363,
         n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371,
         n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379,
         n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387,
         n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395,
         n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403,
         n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411,
         n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419,
         n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427,
         n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435,
         n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443,
         n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451,
         n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459,
         n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467,
         n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475,
         n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483,
         n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491,
         n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499,
         n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507,
         n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515,
         n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523,
         n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531,
         n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539,
         n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547,
         n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555,
         n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563,
         n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571,
         n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579,
         n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587,
         n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595,
         n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603,
         n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611,
         n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619,
         n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627,
         n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635,
         n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643,
         n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651,
         n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659,
         n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667,
         n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675,
         n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683,
         n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691,
         n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699,
         n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707,
         n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715,
         n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723,
         n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731,
         n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739,
         n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747,
         n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755,
         n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763,
         n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771,
         n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779,
         n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787,
         n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795,
         n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803,
         n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811,
         n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819,
         n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827,
         n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835,
         n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843,
         n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851,
         n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859,
         n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867,
         n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875,
         n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883,
         n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891,
         n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899,
         n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907,
         n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915,
         n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923,
         n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931,
         n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939,
         n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947,
         n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955,
         n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963,
         n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971,
         n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979,
         n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987,
         n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995,
         n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003,
         n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011,
         n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019,
         n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027,
         n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035,
         n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043,
         n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051,
         n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059,
         n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067,
         n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075,
         n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083,
         n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091,
         n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099,
         n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107,
         n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115,
         n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123,
         n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131,
         n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139,
         n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147,
         n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155,
         n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163,
         n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171,
         n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179,
         n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187,
         n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195,
         n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203,
         n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211,
         n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219,
         n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227,
         n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235,
         n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243,
         n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251,
         n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259,
         n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267,
         n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275,
         n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283,
         n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291,
         n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299,
         n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307,
         n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315,
         n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323,
         n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331,
         n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339,
         n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347,
         n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355,
         n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363,
         n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371,
         n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379,
         n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387,
         n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395,
         n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403,
         n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411,
         n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419,
         n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427,
         n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435,
         n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443,
         n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451,
         n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459,
         n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467,
         n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475,
         n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483,
         n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491,
         n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499,
         n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507,
         n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515,
         n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523,
         n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531,
         n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539,
         n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547,
         n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555,
         n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563,
         n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571,
         n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579,
         n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587,
         n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595,
         n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603,
         n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611,
         n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619,
         n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627,
         n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635,
         n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643,
         n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651,
         n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659,
         n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667,
         n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675,
         n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683,
         n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691,
         n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699,
         n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707,
         n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715,
         n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723,
         n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731,
         n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739,
         n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747,
         n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755,
         n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763,
         n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771,
         n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779,
         n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787,
         n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795,
         n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803,
         n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811,
         n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819,
         n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827,
         n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835,
         n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843,
         n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851,
         n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859,
         n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867,
         n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875,
         n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883,
         n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891,
         n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899,
         n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907,
         n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915,
         n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923,
         n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931,
         n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939,
         n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947,
         n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955,
         n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963,
         n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971,
         n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979,
         n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987,
         n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995,
         n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003,
         n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011,
         n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019,
         n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027,
         n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035,
         n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043,
         n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051,
         n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059,
         n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067,
         n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075,
         n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083,
         n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091,
         n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099,
         n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107,
         n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115,
         n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123,
         n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131,
         n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139,
         n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147,
         n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155,
         n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163,
         n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171,
         n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179,
         n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187,
         n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195,
         n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203,
         n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211,
         n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219,
         n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227,
         n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235,
         n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243,
         n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251,
         n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259,
         n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267,
         n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275,
         n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283,
         n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291,
         n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299,
         n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307,
         n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315,
         n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323,
         n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331,
         n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339,
         n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347,
         n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355,
         n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363,
         n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371,
         n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379,
         n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387,
         n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395,
         n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403,
         n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411,
         n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419,
         n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427,
         n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435,
         n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443,
         n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451,
         n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459,
         n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467,
         n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475,
         n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483,
         n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491,
         n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499,
         n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507,
         n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515,
         n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523,
         n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531,
         n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539,
         n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547,
         n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555,
         n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563,
         n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571,
         n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579,
         n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587,
         n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595,
         n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603,
         n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611,
         n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619,
         n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627,
         n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635,
         n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643,
         n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651,
         n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659,
         n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667,
         n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675,
         n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683,
         n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691,
         n26692, n26693, n26694, n26695, n26696, n26697, n26698, n26699,
         n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707,
         n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715,
         n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723,
         n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731,
         n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739,
         n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747,
         n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755,
         n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763,
         n26764, n26765, n26766, n26767, n26768, n26769, n26770, n26771,
         n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779,
         n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787,
         n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795,
         n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803,
         n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811,
         n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819,
         n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827,
         n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835,
         n26836, n26837, n26838, n26839, n26840, n26841, n26842, n26843,
         n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851,
         n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859,
         n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867,
         n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875,
         n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883,
         n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891,
         n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899,
         n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907,
         n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915,
         n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923,
         n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931,
         n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939,
         n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947,
         n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955,
         n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963,
         n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971,
         n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979,
         n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987,
         n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995,
         n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003,
         n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011,
         n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019,
         n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027,
         n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035,
         n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043,
         n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051,
         n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059,
         n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067,
         n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075,
         n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083,
         n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091,
         n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099,
         n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107,
         n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115,
         n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123,
         n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131,
         n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139,
         n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147,
         n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155,
         n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163,
         n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171,
         n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179,
         n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187,
         n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195,
         n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203,
         n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211,
         n27212, n27213, n27214, n27215, n27216, n27217, n27218, n27219,
         n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227,
         n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235,
         n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243,
         n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251,
         n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259,
         n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267,
         n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275,
         n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283,
         n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291,
         n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299,
         n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307,
         n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315,
         n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323,
         n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331,
         n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339,
         n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347,
         n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355,
         n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363,
         n27364, n27365, n27366, n27367, n27368, n27369, n27370, n27371,
         n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379,
         n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387,
         n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395,
         n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403,
         n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411,
         n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419,
         n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427,
         n27428, n27429, n27430, n27431, n27432, n27433, n27434, n27435,
         n27436, n27437, n27438, n27439, n27440, n27441, n27442, n27443,
         n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451,
         n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459,
         n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467,
         n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475,
         n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483,
         n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491,
         n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499,
         n27500, n27501, n27502, n27503, n27504, n27505, n27506, n27507,
         n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515,
         n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523,
         n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531,
         n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539,
         n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547,
         n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555,
         n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563,
         n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571,
         n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579,
         n27580, n27581, n27582, n27583, n27584, n27585, n27586, n27587,
         n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595,
         n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603,
         n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611,
         n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619,
         n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627,
         n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635,
         n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643,
         n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651,
         n27652, n27653, n27654, n27655, n27656, n27657, n27658, n27659,
         n27660, n27661, n27662, n27663, n27664, n27665, n27666, n27667,
         n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675,
         n27676, n27677, n27678, n27679, n27680, n27681, n27682, n27683,
         n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691,
         n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699,
         n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707,
         n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715,
         n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723,
         n27724, n27725, n27726, n27727, n27728, n27729, n27730, n27731,
         n27732, n27733, n27734, n27735, n27736, n27737, n27738, n27739,
         n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747,
         n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755,
         n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763,
         n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771,
         n27772, n27773, n27774, n27775, n27776, n27777, n27778, n27779,
         n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787,
         n27788, n27789, n27790, n27791, n27792, n27793, n27794, n27795,
         n27796, n27797, n27798, n27799, n27800, n27801, n27802, n27803,
         n27804, n27805, n27806, n27807, n27808, n27809, n27810, n27811,
         n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819,
         n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827,
         n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835,
         n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843,
         n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851,
         n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859,
         n27860, n27861, n27862, n27863, n27864, n27865, n27866, n27867,
         n27868, n27869, n27870, n27871, n27872, n27873, n27874, n27875,
         n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883,
         n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891,
         n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899,
         n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907,
         n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915,
         n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923,
         n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931,
         n27932, n27933, n27934, n27935, n27936, n27937, n27938, n27939,
         n27940, n27941, n27942, n27943, n27944, n27945, n27946, n27947,
         n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955,
         n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963,
         n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971,
         n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979,
         n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987,
         n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995,
         n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003,
         n28004, n28005, n28006, n28007, n28008, n28009, n28010, n28011,
         n28012, n28013, n28014, n28015, n28016, n28017, n28018, n28019,
         n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027,
         n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035,
         n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043,
         n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051,
         n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059,
         n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067,
         n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075,
         n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083,
         n28084, n28085, n28086, n28087, n28088, n28089, n28090, n28091,
         n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099,
         n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107,
         n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115,
         n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123,
         n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131,
         n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139,
         n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147,
         n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155,
         n28156, n28157, n28158, n28159, n28160, n28161, n28162, n28163,
         n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171,
         n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179,
         n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187,
         n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195,
         n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203,
         n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211,
         n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219,
         n28220, n28221, n28222, n28223, n28224, n28225, n28226, n28227,
         n28228, n28229, n28230, n28231, n28232, n28233, n28234, n28235,
         n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243,
         n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251,
         n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259,
         n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267,
         n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275,
         n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283,
         n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291,
         n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299,
         n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307,
         n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315,
         n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323,
         n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331,
         n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339,
         n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347,
         n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355,
         n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363,
         n28364, n28365, n28366, n28367, n28368, n28369, n28370, n28371,
         n28372, n28373, n28374, n28375, n28376, n28377, n28378, n28379,
         n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387,
         n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395,
         n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403,
         n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411,
         n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419,
         n28420, n28421, n28422, n28423, n28424, n28425, n28426, n28427,
         n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435,
         n28436, n28437, n28438, n28439, n28440, n28441, n28442, n28443,
         n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451,
         n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459,
         n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467,
         n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475,
         n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483,
         n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491,
         n28492, n28493, n28494, n28495, n28496, n28497, n28498, n28499,
         n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507,
         n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515,
         n28516, n28517, n28518, n28519, n28520, n28521, n28522, n28523,
         n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531,
         n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539,
         n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547,
         n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555,
         n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563,
         n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571,
         n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579,
         n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587,
         n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595,
         n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603,
         n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611,
         n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619,
         n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627,
         n28628, n28629, n28630, n28631, n28632, n28633, n28634, n28635,
         n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643,
         n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651,
         n28652, n28653, n28654, n28655, n28656, n28657, n28658, n28659,
         n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667,
         n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675,
         n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683,
         n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691,
         n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699,
         n28700, n28701, n28702, n28703, n28704, n28705, n28706, n28707,
         n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715,
         n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723,
         n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731,
         n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28739,
         n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747,
         n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755,
         n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763,
         n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771,
         n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779,
         n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787,
         n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795,
         n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803,
         n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811,
         n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819,
         n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827,
         n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835,
         n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843,
         n28844, n28845, n28846, n28847, n28848, n28849, n28850, n28851,
         n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859,
         n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867,
         n28868, n28869, n28870, n28871, n28872, n28873, n28874, n28875,
         n28876, n28877, n28878, n28879, n28880, n28881, n28882, n28883,
         n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891,
         n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899,
         n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907,
         n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915,
         n28916, n28917, n28918, n28919, n28920, n28921, n28922, n28923,
         n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931,
         n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939,
         n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947,
         n28948, n28949, n28950, n28951, n28952, n28953, n28954, n28955,
         n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963,
         n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971,
         n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979,
         n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987,
         n28988, n28989, n28990, n28991, n28992, n28993, n28994, n28995,
         n28996, n28997, n28998, n28999, n29000, n29001, n29002, n29003,
         n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011,
         n29012, n29013, n29014, n29015, n29016, n29017, n29018, n29019,
         n29020, n29021, n29022, n29023, n29024, n29025, n29026, n29027,
         n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035,
         n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043,
         n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051,
         n29052, n29053, n29054, n29055, n29056, n29057, n29058, n29059,
         n29060, n29061, n29062, n29063, n29064, n29065, n29066, n29067,
         n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075,
         n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083,
         n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091,
         n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099,
         n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107,
         n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115,
         n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123,
         n29124, n29125, n29126, n29127, n29128, n29129, n29130, n29131,
         n29132, n29133, n29134, n29135, n29136, n29137, n29138, n29139,
         n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147,
         n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155,
         n29156, n29157, n29158, n29159, n29160, n29161, n29162, n29163,
         n29164, n29165, n29166, n29167, n29168, n29169, n29170, n29171,
         n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179,
         n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187,
         n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195,
         n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203,
         n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211,
         n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219,
         n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227,
         n29228, n29229, n29230, n29231, n29232, n29233, n29234, n29235,
         n29236, n29237, n29238, n29239, n29240, n29241, n29242, n29243,
         n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251,
         n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259,
         n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267,
         n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275,
         n29276, n29277, n29278, n29279, n29280, n29281, n29282, n29283,
         n29284, n29285, n29286, n29287, n29288, n29289, n29290, n29291,
         n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299,
         n29300, n29301, n29302, n29303, n29304, n29305, n29306, n29307,
         n29308, n29309, n29310, n29311, n29312, n29313, n29314, n29315,
         n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323,
         n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331,
         n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339,
         n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347,
         n29348, n29349, n29350, n29351, n29352, n29353, n29354, n29355,
         n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363,
         n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371,
         n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379,
         n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387,
         n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395,
         n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403,
         n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411,
         n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29419,
         n29420, n29421, n29422, n29423, n29424, n29425, n29426, n29427,
         n29428, n29429, n29430, n29431, n29432, n29433, n29434, n29435,
         n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443,
         n29444, n29445, n29446, n29447, n29448, n29449, n29450, n29451,
         n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459,
         n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467,
         n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475,
         n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483,
         n29484, n29485, n29486, n29487, n29488, n29489, n29490, n29491,
         n29492, n29493, n29494, n29495, n29496, n29497, n29498, n29499,
         n29500, n29501, n29502, n29503, n29504, n29505, n29506, n29507,
         n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515,
         n29516, n29517, n29518, n29519, n29520, n29521, n29522, n29523,
         n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531,
         n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539,
         n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547,
         n29548, n29549, n29550, n29551, n29552, n29553, n29554, n29555,
         n29556, n29557, n29558, n29559, n29560, n29561, n29562, n29563,
         n29564, n29565, n29566, n29567, n29568, n29569, n29570, n29571,
         n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29579,
         n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587,
         n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595,
         n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603,
         n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611,
         n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619,
         n29620, n29621, n29622, n29623, n29624, n29625, n29626, n29627,
         n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635,
         n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643,
         n29644, n29645, n29646, n29647, n29648, n29649, n29650, n29651,
         n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659,
         n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667,
         n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675,
         n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683,
         n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691,
         n29692, n29693, n29694, n29695, n29696, n29697, n29698, n29699,
         n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707,
         n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715,
         n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723,
         n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731,
         n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739,
         n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747,
         n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755,
         n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763,
         n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771,
         n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779,
         n29780, n29781, n29782, n29783, n29784, n29785, n29786, n29787,
         n29788, n29789, n29790, n29791, n29792, n29793, n29794, n29795,
         n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803,
         n29804, n29805, n29806, n29807, n29808, n29809, n29810, n29811,
         n29812, n29813, n29814, n29815, n29816, n29817, n29818, n29819,
         n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827,
         n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835,
         n29836, n29837, n29838, n29839, n29840, n29841, n29842, n29843,
         n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851,
         n29852, n29853, n29854, n29855, n29856, n29857, n29858, n29859,
         n29860, n29861, n29862, n29863, n29864, n29865, n29866, n29867,
         n29868, n29869, n29870, n29871, n29872, n29873, n29874, n29875,
         n29876, n29877, n29878, n29879, n29880, n29881, n29882, n29883,
         n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891,
         n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899,
         n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907,
         n29908, n29909, n29910, n29911, n29912, n29913, n29914, n29915,
         n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923,
         n29924, n29925, n29926, n29927, n29928, n29929, n29930, n29931,
         n29932, n29933, n29934, n29935, n29936, n29937, n29938, n29939,
         n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947,
         n29948, n29949, n29950, n29951, n29952, n29953, n29954, n29955,
         n29956, n29957, n29958, n29959, n29960, n29961, n29962, n29963,
         n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971,
         n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979,
         n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987,
         n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995,
         n29996, n29997, n29998, n29999, n30000, n30001, n30002, n30003,
         n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011,
         n30012, n30013, n30014, n30015, n30016, n30017, n30018, n30019,
         n30020, n30021, n30022, n30023, n30024, n30025, n30026, n30027,
         n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035,
         n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043,
         n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051,
         n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059,
         n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067,
         n30068, n30069, n30070, n30071, n30072, n30073, n30074, n30075,
         n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083,
         n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091,
         n30092, n30093, n30094, n30095, n30096, n30097, n30098, n30099,
         n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107,
         n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115,
         n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123,
         n30124, n30125, n30126, n30127, n30128, n30129, n30130, n30131,
         n30132, n30133, n30134, n30135, n30136, n30137, n30138, n30139,
         n30140, n30141, n30142, n30143, n30144, n30145, n30146, n30147,
         n30148, n30149, n30150, n30151, n30152, n30153, n30154, n30155,
         n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163,
         n30164, n30165, n30166, n30167, n30168, n30169, n30170, n30171,
         n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179,
         n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187,
         n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195,
         n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203,
         n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211,
         n30212, n30213, n30214, n30215, n30216, n30217, n30218, n30219,
         n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227,
         n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235,
         n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243,
         n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251,
         n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259,
         n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267,
         n30268, n30269, n30270, n30271, n30272, n30273, n30274, n30275,
         n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283,
         n30284, n30285, n30286, n30287, n30288, n30289, n30290, n30291,
         n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299,
         n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307,
         n30308, n30309, n30310, n30311, n30312, n30313, n30314, n30315,
         n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323,
         n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331,
         n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339,
         n30340, n30341, n30342, n30343, n30344, n30345, n30346, n30347,
         n30348, n30349, n30350, n30351, n30352, n30353, n30354, n30355,
         n30356, n30357, n30358, n30359, n30360, n30361, n30362, n30363,
         n30364, n30365, n30366, n30367, n30368, n30369, n30370, n30371,
         n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379,
         n30380, n30381, n30382, n30383, n30384, n30385, n30386, n30387,
         n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395,
         n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403,
         n30404, n30405, n30406, n30407, n30408, n30409, n30410, n30411,
         n30412, n30413, n30414, n30415, n30416, n30417, n30418, n30419,
         n30420, n30421, n30422, n30423, n30424, n30425, n30426, n30427,
         n30428, n30429, n30430, n30431, n30432, n30433, n30434, n30435,
         n30436, n30437, n30438, n30439, n30440, n30441, n30442, n30443,
         n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451,
         n30452, n30453, n30454, n30455, n30456, n30457, n30458, n30459,
         n30460, n30461, n30462, n30463, n30464, n30465, n30466, n30467,
         n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475,
         n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483,
         n30484, n30485, n30486, n30487, n30488, n30489, n30490, n30491,
         n30492, n30493, n30494, n30495, n30496, n30497, n30498, n30499,
         n30500, n30501, n30502, n30503, n30504, n30505, n30506, n30507,
         n30508, n30509, n30510, n30511, n30512, n30513, n30514, n30515,
         n30516, n30517, n30518, n30519, n30520, n30521, n30522, n30523,
         n30524, n30525, n30526, n30527, n30528, n30529, n30530, n30531,
         n30532, n30533, n30534, n30535, n30536, n30537, n30538, n30539,
         n30540, n30541, n30542, n30543, n30544, n30545, n30546, n30547,
         n30548, n30549, n30550, n30551, n30552, n30553, n30554, n30555,
         n30556, n30557, n30558, n30559, n30560, n30561, n30562, n30563,
         n30564, n30565, n30566, n30567, n30568, n30569, n30570, n30571,
         n30572, n30573, n30574, n30575, n30576, n30577, n30578, n30579,
         n30580, n30581, n30582, n30583, n30584, n30585, n30586, n30587,
         n30588, n30589, n30590, n30591, n30592, n30593, n30594, n30595,
         n30596, n30597, n30598, n30599, n30600, n30601, n30602, n30603,
         n30604, n30605, n30606, n30607, n30608, n30609, n30610, n30611,
         n30612, n30613, n30614, n30615, n30616, n30617, n30618, n30619,
         n30620, n30621, n30622, n30623, n30624, n30625, n30626, n30627,
         n30628, n30629, n30630, n30631, n30632, n30633, n30634, n30635,
         n30636, n30637, n30638, n30639, n30640, n30641, n30642, n30643,
         n30644, n30645, n30646, n30647, n30648, n30649, n30650, n30651,
         n30652, n30653, n30654, n30655, n30656, n30657, n30658, n30659,
         n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667,
         n30668, n30669, n30670, n30671, n30672, n30673, n30674, n30675,
         n30676, n30677, n30678, n30679, n30680, n30681, n30682, n30683,
         n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691,
         n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699,
         n30700, n30701, n30702, n30703, n30704, n30705, n30706, n30707,
         n30708, n30709, n30710, n30711, n30712, n30713, n30714, n30715,
         n30716, n30717, n30718, n30719, n30720, n30721, n30722, n30723,
         n30724, n30725, n30726, n30727, n30728, n30729, n30730, n30731,
         n30732, n30733, n30734, n30735, n30736, n30737, n30738, n30739,
         n30740, n30741, n30742, n30743, n30744, n30745, n30746, n30747,
         n30748, n30749, n30750, n30751, n30752, n30753, n30754, n30755,
         n30756, n30757, n30758, n30759, n30760, n30761, n30762, n30763,
         n30764, n30765, n30766, n30767, n30768, n30769, n30770, n30771,
         n30772, n30773, n30774, n30775, n30776, n30777, n30778, n30779,
         n30780, n30781, n30782, n30783, n30784, n30785, n30786, n30787,
         n30788, n30789, n30790, n30791, n30792, n30793, n30794, n30795,
         n30796, n30797, n30798, n30799, n30800, n30801, n30802, n30803,
         n30804, n30805, n30806, n30807, n30808, n30809, n30810, n30811,
         n30812, n30813, n30814, n30815, n30816, n30817, n30818, n30819,
         n30820, n30821, n30822, n30823, n30824, n30825, n30826, n30827,
         n30828, n30829, n30830, n30831, n30832, n30833, n30834, n30835,
         n30836, n30837, n30838, n30839, n30840, n30841, n30842, n30843,
         n30844, n30845, n30846, n30847, n30848, n30849, n30850, n30851,
         n30852, n30853, n30854, n30855, n30856, n30857, n30858, n30859,
         n30860, n30861, n30862, n30863, n30864, n30865, n30866, n30867,
         n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30875,
         n30876, n30877, n30878, n30879, n30880, n30881, n30882, n30883,
         n30884, n30885, n30886, n30887, n30888, n30889, n30890, n30891,
         n30892, n30893, n30894, n30895, n30896, n30897, n30898, n30899,
         n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907,
         n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915,
         n30916, n30917, n30918, n30919, n30920, n30921, n30922, n30923,
         n30924, n30925, n30926, n30927, n30928, n30929, n30930, n30931,
         n30932, n30933, n30934, n30935, n30936, n30937, n30938, n30939,
         n30940, n30941, n30942, n30943, n30944, n30945, n30946, n30947,
         n30948, n30949, n30950, n30951, n30952, n30953, n30954, n30955,
         n30956, n30957, n30958, n30959, n30960, n30961, n30962, n30963,
         n30964, n30965, n30966, n30967, n30968, n30969, n30970, n30971,
         n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979,
         n30980, n30981, n30982, n30983, n30984, n30985, n30986, n30987,
         n30988, n30989, n30990, n30991, n30992, n30993, n30994, n30995,
         n30996, n30997, n30998, n30999, n31000, n31001, n31002, n31003,
         n31004, n31005, n31006, n31007, n31008, n31009, n31010, n31011,
         n31012, n31013, n31014, n31015, n31016, n31017, n31018, n31019,
         n31020, n31021, n31022, n31023, n31024, n31025, n31026, n31027,
         n31028, n31029, n31030, n31031, n31032, n31033, n31034, n31035,
         n31036, n31037, n31038, n31039, n31040, n31041, n31042, n31043,
         n31044, n31045, n31046, n31047, n31048, n31049, n31050, n31051,
         n31052, n31053, n31054, n31055, n31056, n31057, n31058, n31059,
         n31060, n31061, n31062, n31063, n31064, n31065, n31066, n31067,
         n31068, n31069, n31070, n31071, n31072, n31073, n31074, n31075,
         n31076, n31077, n31078, n31079, n31080, n31081, n31082, n31083,
         n31084, n31085, n31086, n31087, n31088, n31089, n31090, n31091,
         n31092, n31093, n31094, n31095, n31096, n31097, n31098, n31099,
         n31100, n31101, n31102, n31103, n31104, n31105, n31106, n31107,
         n31108, n31109, n31110, n31111, n31112, n31113, n31114, n31115,
         n31116, n31117, n31118, n31119, n31120, n31121, n31122, n31123,
         n31124, n31125, n31126, n31127, n31128, n31129, n31130, n31131,
         n31132, n31133, n31134, n31135, n31136, n31137, n31138, n31139,
         n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147,
         n31148, n31149, n31150, n31151, n31152, n31153, n31154, n31155,
         n31156, n31157, n31158, n31159, n31160, n31161, n31162, n31163,
         n31164, n31165, n31166, n31167, n31168, n31169, n31170, n31171,
         n31172, n31173, n31174, n31175, n31176, n31177, n31178, n31179,
         n31180, n31181, n31182, n31183, n31184, n31185, n31186, n31187,
         n31188, n31189, n31190, n31191, n31192, n31193, n31194, n31195,
         n31196, n31197, n31198, n31199, n31200, n31201, n31202, n31203,
         n31204, n31205, n31206, n31207, n31208, n31209, n31210, n31211,
         n31212, n31213, n31214, n31215, n31216, n31217, n31218, n31219,
         n31220, n31221, n31222, n31223, n31224, n31225, n31226, n31227,
         n31228, n31229, n31230, n31231, n31232, n31233, n31234, n31235,
         n31236, n31237, n31238, n31239, n31240, n31241, n31242, n31243,
         n31244, n31245, n31246, n31247, n31248, n31249, n31250, n31251,
         n31252, n31253, n31254, n31255, n31256, n31257, n31258, n31259,
         n31260, n31261, n31262, n31263, n31264, n31265, n31266, n31267,
         n31268, n31269, n31270, n31271, n31272, n31273, n31274, n31275,
         n31276, n31277, n31278, n31279, n31280, n31281, n31282, n31283,
         n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291,
         n31292, n31293, n31294, n31295, n31296, n31297, n31298, n31299,
         n31300, n31301, n31302, n31303, n31304, n31305, n31306, n31307,
         n31308, n31309, n31310, n31311, n31312, n31313, n31314, n31315,
         n31316, n31317, n31318, n31319, n31320, n31321, n31322, n31323,
         n31324, n31325, n31326, n31327, n31328, n31329, n31330, n31331,
         n31332, n31333, n31334, n31335, n31336, n31337, n31338, n31339,
         n31340, n31341, n31342, n31343, n31344, n31345, n31346, n31347,
         n31348, n31349, n31350, n31351, n31352, n31353, n31354, n31355,
         n31356, n31357, n31358, n31359, n31360, n31361, n31362, n31363,
         n31364, n31365, n31366, n31367, n31368, n31369, n31370, n31371,
         n31372, n31373, n31374, n31375, n31376, n31377, n31378, n31379,
         n31380, n31381, n31382, n31383, n31384, n31385, n31386, n31387,
         n31388, n31389, n31390, n31391, n31392, n31393, n31394, n31395,
         n31396, n31397, n31398, n31399, n31400, n31401, n31402, n31403,
         n31404, n31405, n31406, n31407, n31408, n31409, n31410, n31411,
         n31412, n31413, n31414, n31415, n31416, n31417, n31418, n31419,
         n31420, n31421, n31422, n31423, n31424, n31425, n31426, n31427,
         n31428, n31429, n31430, n31431, n31432, n31433, n31434, n31435,
         n31436, n31437, n31438, n31439, n31440, n31441, n31442, n31443,
         n31444, n31445, n31446, n31447, n31448, n31449, n31450, n31451,
         n31452, n31453, n31454, n31455, n31456, n31457, n31458, n31459,
         n31460, n31461, n31462, n31463, n31464, n31465, n31466, n31467,
         n31468, n31469, n31470, n31471, n31472, n31473, n31474, n31475,
         n31476, n31477, n31478, n31479, n31480, n31481, n31482, n31483,
         n31484, n31485, n31486, n31487, n31488, n31489, n31490, n31491,
         n31492, n31493, n31494, n31495, n31496, n31497, n31498, n31499,
         n31500, n31501, n31502, n31503, n31504, n31505, n31506, n31507,
         n31508, n31509, n31510, n31511, n31512, n31513, n31514, n31515,
         n31516, n31517, n31518, n31519, n31520, n31521, n31522, n31523,
         n31524, n31525, n31526, n31527, n31528, n31529, n31530, n31531,
         n31532, n31533, n31534, n31535, n31536, n31537, n31538, n31539,
         n31540, n31541, n31542, n31543, n31544, n31545, n31546, n31547,
         n31548, n31549, n31550, n31551, n31552, n31553, n31554, n31555,
         n31556, n31557, n31558, n31559, n31560, n31561, n31562, n31563,
         n31564, n31565, n31566, n31567, n31568, n31569, n31570, n31571,
         n31572, n31573, n31574, n31575, n31576, n31577, n31578, n31579,
         n31580, n31581, n31582, n31583, n31584, n31585, n31586, n31587,
         n31588, n31589, n31590, n31591, n31592, n31593, n31594, n31595,
         n31596, n31597, n31598, n31599, n31600, n31601, n31602, n31603,
         n31604, n31605, n31606, n31607, n31608, n31609, n31610, n31611,
         n31612, n31613, n31614, n31615, n31616, n31617, n31618, n31619,
         n31620, n31621, n31622, n31623, n31624, n31625, n31626, n31627,
         n31628, n31629, n31630, n31631, n31632, n31633, n31634, n31635,
         n31636, n31637, n31638, n31639, n31640, n31641, n31642, n31643,
         n31644, n31645, n31646, n31647, n31648, n31649, n31650, n31651,
         n31652, n31653, n31654, n31655, n31656, n31657, n31658, n31659,
         n31660, n31661, n31662, n31663, n31664, n31665, n31666, n31667,
         n31668, n31669, n31670, n31671, n31672, n31673, n31674, n31675,
         n31676, n31677, n31678, n31679, n31680, n31681, n31682, n31683,
         n31684, n31685, n31686, n31687, n31688, n31689, n31690, n31691,
         n31692, n31693, n31694, n31695, n31696, n31697, n31698, n31699,
         n31700, n31701, n31702, n31703, n31704, n31705, n31706, n31707,
         n31708, n31709, n31710, n31711, n31712, n31713, n31714, n31715,
         n31716, n31717, n31718, n31719, n31720, n31721, n31722, n31723,
         n31724, n31725, n31726, n31727, n31728, n31729, n31730, n31731,
         n31732, n31733, n31734, n31735, n31736, n31737, n31738, n31739,
         n31740, n31741, n31742, n31743, n31744, n31745, n31746, n31747,
         n31748, n31749, n31750, n31751, n31752, n31753, n31754, n31755,
         n31756, n31757, n31758, n31759, n31760, n31761, n31762, n31763,
         n31764, n31765, n31766, n31767, n31768, n31769, n31770, n31771,
         n31772, n31773, n31774, n31775, n31776, n31777, n31778, n31779,
         n31780, n31781, n31782, n31783, n31784, n31785, n31786, n31787,
         n31788, n31789, n31790, n31791, n31792, n31793, n31794, n31795,
         n31796, n31797, n31798, n31799, n31800, n31801, n31802, n31803,
         n31804, n31805, n31806, n31807, n31808, n31809, n31810, n31811,
         n31812, n31813, n31814, n31815, n31816, n31817, n31818, n31819,
         n31820, n31821, n31822, n31823, n31824, n31825, n31826, n31827,
         n31828, n31829, n31830, n31831, n31832, n31833, n31834, n31835,
         n31836, n31837, n31838, n31839, n31840, n31841, n31842, n31843,
         n31844, n31845, n31846, n31847, n31848, n31849, n31850, n31851,
         n31852, n31853, n31854, n31855, n31856, n31857, n31858, n31859,
         n31860, n31861, n31862, n31863, n31864, n31865, n31866, n31867,
         n31868, n31869, n31870, n31871, n31872, n31873, n31874, n31875,
         n31876, n31877, n31878, n31879, n31880, n31881, n31882, n31883,
         n31884, n31885, n31886, n31887, n31888, n31889, n31890, n31891,
         n31892, n31893, n31894, n31895, n31896, n31897, n31898, n31899,
         n31900, n31901, n31902, n31903, n31904, n31905, n31906, n31907,
         n31908, n31909, n31910, n31911, n31912, n31913, n31914, n31915,
         n31916, n31917, n31918, n31919, n31920, n31921, n31922, n31923,
         n31924, n31925, n31926, n31927, n31928, n31929, n31930, n31931,
         n31932, n31933, n31934, n31935, n31936, n31937, n31938, n31939,
         n31940, n31941, n31942, n31943, n31944, n31945, n31946, n31947,
         n31948, n31949, n31950, n31951, n31952, n31953, n31954, n31955,
         n31956, n31957, n31958, n31959, n31960, n31961, n31962, n31963,
         n31964, n31965, n31966, n31967, n31968, n31969, n31970, n31971,
         n31972, n31973, n31974, n31975, n31976, n31977, n31978, n31979,
         n31980, n31981, n31982, n31983, n31984, n31985, n31986, n31987,
         n31988, n31989, n31990, n31991, n31992, n31993, n31994, n31995,
         n31996, n31997, n31998, n31999, n32000, n32001, n32002, n32003,
         n32004, n32005, n32006, n32007, n32008, n32009, n32010, n32011,
         n32012, n32013, n32014, n32015, n32016, n32017, n32018, n32019,
         n32020, n32021, n32022, n32023, n32024, n32025, n32026, n32027,
         n32028, n32029, n32030, n32031, n32032, n32033, n32034, n32035,
         n32036, n32037, n32038, n32039, n32040, n32041, n32042, n32043,
         n32044, n32045, n32046, n32047, n32048, n32049, n32050, n32051,
         n32052, n32053, n32054, n32055, n32056, n32057, n32058, n32059,
         n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067,
         n32068, n32069, n32070, n32071, n32072, n32073, n32074, n32075,
         n32076, n32077, n32078, n32079, n32080, n32081, n32082, n32083,
         n32084, n32085, n32086, n32087, n32088, n32089, n32090, n32091,
         n32092, n32093, n32094, n32095, n32096, n32097, n32098, n32099,
         n32100, n32101, n32102, n32103, n32104, n32105, n32106, n32107,
         n32108, n32109, n32110, n32111, n32112, n32113, n32114, n32115,
         n32116, n32117, n32118, n32119, n32120, n32121, n32122, n32123,
         n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131,
         n32132, n32133, n32134, n32135, n32136, n32137, n32138, n32139,
         n32140, n32141, n32142, n32143, n32144, n32145, n32146, n32147,
         n32148, n32149, n32150, n32151, n32152, n32153, n32154, n32155,
         n32156, n32157, n32158, n32159, n32160, n32161, n32162, n32163,
         n32164, n32165, n32166, n32167, n32168, n32169, n32170, n32171,
         n32172, n32173, n32174, n32175, n32176, n32177, n32178, n32179,
         n32180, n32181, n32182, n32183, n32184, n32185, n32186, n32187,
         n32188, n32189, n32190, n32191, n32192, n32193, n32194, n32195,
         n32196, n32197, n32198, n32199, n32200, n32201, n32202, n32203,
         n32204, n32205, n32206, n32207, n32208, n32209, n32210, n32211,
         n32212, n32213, n32214, n32215, n32216, n32217, n32218, n32219,
         n32220, n32221, n32222, n32223, n32224, n32225, n32226, n32227,
         n32228, n32229, n32230, n32231, n32232, n32233, n32234, n32235,
         n32236, n32237, n32238, n32239, n32240, n32241, n32242, n32243,
         n32244, n32245, n32246, n32247, n32248, n32249, n32250, n32251,
         n32252, n32253, n32254, n32255, n32256, n32257, n32258, n32259,
         n32260, n32261, n32262, n32263, n32264, n32265, n32266, n32267,
         n32268, n32269, n32270, n32271, n32272, n32273, n32274, n32275,
         n32276, n32277, n32278, n32279, n32280, n32281, n32282, n32283,
         n32284, n32285, n32286, n32287, n32288, n32289, n32290, n32291,
         n32292, n32293, n32294, n32295, n32296, n32297, n32298, n32299,
         n32300, n32301, n32302, n32303, n32304, n32305, n32306, n32307,
         n32308, n32309, n32310, n32311, n32312, n32313, n32314, n32315,
         n32316, n32317, n32318, n32319, n32320, n32321, n32322, n32323,
         n32324, n32325, n32326, n32327, n32328, n32329, n32330, n32331,
         n32332, n32333, n32334, n32335, n32336, n32337, n32338, n32339,
         n32340, n32341, n32342, n32343, n32344, n32345, n32346, n32347,
         n32348, n32349, n32350, n32351, n32352, n32353, n32354, n32355,
         n32356, n32357, n32358, n32359, n32360, n32361, n32362, n32363,
         n32364, n32365, n32366, n32367, n32368, n32369, n32370, n32371,
         n32372, n32373, n32374, n32375, n32376, n32377, n32378, n32379,
         n32380, n32381, n32382, n32383, n32384, n32385, n32386, n32387,
         n32388, n32389, n32390, n32391, n32392, n32393, n32394, n32395,
         n32396, n32397, n32398, n32399, n32400, n32401, n32402, n32403,
         n32404, n32405, n32406, n32407, n32408, n32409, n32410, n32411,
         n32412, n32413, n32414, n32415, n32416, n32417, n32418, n32419,
         n32420, n32421, n32422, n32423, n32424, n32425, n32426, n32427,
         n32428, n32429, n32430, n32431, n32432, n32433, n32434, n32435,
         n32436, n32437, n32438, n32439, n32440, n32441, n32442, n32443,
         n32444, n32445, n32446, n32447, n32448, n32449, n32450, n32451,
         n32452, n32453, n32454, n32455, n32456, n32457, n32458, n32459,
         n32460, n32461, n32462, n32463, n32464, n32465, n32466, n32467,
         n32468, n32469, n32470, n32471, n32472, n32473, n32474, n32475,
         n32476, n32477, n32478, n32479, n32480, n32481, n32482, n32483,
         n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491,
         n32492, n32493, n32494, n32495, n32496, n32497, n32498, n32499,
         n32500, n32501, n32502, n32503, n32504, n32505, n32506, n32507,
         n32508, n32509, n32510, n32511, n32512, n32513, n32514, n32515,
         n32516, n32517, n32518, n32519, n32520, n32521, n32522, n32523,
         n32524, n32525, n32526, n32527, n32528, n32529, n32530, n32531,
         n32532, n32533, n32534, n32535, n32536, n32537, n32538, n32539,
         n32540, n32541, n32542, n32543, n32544, n32545, n32546, n32547,
         n32548, n32549, n32550, n32551, n32552, n32553, n32554, n32555,
         n32556, n32557, n32558, n32559, n32560, n32561, n32562, n32563,
         n32564, n32565, n32566, n32567, n32568, n32569, n32570, n32571,
         n32572, n32573, n32574, n32575, n32576, n32577, n32578, n32579,
         n32580, n32581, n32582, n32583, n32584, n32585, n32586, n32587,
         n32588, n32589, n32590, n32591, n32592, n32593, n32594, n32595,
         n32596, n32597, n32598, n32599, n32600, n32601, n32602, n32603,
         n32604, n32605, n32606, n32607, n32608, n32609, n32610, n32611,
         n32612, n32613, n32614, n32615, n32616, n32617, n32618, n32619,
         n32620, n32621, n32622, n32623, n32624, n32625, n32626, n32627,
         n32628, n32629, n32630, n32631, n32632, n32633, n32634, n32635,
         n32636, n32637, n32638, n32639, n32640, n32641, n32642, n32643,
         n32644, n32645, n32646, n32647, n32648, n32649, n32650, n32651,
         n32652, n32653, n32654, n32655, n32656, n32657, n32658, n32659,
         n32660, n32661, n32662, n32663, n32664, n32665, n32666, n32667,
         n32668, n32669, n32670, n32671, n32672, n32673, n32674, n32675,
         n32676, n32677, n32678, n32679, n32680, n32681, n32682, n32683,
         n32684, n32685, n32686, n32687, n32688, n32689, n32690, n32691,
         n32692, n32693, n32694, n32695, n32696, n32697, n32698, n32699,
         n32700, n32701, n32702, n32703, n32704, n32705, n32706, n32707,
         n32708, n32709, n32710, n32711, n32712, n32713, n32714, n32715,
         n32716, n32717, n32718, n32719, n32720, n32721, n32722, n32723,
         n32724, n32725, n32726, n32727, n32728, n32729, n32730, n32731,
         n32732, n32733, n32734, n32735, n32736, n32737, n32738, n32739,
         n32740, n32741, n32742, n32743, n32744, n32745, n32746, n32747,
         n32748, n32749, n32750, n32751, n32752, n32753, n32754, n32755,
         n32756, n32757, n32758, n32759, n32760, n32761, n32762, n32763,
         n32764, n32765, n32766, n32767, n32768, n32769, n32770, n32771,
         n32772, n32773, n32774, n32775, n32776, n32777, n32778, n32779,
         n32780, n32781, n32782, n32783, n32784, n32785, n32786, n32787,
         n32788, n32789, n32790, n32791, n32792, n32793, n32794, n32795,
         n32796, n32797, n32798, n32799, n32800, n32801, n32802, n32803,
         n32804, n32805, n32806, n32807, n32808, n32809, n32810, n32811,
         n32812, n32813, n32814, n32815, n32816, n32817, n32818, n32819,
         n32820, n32821, n32822, n32823, n32824, n32825, n32826, n32827,
         n32828, n32829, n32830, n32831, n32832, n32833, n32834, n32835,
         n32836, n32837, n32838, n32839, n32840, n32841, n32842, n32843,
         n32844, n32845, n32846, n32847, n32848, n32849, n32850, n32851,
         n32852, n32853, n32854, n32855, n32856, n32857, n32858, n32859,
         n32860, n32861, n32862, n32863, n32864, n32865, n32866, n32867,
         n32868, n32869, n32870, n32871, n32872, n32873, n32874, n32875,
         n32876, n32877, n32878, n32879, n32880, n32881, n32882, n32883,
         n32884, n32885, n32886, n32887, n32888, n32889, n32890, n32891,
         n32892, n32893, n32894, n32895, n32896, n32897, n32898, n32899,
         n32900, n32901, n32902, n32903, n32904, n32905, n32906, n32907,
         n32908, n32909, n32910, n32911, n32912, n32913, n32914, n32915,
         n32916, n32917, n32918, n32919, n32920, n32921, n32922, n32923,
         n32924, n32925, n32926, n32927, n32928, n32929, n32930, n32931,
         n32932, n32933, n32934, n32935, n32936, n32937, n32938, n32939,
         n32940, n32941, n32942, n32943, n32944, n32945, n32946, n32947,
         n32948, n32949, n32950, n32951, n32952, n32953, n32954, n32955,
         n32956, n32957, n32958, n32959, n32960, n32961, n32962, n32963,
         n32964, n32965, n32966, n32967, n32968, n32969, n32970, n32971,
         n32972, n32973, n32974, n32975, n32976, n32977, n32978, n32979,
         n32980, n32981, n32982, n32983, n32984, n32985, n32986, n32987,
         n32988, n32989, n32990, n32991, n32992, n32993, n32994, n32995,
         n32996, n32997, n32998, n32999, n33000, n33001, n33002, n33003,
         n33004, n33005, n33006, n33007, n33008, n33009, n33010, n33011,
         n33012, n33013, n33014, n33015, n33016, n33017, n33018, n33019,
         n33020, n33021, n33022, n33023, n33024, n33025, n33026, n33027,
         n33028, n33029, n33030, n33031, n33032, n33033, n33034, n33035,
         n33036, n33037, n33038, n33039, n33040, n33041, n33042, n33043,
         n33044, n33045, n33046, n33047, n33048, n33049, n33050, n33051,
         n33052, n33053, n33054, n33055, n33056, n33057, n33058, n33059,
         n33060, n33061, n33062, n33063, n33064, n33065, n33066, n33067,
         n33068, n33069, n33070, n33071, n33072, n33073, n33074, n33075,
         n33076, n33077, n33078, n33079, n33080, n33081, n33082, n33083,
         n33084, n33085, n33086, n33087, n33088, n33089, n33090, n33091,
         n33092, n33093, n33094, n33095, n33096, n33097, n33098, n33099,
         n33100, n33101, n33102, n33103, n33104, n33105, n33106, n33107,
         n33108, n33109, n33110, n33111, n33112, n33113, n33114, n33115,
         n33116, n33117, n33118, n33119, n33120, n33121, n33122, n33123,
         n33124, n33125, n33126, n33127, n33128, n33129, n33130, n33131,
         n33132, n33133, n33134, n33135, n33136, n33137, n33138, n33139,
         n33140, n33141, n33142, n33143, n33144, n33145, n33146, n33147,
         n33148, n33149, n33150, n33151, n33152, n33153, n33154, n33155,
         n33156, n33157, n33158, n33159, n33160, n33161, n33162, n33163,
         n33164, n33165, n33166, n33167, n33168, n33169, n33170, n33171,
         n33172, n33173, n33174, n33175, n33176, n33177, n33178, n33179,
         n33180, n33181, n33182, n33183, n33184, n33185, n33186, n33187,
         n33188, n33189, n33190, n33191, n33192, n33193, n33194, n33195,
         n33196, n33197, n33198, n33199, n33200, n33201, n33202, n33203,
         n33204, n33205, n33206, n33207, n33208, n33209, n33210, n33211,
         n33212, n33213, n33214, n33215, n33216, n33217, n33218, n33219,
         n33220, n33221, n33222, n33223, n33224, n33225, n33226, n33227,
         n33228, n33229, n33230, n33231, n33232, n33233, n33234, n33235,
         n33236, n33237, n33238, n33239, n33240, n33241, n33242, n33243,
         n33244, n33245, n33246, n33247, n33248, n33249, n33250, n33251,
         n33252, n33253, n33254, n33255, n33256, n33257, n33258, n33259,
         n33260, n33261, n33262, n33263, n33264, n33265, n33266, n33267,
         n33268, n33269, n33270, n33271, n33272, n33273, n33274, n33275,
         n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283,
         n33284, n33285, n33286, n33287, n33288, n33289, n33290, n33291,
         n33292, n33293, n33294, n33295, n33296, n33297, n33298, n33299,
         n33300, n33301, n33302, n33303, n33304, n33305, n33306, n33307,
         n33308, n33309, n33310, n33311, n33312, n33313, n33314, n33315,
         n33316, n33317, n33318, n33319, n33320, n33321, n33322, n33323,
         n33324, n33325, n33326, n33327, n33328, n33329, n33330, n33331,
         n33332, n33333, n33334, n33335, n33336, n33337, n33338, n33339,
         n33340, n33341, n33342, n33343, n33344, n33345, n33346, n33347,
         n33348, n33349, n33350, n33351, n33352, n33353, n33354, n33355,
         n33356, n33357, n33358, n33359, n33360, n33361, n33362, n33363,
         n33364, n33365, n33366, n33367, n33368, n33369, n33370, n33371,
         n33372, n33373, n33374, n33375, n33376, n33377, n33378, n33379,
         n33380, n33381, n33382, n33383, n33384, n33385, n33386, n33387,
         n33388, n33389, n33390, n33391, n33392, n33393, n33394, n33395,
         n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403,
         n33404, n33405, n33406, n33407, n33408, n33409, n33410, n33411,
         n33412, n33413, n33414, n33415, n33416, n33417, n33418, n33419,
         n33420, n33421, n33422, n33423, n33424, n33425, n33426, n33427,
         n33428, n33429, n33430, n33431, n33432, n33433, n33434, n33435,
         n33436, n33437, n33438, n33439, n33440, n33441, n33442, n33443,
         n33444, n33445, n33446, n33447, n33448, n33449, n33450, n33451,
         n33452, n33453, n33454, n33455, n33456, n33457, n33458, n33459,
         n33460, n33461, n33462, n33463, n33464, n33465, n33466, n33467,
         n33468, n33469, n33470, n33471, n33472, n33473, n33474, n33475,
         n33476, n33477, n33478, n33479, n33480, n33481, n33482, n33483,
         n33484, n33485, n33486, n33487, n33488, n33489, n33490, n33491,
         n33492, n33493, n33494, n33495, n33496, n33497, n33498, n33499,
         n33500, n33501, n33502, n33503, n33504, n33505, n33506, n33507,
         n33508, n33509, n33510, n33511, n33512, n33513, n33514, n33515,
         n33516, n33517, n33518, n33519, n33520, n33521, n33522, n33523,
         n33524, n33525, n33526, n33527, n33528, n33529, n33530, n33531,
         n33532, n33533, n33534, n33535, n33536, n33537, n33538, n33539,
         n33540, n33541, n33542, n33543, n33544, n33545, n33546, n33547,
         n33548, n33549, n33550, n33551, n33552, n33553, n33554, n33555,
         n33556, n33557, n33558, n33559, n33560, n33561, n33562, n33563,
         n33564, n33565, n33566, n33567, n33568, n33569, n33570, n33571,
         n33572, n33573, n33574, n33575, n33576, n33577, n33578, n33579,
         n33580, n33581, n33582, n33583, n33584, n33585, n33586, n33587,
         n33588, n33589, n33590, n33591, n33592, n33593, n33594, n33595,
         n33596, n33597, n33598, n33599, n33600, n33601, n33602, n33603,
         n33604, n33605, n33606, n33607, n33608, n33609, n33610, n33611,
         n33612, n33613, n33614, n33615, n33616, n33617, n33618, n33619,
         n33620, n33621, n33622, n33623, n33624, n33625, n33626, n33627,
         n33628, n33629, n33630, n33631, n33632, n33633, n33634, n33635,
         n33636, n33637, n33638, n33639, n33640, n33641, n33642, n33643,
         n33644, n33645, n33646, n33647, n33648, n33649, n33650, n33651,
         n33652, n33653, n33654, n33655, n33656, n33657, n33658, n33659,
         n33660, n33661, n33662, n33663, n33664, n33665, n33666, n33667,
         n33668, n33669, n33670, n33671, n33672, n33673, n33674, n33675,
         n33676, n33677, n33678, n33679, n33680, n33681, n33682, n33683,
         n33684, n33685, n33686, n33687, n33688, n33689, n33690, n33691,
         n33692, n33693, n33694, n33695, n33696, n33697, n33698, n33699,
         n33700, n33701, n33702, n33703, n33704, n33705, n33706, n33707,
         n33708, n33709, n33710, n33711, n33712, n33713, n33714, n33715,
         n33716, n33717, n33718, n33719, n33720, n33721, n33722, n33723,
         n33724, n33725, n33726, n33727, n33728, n33729, n33730, n33731,
         n33732, n33733, n33734, n33735, n33736, n33737, n33738, n33739,
         n33740, n33741, n33742, n33743, n33744, n33745, n33746, n33747,
         n33748, n33749, n33750, n33751, n33752, n33753, n33754, n33755,
         n33756, n33757, n33758, n33759, n33760, n33761, n33762, n33763,
         n33764, n33765, n33766, n33767, n33768, n33769, n33770, n33771,
         n33772, n33773, n33774, n33775, n33776, n33777, n33778, n33779,
         n33780, n33781, n33782, n33783, n33784, n33785, n33786, n33787,
         n33788, n33789, n33790, n33791, n33792, n33793, n33794, n33795,
         n33796, n33797, n33798, n33799, n33800, n33801, n33802, n33803,
         n33804, n33805, n33806, n33807, n33808, n33809, n33810, n33811,
         n33812, n33813, n33814, n33815, n33816, n33817, n33818, n33819,
         n33820, n33821, n33822, n33823, n33824, n33825, n33826, n33827,
         n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835,
         n33836, n33837, n33838, n33839, n33840, n33841, n33842, n33843,
         n33844, n33845, n33846, n33847, n33848, n33849, n33850, n33851,
         n33852, n33853, n33854, n33855, n33856, n33857, n33858, n33859,
         n33860, n33861, n33862, n33863, n33864, n33865, n33866, n33867,
         n33868, n33869, n33870, n33871, n33872, n33873, n33874, n33875,
         n33876, n33877, n33878, n33879, n33880, n33881, n33882, n33883,
         n33884, n33885, n33886, n33887, n33888, n33889, n33890, n33891,
         n33892, n33893, n33894, n33895, n33896, n33897, n33898, n33899,
         n33900, n33901, n33902, n33903, n33904, n33905, n33906, n33907,
         n33908, n33909, n33910, n33911, n33912, n33913, n33914, n33915,
         n33916, n33917, n33918, n33919, n33920, n33921, n33922, n33923,
         n33924, n33925, n33926, n33927, n33928, n33929, n33930, n33931,
         n33932, n33933, n33934, n33935, n33936, n33937, n33938, n33939,
         n33940, n33941, n33942, n33943, n33944, n33945, n33946, n33947,
         n33948, n33949, n33950, n33951, n33952, n33953, n33954, n33955,
         n33956, n33957, n33958, n33959, n33960, n33961, n33962, n33963,
         n33964, n33965, n33966, n33967, n33968, n33969, n33970, n33971,
         n33972, n33973, n33974, n33975, n33976, n33977, n33978, n33979,
         n33980, n33981, n33982, n33983, n33984, n33985, n33986, n33987,
         n33988, n33989, n33990, n33991, n33992, n33993, n33994, n33995,
         n33996, n33997, n33998, n33999, n34000, n34001, n34002, n34003,
         n34004, n34005, n34006, n34007, n34008, n34009, n34010, n34011,
         n34012, n34013, n34014, n34015, n34016, n34017, n34018, n34019,
         n34020, n34021, n34022, n34023, n34024, n34025, n34026, n34027,
         n34028, n34029, n34030, n34031, n34032, n34033, n34034, n34035,
         n34036, n34037, n34038, n34039, n34040, n34041, n34042, n34043,
         n34044, n34045, n34046, n34047, n34048, n34049, n34050, n34051,
         n34052, n34053, n34054, n34055, n34056, n34057, n34058, n34059,
         n34060, n34061, n34062, n34063, n34064, n34065, n34066, n34067,
         n34068, n34069, n34070, n34071, n34072, n34073, n34074, n34075,
         n34076, n34077, n34078, n34079, n34080, n34081, n34082, n34083,
         n34084, n34085, n34086, n34087, n34088, n34089, n34090, n34091,
         n34092, n34093, n34094, n34095, n34096, n34097, n34098, n34099,
         n34100, n34101, n34102, n34103, n34104, n34105, n34106, n34107,
         n34108, n34109, n34110, n34111, n34112, n34113, n34114, n34115,
         n34116, n34117, n34118, n34119, n34120, n34121, n34122, n34123,
         n34124, n34125, n34126, n34127, n34128, n34129, n34130, n34131,
         n34132, n34133, n34134, n34135, n34136, n34137, n34138, n34139,
         n34140, n34141, n34142, n34143, n34144, n34145, n34146, n34147,
         n34148, n34149, n34150, n34151, n34152, n34153, n34154, n34155,
         n34156, n34157, n34158, n34159, n34160, n34161, n34162, n34163,
         n34164, n34165, n34166, n34167, n34168, n34169, n34170, n34171,
         n34172, n34173, n34174, n34175, n34176, n34177, n34178, n34179,
         n34180, n34181, n34182, n34183, n34184, n34185, n34186, n34187,
         n34188, n34189, n34190, n34191, n34192, n34193, n34194, n34195,
         n34196, n34197, n34198, n34199, n34200, n34201, n34202, n34203,
         n34204, n34205, n34206, n34207, n34208, n34209, n34210, n34211,
         n34212, n34213, n34214, n34215, n34216, n34217, n34218, n34219,
         n34220, n34221, n34222, n34223, n34224, n34225, n34226, n34227,
         n34228, n34229, n34230, n34231, n34232, n34233, n34234, n34235,
         n34236, n34237, n34238, n34239, n34240, n34241, n34242, n34243,
         n34244, n34245, n34246, n34247, n34248, n34249, n34250, n34251,
         n34252, n34253, n34254, n34255, n34256, n34257, n34258, n34259,
         n34260, n34261, n34262, n34263, n34264, n34265, n34266, n34267,
         n34268, n34269, n34270, n34271, n34272, n34273, n34274, n34275,
         n34276, n34277, n34278, n34279, n34280, n34281, n34282, n34283,
         n34284, n34285, n34286, n34287, n34288, n34289, n34290, n34291,
         n34292, n34293, n34294, n34295, n34296, n34297, n34298, n34299,
         n34300, n34301, n34302, n34303, n34304, n34305, n34306, n34307,
         n34308, n34309, n34310, n34311, n34312, n34313, n34314, n34315,
         n34316, n34317, n34318, n34319, n34320, n34321, n34322, n34323,
         n34324, n34325, n34326, n34327, n34328, n34329, n34330, n34331,
         n34332, n34333, n34334, n34335, n34336, n34337, n34338, n34339,
         n34340, n34341, n34342, n34343, n34344, n34345, n34346, n34347,
         n34348, n34349, n34350, n34351, n34352, n34353, n34354, n34355,
         n34356, n34357, n34358, n34359, n34360, n34361, n34362, n34363,
         n34364, n34365, n34366, n34367, n34368, n34369, n34370, n34371,
         n34372, n34373, n34374, n34375, n34376, n34377, n34378, n34379,
         n34380, n34381, n34382, n34383, n34384, n34385, n34386, n34387,
         n34388, n34389, n34390, n34391, n34392, n34393, n34394, n34395,
         n34396, n34397, n34398, n34399, n34400, n34401, n34402, n34403,
         n34404, n34405, n34406, n34407, n34408, n34409, n34410, n34411,
         n34412, n34413, n34414, n34415, n34416, n34417, n34418, n34419,
         n34420, n34421, n34422, n34423, n34424, n34425, n34426, n34427,
         n34428, n34429, n34430, n34431, n34432, n34433, n34434, n34435,
         n34436, n34437, n34438, n34439, n34440, n34441, n34442, n34443,
         n34444, n34445, n34446, n34447, n34448, n34449, n34450, n34451,
         n34452, n34453, n34454, n34455, n34456, n34457, n34458, n34459,
         n34460, n34461, n34462, n34463, n34464, n34465, n34466, n34467,
         n34468, n34469, n34470, n34471, n34472, n34473, n34474, n34475,
         n34476, n34477, n34478, n34479, n34480, n34481, n34482, n34483,
         n34484, n34485, n34486, n34487, n34488, n34489, n34490, n34491,
         n34492, n34493, n34494, n34495, n34496, n34497, n34498, n34499,
         n34500, n34501, n34502, n34503, n34504, n34505, n34506, n34507,
         n34508, n34509, n34510, n34511, n34512, n34513, n34514, n34515,
         n34516, n34517, n34518, n34519, n34520, n34521, n34522, n34523,
         n34524, n34525, n34526, n34527, n34528, n34529, n34530, n34531,
         n34532, n34533, n34534, n34535, n34536, n34537, n34538, n34539,
         n34540, n34541, n34542, n34543, n34544, n34545, n34546, n34547,
         n34548, n34549, n34550, n34551, n34552, n34553, n34554, n34555,
         n34556, n34557, n34558, n34559, n34560, n34561, n34562, n34563,
         n34564, n34565, n34566, n34567, n34568, n34569, n34570, n34571,
         n34572, n34573, n34574, n34575, n34576, n34577, n34578, n34579,
         n34580, n34581, n34582, n34583, n34584, n34585, n34586, n34587,
         n34588, n34589, n34590, n34591, n34592, n34593, n34594, n34595,
         n34596, n34597, n34598, n34599, n34600, n34601, n34602, n34603,
         n34604, n34605, n34606, n34607, n34608, n34609, n34610, n34611,
         n34612, n34613, n34614, n34615, n34616, n34617, n34618, n34619,
         n34620, n34621, n34622, n34623, n34624, n34625, n34626, n34627,
         n34628, n34629, n34630, n34631, n34632, n34633, n34634, n34635,
         n34636, n34637, n34638, n34639, n34640, n34641, n34642, n34643,
         n34644, n34645, n34646, n34647, n34648, n34649, n34650, n34651,
         n34652, n34653, n34654, n34655, n34656, n34657, n34658, n34659,
         n34660, n34661, n34662, n34663, n34664, n34665, n34666, n34667,
         n34668, n34669, n34670, n34671, n34672, n34673, n34674, n34675,
         n34676, n34677, n34678, n34679, n34680, n34681, n34682, n34683,
         n34684, n34685, n34686, n34687, n34688, n34689, n34690, n34691,
         n34692, n34693, n34694, n34695, n34696, n34697, n34698, n34699,
         n34700, n34701, n34702, n34703, n34704, n34705, n34706, n34707,
         n34708, n34709, n34710, n34711, n34712, n34713, n34714, n34715,
         n34716, n34717, n34718, n34719, n34720, n34721, n34722, n34723,
         n34724, n34725, n34726, n34727, n34728, n34729, n34730, n34731,
         n34732, n34733, n34734, n34735, n34736, n34737, n34738, n34739,
         n34740, n34741, n34742, n34743, n34744, n34745, n34746, n34747,
         n34748, n34749, n34750, n34751, n34752, n34753, n34754, n34755,
         n34756, n34757, n34758, n34759, n34760, n34761, n34762, n34763,
         n34764, n34765, n34766, n34767, n34768, n34769, n34770, n34771,
         n34772, n34773, n34774, n34775, n34776, n34777, n34778, n34779,
         n34780, n34781, n34782, n34783, n34784, n34785, n34786, n34787,
         n34788, n34789, n34790, n34791, n34792, n34793, n34794, n34795,
         n34796, n34797, n34798, n34799, n34800, n34801, n34802, n34803,
         n34804, n34805, n34806, n34807, n34808, n34809, n34810, n34811,
         n34812, n34813, n34814, n34815, n34816, n34817, n34818, n34819,
         n34820, n34821, n34822, n34823, n34824, n34825, n34826, n34827,
         n34828, n34829, n34830, n34831, n34832, n34833, n34834, n34835,
         n34836, n34837, n34838, n34839, n34840, n34841, n34842, n34843,
         n34844, n34845, n34846, n34847, n34848, n34849, n34850, n34851,
         n34852, n34853, n34854, n34855, n34856, n34857, n34858, n34859,
         n34860, n34861, n34862, n34863, n34864, n34865, n34866, n34867,
         n34868, n34869, n34870, n34871, n34872, n34873, n34874, n34875,
         n34876, n34877, n34878, n34879, n34880, n34881, n34882, n34883,
         n34884, n34885, n34886, n34887, n34888, n34889, n34890, n34891,
         n34892, n34893, n34894, n34895, n34896, n34897, n34898, n34899,
         n34900, n34901, n34902, n34903, n34904, n34905, n34906, n34907,
         n34908, n34909, n34910, n34911, n34912, n34913, n34914, n34915,
         n34916, n34917, n34918, n34919, n34920, n34921, n34922, n34923,
         n34924, n34925, n34926, n34927, n34928, n34929, n34930, n34931,
         n34932, n34933, n34934, n34935, n34936, n34937, n34938, n34939,
         n34940, n34941, n34942, n34943, n34944, n34945, n34946, n34947,
         n34948, n34949, n34950, n34951, n34952, n34953, n34954, n34955,
         n34956, n34957, n34958, n34959, n34960, n34961, n34962, n34963,
         n34964, n34965, n34966, n34967, n34968, n34969, n34970, n34971,
         n34972, n34973, n34974, n34975, n34976, n34977, n34978, n34979,
         n34980, n34981, n34982, n34983, n34984, n34985, n34986, n34987,
         n34988, n34989, n34990, n34991, n34992, n34993, n34994, n34995,
         n34996, n34997, n34998, n34999, n35000, n35001, n35002, n35003,
         n35004, n35005, n35006, n35007, n35008, n35009, n35010, n35011,
         n35012, n35013, n35014, n35015, n35016, n35017, n35018, n35019,
         n35020, n35021, n35022, n35023, n35024, n35025, n35026, n35027,
         n35028, n35029, n35030, n35031, n35032, n35033, n35034, n35035,
         n35036, n35037, n35038, n35039, n35040, n35041, n35042, n35043,
         n35044, n35045, n35046, n35047, n35048, n35049, n35050, n35051,
         n35052, n35053, n35054, n35055, n35056, n35057, n35058, n35059,
         n35060, n35061, n35062, n35063, n35064, n35065, n35066, n35067,
         n35068, n35069, n35070, n35071, n35072, n35073, n35074, n35075,
         n35076, n35077, n35078, n35079, n35080, n35081, n35082, n35083,
         n35084, n35085, n35086, n35087, n35088, n35089, n35090, n35091,
         n35092, n35093, n35094, n35095, n35096, n35097, n35098, n35099,
         n35100, n35101, n35102, n35103, n35104, n35105, n35106, n35107,
         n35108, n35109, n35110, n35111, n35112, n35113, n35114, n35115,
         n35116, n35117, n35118, n35119, n35120, n35121, n35122, n35123,
         n35124, n35125, n35126, n35127, n35128, n35129, n35130, n35131,
         n35132, n35133, n35134, n35135, n35136, n35137, n35138, n35139,
         n35140, n35141, n35142, n35143, n35144, n35145, n35146, n35147,
         n35148, n35149, n35150, n35151, n35152, n35153, n35154, n35155,
         n35156, n35157, n35158, n35159, n35160, n35161, n35162, n35163,
         n35164, n35165, n35166, n35167, n35168, n35169, n35170, n35171,
         n35172, n35173, n35174, n35175, n35176, n35177, n35178, n35179,
         n35180, n35181, n35182, n35183, n35184, n35185, n35186, n35187,
         n35188, n35189, n35190, n35191, n35192, n35193, n35194, n35195,
         n35196, n35197, n35198, n35199, n35200, n35201, n35202, n35203,
         n35204, n35205, n35206, n35207, n35208, n35209, n35210, n35211,
         n35212, n35213, n35214, n35215, n35216, n35217, n35218, n35219,
         n35220, n35221, n35222, n35223, n35224, n35225, n35226, n35227,
         n35228, n35229, n35230, n35231, n35232, n35233, n35234, n35235,
         n35236, n35237, n35238, n35239, n35240, n35241, n35242, n35243,
         n35244, n35245, n35246, n35247, n35248, n35249, n35250, n35251,
         n35252, n35253, n35254, n35255, n35256, n35257, n35258, n35259,
         n35260, n35261, n35262, n35263, n35264, n35265, n35266, n35267,
         n35268, n35269, n35270, n35271, n35272, n35273, n35274, n35275,
         n35276, n35277, n35278, n35279, n35280, n35281, n35282, n35283,
         n35284, n35285, n35286, n35287, n35288, n35289, n35290, n35291,
         n35292, n35293, n35294, n35295, n35296, n35297, n35298, n35299,
         n35300, n35301, n35302, n35303, n35304, n35305, n35306, n35307,
         n35308, n35309, n35310, n35311, n35312, n35313, n35314, n35315,
         n35316, n35317, n35318, n35319, n35320, n35321, n35322, n35323,
         n35324, n35325, n35326, n35327, n35328, n35329, n35330, n35331,
         n35332, n35333, n35334, n35335, n35336, n35337, n35338, n35339,
         n35340, n35341, n35342, n35343, n35344, n35345, n35346, n35347,
         n35348, n35349, n35350, n35351, n35352, n35353, n35354, n35355,
         n35356, n35357, n35358, n35359, n35360, n35361, n35362, n35363,
         n35364, n35365, n35366, n35367, n35368, n35369, n35370, n35371,
         n35372, n35373, n35374, n35375, n35376, n35377, n35378, n35379,
         n35380, n35381, n35382, n35383, n35384, n35385, n35386, n35387,
         n35388, n35389, n35390, n35391, n35392, n35393, n35394, n35395,
         n35396, n35397, n35398, n35399, n35400, n35401, n35402, n35403,
         n35404, n35405, n35406, n35407, n35408, n35409, n35410, n35411,
         n35412, n35413, n35414, n35415, n35416, n35417, n35418, n35419,
         n35420, n35421, n35422, n35423, n35424, n35425, n35426, n35427,
         n35428, n35429, n35430, n35431, n35432, n35433, n35434, n35435,
         n35436, n35437, n35438, n35439, n35440, n35441, n35442, n35443,
         n35444, n35445, n35446, n35447, n35448, n35449, n35450, n35451,
         n35452, n35453, n35454, n35455, n35456, n35457, n35458, n35459,
         n35460, n35461, n35462, n35463, n35464, n35465, n35466, n35467,
         n35468, n35469, n35470, n35471, n35472, n35473, n35474, n35475,
         n35476, n35477, n35478, n35479, n35480, n35481, n35482, n35483,
         n35484, n35485, n35486, n35487, n35488, n35489, n35490, n35491,
         n35492, n35493, n35494, n35495, n35496, n35497, n35498, n35499,
         n35500, n35501, n35502, n35503, n35504, n35505, n35506, n35507,
         n35508, n35509, n35510, n35511, n35512, n35513, n35514, n35515,
         n35516, n35517, n35518, n35519, n35520, n35521, n35522, n35523,
         n35524, n35525, n35526, n35527, n35528, n35529, n35530, n35531,
         n35532, n35533, n35534, n35535, n35536, n35537, n35538, n35539,
         n35540, n35541, n35542, n35543, n35544, n35545, n35546, n35547,
         n35548, n35549, n35550, n35551, n35552, n35553, n35554, n35555,
         n35556, n35557, n35558, n35559, n35560, n35561, n35562, n35563,
         n35564, n35565, n35566, n35567, n35568, n35569, n35570, n35571,
         n35572, n35573, n35574, n35575, n35576, n35577, n35578, n35579,
         n35580, n35581, n35582, n35583, n35584, n35585, n35586, n35587,
         n35588, n35589, n35590, n35591, n35592, n35593, n35594, n35595,
         n35596, n35597, n35598, n35599, n35600, n35601, n35602, n35603,
         n35604, n35605, n35606, n35607, n35608, n35609, n35610, n35611,
         n35612, n35613, n35614, n35615, n35616, n35617, n35618, n35619,
         n35620, n35621, n35622, n35623, n35624, n35625, n35626, n35627,
         n35628, n35629, n35630, n35631, n35632, n35633, n35634, n35635,
         n35636, n35637, n35638, n35639, n35640, n35641, n35642, n35643,
         n35644, n35645, n35646, n35647, n35648, n35649, n35650, n35651,
         n35652, n35653, n35654, n35655, n35656, n35657, n35658, n35659,
         n35660, n35661, n35662, n35663, n35664, n35665, n35666, n35667,
         n35668, n35669, n35670, n35671, n35672, n35673, n35674, n35675,
         n35676, n35677, n35678, n35679, n35680, n35681, n35682, n35683,
         n35684, n35685, n35686, n35687, n35688, n35689, n35690, n35691,
         n35692, n35693, n35694, n35695, n35696, n35697, n35698, n35699,
         n35700, n35701, n35702, n35703, n35704, n35705, n35706, n35707,
         n35708, n35709, n35710, n35711, n35712, n35713, n35714, n35715,
         n35716, n35717, n35718, n35719, n35720, n35721, n35722, n35723,
         n35724, n35725, n35726, n35727, n35728, n35729, n35730, n35731,
         n35732, n35733, n35734, n35735, n35736, n35737, n35738, n35739,
         n35740, n35741, n35742, n35743, n35744, n35745, n35746, n35747,
         n35748, n35749, n35750, n35751, n35752, n35753, n35754, n35755,
         n35756, n35757, n35758, n35759, n35760, n35761, n35762, n35763,
         n35764, n35765, n35766, n35767, n35768, n35769, n35770, n35771,
         n35772, n35773, n35774, n35775, n35776, n35777, n35778, n35779,
         n35780, n35781, n35782, n35783, n35784, n35785, n35786, n35787,
         n35788, n35789, n35790, n35791, n35792, n35793, n35794, n35795,
         n35796, n35797, n35798, n35799, n35800, n35801, n35802, n35803,
         n35804, n35805, n35806, n35807, n35808, n35809, n35810, n35811,
         n35812, n35813, n35814, n35815, n35816, n35817, n35818, n35819,
         n35820, n35821, n35822, n35823, n35824, n35825, n35826, n35827,
         n35828, n35829, n35830, n35831, n35832, n35833, n35834, n35835,
         n35836, n35837, n35838, n35839, n35840, n35841, n35842, n35843,
         n35844, n35845, n35846, n35847, n35848, n35849, n35850, n35851,
         n35852, n35853, n35854, n35855, n35856, n35857, n35858, n35859,
         n35860, n35861, n35862, n35863, n35864, n35865, n35866, n35867,
         n35868, n35869, n35870, n35871, n35872, n35873, n35874, n35875,
         n35876, n35877, n35878, n35879, n35880, n35881, n35882, n35883,
         n35884, n35885, n35886, n35887, n35888, n35889, n35890, n35891,
         n35892, n35893, n35894, n35895, n35896, n35897, n35898, n35899,
         n35900, n35901, n35902, n35903, n35904, n35905, n35906, n35907,
         n35908, n35909, n35910, n35911, n35912, n35913, n35914, n35915,
         n35916, n35917, n35918, n35919, n35920, n35921, n35922, n35923,
         n35924, n35925, n35926, n35927, n35928, n35929, n35930, n35931,
         n35932, n35933, n35934, n35935, n35936, n35937, n35938, n35939,
         n35940, n35941, n35942, n35943, n35944, n35945, n35946, n35947,
         n35948, n35949, n35950, n35951, n35952, n35953, n35954, n35955,
         n35956, n35957, n35958, n35959, n35960, n35961, n35962, n35963,
         n35964, n35965, n35966, n35967, n35968, n35969, n35970, n35971,
         n35972, n35973, n35974, n35975, n35976, n35977, n35978, n35979,
         n35980, n35981, n35982, n35983, n35984, n35985, n35986, n35987,
         n35988, n35989, n35990, n35991, n35992, n35993, n35994, n35995,
         n35996, n35997, n35998, n35999, n36000, n36001, n36002, n36003,
         n36004, n36005, n36006, n36007, n36008, n36009, n36010, n36011,
         n36012, n36013, n36014, n36015, n36016, n36017, n36018, n36019,
         n36020, n36021, n36022, n36023, n36024, n36025, n36026, n36027,
         n36028, n36029, n36030, n36031, n36032, n36033, n36034, n36035,
         n36036, n36037, n36038, n36039, n36040, n36041, n36042, n36043,
         n36044, n36045, n36046, n36047, n36048, n36049, n36050, n36051,
         n36052, n36053, n36054, n36055, n36056, n36057, n36058, n36059,
         n36060, n36061, n36062, n36063, n36064, n36065, n36066, n36067,
         n36068, n36069, n36070, n36071, n36072, n36073, n36074, n36075,
         n36076, n36077, n36078, n36079, n36080, n36081, n36082, n36083,
         n36084, n36085, n36086, n36087, n36088, n36089, n36090, n36091,
         n36092, n36093, n36094, n36095, n36096, n36097, n36098, n36099,
         n36100, n36101, n36102, n36103, n36104, n36105, n36106, n36107,
         n36108, n36109, n36110, n36111, n36112, n36113, n36114, n36115,
         n36116, n36117, n36118, n36119, n36120, n36121, n36122, n36123,
         n36124, n36125, n36126, n36127, n36128, n36129, n36130, n36131,
         n36132, n36133, n36134, n36135, n36136, n36137, n36138, n36139,
         n36140, n36141, n36142, n36143, n36144, n36145, n36146, n36147,
         n36148, n36149, n36150, n36151, n36152, n36153, n36154, n36155,
         n36156, n36157, n36158, n36159, n36160, n36161, n36162, n36163,
         n36164, n36165, n36166, n36167, n36168, n36169, n36170, n36171,
         n36172, n36173, n36174, n36175, n36176, n36177, n36178, n36179,
         n36180, n36181, n36182, n36183, n36184, n36185, n36186, n36187,
         n36188, n36189, n36190, n36191, n36192, n36193, n36194, n36195,
         n36196, n36197, n36198, n36199, n36200, n36201, n36202, n36203,
         n36204, n36205, n36206, n36207, n36208, n36209, n36210, n36211,
         n36212, n36213, n36214, n36215, n36216, n36217, n36218, n36219,
         n36220, n36221, n36222, n36223, n36224, n36225, n36226, n36227,
         n36228, n36229, n36230, n36231, n36232, n36233, n36234, n36235,
         n36236, n36237, n36238, n36239, n36240, n36241, n36242, n36243,
         n36244, n36245, n36246, n36247, n36248, n36249, n36250, n36251,
         n36252, n36253, n36254, n36255, n36256, n36257, n36258, n36259,
         n36260, n36261, n36262, n36263, n36264, n36265, n36266, n36267,
         n36268, n36269, n36270, n36271, n36272, n36273, n36274, n36275,
         n36276, n36277, n36278, n36279, n36280, n36281, n36282, n36283,
         n36284, n36285, n36286, n36287, n36288, n36289, n36290, n36291,
         n36292, n36293, n36294, n36295, n36296, n36297, n36298, n36299,
         n36300, n36301, n36302, n36303, n36304, n36305, n36306, n36307,
         n36308, n36309, n36310, n36311, n36312, n36313, n36314, n36315,
         n36316, n36317, n36318, n36319, n36320, n36321, n36322, n36323,
         n36324, n36325, n36326, n36327, n36328, n36329, n36330, n36331,
         n36332, n36333, n36334, n36335, n36336, n36337, n36338, n36339,
         n36340, n36341, n36342, n36343, n36344, n36345, n36346, n36347,
         n36348, n36349, n36350, n36351, n36352, n36353, n36354, n36355,
         n36356, n36357, n36358, n36359, n36360, n36361, n36362, n36363,
         n36364, n36365, n36366, n36367, n36368, n36369, n36370, n36371,
         n36372, n36373, n36374, n36375, n36376, n36377, n36378, n36379,
         n36380, n36381, n36382, n36383, n36384, n36385, n36386, n36387,
         n36388, n36389, n36390, n36391, n36392, n36393, n36394, n36395,
         n36396, n36397, n36398, n36399, n36400, n36401, n36402, n36403,
         n36404, n36405, n36406, n36407, n36408, n36409, n36410, n36411,
         n36412, n36413, n36414, n36415, n36416, n36417, n36418, n36419,
         n36420, n36421, n36422, n36423, n36424, n36425, n36426, n36427,
         n36428, n36429, n36430, n36431, n36432, n36433, n36434, n36435,
         n36436, n36437, n36438, n36439, n36440, n36441, n36442, n36443,
         n36444, n36445, n36446, n36447, n36448, n36449, n36450, n36451,
         n36452, n36453, n36454, n36455, n36456, n36457, n36458, n36459,
         n36460, n36461, n36462, n36463, n36464, n36465, n36466, n36467,
         n36468, n36469, n36470, n36471, n36472, n36473, n36474, n36475,
         n36476, n36477, n36478, n36479, n36480, n36481, n36482, n36483,
         n36484, n36485, n36486, n36487, n36488, n36489, n36490, n36491,
         n36492, n36493, n36494, n36495, n36496, n36497, n36498, n36499,
         n36500, n36501, n36502, n36503, n36504, n36505, n36506, n36507,
         n36508, n36509, n36510, n36511, n36512, n36513, n36514, n36515,
         n36516, n36517, n36518, n36519, n36520, n36521, n36522, n36523,
         n36524, n36525, n36526, n36527, n36528, n36529, n36530, n36531,
         n36532, n36533, n36534, n36535, n36536, n36537, n36538, n36539,
         n36540, n36541, n36542, n36543, n36544, n36545, n36546, n36547,
         n36548, n36549, n36550, n36551, n36552, n36553, n36554, n36555,
         n36556, n36557, n36558, n36559, n36560, n36561, n36562, n36563,
         n36564, n36565, n36566, n36567, n36568, n36569, n36570, n36571,
         n36572, n36573, n36574, n36575, n36576, n36577, n36578, n36579,
         n36580, n36581, n36582, n36583, n36584, n36585, n36586, n36587,
         n36588, n36589, n36590, n36591, n36592, n36593, n36594, n36595,
         n36596, n36597, n36598, n36599, n36600, n36601, n36602, n36603,
         n36604, n36605, n36606, n36607, n36608, n36609, n36610, n36611,
         n36612, n36613, n36614, n36615, n36616, n36617, n36618, n36619,
         n36620, n36621, n36622, n36623, n36624, n36625, n36626, n36627,
         n36628, n36629, n36630, n36631, n36632, n36633, n36634, n36635,
         n36636, n36637, n36638, n36639, n36640, n36641, n36642, n36643,
         n36644, n36645, n36646, n36647, n36648, n36649, n36650, n36651,
         n36652, n36653, n36654, n36655, n36656, n36657, n36658, n36659,
         n36660, n36661, n36662, n36663, n36664, n36665, n36666, n36667,
         n36668, n36669, n36670, n36671, n36672, n36673, n36674, n36675,
         n36676, n36677, n36678, n36679, n36680, n36681, n36682, n36683,
         n36684, n36685, n36686, n36687, n36688, n36689, n36690, n36691,
         n36692, n36693, n36694, n36695, n36696, n36697, n36698, n36699,
         n36700, n36701, n36702, n36703, n36704, n36705, n36706, n36707,
         n36708, n36709, n36710, n36711, n36712, n36713, n36714, n36715,
         n36716, n36717, n36718, n36719, n36720, n36721, n36722, n36723,
         n36724, n36725, n36726, n36727, n36728, n36729, n36730, n36731,
         n36732, n36733, n36734, n36735, n36736, n36737, n36738, n36739,
         n36740, n36741, n36742, n36743, n36744, n36745, n36746, n36747,
         n36748, n36749, n36750, n36751, n36752, n36753, n36754, n36755,
         n36756, n36757, n36758, n36759, n36760, n36761, n36762, n36763,
         n36764, n36765, n36766, n36767, n36768, n36769, n36770, n36771,
         n36772, n36773, n36774, n36775, n36776, n36777, n36778, n36779,
         n36780, n36781, n36782, n36783, n36784, n36785, n36786, n36787,
         n36788, n36789, n36790, n36791, n36792, n36793, n36794, n36795,
         n36796, n36797, n36798, n36799, n36800, n36801, n36802, n36803,
         n36804, n36805, n36806, n36807, n36808, n36809, n36810, n36811,
         n36812, n36813, n36814, n36815, n36816, n36817, n36818, n36819,
         n36820, n36821, n36822, n36823, n36824, n36825, n36826, n36827,
         n36828, n36829, n36830, n36831, n36832, n36833, n36834, n36835,
         n36836, n36837, n36838, n36839, n36840, n36841, n36842, n36843,
         n36844, n36845, n36846, n36847, n36848, n36849, n36850, n36851,
         n36852, n36853, n36854, n36855, n36856, n36857, n36858, n36859,
         n36860, n36861, n36862, n36863, n36864, n36865, n36866, n36867,
         n36868, n36869, n36870, n36871, n36872, n36873, n36874, n36875,
         n36876, n36877, n36878, n36879, n36880, n36881, n36882, n36883,
         n36884, n36885, n36886, n36887, n36888, n36889, n36890, n36891,
         n36892, n36893, n36894, n36895, n36896, n36897, n36898, n36899,
         n36900, n36901, n36902, n36903, n36904, n36905, n36906, n36907,
         n36908, n36909, n36910, n36911, n36912, n36913, n36914, n36915,
         n36916, n36917, n36918, n36919, n36920, n36921, n36922, n36923,
         n36924, n36925, n36926, n36927, n36928, n36929, n36930, n36931,
         n36932, n36933, n36934, n36935, n36936, n36937, n36938, n36939,
         n36940, n36941, n36942, n36943, n36944, n36945, n36946, n36947,
         n36948, n36949, n36950, n36951, n36952, n36953, n36954, n36955,
         n36956, n36957, n36958, n36959, n36960, n36961, n36962, n36963,
         n36964, n36965, n36966, n36967, n36968, n36969, n36970, n36971,
         n36972, n36973, n36974, n36975, n36976, n36977, n36978, n36979,
         n36980, n36981, n36982, n36983, n36984, n36985, n36986, n36987,
         n36988, n36989, n36990, n36991, n36992, n36993, n36994, n36995,
         n36996, n36997, n36998, n36999, n37000, n37001, n37002, n37003,
         n37004, n37005, n37006, n37007, n37008, n37009, n37010, n37011,
         n37012, n37013, n37014, n37015, n37016, n37017, n37018, n37019,
         n37020, n37021, n37022, n37023, n37024, n37025, n37026, n37027,
         n37028, n37029, n37030, n37031, n37032, n37033, n37034, n37035,
         n37036, n37037, n37038, n37039, n37040, n37041, n37042, n37043,
         n37044, n37045, n37046, n37047, n37048, n37049, n37050, n37051,
         n37052, n37053, n37054, n37055, n37056, n37057, n37058, n37059,
         n37060, n37061, n37062, n37063, n37064, n37065, n37066, n37067,
         n37068, n37069, n37070, n37071, n37072, n37073, n37074, n37075,
         n37076, n37077, n37078, n37079, n37080, n37081, n37082, n37083,
         n37084, n37085, n37086, n37087, n37088, n37089, n37090, n37091,
         n37092, n37093, n37094, n37095, n37096, n37097, n37098, n37099,
         n37100, n37101, n37102, n37103, n37104, n37105, n37106, n37107,
         n37108, n37109, n37110, n37111, n37112, n37113, n37114, n37115,
         n37116, n37117, n37118, n37119, n37120, n37121, n37122, n37123,
         n37124, n37125, n37126, n37127, n37128, n37129, n37130, n37131,
         n37132, n37133, n37134, n37135, n37136, n37137, n37138, n37139,
         n37140, n37141, n37142, n37143, n37144, n37145, n37146, n37147,
         n37148, n37149, n37150, n37151, n37152, n37153, n37154, n37155,
         n37156, n37157, n37158, n37159, n37160, n37161, n37162, n37163,
         n37164, n37165, n37166, n37167, n37168, n37169, n37170, n37171,
         n37172, n37173, n37174, n37175, n37176, n37177, n37178, n37179,
         n37180, n37181, n37182, n37183, n37184, n37185, n37186, n37187,
         n37188, n37189, n37190, n37191, n37192, n37193, n37194, n37195,
         n37196, n37197, n37198, n37199, n37200, n37201, n37202, n37203,
         n37204, n37205, n37206, n37207, n37208, n37209, n37210, n37211,
         n37212, n37213, n37214, n37215, n37216, n37217, n37218, n37219,
         n37220, n37221, n37222, n37223, n37224, n37225, n37226, n37227,
         n37228, n37229, n37230, n37231, n37232, n37233, n37234, n37235,
         n37236, n37237, n37238, n37239, n37240, n37241, n37242, n37243,
         n37244, n37245, n37246, n37247, n37248, n37249, n37250, n37251,
         n37252, n37253, n37254, n37255, n37256, n37257, n37258, n37259,
         n37260, n37261, n37262, n37263, n37264, n37265, n37266, n37267,
         n37268, n37269, n37270, n37271, n37272, n37273, n37274, n37275,
         n37276, n37277, n37278, n37279, n37280, n37281, n37282, n37283,
         n37284, n37285, n37286, n37287, n37288, n37289, n37290, n37291,
         n37292, n37293, n37294, n37295, n37296, n37297, n37298, n37299,
         n37300, n37301, n37302, n37303, n37304, n37305, n37306, n37307,
         n37308, n37309, n37310, n37311, n37312, n37313, n37314, n37315,
         n37316, n37317, n37318, n37319, n37320, n37321, n37322, n37323,
         n37324, n37325, n37326, n37327, n37328, n37329, n37330, n37331,
         n37332, n37333, n37334, n37335, n37336, n37337, n37338, n37339,
         n37340, n37341, n37342, n37343, n37344, n37345, n37346, n37347,
         n37348, n37349, n37350, n37351, n37352, n37353, n37354, n37355,
         n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363,
         n37364, n37365, n37366, n37367, n37368, n37369, n37370, n37371;
  assign \knn_comb_/min_val_out[0][0]  = p_input[2032];
  assign \knn_comb_/min_val_out[0][1]  = p_input[2033];
  assign \knn_comb_/min_val_out[0][2]  = p_input[2034];
  assign \knn_comb_/min_val_out[0][3]  = p_input[2035];
  assign \knn_comb_/min_val_out[0][4]  = p_input[2036];
  assign \knn_comb_/min_val_out[0][5]  = p_input[2037];
  assign \knn_comb_/min_val_out[0][6]  = p_input[2038];
  assign \knn_comb_/min_val_out[0][7]  = p_input[2039];
  assign \knn_comb_/min_val_out[0][8]  = p_input[2040];
  assign \knn_comb_/min_val_out[0][9]  = p_input[2041];
  assign \knn_comb_/min_val_out[0][10]  = p_input[2042];
  assign \knn_comb_/min_val_out[0][11]  = p_input[2043];
  assign \knn_comb_/min_val_out[0][12]  = p_input[2044];
  assign \knn_comb_/min_val_out[0][13]  = p_input[2045];
  assign \knn_comb_/min_val_out[0][14]  = p_input[2046];
  assign \knn_comb_/min_val_out[0][15]  = p_input[2047];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][0]  = p_input[2016];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][1]  = p_input[2017];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][2]  = p_input[2018];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][3]  = p_input[2019];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][4]  = p_input[2020];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][5]  = p_input[2021];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][6]  = p_input[2022];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][7]  = p_input[2023];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][8]  = p_input[2024];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][9]  = p_input[2025];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][10]  = p_input[2026];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][11]  = p_input[2027];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][12]  = p_input[2028];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][13]  = p_input[2029];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][14]  = p_input[2030];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][15]  = p_input[2031];

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  XOR U2 ( .A(n3), .B(n4), .Z(o[8]) );
  XOR U3 ( .A(n5), .B(n6), .Z(o[7]) );
  XOR U4 ( .A(n7), .B(n8), .Z(o[6]) );
  XOR U5 ( .A(n9), .B(n10), .Z(o[5]) );
  XOR U6 ( .A(n11), .B(n12), .Z(o[4]) );
  XOR U7 ( .A(n13), .B(n14), .Z(o[3]) );
  XOR U8 ( .A(n15), .B(n16), .Z(o[31]) );
  XOR U9 ( .A(n17), .B(n18), .Z(o[30]) );
  XOR U10 ( .A(n19), .B(n20), .Z(o[2]) );
  XOR U11 ( .A(n21), .B(n22), .Z(o[29]) );
  XOR U12 ( .A(n23), .B(n24), .Z(o[28]) );
  XOR U13 ( .A(n25), .B(n26), .Z(o[27]) );
  XOR U14 ( .A(n27), .B(n28), .Z(o[26]) );
  XOR U15 ( .A(n1), .B(n29), .Z(o[25]) );
  AND U16 ( .A(n30), .B(n31), .Z(n1) );
  XOR U17 ( .A(n2), .B(n29), .Z(n31) );
  XOR U18 ( .A(n32), .B(n33), .Z(n29) );
  AND U19 ( .A(n34), .B(n35), .Z(n33) );
  XOR U20 ( .A(p_input[9]), .B(n32), .Z(n35) );
  XOR U21 ( .A(n36), .B(n37), .Z(n32) );
  AND U22 ( .A(n38), .B(n39), .Z(n37) );
  XOR U23 ( .A(n40), .B(n41), .Z(n2) );
  AND U24 ( .A(n42), .B(n39), .Z(n41) );
  XNOR U25 ( .A(n43), .B(n36), .Z(n39) );
  XOR U26 ( .A(n44), .B(n45), .Z(n36) );
  AND U27 ( .A(n46), .B(n47), .Z(n45) );
  XOR U28 ( .A(p_input[25]), .B(n44), .Z(n47) );
  XOR U29 ( .A(n48), .B(n49), .Z(n44) );
  AND U30 ( .A(n50), .B(n51), .Z(n49) );
  IV U31 ( .A(n40), .Z(n43) );
  XNOR U32 ( .A(n52), .B(n53), .Z(n40) );
  AND U33 ( .A(n54), .B(n51), .Z(n53) );
  XNOR U34 ( .A(n52), .B(n48), .Z(n51) );
  XOR U35 ( .A(n55), .B(n56), .Z(n48) );
  AND U36 ( .A(n57), .B(n58), .Z(n56) );
  XOR U37 ( .A(p_input[41]), .B(n55), .Z(n58) );
  XOR U38 ( .A(n59), .B(n60), .Z(n55) );
  AND U39 ( .A(n61), .B(n62), .Z(n60) );
  XOR U40 ( .A(n63), .B(n64), .Z(n52) );
  AND U41 ( .A(n65), .B(n62), .Z(n64) );
  XNOR U42 ( .A(n63), .B(n59), .Z(n62) );
  XOR U43 ( .A(n66), .B(n67), .Z(n59) );
  AND U44 ( .A(n68), .B(n69), .Z(n67) );
  XOR U45 ( .A(p_input[57]), .B(n66), .Z(n69) );
  XOR U46 ( .A(n70), .B(n71), .Z(n66) );
  AND U47 ( .A(n72), .B(n73), .Z(n71) );
  XOR U48 ( .A(n74), .B(n75), .Z(n63) );
  AND U49 ( .A(n76), .B(n73), .Z(n75) );
  XNOR U50 ( .A(n74), .B(n70), .Z(n73) );
  XOR U51 ( .A(n77), .B(n78), .Z(n70) );
  AND U52 ( .A(n79), .B(n80), .Z(n78) );
  XOR U53 ( .A(p_input[73]), .B(n77), .Z(n80) );
  XOR U54 ( .A(n81), .B(n82), .Z(n77) );
  AND U55 ( .A(n83), .B(n84), .Z(n82) );
  XOR U56 ( .A(n85), .B(n86), .Z(n74) );
  AND U57 ( .A(n87), .B(n84), .Z(n86) );
  XNOR U58 ( .A(n85), .B(n81), .Z(n84) );
  XOR U59 ( .A(n88), .B(n89), .Z(n81) );
  AND U60 ( .A(n90), .B(n91), .Z(n89) );
  XOR U61 ( .A(p_input[89]), .B(n88), .Z(n91) );
  XOR U62 ( .A(n92), .B(n93), .Z(n88) );
  AND U63 ( .A(n94), .B(n95), .Z(n93) );
  XOR U64 ( .A(n96), .B(n97), .Z(n85) );
  AND U65 ( .A(n98), .B(n95), .Z(n97) );
  XNOR U66 ( .A(n96), .B(n92), .Z(n95) );
  XOR U67 ( .A(n99), .B(n100), .Z(n92) );
  AND U68 ( .A(n101), .B(n102), .Z(n100) );
  XOR U69 ( .A(p_input[105]), .B(n99), .Z(n102) );
  XOR U70 ( .A(n103), .B(n104), .Z(n99) );
  AND U71 ( .A(n105), .B(n106), .Z(n104) );
  XOR U72 ( .A(n107), .B(n108), .Z(n96) );
  AND U73 ( .A(n109), .B(n106), .Z(n108) );
  XNOR U74 ( .A(n107), .B(n103), .Z(n106) );
  XOR U75 ( .A(n110), .B(n111), .Z(n103) );
  AND U76 ( .A(n112), .B(n113), .Z(n111) );
  XOR U77 ( .A(p_input[121]), .B(n110), .Z(n113) );
  XOR U78 ( .A(n114), .B(n115), .Z(n110) );
  AND U79 ( .A(n116), .B(n117), .Z(n115) );
  XOR U80 ( .A(n118), .B(n119), .Z(n107) );
  AND U81 ( .A(n120), .B(n117), .Z(n119) );
  XNOR U82 ( .A(n118), .B(n114), .Z(n117) );
  XOR U83 ( .A(n121), .B(n122), .Z(n114) );
  AND U84 ( .A(n123), .B(n124), .Z(n122) );
  XOR U85 ( .A(p_input[137]), .B(n121), .Z(n124) );
  XOR U86 ( .A(n125), .B(n126), .Z(n121) );
  AND U87 ( .A(n127), .B(n128), .Z(n126) );
  XOR U88 ( .A(n129), .B(n130), .Z(n118) );
  AND U89 ( .A(n131), .B(n128), .Z(n130) );
  XNOR U90 ( .A(n129), .B(n125), .Z(n128) );
  XOR U91 ( .A(n132), .B(n133), .Z(n125) );
  AND U92 ( .A(n134), .B(n135), .Z(n133) );
  XOR U93 ( .A(p_input[153]), .B(n132), .Z(n135) );
  XOR U94 ( .A(n136), .B(n137), .Z(n132) );
  AND U95 ( .A(n138), .B(n139), .Z(n137) );
  XOR U96 ( .A(n140), .B(n141), .Z(n129) );
  AND U97 ( .A(n142), .B(n139), .Z(n141) );
  XNOR U98 ( .A(n140), .B(n136), .Z(n139) );
  XOR U99 ( .A(n143), .B(n144), .Z(n136) );
  AND U100 ( .A(n145), .B(n146), .Z(n144) );
  XOR U101 ( .A(p_input[169]), .B(n143), .Z(n146) );
  XOR U102 ( .A(n147), .B(n148), .Z(n143) );
  AND U103 ( .A(n149), .B(n150), .Z(n148) );
  XOR U104 ( .A(n151), .B(n152), .Z(n140) );
  AND U105 ( .A(n153), .B(n150), .Z(n152) );
  XNOR U106 ( .A(n151), .B(n147), .Z(n150) );
  XOR U107 ( .A(n154), .B(n155), .Z(n147) );
  AND U108 ( .A(n156), .B(n157), .Z(n155) );
  XOR U109 ( .A(p_input[185]), .B(n154), .Z(n157) );
  XOR U110 ( .A(n158), .B(n159), .Z(n154) );
  AND U111 ( .A(n160), .B(n161), .Z(n159) );
  XOR U112 ( .A(n162), .B(n163), .Z(n151) );
  AND U113 ( .A(n164), .B(n161), .Z(n163) );
  XNOR U114 ( .A(n162), .B(n158), .Z(n161) );
  XOR U115 ( .A(n165), .B(n166), .Z(n158) );
  AND U116 ( .A(n167), .B(n168), .Z(n166) );
  XOR U117 ( .A(p_input[201]), .B(n165), .Z(n168) );
  XOR U118 ( .A(n169), .B(n170), .Z(n165) );
  AND U119 ( .A(n171), .B(n172), .Z(n170) );
  XOR U120 ( .A(n173), .B(n174), .Z(n162) );
  AND U121 ( .A(n175), .B(n172), .Z(n174) );
  XNOR U122 ( .A(n173), .B(n169), .Z(n172) );
  XOR U123 ( .A(n176), .B(n177), .Z(n169) );
  AND U124 ( .A(n178), .B(n179), .Z(n177) );
  XOR U125 ( .A(p_input[217]), .B(n176), .Z(n179) );
  XOR U126 ( .A(n180), .B(n181), .Z(n176) );
  AND U127 ( .A(n182), .B(n183), .Z(n181) );
  XOR U128 ( .A(n184), .B(n185), .Z(n173) );
  AND U129 ( .A(n186), .B(n183), .Z(n185) );
  XNOR U130 ( .A(n184), .B(n180), .Z(n183) );
  XOR U131 ( .A(n187), .B(n188), .Z(n180) );
  AND U132 ( .A(n189), .B(n190), .Z(n188) );
  XOR U133 ( .A(p_input[233]), .B(n187), .Z(n190) );
  XOR U134 ( .A(n191), .B(n192), .Z(n187) );
  AND U135 ( .A(n193), .B(n194), .Z(n192) );
  XOR U136 ( .A(n195), .B(n196), .Z(n184) );
  AND U137 ( .A(n197), .B(n194), .Z(n196) );
  XNOR U138 ( .A(n195), .B(n191), .Z(n194) );
  XOR U139 ( .A(n198), .B(n199), .Z(n191) );
  AND U140 ( .A(n200), .B(n201), .Z(n199) );
  XOR U141 ( .A(p_input[249]), .B(n198), .Z(n201) );
  XOR U142 ( .A(n202), .B(n203), .Z(n198) );
  AND U143 ( .A(n204), .B(n205), .Z(n203) );
  XOR U144 ( .A(n206), .B(n207), .Z(n195) );
  AND U145 ( .A(n208), .B(n205), .Z(n207) );
  XNOR U146 ( .A(n206), .B(n202), .Z(n205) );
  XOR U147 ( .A(n209), .B(n210), .Z(n202) );
  AND U148 ( .A(n211), .B(n212), .Z(n210) );
  XOR U149 ( .A(p_input[265]), .B(n209), .Z(n212) );
  XOR U150 ( .A(n213), .B(n214), .Z(n209) );
  AND U151 ( .A(n215), .B(n216), .Z(n214) );
  XOR U152 ( .A(n217), .B(n218), .Z(n206) );
  AND U153 ( .A(n219), .B(n216), .Z(n218) );
  XNOR U154 ( .A(n217), .B(n213), .Z(n216) );
  XOR U155 ( .A(n220), .B(n221), .Z(n213) );
  AND U156 ( .A(n222), .B(n223), .Z(n221) );
  XOR U157 ( .A(p_input[281]), .B(n220), .Z(n223) );
  XOR U158 ( .A(n224), .B(n225), .Z(n220) );
  AND U159 ( .A(n226), .B(n227), .Z(n225) );
  XOR U160 ( .A(n228), .B(n229), .Z(n217) );
  AND U161 ( .A(n230), .B(n227), .Z(n229) );
  XNOR U162 ( .A(n228), .B(n224), .Z(n227) );
  XOR U163 ( .A(n231), .B(n232), .Z(n224) );
  AND U164 ( .A(n233), .B(n234), .Z(n232) );
  XOR U165 ( .A(p_input[297]), .B(n231), .Z(n234) );
  XOR U166 ( .A(n235), .B(n236), .Z(n231) );
  AND U167 ( .A(n237), .B(n238), .Z(n236) );
  XOR U168 ( .A(n239), .B(n240), .Z(n228) );
  AND U169 ( .A(n241), .B(n238), .Z(n240) );
  XNOR U170 ( .A(n239), .B(n235), .Z(n238) );
  XOR U171 ( .A(n242), .B(n243), .Z(n235) );
  AND U172 ( .A(n244), .B(n245), .Z(n243) );
  XOR U173 ( .A(p_input[313]), .B(n242), .Z(n245) );
  XOR U174 ( .A(n246), .B(n247), .Z(n242) );
  AND U175 ( .A(n248), .B(n249), .Z(n247) );
  XOR U176 ( .A(n250), .B(n251), .Z(n239) );
  AND U177 ( .A(n252), .B(n249), .Z(n251) );
  XNOR U178 ( .A(n250), .B(n246), .Z(n249) );
  XOR U179 ( .A(n253), .B(n254), .Z(n246) );
  AND U180 ( .A(n255), .B(n256), .Z(n254) );
  XOR U181 ( .A(p_input[329]), .B(n253), .Z(n256) );
  XOR U182 ( .A(n257), .B(n258), .Z(n253) );
  AND U183 ( .A(n259), .B(n260), .Z(n258) );
  XOR U184 ( .A(n261), .B(n262), .Z(n250) );
  AND U185 ( .A(n263), .B(n260), .Z(n262) );
  XNOR U186 ( .A(n261), .B(n257), .Z(n260) );
  XOR U187 ( .A(n264), .B(n265), .Z(n257) );
  AND U188 ( .A(n266), .B(n267), .Z(n265) );
  XOR U189 ( .A(p_input[345]), .B(n264), .Z(n267) );
  XOR U190 ( .A(n268), .B(n269), .Z(n264) );
  AND U191 ( .A(n270), .B(n271), .Z(n269) );
  XOR U192 ( .A(n272), .B(n273), .Z(n261) );
  AND U193 ( .A(n274), .B(n271), .Z(n273) );
  XNOR U194 ( .A(n272), .B(n268), .Z(n271) );
  XOR U195 ( .A(n275), .B(n276), .Z(n268) );
  AND U196 ( .A(n277), .B(n278), .Z(n276) );
  XOR U197 ( .A(p_input[361]), .B(n275), .Z(n278) );
  XOR U198 ( .A(n279), .B(n280), .Z(n275) );
  AND U199 ( .A(n281), .B(n282), .Z(n280) );
  XOR U200 ( .A(n283), .B(n284), .Z(n272) );
  AND U201 ( .A(n285), .B(n282), .Z(n284) );
  XNOR U202 ( .A(n283), .B(n279), .Z(n282) );
  XOR U203 ( .A(n286), .B(n287), .Z(n279) );
  AND U204 ( .A(n288), .B(n289), .Z(n287) );
  XOR U205 ( .A(p_input[377]), .B(n286), .Z(n289) );
  XOR U206 ( .A(n290), .B(n291), .Z(n286) );
  AND U207 ( .A(n292), .B(n293), .Z(n291) );
  XOR U208 ( .A(n294), .B(n295), .Z(n283) );
  AND U209 ( .A(n296), .B(n293), .Z(n295) );
  XNOR U210 ( .A(n294), .B(n290), .Z(n293) );
  XOR U211 ( .A(n297), .B(n298), .Z(n290) );
  AND U212 ( .A(n299), .B(n300), .Z(n298) );
  XOR U213 ( .A(p_input[393]), .B(n297), .Z(n300) );
  XOR U214 ( .A(n301), .B(n302), .Z(n297) );
  AND U215 ( .A(n303), .B(n304), .Z(n302) );
  XOR U216 ( .A(n305), .B(n306), .Z(n294) );
  AND U217 ( .A(n307), .B(n304), .Z(n306) );
  XNOR U218 ( .A(n305), .B(n301), .Z(n304) );
  XOR U219 ( .A(n308), .B(n309), .Z(n301) );
  AND U220 ( .A(n310), .B(n311), .Z(n309) );
  XOR U221 ( .A(p_input[409]), .B(n308), .Z(n311) );
  XOR U222 ( .A(n312), .B(n313), .Z(n308) );
  AND U223 ( .A(n314), .B(n315), .Z(n313) );
  XOR U224 ( .A(n316), .B(n317), .Z(n305) );
  AND U225 ( .A(n318), .B(n315), .Z(n317) );
  XNOR U226 ( .A(n316), .B(n312), .Z(n315) );
  XOR U227 ( .A(n319), .B(n320), .Z(n312) );
  AND U228 ( .A(n321), .B(n322), .Z(n320) );
  XOR U229 ( .A(p_input[425]), .B(n319), .Z(n322) );
  XOR U230 ( .A(n323), .B(n324), .Z(n319) );
  AND U231 ( .A(n325), .B(n326), .Z(n324) );
  XOR U232 ( .A(n327), .B(n328), .Z(n316) );
  AND U233 ( .A(n329), .B(n326), .Z(n328) );
  XNOR U234 ( .A(n327), .B(n323), .Z(n326) );
  XOR U235 ( .A(n330), .B(n331), .Z(n323) );
  AND U236 ( .A(n332), .B(n333), .Z(n331) );
  XOR U237 ( .A(p_input[441]), .B(n330), .Z(n333) );
  XOR U238 ( .A(n334), .B(n335), .Z(n330) );
  AND U239 ( .A(n336), .B(n337), .Z(n335) );
  XOR U240 ( .A(n338), .B(n339), .Z(n327) );
  AND U241 ( .A(n340), .B(n337), .Z(n339) );
  XNOR U242 ( .A(n338), .B(n334), .Z(n337) );
  XOR U243 ( .A(n341), .B(n342), .Z(n334) );
  AND U244 ( .A(n343), .B(n344), .Z(n342) );
  XOR U245 ( .A(p_input[457]), .B(n341), .Z(n344) );
  XOR U246 ( .A(n345), .B(n346), .Z(n341) );
  AND U247 ( .A(n347), .B(n348), .Z(n346) );
  XOR U248 ( .A(n349), .B(n350), .Z(n338) );
  AND U249 ( .A(n351), .B(n348), .Z(n350) );
  XNOR U250 ( .A(n349), .B(n345), .Z(n348) );
  XOR U251 ( .A(n352), .B(n353), .Z(n345) );
  AND U252 ( .A(n354), .B(n355), .Z(n353) );
  XOR U253 ( .A(p_input[473]), .B(n352), .Z(n355) );
  XOR U254 ( .A(n356), .B(n357), .Z(n352) );
  AND U255 ( .A(n358), .B(n359), .Z(n357) );
  XOR U256 ( .A(n360), .B(n361), .Z(n349) );
  AND U257 ( .A(n362), .B(n359), .Z(n361) );
  XNOR U258 ( .A(n360), .B(n356), .Z(n359) );
  XOR U259 ( .A(n363), .B(n364), .Z(n356) );
  AND U260 ( .A(n365), .B(n366), .Z(n364) );
  XOR U261 ( .A(p_input[489]), .B(n363), .Z(n366) );
  XOR U262 ( .A(n367), .B(n368), .Z(n363) );
  AND U263 ( .A(n369), .B(n370), .Z(n368) );
  XOR U264 ( .A(n371), .B(n372), .Z(n360) );
  AND U265 ( .A(n373), .B(n370), .Z(n372) );
  XNOR U266 ( .A(n371), .B(n367), .Z(n370) );
  XOR U267 ( .A(n374), .B(n375), .Z(n367) );
  AND U268 ( .A(n376), .B(n377), .Z(n375) );
  XOR U269 ( .A(p_input[505]), .B(n374), .Z(n377) );
  XOR U270 ( .A(n378), .B(n379), .Z(n374) );
  AND U271 ( .A(n380), .B(n381), .Z(n379) );
  XOR U272 ( .A(n382), .B(n383), .Z(n371) );
  AND U273 ( .A(n384), .B(n381), .Z(n383) );
  XNOR U274 ( .A(n382), .B(n378), .Z(n381) );
  XOR U275 ( .A(n385), .B(n386), .Z(n378) );
  AND U276 ( .A(n387), .B(n388), .Z(n386) );
  XOR U277 ( .A(p_input[521]), .B(n385), .Z(n388) );
  XOR U278 ( .A(n389), .B(n390), .Z(n385) );
  AND U279 ( .A(n391), .B(n392), .Z(n390) );
  XOR U280 ( .A(n393), .B(n394), .Z(n382) );
  AND U281 ( .A(n395), .B(n392), .Z(n394) );
  XNOR U282 ( .A(n393), .B(n389), .Z(n392) );
  XOR U283 ( .A(n396), .B(n397), .Z(n389) );
  AND U284 ( .A(n398), .B(n399), .Z(n397) );
  XOR U285 ( .A(p_input[537]), .B(n396), .Z(n399) );
  XOR U286 ( .A(n400), .B(n401), .Z(n396) );
  AND U287 ( .A(n402), .B(n403), .Z(n401) );
  XOR U288 ( .A(n404), .B(n405), .Z(n393) );
  AND U289 ( .A(n406), .B(n403), .Z(n405) );
  XNOR U290 ( .A(n404), .B(n400), .Z(n403) );
  XOR U291 ( .A(n407), .B(n408), .Z(n400) );
  AND U292 ( .A(n409), .B(n410), .Z(n408) );
  XOR U293 ( .A(p_input[553]), .B(n407), .Z(n410) );
  XOR U294 ( .A(n411), .B(n412), .Z(n407) );
  AND U295 ( .A(n413), .B(n414), .Z(n412) );
  XOR U296 ( .A(n415), .B(n416), .Z(n404) );
  AND U297 ( .A(n417), .B(n414), .Z(n416) );
  XNOR U298 ( .A(n415), .B(n411), .Z(n414) );
  XOR U299 ( .A(n418), .B(n419), .Z(n411) );
  AND U300 ( .A(n420), .B(n421), .Z(n419) );
  XOR U301 ( .A(p_input[569]), .B(n418), .Z(n421) );
  XOR U302 ( .A(n422), .B(n423), .Z(n418) );
  AND U303 ( .A(n424), .B(n425), .Z(n423) );
  XOR U304 ( .A(n426), .B(n427), .Z(n415) );
  AND U305 ( .A(n428), .B(n425), .Z(n427) );
  XNOR U306 ( .A(n426), .B(n422), .Z(n425) );
  XOR U307 ( .A(n429), .B(n430), .Z(n422) );
  AND U308 ( .A(n431), .B(n432), .Z(n430) );
  XOR U309 ( .A(p_input[585]), .B(n429), .Z(n432) );
  XOR U310 ( .A(n433), .B(n434), .Z(n429) );
  AND U311 ( .A(n435), .B(n436), .Z(n434) );
  XOR U312 ( .A(n437), .B(n438), .Z(n426) );
  AND U313 ( .A(n439), .B(n436), .Z(n438) );
  XNOR U314 ( .A(n437), .B(n433), .Z(n436) );
  XOR U315 ( .A(n440), .B(n441), .Z(n433) );
  AND U316 ( .A(n442), .B(n443), .Z(n441) );
  XOR U317 ( .A(p_input[601]), .B(n440), .Z(n443) );
  XOR U318 ( .A(n444), .B(n445), .Z(n440) );
  AND U319 ( .A(n446), .B(n447), .Z(n445) );
  XOR U320 ( .A(n448), .B(n449), .Z(n437) );
  AND U321 ( .A(n450), .B(n447), .Z(n449) );
  XNOR U322 ( .A(n448), .B(n444), .Z(n447) );
  XOR U323 ( .A(n451), .B(n452), .Z(n444) );
  AND U324 ( .A(n453), .B(n454), .Z(n452) );
  XOR U325 ( .A(p_input[617]), .B(n451), .Z(n454) );
  XOR U326 ( .A(n455), .B(n456), .Z(n451) );
  AND U327 ( .A(n457), .B(n458), .Z(n456) );
  XOR U328 ( .A(n459), .B(n460), .Z(n448) );
  AND U329 ( .A(n461), .B(n458), .Z(n460) );
  XNOR U330 ( .A(n459), .B(n455), .Z(n458) );
  XOR U331 ( .A(n462), .B(n463), .Z(n455) );
  AND U332 ( .A(n464), .B(n465), .Z(n463) );
  XOR U333 ( .A(p_input[633]), .B(n462), .Z(n465) );
  XOR U334 ( .A(n466), .B(n467), .Z(n462) );
  AND U335 ( .A(n468), .B(n469), .Z(n467) );
  XOR U336 ( .A(n470), .B(n471), .Z(n459) );
  AND U337 ( .A(n472), .B(n469), .Z(n471) );
  XNOR U338 ( .A(n470), .B(n466), .Z(n469) );
  XOR U339 ( .A(n473), .B(n474), .Z(n466) );
  AND U340 ( .A(n475), .B(n476), .Z(n474) );
  XOR U341 ( .A(p_input[649]), .B(n473), .Z(n476) );
  XOR U342 ( .A(n477), .B(n478), .Z(n473) );
  AND U343 ( .A(n479), .B(n480), .Z(n478) );
  XOR U344 ( .A(n481), .B(n482), .Z(n470) );
  AND U345 ( .A(n483), .B(n480), .Z(n482) );
  XNOR U346 ( .A(n481), .B(n477), .Z(n480) );
  XOR U347 ( .A(n484), .B(n485), .Z(n477) );
  AND U348 ( .A(n486), .B(n487), .Z(n485) );
  XOR U349 ( .A(p_input[665]), .B(n484), .Z(n487) );
  XOR U350 ( .A(n488), .B(n489), .Z(n484) );
  AND U351 ( .A(n490), .B(n491), .Z(n489) );
  XOR U352 ( .A(n492), .B(n493), .Z(n481) );
  AND U353 ( .A(n494), .B(n491), .Z(n493) );
  XNOR U354 ( .A(n492), .B(n488), .Z(n491) );
  XOR U355 ( .A(n495), .B(n496), .Z(n488) );
  AND U356 ( .A(n497), .B(n498), .Z(n496) );
  XOR U357 ( .A(p_input[681]), .B(n495), .Z(n498) );
  XOR U358 ( .A(n499), .B(n500), .Z(n495) );
  AND U359 ( .A(n501), .B(n502), .Z(n500) );
  XOR U360 ( .A(n503), .B(n504), .Z(n492) );
  AND U361 ( .A(n505), .B(n502), .Z(n504) );
  XNOR U362 ( .A(n503), .B(n499), .Z(n502) );
  XOR U363 ( .A(n506), .B(n507), .Z(n499) );
  AND U364 ( .A(n508), .B(n509), .Z(n507) );
  XOR U365 ( .A(p_input[697]), .B(n506), .Z(n509) );
  XOR U366 ( .A(n510), .B(n511), .Z(n506) );
  AND U367 ( .A(n512), .B(n513), .Z(n511) );
  XOR U368 ( .A(n514), .B(n515), .Z(n503) );
  AND U369 ( .A(n516), .B(n513), .Z(n515) );
  XNOR U370 ( .A(n514), .B(n510), .Z(n513) );
  XOR U371 ( .A(n517), .B(n518), .Z(n510) );
  AND U372 ( .A(n519), .B(n520), .Z(n518) );
  XOR U373 ( .A(p_input[713]), .B(n517), .Z(n520) );
  XOR U374 ( .A(n521), .B(n522), .Z(n517) );
  AND U375 ( .A(n523), .B(n524), .Z(n522) );
  XOR U376 ( .A(n525), .B(n526), .Z(n514) );
  AND U377 ( .A(n527), .B(n524), .Z(n526) );
  XNOR U378 ( .A(n525), .B(n521), .Z(n524) );
  XOR U379 ( .A(n528), .B(n529), .Z(n521) );
  AND U380 ( .A(n530), .B(n531), .Z(n529) );
  XOR U381 ( .A(p_input[729]), .B(n528), .Z(n531) );
  XOR U382 ( .A(n532), .B(n533), .Z(n528) );
  AND U383 ( .A(n534), .B(n535), .Z(n533) );
  XOR U384 ( .A(n536), .B(n537), .Z(n525) );
  AND U385 ( .A(n538), .B(n535), .Z(n537) );
  XNOR U386 ( .A(n536), .B(n532), .Z(n535) );
  XOR U387 ( .A(n539), .B(n540), .Z(n532) );
  AND U388 ( .A(n541), .B(n542), .Z(n540) );
  XOR U389 ( .A(p_input[745]), .B(n539), .Z(n542) );
  XOR U390 ( .A(n543), .B(n544), .Z(n539) );
  AND U391 ( .A(n545), .B(n546), .Z(n544) );
  XOR U392 ( .A(n547), .B(n548), .Z(n536) );
  AND U393 ( .A(n549), .B(n546), .Z(n548) );
  XNOR U394 ( .A(n547), .B(n543), .Z(n546) );
  XOR U395 ( .A(n550), .B(n551), .Z(n543) );
  AND U396 ( .A(n552), .B(n553), .Z(n551) );
  XOR U397 ( .A(p_input[761]), .B(n550), .Z(n553) );
  XOR U398 ( .A(n554), .B(n555), .Z(n550) );
  AND U399 ( .A(n556), .B(n557), .Z(n555) );
  XOR U400 ( .A(n558), .B(n559), .Z(n547) );
  AND U401 ( .A(n560), .B(n557), .Z(n559) );
  XNOR U402 ( .A(n558), .B(n554), .Z(n557) );
  XOR U403 ( .A(n561), .B(n562), .Z(n554) );
  AND U404 ( .A(n563), .B(n564), .Z(n562) );
  XOR U405 ( .A(p_input[777]), .B(n561), .Z(n564) );
  XOR U406 ( .A(n565), .B(n566), .Z(n561) );
  AND U407 ( .A(n567), .B(n568), .Z(n566) );
  XOR U408 ( .A(n569), .B(n570), .Z(n558) );
  AND U409 ( .A(n571), .B(n568), .Z(n570) );
  XNOR U410 ( .A(n569), .B(n565), .Z(n568) );
  XOR U411 ( .A(n572), .B(n573), .Z(n565) );
  AND U412 ( .A(n574), .B(n575), .Z(n573) );
  XOR U413 ( .A(p_input[793]), .B(n572), .Z(n575) );
  XOR U414 ( .A(n576), .B(n577), .Z(n572) );
  AND U415 ( .A(n578), .B(n579), .Z(n577) );
  XOR U416 ( .A(n580), .B(n581), .Z(n569) );
  AND U417 ( .A(n582), .B(n579), .Z(n581) );
  XNOR U418 ( .A(n580), .B(n576), .Z(n579) );
  XOR U419 ( .A(n583), .B(n584), .Z(n576) );
  AND U420 ( .A(n585), .B(n586), .Z(n584) );
  XOR U421 ( .A(p_input[809]), .B(n583), .Z(n586) );
  XOR U422 ( .A(n587), .B(n588), .Z(n583) );
  AND U423 ( .A(n589), .B(n590), .Z(n588) );
  XOR U424 ( .A(n591), .B(n592), .Z(n580) );
  AND U425 ( .A(n593), .B(n590), .Z(n592) );
  XNOR U426 ( .A(n591), .B(n587), .Z(n590) );
  XOR U427 ( .A(n594), .B(n595), .Z(n587) );
  AND U428 ( .A(n596), .B(n597), .Z(n595) );
  XOR U429 ( .A(p_input[825]), .B(n594), .Z(n597) );
  XOR U430 ( .A(n598), .B(n599), .Z(n594) );
  AND U431 ( .A(n600), .B(n601), .Z(n599) );
  XOR U432 ( .A(n602), .B(n603), .Z(n591) );
  AND U433 ( .A(n604), .B(n601), .Z(n603) );
  XNOR U434 ( .A(n602), .B(n598), .Z(n601) );
  XOR U435 ( .A(n605), .B(n606), .Z(n598) );
  AND U436 ( .A(n607), .B(n608), .Z(n606) );
  XOR U437 ( .A(p_input[841]), .B(n605), .Z(n608) );
  XOR U438 ( .A(n609), .B(n610), .Z(n605) );
  AND U439 ( .A(n611), .B(n612), .Z(n610) );
  XOR U440 ( .A(n613), .B(n614), .Z(n602) );
  AND U441 ( .A(n615), .B(n612), .Z(n614) );
  XNOR U442 ( .A(n613), .B(n609), .Z(n612) );
  XOR U443 ( .A(n616), .B(n617), .Z(n609) );
  AND U444 ( .A(n618), .B(n619), .Z(n617) );
  XOR U445 ( .A(p_input[857]), .B(n616), .Z(n619) );
  XOR U446 ( .A(n620), .B(n621), .Z(n616) );
  AND U447 ( .A(n622), .B(n623), .Z(n621) );
  XOR U448 ( .A(n624), .B(n625), .Z(n613) );
  AND U449 ( .A(n626), .B(n623), .Z(n625) );
  XNOR U450 ( .A(n624), .B(n620), .Z(n623) );
  XOR U451 ( .A(n627), .B(n628), .Z(n620) );
  AND U452 ( .A(n629), .B(n630), .Z(n628) );
  XOR U453 ( .A(p_input[873]), .B(n627), .Z(n630) );
  XOR U454 ( .A(n631), .B(n632), .Z(n627) );
  AND U455 ( .A(n633), .B(n634), .Z(n632) );
  XOR U456 ( .A(n635), .B(n636), .Z(n624) );
  AND U457 ( .A(n637), .B(n634), .Z(n636) );
  XNOR U458 ( .A(n635), .B(n631), .Z(n634) );
  XOR U459 ( .A(n638), .B(n639), .Z(n631) );
  AND U460 ( .A(n640), .B(n641), .Z(n639) );
  XOR U461 ( .A(p_input[889]), .B(n638), .Z(n641) );
  XOR U462 ( .A(n642), .B(n643), .Z(n638) );
  AND U463 ( .A(n644), .B(n645), .Z(n643) );
  XOR U464 ( .A(n646), .B(n647), .Z(n635) );
  AND U465 ( .A(n648), .B(n645), .Z(n647) );
  XNOR U466 ( .A(n646), .B(n642), .Z(n645) );
  XOR U467 ( .A(n649), .B(n650), .Z(n642) );
  AND U468 ( .A(n651), .B(n652), .Z(n650) );
  XOR U469 ( .A(p_input[905]), .B(n649), .Z(n652) );
  XOR U470 ( .A(n653), .B(n654), .Z(n649) );
  AND U471 ( .A(n655), .B(n656), .Z(n654) );
  XOR U472 ( .A(n657), .B(n658), .Z(n646) );
  AND U473 ( .A(n659), .B(n656), .Z(n658) );
  XNOR U474 ( .A(n657), .B(n653), .Z(n656) );
  XOR U475 ( .A(n660), .B(n661), .Z(n653) );
  AND U476 ( .A(n662), .B(n663), .Z(n661) );
  XOR U477 ( .A(p_input[921]), .B(n660), .Z(n663) );
  XOR U478 ( .A(n664), .B(n665), .Z(n660) );
  AND U479 ( .A(n666), .B(n667), .Z(n665) );
  XOR U480 ( .A(n668), .B(n669), .Z(n657) );
  AND U481 ( .A(n670), .B(n667), .Z(n669) );
  XNOR U482 ( .A(n668), .B(n664), .Z(n667) );
  XOR U483 ( .A(n671), .B(n672), .Z(n664) );
  AND U484 ( .A(n673), .B(n674), .Z(n672) );
  XOR U485 ( .A(p_input[937]), .B(n671), .Z(n674) );
  XOR U486 ( .A(n675), .B(n676), .Z(n671) );
  AND U487 ( .A(n677), .B(n678), .Z(n676) );
  XOR U488 ( .A(n679), .B(n680), .Z(n668) );
  AND U489 ( .A(n681), .B(n678), .Z(n680) );
  XNOR U490 ( .A(n679), .B(n675), .Z(n678) );
  XOR U491 ( .A(n682), .B(n683), .Z(n675) );
  AND U492 ( .A(n684), .B(n685), .Z(n683) );
  XOR U493 ( .A(p_input[953]), .B(n682), .Z(n685) );
  XOR U494 ( .A(n686), .B(n687), .Z(n682) );
  AND U495 ( .A(n688), .B(n689), .Z(n687) );
  XOR U496 ( .A(n690), .B(n691), .Z(n679) );
  AND U497 ( .A(n692), .B(n689), .Z(n691) );
  XNOR U498 ( .A(n690), .B(n686), .Z(n689) );
  XOR U499 ( .A(n693), .B(n694), .Z(n686) );
  AND U500 ( .A(n695), .B(n696), .Z(n694) );
  XOR U501 ( .A(p_input[969]), .B(n693), .Z(n696) );
  XOR U502 ( .A(n697), .B(n698), .Z(n693) );
  AND U503 ( .A(n699), .B(n700), .Z(n698) );
  XOR U504 ( .A(n701), .B(n702), .Z(n690) );
  AND U505 ( .A(n703), .B(n700), .Z(n702) );
  XNOR U506 ( .A(n701), .B(n697), .Z(n700) );
  XOR U507 ( .A(n704), .B(n705), .Z(n697) );
  AND U508 ( .A(n706), .B(n707), .Z(n705) );
  XOR U509 ( .A(p_input[985]), .B(n704), .Z(n707) );
  XOR U510 ( .A(n708), .B(n709), .Z(n704) );
  AND U511 ( .A(n710), .B(n711), .Z(n709) );
  XOR U512 ( .A(n712), .B(n713), .Z(n701) );
  AND U513 ( .A(n714), .B(n711), .Z(n713) );
  XNOR U514 ( .A(n712), .B(n708), .Z(n711) );
  XOR U515 ( .A(n715), .B(n716), .Z(n708) );
  AND U516 ( .A(n717), .B(n718), .Z(n716) );
  XOR U517 ( .A(p_input[1001]), .B(n715), .Z(n718) );
  XOR U518 ( .A(n719), .B(n720), .Z(n715) );
  AND U519 ( .A(n721), .B(n722), .Z(n720) );
  XOR U520 ( .A(n723), .B(n724), .Z(n712) );
  AND U521 ( .A(n725), .B(n722), .Z(n724) );
  XNOR U522 ( .A(n723), .B(n719), .Z(n722) );
  XOR U523 ( .A(n726), .B(n727), .Z(n719) );
  AND U524 ( .A(n728), .B(n729), .Z(n727) );
  XOR U525 ( .A(p_input[1017]), .B(n726), .Z(n729) );
  XOR U526 ( .A(n730), .B(n731), .Z(n726) );
  AND U527 ( .A(n732), .B(n733), .Z(n731) );
  XOR U528 ( .A(n734), .B(n735), .Z(n723) );
  AND U529 ( .A(n736), .B(n733), .Z(n735) );
  XNOR U530 ( .A(n734), .B(n730), .Z(n733) );
  XOR U531 ( .A(n737), .B(n738), .Z(n730) );
  AND U532 ( .A(n739), .B(n740), .Z(n738) );
  XOR U533 ( .A(p_input[1033]), .B(n737), .Z(n740) );
  XOR U534 ( .A(n741), .B(n742), .Z(n737) );
  AND U535 ( .A(n743), .B(n744), .Z(n742) );
  XOR U536 ( .A(n745), .B(n746), .Z(n734) );
  AND U537 ( .A(n747), .B(n744), .Z(n746) );
  XNOR U538 ( .A(n745), .B(n741), .Z(n744) );
  XOR U539 ( .A(n748), .B(n749), .Z(n741) );
  AND U540 ( .A(n750), .B(n751), .Z(n749) );
  XOR U541 ( .A(p_input[1049]), .B(n748), .Z(n751) );
  XOR U542 ( .A(n752), .B(n753), .Z(n748) );
  AND U543 ( .A(n754), .B(n755), .Z(n753) );
  XOR U544 ( .A(n756), .B(n757), .Z(n745) );
  AND U545 ( .A(n758), .B(n755), .Z(n757) );
  XNOR U546 ( .A(n756), .B(n752), .Z(n755) );
  XOR U547 ( .A(n759), .B(n760), .Z(n752) );
  AND U548 ( .A(n761), .B(n762), .Z(n760) );
  XOR U549 ( .A(p_input[1065]), .B(n759), .Z(n762) );
  XOR U550 ( .A(n763), .B(n764), .Z(n759) );
  AND U551 ( .A(n765), .B(n766), .Z(n764) );
  XOR U552 ( .A(n767), .B(n768), .Z(n756) );
  AND U553 ( .A(n769), .B(n766), .Z(n768) );
  XNOR U554 ( .A(n767), .B(n763), .Z(n766) );
  XOR U555 ( .A(n770), .B(n771), .Z(n763) );
  AND U556 ( .A(n772), .B(n773), .Z(n771) );
  XOR U557 ( .A(p_input[1081]), .B(n770), .Z(n773) );
  XOR U558 ( .A(n774), .B(n775), .Z(n770) );
  AND U559 ( .A(n776), .B(n777), .Z(n775) );
  XOR U560 ( .A(n778), .B(n779), .Z(n767) );
  AND U561 ( .A(n780), .B(n777), .Z(n779) );
  XNOR U562 ( .A(n778), .B(n774), .Z(n777) );
  XOR U563 ( .A(n781), .B(n782), .Z(n774) );
  AND U564 ( .A(n783), .B(n784), .Z(n782) );
  XOR U565 ( .A(p_input[1097]), .B(n781), .Z(n784) );
  XOR U566 ( .A(n785), .B(n786), .Z(n781) );
  AND U567 ( .A(n787), .B(n788), .Z(n786) );
  XOR U568 ( .A(n789), .B(n790), .Z(n778) );
  AND U569 ( .A(n791), .B(n788), .Z(n790) );
  XNOR U570 ( .A(n789), .B(n785), .Z(n788) );
  XOR U571 ( .A(n792), .B(n793), .Z(n785) );
  AND U572 ( .A(n794), .B(n795), .Z(n793) );
  XOR U573 ( .A(p_input[1113]), .B(n792), .Z(n795) );
  XOR U574 ( .A(n796), .B(n797), .Z(n792) );
  AND U575 ( .A(n798), .B(n799), .Z(n797) );
  XOR U576 ( .A(n800), .B(n801), .Z(n789) );
  AND U577 ( .A(n802), .B(n799), .Z(n801) );
  XNOR U578 ( .A(n800), .B(n796), .Z(n799) );
  XOR U579 ( .A(n803), .B(n804), .Z(n796) );
  AND U580 ( .A(n805), .B(n806), .Z(n804) );
  XOR U581 ( .A(p_input[1129]), .B(n803), .Z(n806) );
  XOR U582 ( .A(n807), .B(n808), .Z(n803) );
  AND U583 ( .A(n809), .B(n810), .Z(n808) );
  XOR U584 ( .A(n811), .B(n812), .Z(n800) );
  AND U585 ( .A(n813), .B(n810), .Z(n812) );
  XNOR U586 ( .A(n811), .B(n807), .Z(n810) );
  XOR U587 ( .A(n814), .B(n815), .Z(n807) );
  AND U588 ( .A(n816), .B(n817), .Z(n815) );
  XOR U589 ( .A(p_input[1145]), .B(n814), .Z(n817) );
  XOR U590 ( .A(n818), .B(n819), .Z(n814) );
  AND U591 ( .A(n820), .B(n821), .Z(n819) );
  XOR U592 ( .A(n822), .B(n823), .Z(n811) );
  AND U593 ( .A(n824), .B(n821), .Z(n823) );
  XNOR U594 ( .A(n822), .B(n818), .Z(n821) );
  XOR U595 ( .A(n825), .B(n826), .Z(n818) );
  AND U596 ( .A(n827), .B(n828), .Z(n826) );
  XOR U597 ( .A(p_input[1161]), .B(n825), .Z(n828) );
  XOR U598 ( .A(n829), .B(n830), .Z(n825) );
  AND U599 ( .A(n831), .B(n832), .Z(n830) );
  XOR U600 ( .A(n833), .B(n834), .Z(n822) );
  AND U601 ( .A(n835), .B(n832), .Z(n834) );
  XNOR U602 ( .A(n833), .B(n829), .Z(n832) );
  XOR U603 ( .A(n836), .B(n837), .Z(n829) );
  AND U604 ( .A(n838), .B(n839), .Z(n837) );
  XOR U605 ( .A(p_input[1177]), .B(n836), .Z(n839) );
  XOR U606 ( .A(n840), .B(n841), .Z(n836) );
  AND U607 ( .A(n842), .B(n843), .Z(n841) );
  XOR U608 ( .A(n844), .B(n845), .Z(n833) );
  AND U609 ( .A(n846), .B(n843), .Z(n845) );
  XNOR U610 ( .A(n844), .B(n840), .Z(n843) );
  XOR U611 ( .A(n847), .B(n848), .Z(n840) );
  AND U612 ( .A(n849), .B(n850), .Z(n848) );
  XOR U613 ( .A(p_input[1193]), .B(n847), .Z(n850) );
  XOR U614 ( .A(n851), .B(n852), .Z(n847) );
  AND U615 ( .A(n853), .B(n854), .Z(n852) );
  XOR U616 ( .A(n855), .B(n856), .Z(n844) );
  AND U617 ( .A(n857), .B(n854), .Z(n856) );
  XNOR U618 ( .A(n855), .B(n851), .Z(n854) );
  XOR U619 ( .A(n858), .B(n859), .Z(n851) );
  AND U620 ( .A(n860), .B(n861), .Z(n859) );
  XOR U621 ( .A(p_input[1209]), .B(n858), .Z(n861) );
  XOR U622 ( .A(n862), .B(n863), .Z(n858) );
  AND U623 ( .A(n864), .B(n865), .Z(n863) );
  XOR U624 ( .A(n866), .B(n867), .Z(n855) );
  AND U625 ( .A(n868), .B(n865), .Z(n867) );
  XNOR U626 ( .A(n866), .B(n862), .Z(n865) );
  XOR U627 ( .A(n869), .B(n870), .Z(n862) );
  AND U628 ( .A(n871), .B(n872), .Z(n870) );
  XOR U629 ( .A(p_input[1225]), .B(n869), .Z(n872) );
  XOR U630 ( .A(n873), .B(n874), .Z(n869) );
  AND U631 ( .A(n875), .B(n876), .Z(n874) );
  XOR U632 ( .A(n877), .B(n878), .Z(n866) );
  AND U633 ( .A(n879), .B(n876), .Z(n878) );
  XNOR U634 ( .A(n877), .B(n873), .Z(n876) );
  XOR U635 ( .A(n880), .B(n881), .Z(n873) );
  AND U636 ( .A(n882), .B(n883), .Z(n881) );
  XOR U637 ( .A(p_input[1241]), .B(n880), .Z(n883) );
  XOR U638 ( .A(n884), .B(n885), .Z(n880) );
  AND U639 ( .A(n886), .B(n887), .Z(n885) );
  XOR U640 ( .A(n888), .B(n889), .Z(n877) );
  AND U641 ( .A(n890), .B(n887), .Z(n889) );
  XNOR U642 ( .A(n888), .B(n884), .Z(n887) );
  XOR U643 ( .A(n891), .B(n892), .Z(n884) );
  AND U644 ( .A(n893), .B(n894), .Z(n892) );
  XOR U645 ( .A(p_input[1257]), .B(n891), .Z(n894) );
  XOR U646 ( .A(n895), .B(n896), .Z(n891) );
  AND U647 ( .A(n897), .B(n898), .Z(n896) );
  XOR U648 ( .A(n899), .B(n900), .Z(n888) );
  AND U649 ( .A(n901), .B(n898), .Z(n900) );
  XNOR U650 ( .A(n899), .B(n895), .Z(n898) );
  XOR U651 ( .A(n902), .B(n903), .Z(n895) );
  AND U652 ( .A(n904), .B(n905), .Z(n903) );
  XOR U653 ( .A(p_input[1273]), .B(n902), .Z(n905) );
  XOR U654 ( .A(n906), .B(n907), .Z(n902) );
  AND U655 ( .A(n908), .B(n909), .Z(n907) );
  XOR U656 ( .A(n910), .B(n911), .Z(n899) );
  AND U657 ( .A(n912), .B(n909), .Z(n911) );
  XNOR U658 ( .A(n910), .B(n906), .Z(n909) );
  XOR U659 ( .A(n913), .B(n914), .Z(n906) );
  AND U660 ( .A(n915), .B(n916), .Z(n914) );
  XOR U661 ( .A(p_input[1289]), .B(n913), .Z(n916) );
  XOR U662 ( .A(n917), .B(n918), .Z(n913) );
  AND U663 ( .A(n919), .B(n920), .Z(n918) );
  XOR U664 ( .A(n921), .B(n922), .Z(n910) );
  AND U665 ( .A(n923), .B(n920), .Z(n922) );
  XNOR U666 ( .A(n921), .B(n917), .Z(n920) );
  XOR U667 ( .A(n924), .B(n925), .Z(n917) );
  AND U668 ( .A(n926), .B(n927), .Z(n925) );
  XOR U669 ( .A(p_input[1305]), .B(n924), .Z(n927) );
  XOR U670 ( .A(n928), .B(n929), .Z(n924) );
  AND U671 ( .A(n930), .B(n931), .Z(n929) );
  XOR U672 ( .A(n932), .B(n933), .Z(n921) );
  AND U673 ( .A(n934), .B(n931), .Z(n933) );
  XNOR U674 ( .A(n932), .B(n928), .Z(n931) );
  XOR U675 ( .A(n935), .B(n936), .Z(n928) );
  AND U676 ( .A(n937), .B(n938), .Z(n936) );
  XOR U677 ( .A(p_input[1321]), .B(n935), .Z(n938) );
  XOR U678 ( .A(n939), .B(n940), .Z(n935) );
  AND U679 ( .A(n941), .B(n942), .Z(n940) );
  XOR U680 ( .A(n943), .B(n944), .Z(n932) );
  AND U681 ( .A(n945), .B(n942), .Z(n944) );
  XNOR U682 ( .A(n943), .B(n939), .Z(n942) );
  XOR U683 ( .A(n946), .B(n947), .Z(n939) );
  AND U684 ( .A(n948), .B(n949), .Z(n947) );
  XOR U685 ( .A(p_input[1337]), .B(n946), .Z(n949) );
  XOR U686 ( .A(n950), .B(n951), .Z(n946) );
  AND U687 ( .A(n952), .B(n953), .Z(n951) );
  XOR U688 ( .A(n954), .B(n955), .Z(n943) );
  AND U689 ( .A(n956), .B(n953), .Z(n955) );
  XNOR U690 ( .A(n954), .B(n950), .Z(n953) );
  XOR U691 ( .A(n957), .B(n958), .Z(n950) );
  AND U692 ( .A(n959), .B(n960), .Z(n958) );
  XOR U693 ( .A(p_input[1353]), .B(n957), .Z(n960) );
  XOR U694 ( .A(n961), .B(n962), .Z(n957) );
  AND U695 ( .A(n963), .B(n964), .Z(n962) );
  XOR U696 ( .A(n965), .B(n966), .Z(n954) );
  AND U697 ( .A(n967), .B(n964), .Z(n966) );
  XNOR U698 ( .A(n965), .B(n961), .Z(n964) );
  XOR U699 ( .A(n968), .B(n969), .Z(n961) );
  AND U700 ( .A(n970), .B(n971), .Z(n969) );
  XOR U701 ( .A(p_input[1369]), .B(n968), .Z(n971) );
  XOR U702 ( .A(n972), .B(n973), .Z(n968) );
  AND U703 ( .A(n974), .B(n975), .Z(n973) );
  XOR U704 ( .A(n976), .B(n977), .Z(n965) );
  AND U705 ( .A(n978), .B(n975), .Z(n977) );
  XNOR U706 ( .A(n976), .B(n972), .Z(n975) );
  XOR U707 ( .A(n979), .B(n980), .Z(n972) );
  AND U708 ( .A(n981), .B(n982), .Z(n980) );
  XOR U709 ( .A(p_input[1385]), .B(n979), .Z(n982) );
  XOR U710 ( .A(n983), .B(n984), .Z(n979) );
  AND U711 ( .A(n985), .B(n986), .Z(n984) );
  XOR U712 ( .A(n987), .B(n988), .Z(n976) );
  AND U713 ( .A(n989), .B(n986), .Z(n988) );
  XNOR U714 ( .A(n987), .B(n983), .Z(n986) );
  XOR U715 ( .A(n990), .B(n991), .Z(n983) );
  AND U716 ( .A(n992), .B(n993), .Z(n991) );
  XOR U717 ( .A(p_input[1401]), .B(n990), .Z(n993) );
  XOR U718 ( .A(n994), .B(n995), .Z(n990) );
  AND U719 ( .A(n996), .B(n997), .Z(n995) );
  XOR U720 ( .A(n998), .B(n999), .Z(n987) );
  AND U721 ( .A(n1000), .B(n997), .Z(n999) );
  XNOR U722 ( .A(n998), .B(n994), .Z(n997) );
  XOR U723 ( .A(n1001), .B(n1002), .Z(n994) );
  AND U724 ( .A(n1003), .B(n1004), .Z(n1002) );
  XOR U725 ( .A(p_input[1417]), .B(n1001), .Z(n1004) );
  XOR U726 ( .A(n1005), .B(n1006), .Z(n1001) );
  AND U727 ( .A(n1007), .B(n1008), .Z(n1006) );
  XOR U728 ( .A(n1009), .B(n1010), .Z(n998) );
  AND U729 ( .A(n1011), .B(n1008), .Z(n1010) );
  XNOR U730 ( .A(n1009), .B(n1005), .Z(n1008) );
  XOR U731 ( .A(n1012), .B(n1013), .Z(n1005) );
  AND U732 ( .A(n1014), .B(n1015), .Z(n1013) );
  XOR U733 ( .A(p_input[1433]), .B(n1012), .Z(n1015) );
  XOR U734 ( .A(n1016), .B(n1017), .Z(n1012) );
  AND U735 ( .A(n1018), .B(n1019), .Z(n1017) );
  XOR U736 ( .A(n1020), .B(n1021), .Z(n1009) );
  AND U737 ( .A(n1022), .B(n1019), .Z(n1021) );
  XNOR U738 ( .A(n1020), .B(n1016), .Z(n1019) );
  XOR U739 ( .A(n1023), .B(n1024), .Z(n1016) );
  AND U740 ( .A(n1025), .B(n1026), .Z(n1024) );
  XOR U741 ( .A(p_input[1449]), .B(n1023), .Z(n1026) );
  XOR U742 ( .A(n1027), .B(n1028), .Z(n1023) );
  AND U743 ( .A(n1029), .B(n1030), .Z(n1028) );
  XOR U744 ( .A(n1031), .B(n1032), .Z(n1020) );
  AND U745 ( .A(n1033), .B(n1030), .Z(n1032) );
  XNOR U746 ( .A(n1031), .B(n1027), .Z(n1030) );
  XOR U747 ( .A(n1034), .B(n1035), .Z(n1027) );
  AND U748 ( .A(n1036), .B(n1037), .Z(n1035) );
  XOR U749 ( .A(p_input[1465]), .B(n1034), .Z(n1037) );
  XOR U750 ( .A(n1038), .B(n1039), .Z(n1034) );
  AND U751 ( .A(n1040), .B(n1041), .Z(n1039) );
  XOR U752 ( .A(n1042), .B(n1043), .Z(n1031) );
  AND U753 ( .A(n1044), .B(n1041), .Z(n1043) );
  XNOR U754 ( .A(n1042), .B(n1038), .Z(n1041) );
  XOR U755 ( .A(n1045), .B(n1046), .Z(n1038) );
  AND U756 ( .A(n1047), .B(n1048), .Z(n1046) );
  XOR U757 ( .A(p_input[1481]), .B(n1045), .Z(n1048) );
  XOR U758 ( .A(n1049), .B(n1050), .Z(n1045) );
  AND U759 ( .A(n1051), .B(n1052), .Z(n1050) );
  XOR U760 ( .A(n1053), .B(n1054), .Z(n1042) );
  AND U761 ( .A(n1055), .B(n1052), .Z(n1054) );
  XNOR U762 ( .A(n1053), .B(n1049), .Z(n1052) );
  XOR U763 ( .A(n1056), .B(n1057), .Z(n1049) );
  AND U764 ( .A(n1058), .B(n1059), .Z(n1057) );
  XOR U765 ( .A(p_input[1497]), .B(n1056), .Z(n1059) );
  XOR U766 ( .A(n1060), .B(n1061), .Z(n1056) );
  AND U767 ( .A(n1062), .B(n1063), .Z(n1061) );
  XOR U768 ( .A(n1064), .B(n1065), .Z(n1053) );
  AND U769 ( .A(n1066), .B(n1063), .Z(n1065) );
  XNOR U770 ( .A(n1064), .B(n1060), .Z(n1063) );
  XOR U771 ( .A(n1067), .B(n1068), .Z(n1060) );
  AND U772 ( .A(n1069), .B(n1070), .Z(n1068) );
  XOR U773 ( .A(p_input[1513]), .B(n1067), .Z(n1070) );
  XOR U774 ( .A(n1071), .B(n1072), .Z(n1067) );
  AND U775 ( .A(n1073), .B(n1074), .Z(n1072) );
  XOR U776 ( .A(n1075), .B(n1076), .Z(n1064) );
  AND U777 ( .A(n1077), .B(n1074), .Z(n1076) );
  XNOR U778 ( .A(n1075), .B(n1071), .Z(n1074) );
  XOR U779 ( .A(n1078), .B(n1079), .Z(n1071) );
  AND U780 ( .A(n1080), .B(n1081), .Z(n1079) );
  XOR U781 ( .A(p_input[1529]), .B(n1078), .Z(n1081) );
  XOR U782 ( .A(n1082), .B(n1083), .Z(n1078) );
  AND U783 ( .A(n1084), .B(n1085), .Z(n1083) );
  XOR U784 ( .A(n1086), .B(n1087), .Z(n1075) );
  AND U785 ( .A(n1088), .B(n1085), .Z(n1087) );
  XNOR U786 ( .A(n1086), .B(n1082), .Z(n1085) );
  XOR U787 ( .A(n1089), .B(n1090), .Z(n1082) );
  AND U788 ( .A(n1091), .B(n1092), .Z(n1090) );
  XOR U789 ( .A(p_input[1545]), .B(n1089), .Z(n1092) );
  XOR U790 ( .A(n1093), .B(n1094), .Z(n1089) );
  AND U791 ( .A(n1095), .B(n1096), .Z(n1094) );
  XOR U792 ( .A(n1097), .B(n1098), .Z(n1086) );
  AND U793 ( .A(n1099), .B(n1096), .Z(n1098) );
  XNOR U794 ( .A(n1097), .B(n1093), .Z(n1096) );
  XOR U795 ( .A(n1100), .B(n1101), .Z(n1093) );
  AND U796 ( .A(n1102), .B(n1103), .Z(n1101) );
  XOR U797 ( .A(p_input[1561]), .B(n1100), .Z(n1103) );
  XOR U798 ( .A(n1104), .B(n1105), .Z(n1100) );
  AND U799 ( .A(n1106), .B(n1107), .Z(n1105) );
  XOR U800 ( .A(n1108), .B(n1109), .Z(n1097) );
  AND U801 ( .A(n1110), .B(n1107), .Z(n1109) );
  XNOR U802 ( .A(n1108), .B(n1104), .Z(n1107) );
  XOR U803 ( .A(n1111), .B(n1112), .Z(n1104) );
  AND U804 ( .A(n1113), .B(n1114), .Z(n1112) );
  XOR U805 ( .A(p_input[1577]), .B(n1111), .Z(n1114) );
  XOR U806 ( .A(n1115), .B(n1116), .Z(n1111) );
  AND U807 ( .A(n1117), .B(n1118), .Z(n1116) );
  XOR U808 ( .A(n1119), .B(n1120), .Z(n1108) );
  AND U809 ( .A(n1121), .B(n1118), .Z(n1120) );
  XNOR U810 ( .A(n1119), .B(n1115), .Z(n1118) );
  XOR U811 ( .A(n1122), .B(n1123), .Z(n1115) );
  AND U812 ( .A(n1124), .B(n1125), .Z(n1123) );
  XOR U813 ( .A(p_input[1593]), .B(n1122), .Z(n1125) );
  XOR U814 ( .A(n1126), .B(n1127), .Z(n1122) );
  AND U815 ( .A(n1128), .B(n1129), .Z(n1127) );
  XOR U816 ( .A(n1130), .B(n1131), .Z(n1119) );
  AND U817 ( .A(n1132), .B(n1129), .Z(n1131) );
  XNOR U818 ( .A(n1130), .B(n1126), .Z(n1129) );
  XOR U819 ( .A(n1133), .B(n1134), .Z(n1126) );
  AND U820 ( .A(n1135), .B(n1136), .Z(n1134) );
  XOR U821 ( .A(p_input[1609]), .B(n1133), .Z(n1136) );
  XOR U822 ( .A(n1137), .B(n1138), .Z(n1133) );
  AND U823 ( .A(n1139), .B(n1140), .Z(n1138) );
  XOR U824 ( .A(n1141), .B(n1142), .Z(n1130) );
  AND U825 ( .A(n1143), .B(n1140), .Z(n1142) );
  XNOR U826 ( .A(n1141), .B(n1137), .Z(n1140) );
  XOR U827 ( .A(n1144), .B(n1145), .Z(n1137) );
  AND U828 ( .A(n1146), .B(n1147), .Z(n1145) );
  XOR U829 ( .A(p_input[1625]), .B(n1144), .Z(n1147) );
  XOR U830 ( .A(n1148), .B(n1149), .Z(n1144) );
  AND U831 ( .A(n1150), .B(n1151), .Z(n1149) );
  XOR U832 ( .A(n1152), .B(n1153), .Z(n1141) );
  AND U833 ( .A(n1154), .B(n1151), .Z(n1153) );
  XNOR U834 ( .A(n1152), .B(n1148), .Z(n1151) );
  XOR U835 ( .A(n1155), .B(n1156), .Z(n1148) );
  AND U836 ( .A(n1157), .B(n1158), .Z(n1156) );
  XOR U837 ( .A(p_input[1641]), .B(n1155), .Z(n1158) );
  XOR U838 ( .A(n1159), .B(n1160), .Z(n1155) );
  AND U839 ( .A(n1161), .B(n1162), .Z(n1160) );
  XOR U840 ( .A(n1163), .B(n1164), .Z(n1152) );
  AND U841 ( .A(n1165), .B(n1162), .Z(n1164) );
  XNOR U842 ( .A(n1163), .B(n1159), .Z(n1162) );
  XOR U843 ( .A(n1166), .B(n1167), .Z(n1159) );
  AND U844 ( .A(n1168), .B(n1169), .Z(n1167) );
  XOR U845 ( .A(p_input[1657]), .B(n1166), .Z(n1169) );
  XOR U846 ( .A(n1170), .B(n1171), .Z(n1166) );
  AND U847 ( .A(n1172), .B(n1173), .Z(n1171) );
  XOR U848 ( .A(n1174), .B(n1175), .Z(n1163) );
  AND U849 ( .A(n1176), .B(n1173), .Z(n1175) );
  XNOR U850 ( .A(n1174), .B(n1170), .Z(n1173) );
  XOR U851 ( .A(n1177), .B(n1178), .Z(n1170) );
  AND U852 ( .A(n1179), .B(n1180), .Z(n1178) );
  XOR U853 ( .A(p_input[1673]), .B(n1177), .Z(n1180) );
  XOR U854 ( .A(n1181), .B(n1182), .Z(n1177) );
  AND U855 ( .A(n1183), .B(n1184), .Z(n1182) );
  XOR U856 ( .A(n1185), .B(n1186), .Z(n1174) );
  AND U857 ( .A(n1187), .B(n1184), .Z(n1186) );
  XNOR U858 ( .A(n1185), .B(n1181), .Z(n1184) );
  XOR U859 ( .A(n1188), .B(n1189), .Z(n1181) );
  AND U860 ( .A(n1190), .B(n1191), .Z(n1189) );
  XOR U861 ( .A(p_input[1689]), .B(n1188), .Z(n1191) );
  XOR U862 ( .A(n1192), .B(n1193), .Z(n1188) );
  AND U863 ( .A(n1194), .B(n1195), .Z(n1193) );
  XOR U864 ( .A(n1196), .B(n1197), .Z(n1185) );
  AND U865 ( .A(n1198), .B(n1195), .Z(n1197) );
  XNOR U866 ( .A(n1196), .B(n1192), .Z(n1195) );
  XOR U867 ( .A(n1199), .B(n1200), .Z(n1192) );
  AND U868 ( .A(n1201), .B(n1202), .Z(n1200) );
  XOR U869 ( .A(p_input[1705]), .B(n1199), .Z(n1202) );
  XOR U870 ( .A(n1203), .B(n1204), .Z(n1199) );
  AND U871 ( .A(n1205), .B(n1206), .Z(n1204) );
  XOR U872 ( .A(n1207), .B(n1208), .Z(n1196) );
  AND U873 ( .A(n1209), .B(n1206), .Z(n1208) );
  XNOR U874 ( .A(n1207), .B(n1203), .Z(n1206) );
  XOR U875 ( .A(n1210), .B(n1211), .Z(n1203) );
  AND U876 ( .A(n1212), .B(n1213), .Z(n1211) );
  XOR U877 ( .A(p_input[1721]), .B(n1210), .Z(n1213) );
  XOR U878 ( .A(n1214), .B(n1215), .Z(n1210) );
  AND U879 ( .A(n1216), .B(n1217), .Z(n1215) );
  XOR U880 ( .A(n1218), .B(n1219), .Z(n1207) );
  AND U881 ( .A(n1220), .B(n1217), .Z(n1219) );
  XNOR U882 ( .A(n1218), .B(n1214), .Z(n1217) );
  XOR U883 ( .A(n1221), .B(n1222), .Z(n1214) );
  AND U884 ( .A(n1223), .B(n1224), .Z(n1222) );
  XOR U885 ( .A(p_input[1737]), .B(n1221), .Z(n1224) );
  XOR U886 ( .A(n1225), .B(n1226), .Z(n1221) );
  AND U887 ( .A(n1227), .B(n1228), .Z(n1226) );
  XOR U888 ( .A(n1229), .B(n1230), .Z(n1218) );
  AND U889 ( .A(n1231), .B(n1228), .Z(n1230) );
  XNOR U890 ( .A(n1229), .B(n1225), .Z(n1228) );
  XOR U891 ( .A(n1232), .B(n1233), .Z(n1225) );
  AND U892 ( .A(n1234), .B(n1235), .Z(n1233) );
  XOR U893 ( .A(p_input[1753]), .B(n1232), .Z(n1235) );
  XOR U894 ( .A(n1236), .B(n1237), .Z(n1232) );
  AND U895 ( .A(n1238), .B(n1239), .Z(n1237) );
  XOR U896 ( .A(n1240), .B(n1241), .Z(n1229) );
  AND U897 ( .A(n1242), .B(n1239), .Z(n1241) );
  XNOR U898 ( .A(n1240), .B(n1236), .Z(n1239) );
  XOR U899 ( .A(n1243), .B(n1244), .Z(n1236) );
  AND U900 ( .A(n1245), .B(n1246), .Z(n1244) );
  XOR U901 ( .A(p_input[1769]), .B(n1243), .Z(n1246) );
  XOR U902 ( .A(n1247), .B(n1248), .Z(n1243) );
  AND U903 ( .A(n1249), .B(n1250), .Z(n1248) );
  XOR U904 ( .A(n1251), .B(n1252), .Z(n1240) );
  AND U905 ( .A(n1253), .B(n1250), .Z(n1252) );
  XNOR U906 ( .A(n1251), .B(n1247), .Z(n1250) );
  XOR U907 ( .A(n1254), .B(n1255), .Z(n1247) );
  AND U908 ( .A(n1256), .B(n1257), .Z(n1255) );
  XOR U909 ( .A(p_input[1785]), .B(n1254), .Z(n1257) );
  XOR U910 ( .A(n1258), .B(n1259), .Z(n1254) );
  AND U911 ( .A(n1260), .B(n1261), .Z(n1259) );
  XOR U912 ( .A(n1262), .B(n1263), .Z(n1251) );
  AND U913 ( .A(n1264), .B(n1261), .Z(n1263) );
  XNOR U914 ( .A(n1262), .B(n1258), .Z(n1261) );
  XOR U915 ( .A(n1265), .B(n1266), .Z(n1258) );
  AND U916 ( .A(n1267), .B(n1268), .Z(n1266) );
  XOR U917 ( .A(p_input[1801]), .B(n1265), .Z(n1268) );
  XOR U918 ( .A(n1269), .B(n1270), .Z(n1265) );
  AND U919 ( .A(n1271), .B(n1272), .Z(n1270) );
  XOR U920 ( .A(n1273), .B(n1274), .Z(n1262) );
  AND U921 ( .A(n1275), .B(n1272), .Z(n1274) );
  XNOR U922 ( .A(n1273), .B(n1269), .Z(n1272) );
  XOR U923 ( .A(n1276), .B(n1277), .Z(n1269) );
  AND U924 ( .A(n1278), .B(n1279), .Z(n1277) );
  XOR U925 ( .A(p_input[1817]), .B(n1276), .Z(n1279) );
  XOR U926 ( .A(n1280), .B(n1281), .Z(n1276) );
  AND U927 ( .A(n1282), .B(n1283), .Z(n1281) );
  XOR U928 ( .A(n1284), .B(n1285), .Z(n1273) );
  AND U929 ( .A(n1286), .B(n1283), .Z(n1285) );
  XNOR U930 ( .A(n1284), .B(n1280), .Z(n1283) );
  XOR U931 ( .A(n1287), .B(n1288), .Z(n1280) );
  AND U932 ( .A(n1289), .B(n1290), .Z(n1288) );
  XOR U933 ( .A(p_input[1833]), .B(n1287), .Z(n1290) );
  XOR U934 ( .A(n1291), .B(n1292), .Z(n1287) );
  AND U935 ( .A(n1293), .B(n1294), .Z(n1292) );
  XOR U936 ( .A(n1295), .B(n1296), .Z(n1284) );
  AND U937 ( .A(n1297), .B(n1294), .Z(n1296) );
  XNOR U938 ( .A(n1295), .B(n1291), .Z(n1294) );
  XOR U939 ( .A(n1298), .B(n1299), .Z(n1291) );
  AND U940 ( .A(n1300), .B(n1301), .Z(n1299) );
  XOR U941 ( .A(p_input[1849]), .B(n1298), .Z(n1301) );
  XOR U942 ( .A(n1302), .B(n1303), .Z(n1298) );
  AND U943 ( .A(n1304), .B(n1305), .Z(n1303) );
  XOR U944 ( .A(n1306), .B(n1307), .Z(n1295) );
  AND U945 ( .A(n1308), .B(n1305), .Z(n1307) );
  XNOR U946 ( .A(n1306), .B(n1302), .Z(n1305) );
  XOR U947 ( .A(n1309), .B(n1310), .Z(n1302) );
  AND U948 ( .A(n1311), .B(n1312), .Z(n1310) );
  XOR U949 ( .A(p_input[1865]), .B(n1309), .Z(n1312) );
  XOR U950 ( .A(n1313), .B(n1314), .Z(n1309) );
  AND U951 ( .A(n1315), .B(n1316), .Z(n1314) );
  XOR U952 ( .A(n1317), .B(n1318), .Z(n1306) );
  AND U953 ( .A(n1319), .B(n1316), .Z(n1318) );
  XNOR U954 ( .A(n1317), .B(n1313), .Z(n1316) );
  XOR U955 ( .A(n1320), .B(n1321), .Z(n1313) );
  AND U956 ( .A(n1322), .B(n1323), .Z(n1321) );
  XOR U957 ( .A(p_input[1881]), .B(n1320), .Z(n1323) );
  XOR U958 ( .A(n1324), .B(n1325), .Z(n1320) );
  AND U959 ( .A(n1326), .B(n1327), .Z(n1325) );
  XOR U960 ( .A(n1328), .B(n1329), .Z(n1317) );
  AND U961 ( .A(n1330), .B(n1327), .Z(n1329) );
  XNOR U962 ( .A(n1328), .B(n1324), .Z(n1327) );
  XOR U963 ( .A(n1331), .B(n1332), .Z(n1324) );
  AND U964 ( .A(n1333), .B(n1334), .Z(n1332) );
  XOR U965 ( .A(p_input[1897]), .B(n1331), .Z(n1334) );
  XOR U966 ( .A(n1335), .B(n1336), .Z(n1331) );
  AND U967 ( .A(n1337), .B(n1338), .Z(n1336) );
  XOR U968 ( .A(n1339), .B(n1340), .Z(n1328) );
  AND U969 ( .A(n1341), .B(n1338), .Z(n1340) );
  XNOR U970 ( .A(n1339), .B(n1335), .Z(n1338) );
  XOR U971 ( .A(n1342), .B(n1343), .Z(n1335) );
  AND U972 ( .A(n1344), .B(n1345), .Z(n1343) );
  XOR U973 ( .A(p_input[1913]), .B(n1342), .Z(n1345) );
  XOR U974 ( .A(n1346), .B(n1347), .Z(n1342) );
  AND U975 ( .A(n1348), .B(n1349), .Z(n1347) );
  XOR U976 ( .A(n1350), .B(n1351), .Z(n1339) );
  AND U977 ( .A(n1352), .B(n1349), .Z(n1351) );
  XNOR U978 ( .A(n1350), .B(n1346), .Z(n1349) );
  XOR U979 ( .A(n1353), .B(n1354), .Z(n1346) );
  AND U980 ( .A(n1355), .B(n1356), .Z(n1354) );
  XOR U981 ( .A(p_input[1929]), .B(n1353), .Z(n1356) );
  XOR U982 ( .A(n1357), .B(n1358), .Z(n1353) );
  AND U983 ( .A(n1359), .B(n1360), .Z(n1358) );
  XOR U984 ( .A(n1361), .B(n1362), .Z(n1350) );
  AND U985 ( .A(n1363), .B(n1360), .Z(n1362) );
  XNOR U986 ( .A(n1361), .B(n1357), .Z(n1360) );
  XOR U987 ( .A(n1364), .B(n1365), .Z(n1357) );
  AND U988 ( .A(n1366), .B(n1367), .Z(n1365) );
  XOR U989 ( .A(p_input[1945]), .B(n1364), .Z(n1367) );
  XOR U990 ( .A(n1368), .B(n1369), .Z(n1364) );
  AND U991 ( .A(n1370), .B(n1371), .Z(n1369) );
  XOR U992 ( .A(n1372), .B(n1373), .Z(n1361) );
  AND U993 ( .A(n1374), .B(n1371), .Z(n1373) );
  XNOR U994 ( .A(n1372), .B(n1368), .Z(n1371) );
  XOR U995 ( .A(n1375), .B(n1376), .Z(n1368) );
  AND U996 ( .A(n1377), .B(n1378), .Z(n1376) );
  XOR U997 ( .A(p_input[1961]), .B(n1375), .Z(n1378) );
  XOR U998 ( .A(n1379), .B(n1380), .Z(n1375) );
  AND U999 ( .A(n1381), .B(n1382), .Z(n1380) );
  XOR U1000 ( .A(n1383), .B(n1384), .Z(n1372) );
  AND U1001 ( .A(n1385), .B(n1382), .Z(n1384) );
  XNOR U1002 ( .A(n1383), .B(n1379), .Z(n1382) );
  XOR U1003 ( .A(n1386), .B(n1387), .Z(n1379) );
  AND U1004 ( .A(n1388), .B(n1389), .Z(n1387) );
  XOR U1005 ( .A(p_input[1977]), .B(n1386), .Z(n1389) );
  XOR U1006 ( .A(n1390), .B(n1391), .Z(n1386) );
  AND U1007 ( .A(n1392), .B(n1393), .Z(n1391) );
  XOR U1008 ( .A(n1394), .B(n1395), .Z(n1383) );
  AND U1009 ( .A(n1396), .B(n1393), .Z(n1395) );
  XNOR U1010 ( .A(n1394), .B(n1390), .Z(n1393) );
  XOR U1011 ( .A(n1397), .B(n1398), .Z(n1390) );
  AND U1012 ( .A(n1399), .B(n1400), .Z(n1398) );
  XOR U1013 ( .A(p_input[1993]), .B(n1397), .Z(n1400) );
  XOR U1014 ( .A(n1401), .B(n1402), .Z(n1397) );
  AND U1015 ( .A(n1403), .B(n1404), .Z(n1402) );
  XOR U1016 ( .A(n1405), .B(n1406), .Z(n1394) );
  AND U1017 ( .A(n1407), .B(n1404), .Z(n1406) );
  XNOR U1018 ( .A(n1405), .B(n1401), .Z(n1404) );
  XOR U1019 ( .A(n1408), .B(n1409), .Z(n1401) );
  AND U1020 ( .A(n1410), .B(n1411), .Z(n1409) );
  XOR U1021 ( .A(p_input[2009]), .B(n1408), .Z(n1411) );
  XNOR U1022 ( .A(n1412), .B(n1413), .Z(n1408) );
  AND U1023 ( .A(n1414), .B(n1415), .Z(n1413) );
  XNOR U1024 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n1416), .Z(n1405) );
  AND U1025 ( .A(n1417), .B(n1415), .Z(n1416) );
  XOR U1026 ( .A(n1418), .B(n1412), .Z(n1415) );
  XOR U1027 ( .A(n3), .B(n1419), .Z(o[24]) );
  AND U1028 ( .A(n30), .B(n1420), .Z(n3) );
  XOR U1029 ( .A(n4), .B(n1419), .Z(n1420) );
  XOR U1030 ( .A(n1421), .B(n1422), .Z(n1419) );
  AND U1031 ( .A(n34), .B(n1423), .Z(n1422) );
  XOR U1032 ( .A(p_input[8]), .B(n1421), .Z(n1423) );
  XOR U1033 ( .A(n1424), .B(n1425), .Z(n1421) );
  AND U1034 ( .A(n38), .B(n1426), .Z(n1425) );
  XOR U1035 ( .A(n1427), .B(n1428), .Z(n4) );
  AND U1036 ( .A(n42), .B(n1426), .Z(n1428) );
  XNOR U1037 ( .A(n1429), .B(n1424), .Z(n1426) );
  XOR U1038 ( .A(n1430), .B(n1431), .Z(n1424) );
  AND U1039 ( .A(n46), .B(n1432), .Z(n1431) );
  XOR U1040 ( .A(p_input[24]), .B(n1430), .Z(n1432) );
  XOR U1041 ( .A(n1433), .B(n1434), .Z(n1430) );
  AND U1042 ( .A(n50), .B(n1435), .Z(n1434) );
  IV U1043 ( .A(n1427), .Z(n1429) );
  XNOR U1044 ( .A(n1436), .B(n1437), .Z(n1427) );
  AND U1045 ( .A(n54), .B(n1435), .Z(n1437) );
  XNOR U1046 ( .A(n1436), .B(n1433), .Z(n1435) );
  XOR U1047 ( .A(n1438), .B(n1439), .Z(n1433) );
  AND U1048 ( .A(n57), .B(n1440), .Z(n1439) );
  XOR U1049 ( .A(p_input[40]), .B(n1438), .Z(n1440) );
  XOR U1050 ( .A(n1441), .B(n1442), .Z(n1438) );
  AND U1051 ( .A(n61), .B(n1443), .Z(n1442) );
  XOR U1052 ( .A(n1444), .B(n1445), .Z(n1436) );
  AND U1053 ( .A(n65), .B(n1443), .Z(n1445) );
  XNOR U1054 ( .A(n1444), .B(n1441), .Z(n1443) );
  XOR U1055 ( .A(n1446), .B(n1447), .Z(n1441) );
  AND U1056 ( .A(n68), .B(n1448), .Z(n1447) );
  XOR U1057 ( .A(p_input[56]), .B(n1446), .Z(n1448) );
  XOR U1058 ( .A(n1449), .B(n1450), .Z(n1446) );
  AND U1059 ( .A(n72), .B(n1451), .Z(n1450) );
  XOR U1060 ( .A(n1452), .B(n1453), .Z(n1444) );
  AND U1061 ( .A(n76), .B(n1451), .Z(n1453) );
  XNOR U1062 ( .A(n1452), .B(n1449), .Z(n1451) );
  XOR U1063 ( .A(n1454), .B(n1455), .Z(n1449) );
  AND U1064 ( .A(n79), .B(n1456), .Z(n1455) );
  XOR U1065 ( .A(p_input[72]), .B(n1454), .Z(n1456) );
  XOR U1066 ( .A(n1457), .B(n1458), .Z(n1454) );
  AND U1067 ( .A(n83), .B(n1459), .Z(n1458) );
  XOR U1068 ( .A(n1460), .B(n1461), .Z(n1452) );
  AND U1069 ( .A(n87), .B(n1459), .Z(n1461) );
  XNOR U1070 ( .A(n1460), .B(n1457), .Z(n1459) );
  XOR U1071 ( .A(n1462), .B(n1463), .Z(n1457) );
  AND U1072 ( .A(n90), .B(n1464), .Z(n1463) );
  XOR U1073 ( .A(p_input[88]), .B(n1462), .Z(n1464) );
  XOR U1074 ( .A(n1465), .B(n1466), .Z(n1462) );
  AND U1075 ( .A(n94), .B(n1467), .Z(n1466) );
  XOR U1076 ( .A(n1468), .B(n1469), .Z(n1460) );
  AND U1077 ( .A(n98), .B(n1467), .Z(n1469) );
  XNOR U1078 ( .A(n1468), .B(n1465), .Z(n1467) );
  XOR U1079 ( .A(n1470), .B(n1471), .Z(n1465) );
  AND U1080 ( .A(n101), .B(n1472), .Z(n1471) );
  XOR U1081 ( .A(p_input[104]), .B(n1470), .Z(n1472) );
  XOR U1082 ( .A(n1473), .B(n1474), .Z(n1470) );
  AND U1083 ( .A(n105), .B(n1475), .Z(n1474) );
  XOR U1084 ( .A(n1476), .B(n1477), .Z(n1468) );
  AND U1085 ( .A(n109), .B(n1475), .Z(n1477) );
  XNOR U1086 ( .A(n1476), .B(n1473), .Z(n1475) );
  XOR U1087 ( .A(n1478), .B(n1479), .Z(n1473) );
  AND U1088 ( .A(n112), .B(n1480), .Z(n1479) );
  XOR U1089 ( .A(p_input[120]), .B(n1478), .Z(n1480) );
  XOR U1090 ( .A(n1481), .B(n1482), .Z(n1478) );
  AND U1091 ( .A(n116), .B(n1483), .Z(n1482) );
  XOR U1092 ( .A(n1484), .B(n1485), .Z(n1476) );
  AND U1093 ( .A(n120), .B(n1483), .Z(n1485) );
  XNOR U1094 ( .A(n1484), .B(n1481), .Z(n1483) );
  XOR U1095 ( .A(n1486), .B(n1487), .Z(n1481) );
  AND U1096 ( .A(n123), .B(n1488), .Z(n1487) );
  XOR U1097 ( .A(p_input[136]), .B(n1486), .Z(n1488) );
  XOR U1098 ( .A(n1489), .B(n1490), .Z(n1486) );
  AND U1099 ( .A(n127), .B(n1491), .Z(n1490) );
  XOR U1100 ( .A(n1492), .B(n1493), .Z(n1484) );
  AND U1101 ( .A(n131), .B(n1491), .Z(n1493) );
  XNOR U1102 ( .A(n1492), .B(n1489), .Z(n1491) );
  XOR U1103 ( .A(n1494), .B(n1495), .Z(n1489) );
  AND U1104 ( .A(n134), .B(n1496), .Z(n1495) );
  XOR U1105 ( .A(p_input[152]), .B(n1494), .Z(n1496) );
  XOR U1106 ( .A(n1497), .B(n1498), .Z(n1494) );
  AND U1107 ( .A(n138), .B(n1499), .Z(n1498) );
  XOR U1108 ( .A(n1500), .B(n1501), .Z(n1492) );
  AND U1109 ( .A(n142), .B(n1499), .Z(n1501) );
  XNOR U1110 ( .A(n1500), .B(n1497), .Z(n1499) );
  XOR U1111 ( .A(n1502), .B(n1503), .Z(n1497) );
  AND U1112 ( .A(n145), .B(n1504), .Z(n1503) );
  XOR U1113 ( .A(p_input[168]), .B(n1502), .Z(n1504) );
  XOR U1114 ( .A(n1505), .B(n1506), .Z(n1502) );
  AND U1115 ( .A(n149), .B(n1507), .Z(n1506) );
  XOR U1116 ( .A(n1508), .B(n1509), .Z(n1500) );
  AND U1117 ( .A(n153), .B(n1507), .Z(n1509) );
  XNOR U1118 ( .A(n1508), .B(n1505), .Z(n1507) );
  XOR U1119 ( .A(n1510), .B(n1511), .Z(n1505) );
  AND U1120 ( .A(n156), .B(n1512), .Z(n1511) );
  XOR U1121 ( .A(p_input[184]), .B(n1510), .Z(n1512) );
  XOR U1122 ( .A(n1513), .B(n1514), .Z(n1510) );
  AND U1123 ( .A(n160), .B(n1515), .Z(n1514) );
  XOR U1124 ( .A(n1516), .B(n1517), .Z(n1508) );
  AND U1125 ( .A(n164), .B(n1515), .Z(n1517) );
  XNOR U1126 ( .A(n1516), .B(n1513), .Z(n1515) );
  XOR U1127 ( .A(n1518), .B(n1519), .Z(n1513) );
  AND U1128 ( .A(n167), .B(n1520), .Z(n1519) );
  XOR U1129 ( .A(p_input[200]), .B(n1518), .Z(n1520) );
  XOR U1130 ( .A(n1521), .B(n1522), .Z(n1518) );
  AND U1131 ( .A(n171), .B(n1523), .Z(n1522) );
  XOR U1132 ( .A(n1524), .B(n1525), .Z(n1516) );
  AND U1133 ( .A(n175), .B(n1523), .Z(n1525) );
  XNOR U1134 ( .A(n1524), .B(n1521), .Z(n1523) );
  XOR U1135 ( .A(n1526), .B(n1527), .Z(n1521) );
  AND U1136 ( .A(n178), .B(n1528), .Z(n1527) );
  XOR U1137 ( .A(p_input[216]), .B(n1526), .Z(n1528) );
  XOR U1138 ( .A(n1529), .B(n1530), .Z(n1526) );
  AND U1139 ( .A(n182), .B(n1531), .Z(n1530) );
  XOR U1140 ( .A(n1532), .B(n1533), .Z(n1524) );
  AND U1141 ( .A(n186), .B(n1531), .Z(n1533) );
  XNOR U1142 ( .A(n1532), .B(n1529), .Z(n1531) );
  XOR U1143 ( .A(n1534), .B(n1535), .Z(n1529) );
  AND U1144 ( .A(n189), .B(n1536), .Z(n1535) );
  XOR U1145 ( .A(p_input[232]), .B(n1534), .Z(n1536) );
  XOR U1146 ( .A(n1537), .B(n1538), .Z(n1534) );
  AND U1147 ( .A(n193), .B(n1539), .Z(n1538) );
  XOR U1148 ( .A(n1540), .B(n1541), .Z(n1532) );
  AND U1149 ( .A(n197), .B(n1539), .Z(n1541) );
  XNOR U1150 ( .A(n1540), .B(n1537), .Z(n1539) );
  XOR U1151 ( .A(n1542), .B(n1543), .Z(n1537) );
  AND U1152 ( .A(n200), .B(n1544), .Z(n1543) );
  XOR U1153 ( .A(p_input[248]), .B(n1542), .Z(n1544) );
  XOR U1154 ( .A(n1545), .B(n1546), .Z(n1542) );
  AND U1155 ( .A(n204), .B(n1547), .Z(n1546) );
  XOR U1156 ( .A(n1548), .B(n1549), .Z(n1540) );
  AND U1157 ( .A(n208), .B(n1547), .Z(n1549) );
  XNOR U1158 ( .A(n1548), .B(n1545), .Z(n1547) );
  XOR U1159 ( .A(n1550), .B(n1551), .Z(n1545) );
  AND U1160 ( .A(n211), .B(n1552), .Z(n1551) );
  XOR U1161 ( .A(p_input[264]), .B(n1550), .Z(n1552) );
  XOR U1162 ( .A(n1553), .B(n1554), .Z(n1550) );
  AND U1163 ( .A(n215), .B(n1555), .Z(n1554) );
  XOR U1164 ( .A(n1556), .B(n1557), .Z(n1548) );
  AND U1165 ( .A(n219), .B(n1555), .Z(n1557) );
  XNOR U1166 ( .A(n1556), .B(n1553), .Z(n1555) );
  XOR U1167 ( .A(n1558), .B(n1559), .Z(n1553) );
  AND U1168 ( .A(n222), .B(n1560), .Z(n1559) );
  XOR U1169 ( .A(p_input[280]), .B(n1558), .Z(n1560) );
  XOR U1170 ( .A(n1561), .B(n1562), .Z(n1558) );
  AND U1171 ( .A(n226), .B(n1563), .Z(n1562) );
  XOR U1172 ( .A(n1564), .B(n1565), .Z(n1556) );
  AND U1173 ( .A(n230), .B(n1563), .Z(n1565) );
  XNOR U1174 ( .A(n1564), .B(n1561), .Z(n1563) );
  XOR U1175 ( .A(n1566), .B(n1567), .Z(n1561) );
  AND U1176 ( .A(n233), .B(n1568), .Z(n1567) );
  XOR U1177 ( .A(p_input[296]), .B(n1566), .Z(n1568) );
  XOR U1178 ( .A(n1569), .B(n1570), .Z(n1566) );
  AND U1179 ( .A(n237), .B(n1571), .Z(n1570) );
  XOR U1180 ( .A(n1572), .B(n1573), .Z(n1564) );
  AND U1181 ( .A(n241), .B(n1571), .Z(n1573) );
  XNOR U1182 ( .A(n1572), .B(n1569), .Z(n1571) );
  XOR U1183 ( .A(n1574), .B(n1575), .Z(n1569) );
  AND U1184 ( .A(n244), .B(n1576), .Z(n1575) );
  XOR U1185 ( .A(p_input[312]), .B(n1574), .Z(n1576) );
  XOR U1186 ( .A(n1577), .B(n1578), .Z(n1574) );
  AND U1187 ( .A(n248), .B(n1579), .Z(n1578) );
  XOR U1188 ( .A(n1580), .B(n1581), .Z(n1572) );
  AND U1189 ( .A(n252), .B(n1579), .Z(n1581) );
  XNOR U1190 ( .A(n1580), .B(n1577), .Z(n1579) );
  XOR U1191 ( .A(n1582), .B(n1583), .Z(n1577) );
  AND U1192 ( .A(n255), .B(n1584), .Z(n1583) );
  XOR U1193 ( .A(p_input[328]), .B(n1582), .Z(n1584) );
  XOR U1194 ( .A(n1585), .B(n1586), .Z(n1582) );
  AND U1195 ( .A(n259), .B(n1587), .Z(n1586) );
  XOR U1196 ( .A(n1588), .B(n1589), .Z(n1580) );
  AND U1197 ( .A(n263), .B(n1587), .Z(n1589) );
  XNOR U1198 ( .A(n1588), .B(n1585), .Z(n1587) );
  XOR U1199 ( .A(n1590), .B(n1591), .Z(n1585) );
  AND U1200 ( .A(n266), .B(n1592), .Z(n1591) );
  XOR U1201 ( .A(p_input[344]), .B(n1590), .Z(n1592) );
  XOR U1202 ( .A(n1593), .B(n1594), .Z(n1590) );
  AND U1203 ( .A(n270), .B(n1595), .Z(n1594) );
  XOR U1204 ( .A(n1596), .B(n1597), .Z(n1588) );
  AND U1205 ( .A(n274), .B(n1595), .Z(n1597) );
  XNOR U1206 ( .A(n1596), .B(n1593), .Z(n1595) );
  XOR U1207 ( .A(n1598), .B(n1599), .Z(n1593) );
  AND U1208 ( .A(n277), .B(n1600), .Z(n1599) );
  XOR U1209 ( .A(p_input[360]), .B(n1598), .Z(n1600) );
  XOR U1210 ( .A(n1601), .B(n1602), .Z(n1598) );
  AND U1211 ( .A(n281), .B(n1603), .Z(n1602) );
  XOR U1212 ( .A(n1604), .B(n1605), .Z(n1596) );
  AND U1213 ( .A(n285), .B(n1603), .Z(n1605) );
  XNOR U1214 ( .A(n1604), .B(n1601), .Z(n1603) );
  XOR U1215 ( .A(n1606), .B(n1607), .Z(n1601) );
  AND U1216 ( .A(n288), .B(n1608), .Z(n1607) );
  XOR U1217 ( .A(p_input[376]), .B(n1606), .Z(n1608) );
  XOR U1218 ( .A(n1609), .B(n1610), .Z(n1606) );
  AND U1219 ( .A(n292), .B(n1611), .Z(n1610) );
  XOR U1220 ( .A(n1612), .B(n1613), .Z(n1604) );
  AND U1221 ( .A(n296), .B(n1611), .Z(n1613) );
  XNOR U1222 ( .A(n1612), .B(n1609), .Z(n1611) );
  XOR U1223 ( .A(n1614), .B(n1615), .Z(n1609) );
  AND U1224 ( .A(n299), .B(n1616), .Z(n1615) );
  XOR U1225 ( .A(p_input[392]), .B(n1614), .Z(n1616) );
  XOR U1226 ( .A(n1617), .B(n1618), .Z(n1614) );
  AND U1227 ( .A(n303), .B(n1619), .Z(n1618) );
  XOR U1228 ( .A(n1620), .B(n1621), .Z(n1612) );
  AND U1229 ( .A(n307), .B(n1619), .Z(n1621) );
  XNOR U1230 ( .A(n1620), .B(n1617), .Z(n1619) );
  XOR U1231 ( .A(n1622), .B(n1623), .Z(n1617) );
  AND U1232 ( .A(n310), .B(n1624), .Z(n1623) );
  XOR U1233 ( .A(p_input[408]), .B(n1622), .Z(n1624) );
  XOR U1234 ( .A(n1625), .B(n1626), .Z(n1622) );
  AND U1235 ( .A(n314), .B(n1627), .Z(n1626) );
  XOR U1236 ( .A(n1628), .B(n1629), .Z(n1620) );
  AND U1237 ( .A(n318), .B(n1627), .Z(n1629) );
  XNOR U1238 ( .A(n1628), .B(n1625), .Z(n1627) );
  XOR U1239 ( .A(n1630), .B(n1631), .Z(n1625) );
  AND U1240 ( .A(n321), .B(n1632), .Z(n1631) );
  XOR U1241 ( .A(p_input[424]), .B(n1630), .Z(n1632) );
  XOR U1242 ( .A(n1633), .B(n1634), .Z(n1630) );
  AND U1243 ( .A(n325), .B(n1635), .Z(n1634) );
  XOR U1244 ( .A(n1636), .B(n1637), .Z(n1628) );
  AND U1245 ( .A(n329), .B(n1635), .Z(n1637) );
  XNOR U1246 ( .A(n1636), .B(n1633), .Z(n1635) );
  XOR U1247 ( .A(n1638), .B(n1639), .Z(n1633) );
  AND U1248 ( .A(n332), .B(n1640), .Z(n1639) );
  XOR U1249 ( .A(p_input[440]), .B(n1638), .Z(n1640) );
  XOR U1250 ( .A(n1641), .B(n1642), .Z(n1638) );
  AND U1251 ( .A(n336), .B(n1643), .Z(n1642) );
  XOR U1252 ( .A(n1644), .B(n1645), .Z(n1636) );
  AND U1253 ( .A(n340), .B(n1643), .Z(n1645) );
  XNOR U1254 ( .A(n1644), .B(n1641), .Z(n1643) );
  XOR U1255 ( .A(n1646), .B(n1647), .Z(n1641) );
  AND U1256 ( .A(n343), .B(n1648), .Z(n1647) );
  XOR U1257 ( .A(p_input[456]), .B(n1646), .Z(n1648) );
  XOR U1258 ( .A(n1649), .B(n1650), .Z(n1646) );
  AND U1259 ( .A(n347), .B(n1651), .Z(n1650) );
  XOR U1260 ( .A(n1652), .B(n1653), .Z(n1644) );
  AND U1261 ( .A(n351), .B(n1651), .Z(n1653) );
  XNOR U1262 ( .A(n1652), .B(n1649), .Z(n1651) );
  XOR U1263 ( .A(n1654), .B(n1655), .Z(n1649) );
  AND U1264 ( .A(n354), .B(n1656), .Z(n1655) );
  XOR U1265 ( .A(p_input[472]), .B(n1654), .Z(n1656) );
  XOR U1266 ( .A(n1657), .B(n1658), .Z(n1654) );
  AND U1267 ( .A(n358), .B(n1659), .Z(n1658) );
  XOR U1268 ( .A(n1660), .B(n1661), .Z(n1652) );
  AND U1269 ( .A(n362), .B(n1659), .Z(n1661) );
  XNOR U1270 ( .A(n1660), .B(n1657), .Z(n1659) );
  XOR U1271 ( .A(n1662), .B(n1663), .Z(n1657) );
  AND U1272 ( .A(n365), .B(n1664), .Z(n1663) );
  XOR U1273 ( .A(p_input[488]), .B(n1662), .Z(n1664) );
  XOR U1274 ( .A(n1665), .B(n1666), .Z(n1662) );
  AND U1275 ( .A(n369), .B(n1667), .Z(n1666) );
  XOR U1276 ( .A(n1668), .B(n1669), .Z(n1660) );
  AND U1277 ( .A(n373), .B(n1667), .Z(n1669) );
  XNOR U1278 ( .A(n1668), .B(n1665), .Z(n1667) );
  XOR U1279 ( .A(n1670), .B(n1671), .Z(n1665) );
  AND U1280 ( .A(n376), .B(n1672), .Z(n1671) );
  XOR U1281 ( .A(p_input[504]), .B(n1670), .Z(n1672) );
  XOR U1282 ( .A(n1673), .B(n1674), .Z(n1670) );
  AND U1283 ( .A(n380), .B(n1675), .Z(n1674) );
  XOR U1284 ( .A(n1676), .B(n1677), .Z(n1668) );
  AND U1285 ( .A(n384), .B(n1675), .Z(n1677) );
  XNOR U1286 ( .A(n1676), .B(n1673), .Z(n1675) );
  XOR U1287 ( .A(n1678), .B(n1679), .Z(n1673) );
  AND U1288 ( .A(n387), .B(n1680), .Z(n1679) );
  XOR U1289 ( .A(p_input[520]), .B(n1678), .Z(n1680) );
  XOR U1290 ( .A(n1681), .B(n1682), .Z(n1678) );
  AND U1291 ( .A(n391), .B(n1683), .Z(n1682) );
  XOR U1292 ( .A(n1684), .B(n1685), .Z(n1676) );
  AND U1293 ( .A(n395), .B(n1683), .Z(n1685) );
  XNOR U1294 ( .A(n1684), .B(n1681), .Z(n1683) );
  XOR U1295 ( .A(n1686), .B(n1687), .Z(n1681) );
  AND U1296 ( .A(n398), .B(n1688), .Z(n1687) );
  XOR U1297 ( .A(p_input[536]), .B(n1686), .Z(n1688) );
  XOR U1298 ( .A(n1689), .B(n1690), .Z(n1686) );
  AND U1299 ( .A(n402), .B(n1691), .Z(n1690) );
  XOR U1300 ( .A(n1692), .B(n1693), .Z(n1684) );
  AND U1301 ( .A(n406), .B(n1691), .Z(n1693) );
  XNOR U1302 ( .A(n1692), .B(n1689), .Z(n1691) );
  XOR U1303 ( .A(n1694), .B(n1695), .Z(n1689) );
  AND U1304 ( .A(n409), .B(n1696), .Z(n1695) );
  XOR U1305 ( .A(p_input[552]), .B(n1694), .Z(n1696) );
  XOR U1306 ( .A(n1697), .B(n1698), .Z(n1694) );
  AND U1307 ( .A(n413), .B(n1699), .Z(n1698) );
  XOR U1308 ( .A(n1700), .B(n1701), .Z(n1692) );
  AND U1309 ( .A(n417), .B(n1699), .Z(n1701) );
  XNOR U1310 ( .A(n1700), .B(n1697), .Z(n1699) );
  XOR U1311 ( .A(n1702), .B(n1703), .Z(n1697) );
  AND U1312 ( .A(n420), .B(n1704), .Z(n1703) );
  XOR U1313 ( .A(p_input[568]), .B(n1702), .Z(n1704) );
  XOR U1314 ( .A(n1705), .B(n1706), .Z(n1702) );
  AND U1315 ( .A(n424), .B(n1707), .Z(n1706) );
  XOR U1316 ( .A(n1708), .B(n1709), .Z(n1700) );
  AND U1317 ( .A(n428), .B(n1707), .Z(n1709) );
  XNOR U1318 ( .A(n1708), .B(n1705), .Z(n1707) );
  XOR U1319 ( .A(n1710), .B(n1711), .Z(n1705) );
  AND U1320 ( .A(n431), .B(n1712), .Z(n1711) );
  XOR U1321 ( .A(p_input[584]), .B(n1710), .Z(n1712) );
  XOR U1322 ( .A(n1713), .B(n1714), .Z(n1710) );
  AND U1323 ( .A(n435), .B(n1715), .Z(n1714) );
  XOR U1324 ( .A(n1716), .B(n1717), .Z(n1708) );
  AND U1325 ( .A(n439), .B(n1715), .Z(n1717) );
  XNOR U1326 ( .A(n1716), .B(n1713), .Z(n1715) );
  XOR U1327 ( .A(n1718), .B(n1719), .Z(n1713) );
  AND U1328 ( .A(n442), .B(n1720), .Z(n1719) );
  XOR U1329 ( .A(p_input[600]), .B(n1718), .Z(n1720) );
  XOR U1330 ( .A(n1721), .B(n1722), .Z(n1718) );
  AND U1331 ( .A(n446), .B(n1723), .Z(n1722) );
  XOR U1332 ( .A(n1724), .B(n1725), .Z(n1716) );
  AND U1333 ( .A(n450), .B(n1723), .Z(n1725) );
  XNOR U1334 ( .A(n1724), .B(n1721), .Z(n1723) );
  XOR U1335 ( .A(n1726), .B(n1727), .Z(n1721) );
  AND U1336 ( .A(n453), .B(n1728), .Z(n1727) );
  XOR U1337 ( .A(p_input[616]), .B(n1726), .Z(n1728) );
  XOR U1338 ( .A(n1729), .B(n1730), .Z(n1726) );
  AND U1339 ( .A(n457), .B(n1731), .Z(n1730) );
  XOR U1340 ( .A(n1732), .B(n1733), .Z(n1724) );
  AND U1341 ( .A(n461), .B(n1731), .Z(n1733) );
  XNOR U1342 ( .A(n1732), .B(n1729), .Z(n1731) );
  XOR U1343 ( .A(n1734), .B(n1735), .Z(n1729) );
  AND U1344 ( .A(n464), .B(n1736), .Z(n1735) );
  XOR U1345 ( .A(p_input[632]), .B(n1734), .Z(n1736) );
  XOR U1346 ( .A(n1737), .B(n1738), .Z(n1734) );
  AND U1347 ( .A(n468), .B(n1739), .Z(n1738) );
  XOR U1348 ( .A(n1740), .B(n1741), .Z(n1732) );
  AND U1349 ( .A(n472), .B(n1739), .Z(n1741) );
  XNOR U1350 ( .A(n1740), .B(n1737), .Z(n1739) );
  XOR U1351 ( .A(n1742), .B(n1743), .Z(n1737) );
  AND U1352 ( .A(n475), .B(n1744), .Z(n1743) );
  XOR U1353 ( .A(p_input[648]), .B(n1742), .Z(n1744) );
  XOR U1354 ( .A(n1745), .B(n1746), .Z(n1742) );
  AND U1355 ( .A(n479), .B(n1747), .Z(n1746) );
  XOR U1356 ( .A(n1748), .B(n1749), .Z(n1740) );
  AND U1357 ( .A(n483), .B(n1747), .Z(n1749) );
  XNOR U1358 ( .A(n1748), .B(n1745), .Z(n1747) );
  XOR U1359 ( .A(n1750), .B(n1751), .Z(n1745) );
  AND U1360 ( .A(n486), .B(n1752), .Z(n1751) );
  XOR U1361 ( .A(p_input[664]), .B(n1750), .Z(n1752) );
  XOR U1362 ( .A(n1753), .B(n1754), .Z(n1750) );
  AND U1363 ( .A(n490), .B(n1755), .Z(n1754) );
  XOR U1364 ( .A(n1756), .B(n1757), .Z(n1748) );
  AND U1365 ( .A(n494), .B(n1755), .Z(n1757) );
  XNOR U1366 ( .A(n1756), .B(n1753), .Z(n1755) );
  XOR U1367 ( .A(n1758), .B(n1759), .Z(n1753) );
  AND U1368 ( .A(n497), .B(n1760), .Z(n1759) );
  XOR U1369 ( .A(p_input[680]), .B(n1758), .Z(n1760) );
  XOR U1370 ( .A(n1761), .B(n1762), .Z(n1758) );
  AND U1371 ( .A(n501), .B(n1763), .Z(n1762) );
  XOR U1372 ( .A(n1764), .B(n1765), .Z(n1756) );
  AND U1373 ( .A(n505), .B(n1763), .Z(n1765) );
  XNOR U1374 ( .A(n1764), .B(n1761), .Z(n1763) );
  XOR U1375 ( .A(n1766), .B(n1767), .Z(n1761) );
  AND U1376 ( .A(n508), .B(n1768), .Z(n1767) );
  XOR U1377 ( .A(p_input[696]), .B(n1766), .Z(n1768) );
  XOR U1378 ( .A(n1769), .B(n1770), .Z(n1766) );
  AND U1379 ( .A(n512), .B(n1771), .Z(n1770) );
  XOR U1380 ( .A(n1772), .B(n1773), .Z(n1764) );
  AND U1381 ( .A(n516), .B(n1771), .Z(n1773) );
  XNOR U1382 ( .A(n1772), .B(n1769), .Z(n1771) );
  XOR U1383 ( .A(n1774), .B(n1775), .Z(n1769) );
  AND U1384 ( .A(n519), .B(n1776), .Z(n1775) );
  XOR U1385 ( .A(p_input[712]), .B(n1774), .Z(n1776) );
  XOR U1386 ( .A(n1777), .B(n1778), .Z(n1774) );
  AND U1387 ( .A(n523), .B(n1779), .Z(n1778) );
  XOR U1388 ( .A(n1780), .B(n1781), .Z(n1772) );
  AND U1389 ( .A(n527), .B(n1779), .Z(n1781) );
  XNOR U1390 ( .A(n1780), .B(n1777), .Z(n1779) );
  XOR U1391 ( .A(n1782), .B(n1783), .Z(n1777) );
  AND U1392 ( .A(n530), .B(n1784), .Z(n1783) );
  XOR U1393 ( .A(p_input[728]), .B(n1782), .Z(n1784) );
  XOR U1394 ( .A(n1785), .B(n1786), .Z(n1782) );
  AND U1395 ( .A(n534), .B(n1787), .Z(n1786) );
  XOR U1396 ( .A(n1788), .B(n1789), .Z(n1780) );
  AND U1397 ( .A(n538), .B(n1787), .Z(n1789) );
  XNOR U1398 ( .A(n1788), .B(n1785), .Z(n1787) );
  XOR U1399 ( .A(n1790), .B(n1791), .Z(n1785) );
  AND U1400 ( .A(n541), .B(n1792), .Z(n1791) );
  XOR U1401 ( .A(p_input[744]), .B(n1790), .Z(n1792) );
  XOR U1402 ( .A(n1793), .B(n1794), .Z(n1790) );
  AND U1403 ( .A(n545), .B(n1795), .Z(n1794) );
  XOR U1404 ( .A(n1796), .B(n1797), .Z(n1788) );
  AND U1405 ( .A(n549), .B(n1795), .Z(n1797) );
  XNOR U1406 ( .A(n1796), .B(n1793), .Z(n1795) );
  XOR U1407 ( .A(n1798), .B(n1799), .Z(n1793) );
  AND U1408 ( .A(n552), .B(n1800), .Z(n1799) );
  XOR U1409 ( .A(p_input[760]), .B(n1798), .Z(n1800) );
  XOR U1410 ( .A(n1801), .B(n1802), .Z(n1798) );
  AND U1411 ( .A(n556), .B(n1803), .Z(n1802) );
  XOR U1412 ( .A(n1804), .B(n1805), .Z(n1796) );
  AND U1413 ( .A(n560), .B(n1803), .Z(n1805) );
  XNOR U1414 ( .A(n1804), .B(n1801), .Z(n1803) );
  XOR U1415 ( .A(n1806), .B(n1807), .Z(n1801) );
  AND U1416 ( .A(n563), .B(n1808), .Z(n1807) );
  XOR U1417 ( .A(p_input[776]), .B(n1806), .Z(n1808) );
  XOR U1418 ( .A(n1809), .B(n1810), .Z(n1806) );
  AND U1419 ( .A(n567), .B(n1811), .Z(n1810) );
  XOR U1420 ( .A(n1812), .B(n1813), .Z(n1804) );
  AND U1421 ( .A(n571), .B(n1811), .Z(n1813) );
  XNOR U1422 ( .A(n1812), .B(n1809), .Z(n1811) );
  XOR U1423 ( .A(n1814), .B(n1815), .Z(n1809) );
  AND U1424 ( .A(n574), .B(n1816), .Z(n1815) );
  XOR U1425 ( .A(p_input[792]), .B(n1814), .Z(n1816) );
  XOR U1426 ( .A(n1817), .B(n1818), .Z(n1814) );
  AND U1427 ( .A(n578), .B(n1819), .Z(n1818) );
  XOR U1428 ( .A(n1820), .B(n1821), .Z(n1812) );
  AND U1429 ( .A(n582), .B(n1819), .Z(n1821) );
  XNOR U1430 ( .A(n1820), .B(n1817), .Z(n1819) );
  XOR U1431 ( .A(n1822), .B(n1823), .Z(n1817) );
  AND U1432 ( .A(n585), .B(n1824), .Z(n1823) );
  XOR U1433 ( .A(p_input[808]), .B(n1822), .Z(n1824) );
  XOR U1434 ( .A(n1825), .B(n1826), .Z(n1822) );
  AND U1435 ( .A(n589), .B(n1827), .Z(n1826) );
  XOR U1436 ( .A(n1828), .B(n1829), .Z(n1820) );
  AND U1437 ( .A(n593), .B(n1827), .Z(n1829) );
  XNOR U1438 ( .A(n1828), .B(n1825), .Z(n1827) );
  XOR U1439 ( .A(n1830), .B(n1831), .Z(n1825) );
  AND U1440 ( .A(n596), .B(n1832), .Z(n1831) );
  XOR U1441 ( .A(p_input[824]), .B(n1830), .Z(n1832) );
  XOR U1442 ( .A(n1833), .B(n1834), .Z(n1830) );
  AND U1443 ( .A(n600), .B(n1835), .Z(n1834) );
  XOR U1444 ( .A(n1836), .B(n1837), .Z(n1828) );
  AND U1445 ( .A(n604), .B(n1835), .Z(n1837) );
  XNOR U1446 ( .A(n1836), .B(n1833), .Z(n1835) );
  XOR U1447 ( .A(n1838), .B(n1839), .Z(n1833) );
  AND U1448 ( .A(n607), .B(n1840), .Z(n1839) );
  XOR U1449 ( .A(p_input[840]), .B(n1838), .Z(n1840) );
  XOR U1450 ( .A(n1841), .B(n1842), .Z(n1838) );
  AND U1451 ( .A(n611), .B(n1843), .Z(n1842) );
  XOR U1452 ( .A(n1844), .B(n1845), .Z(n1836) );
  AND U1453 ( .A(n615), .B(n1843), .Z(n1845) );
  XNOR U1454 ( .A(n1844), .B(n1841), .Z(n1843) );
  XOR U1455 ( .A(n1846), .B(n1847), .Z(n1841) );
  AND U1456 ( .A(n618), .B(n1848), .Z(n1847) );
  XOR U1457 ( .A(p_input[856]), .B(n1846), .Z(n1848) );
  XOR U1458 ( .A(n1849), .B(n1850), .Z(n1846) );
  AND U1459 ( .A(n622), .B(n1851), .Z(n1850) );
  XOR U1460 ( .A(n1852), .B(n1853), .Z(n1844) );
  AND U1461 ( .A(n626), .B(n1851), .Z(n1853) );
  XNOR U1462 ( .A(n1852), .B(n1849), .Z(n1851) );
  XOR U1463 ( .A(n1854), .B(n1855), .Z(n1849) );
  AND U1464 ( .A(n629), .B(n1856), .Z(n1855) );
  XOR U1465 ( .A(p_input[872]), .B(n1854), .Z(n1856) );
  XOR U1466 ( .A(n1857), .B(n1858), .Z(n1854) );
  AND U1467 ( .A(n633), .B(n1859), .Z(n1858) );
  XOR U1468 ( .A(n1860), .B(n1861), .Z(n1852) );
  AND U1469 ( .A(n637), .B(n1859), .Z(n1861) );
  XNOR U1470 ( .A(n1860), .B(n1857), .Z(n1859) );
  XOR U1471 ( .A(n1862), .B(n1863), .Z(n1857) );
  AND U1472 ( .A(n640), .B(n1864), .Z(n1863) );
  XOR U1473 ( .A(p_input[888]), .B(n1862), .Z(n1864) );
  XOR U1474 ( .A(n1865), .B(n1866), .Z(n1862) );
  AND U1475 ( .A(n644), .B(n1867), .Z(n1866) );
  XOR U1476 ( .A(n1868), .B(n1869), .Z(n1860) );
  AND U1477 ( .A(n648), .B(n1867), .Z(n1869) );
  XNOR U1478 ( .A(n1868), .B(n1865), .Z(n1867) );
  XOR U1479 ( .A(n1870), .B(n1871), .Z(n1865) );
  AND U1480 ( .A(n651), .B(n1872), .Z(n1871) );
  XOR U1481 ( .A(p_input[904]), .B(n1870), .Z(n1872) );
  XOR U1482 ( .A(n1873), .B(n1874), .Z(n1870) );
  AND U1483 ( .A(n655), .B(n1875), .Z(n1874) );
  XOR U1484 ( .A(n1876), .B(n1877), .Z(n1868) );
  AND U1485 ( .A(n659), .B(n1875), .Z(n1877) );
  XNOR U1486 ( .A(n1876), .B(n1873), .Z(n1875) );
  XOR U1487 ( .A(n1878), .B(n1879), .Z(n1873) );
  AND U1488 ( .A(n662), .B(n1880), .Z(n1879) );
  XOR U1489 ( .A(p_input[920]), .B(n1878), .Z(n1880) );
  XOR U1490 ( .A(n1881), .B(n1882), .Z(n1878) );
  AND U1491 ( .A(n666), .B(n1883), .Z(n1882) );
  XOR U1492 ( .A(n1884), .B(n1885), .Z(n1876) );
  AND U1493 ( .A(n670), .B(n1883), .Z(n1885) );
  XNOR U1494 ( .A(n1884), .B(n1881), .Z(n1883) );
  XOR U1495 ( .A(n1886), .B(n1887), .Z(n1881) );
  AND U1496 ( .A(n673), .B(n1888), .Z(n1887) );
  XOR U1497 ( .A(p_input[936]), .B(n1886), .Z(n1888) );
  XOR U1498 ( .A(n1889), .B(n1890), .Z(n1886) );
  AND U1499 ( .A(n677), .B(n1891), .Z(n1890) );
  XOR U1500 ( .A(n1892), .B(n1893), .Z(n1884) );
  AND U1501 ( .A(n681), .B(n1891), .Z(n1893) );
  XNOR U1502 ( .A(n1892), .B(n1889), .Z(n1891) );
  XOR U1503 ( .A(n1894), .B(n1895), .Z(n1889) );
  AND U1504 ( .A(n684), .B(n1896), .Z(n1895) );
  XOR U1505 ( .A(p_input[952]), .B(n1894), .Z(n1896) );
  XOR U1506 ( .A(n1897), .B(n1898), .Z(n1894) );
  AND U1507 ( .A(n688), .B(n1899), .Z(n1898) );
  XOR U1508 ( .A(n1900), .B(n1901), .Z(n1892) );
  AND U1509 ( .A(n692), .B(n1899), .Z(n1901) );
  XNOR U1510 ( .A(n1900), .B(n1897), .Z(n1899) );
  XOR U1511 ( .A(n1902), .B(n1903), .Z(n1897) );
  AND U1512 ( .A(n695), .B(n1904), .Z(n1903) );
  XOR U1513 ( .A(p_input[968]), .B(n1902), .Z(n1904) );
  XOR U1514 ( .A(n1905), .B(n1906), .Z(n1902) );
  AND U1515 ( .A(n699), .B(n1907), .Z(n1906) );
  XOR U1516 ( .A(n1908), .B(n1909), .Z(n1900) );
  AND U1517 ( .A(n703), .B(n1907), .Z(n1909) );
  XNOR U1518 ( .A(n1908), .B(n1905), .Z(n1907) );
  XOR U1519 ( .A(n1910), .B(n1911), .Z(n1905) );
  AND U1520 ( .A(n706), .B(n1912), .Z(n1911) );
  XOR U1521 ( .A(p_input[984]), .B(n1910), .Z(n1912) );
  XOR U1522 ( .A(n1913), .B(n1914), .Z(n1910) );
  AND U1523 ( .A(n710), .B(n1915), .Z(n1914) );
  XOR U1524 ( .A(n1916), .B(n1917), .Z(n1908) );
  AND U1525 ( .A(n714), .B(n1915), .Z(n1917) );
  XNOR U1526 ( .A(n1916), .B(n1913), .Z(n1915) );
  XOR U1527 ( .A(n1918), .B(n1919), .Z(n1913) );
  AND U1528 ( .A(n717), .B(n1920), .Z(n1919) );
  XOR U1529 ( .A(p_input[1000]), .B(n1918), .Z(n1920) );
  XOR U1530 ( .A(n1921), .B(n1922), .Z(n1918) );
  AND U1531 ( .A(n721), .B(n1923), .Z(n1922) );
  XOR U1532 ( .A(n1924), .B(n1925), .Z(n1916) );
  AND U1533 ( .A(n725), .B(n1923), .Z(n1925) );
  XNOR U1534 ( .A(n1924), .B(n1921), .Z(n1923) );
  XOR U1535 ( .A(n1926), .B(n1927), .Z(n1921) );
  AND U1536 ( .A(n728), .B(n1928), .Z(n1927) );
  XOR U1537 ( .A(p_input[1016]), .B(n1926), .Z(n1928) );
  XOR U1538 ( .A(n1929), .B(n1930), .Z(n1926) );
  AND U1539 ( .A(n732), .B(n1931), .Z(n1930) );
  XOR U1540 ( .A(n1932), .B(n1933), .Z(n1924) );
  AND U1541 ( .A(n736), .B(n1931), .Z(n1933) );
  XNOR U1542 ( .A(n1932), .B(n1929), .Z(n1931) );
  XOR U1543 ( .A(n1934), .B(n1935), .Z(n1929) );
  AND U1544 ( .A(n739), .B(n1936), .Z(n1935) );
  XOR U1545 ( .A(p_input[1032]), .B(n1934), .Z(n1936) );
  XOR U1546 ( .A(n1937), .B(n1938), .Z(n1934) );
  AND U1547 ( .A(n743), .B(n1939), .Z(n1938) );
  XOR U1548 ( .A(n1940), .B(n1941), .Z(n1932) );
  AND U1549 ( .A(n747), .B(n1939), .Z(n1941) );
  XNOR U1550 ( .A(n1940), .B(n1937), .Z(n1939) );
  XOR U1551 ( .A(n1942), .B(n1943), .Z(n1937) );
  AND U1552 ( .A(n750), .B(n1944), .Z(n1943) );
  XOR U1553 ( .A(p_input[1048]), .B(n1942), .Z(n1944) );
  XOR U1554 ( .A(n1945), .B(n1946), .Z(n1942) );
  AND U1555 ( .A(n754), .B(n1947), .Z(n1946) );
  XOR U1556 ( .A(n1948), .B(n1949), .Z(n1940) );
  AND U1557 ( .A(n758), .B(n1947), .Z(n1949) );
  XNOR U1558 ( .A(n1948), .B(n1945), .Z(n1947) );
  XOR U1559 ( .A(n1950), .B(n1951), .Z(n1945) );
  AND U1560 ( .A(n761), .B(n1952), .Z(n1951) );
  XOR U1561 ( .A(p_input[1064]), .B(n1950), .Z(n1952) );
  XOR U1562 ( .A(n1953), .B(n1954), .Z(n1950) );
  AND U1563 ( .A(n765), .B(n1955), .Z(n1954) );
  XOR U1564 ( .A(n1956), .B(n1957), .Z(n1948) );
  AND U1565 ( .A(n769), .B(n1955), .Z(n1957) );
  XNOR U1566 ( .A(n1956), .B(n1953), .Z(n1955) );
  XOR U1567 ( .A(n1958), .B(n1959), .Z(n1953) );
  AND U1568 ( .A(n772), .B(n1960), .Z(n1959) );
  XOR U1569 ( .A(p_input[1080]), .B(n1958), .Z(n1960) );
  XOR U1570 ( .A(n1961), .B(n1962), .Z(n1958) );
  AND U1571 ( .A(n776), .B(n1963), .Z(n1962) );
  XOR U1572 ( .A(n1964), .B(n1965), .Z(n1956) );
  AND U1573 ( .A(n780), .B(n1963), .Z(n1965) );
  XNOR U1574 ( .A(n1964), .B(n1961), .Z(n1963) );
  XOR U1575 ( .A(n1966), .B(n1967), .Z(n1961) );
  AND U1576 ( .A(n783), .B(n1968), .Z(n1967) );
  XOR U1577 ( .A(p_input[1096]), .B(n1966), .Z(n1968) );
  XOR U1578 ( .A(n1969), .B(n1970), .Z(n1966) );
  AND U1579 ( .A(n787), .B(n1971), .Z(n1970) );
  XOR U1580 ( .A(n1972), .B(n1973), .Z(n1964) );
  AND U1581 ( .A(n791), .B(n1971), .Z(n1973) );
  XNOR U1582 ( .A(n1972), .B(n1969), .Z(n1971) );
  XOR U1583 ( .A(n1974), .B(n1975), .Z(n1969) );
  AND U1584 ( .A(n794), .B(n1976), .Z(n1975) );
  XOR U1585 ( .A(p_input[1112]), .B(n1974), .Z(n1976) );
  XOR U1586 ( .A(n1977), .B(n1978), .Z(n1974) );
  AND U1587 ( .A(n798), .B(n1979), .Z(n1978) );
  XOR U1588 ( .A(n1980), .B(n1981), .Z(n1972) );
  AND U1589 ( .A(n802), .B(n1979), .Z(n1981) );
  XNOR U1590 ( .A(n1980), .B(n1977), .Z(n1979) );
  XOR U1591 ( .A(n1982), .B(n1983), .Z(n1977) );
  AND U1592 ( .A(n805), .B(n1984), .Z(n1983) );
  XOR U1593 ( .A(p_input[1128]), .B(n1982), .Z(n1984) );
  XOR U1594 ( .A(n1985), .B(n1986), .Z(n1982) );
  AND U1595 ( .A(n809), .B(n1987), .Z(n1986) );
  XOR U1596 ( .A(n1988), .B(n1989), .Z(n1980) );
  AND U1597 ( .A(n813), .B(n1987), .Z(n1989) );
  XNOR U1598 ( .A(n1988), .B(n1985), .Z(n1987) );
  XOR U1599 ( .A(n1990), .B(n1991), .Z(n1985) );
  AND U1600 ( .A(n816), .B(n1992), .Z(n1991) );
  XOR U1601 ( .A(p_input[1144]), .B(n1990), .Z(n1992) );
  XOR U1602 ( .A(n1993), .B(n1994), .Z(n1990) );
  AND U1603 ( .A(n820), .B(n1995), .Z(n1994) );
  XOR U1604 ( .A(n1996), .B(n1997), .Z(n1988) );
  AND U1605 ( .A(n824), .B(n1995), .Z(n1997) );
  XNOR U1606 ( .A(n1996), .B(n1993), .Z(n1995) );
  XOR U1607 ( .A(n1998), .B(n1999), .Z(n1993) );
  AND U1608 ( .A(n827), .B(n2000), .Z(n1999) );
  XOR U1609 ( .A(p_input[1160]), .B(n1998), .Z(n2000) );
  XOR U1610 ( .A(n2001), .B(n2002), .Z(n1998) );
  AND U1611 ( .A(n831), .B(n2003), .Z(n2002) );
  XOR U1612 ( .A(n2004), .B(n2005), .Z(n1996) );
  AND U1613 ( .A(n835), .B(n2003), .Z(n2005) );
  XNOR U1614 ( .A(n2004), .B(n2001), .Z(n2003) );
  XOR U1615 ( .A(n2006), .B(n2007), .Z(n2001) );
  AND U1616 ( .A(n838), .B(n2008), .Z(n2007) );
  XOR U1617 ( .A(p_input[1176]), .B(n2006), .Z(n2008) );
  XOR U1618 ( .A(n2009), .B(n2010), .Z(n2006) );
  AND U1619 ( .A(n842), .B(n2011), .Z(n2010) );
  XOR U1620 ( .A(n2012), .B(n2013), .Z(n2004) );
  AND U1621 ( .A(n846), .B(n2011), .Z(n2013) );
  XNOR U1622 ( .A(n2012), .B(n2009), .Z(n2011) );
  XOR U1623 ( .A(n2014), .B(n2015), .Z(n2009) );
  AND U1624 ( .A(n849), .B(n2016), .Z(n2015) );
  XOR U1625 ( .A(p_input[1192]), .B(n2014), .Z(n2016) );
  XOR U1626 ( .A(n2017), .B(n2018), .Z(n2014) );
  AND U1627 ( .A(n853), .B(n2019), .Z(n2018) );
  XOR U1628 ( .A(n2020), .B(n2021), .Z(n2012) );
  AND U1629 ( .A(n857), .B(n2019), .Z(n2021) );
  XNOR U1630 ( .A(n2020), .B(n2017), .Z(n2019) );
  XOR U1631 ( .A(n2022), .B(n2023), .Z(n2017) );
  AND U1632 ( .A(n860), .B(n2024), .Z(n2023) );
  XOR U1633 ( .A(p_input[1208]), .B(n2022), .Z(n2024) );
  XOR U1634 ( .A(n2025), .B(n2026), .Z(n2022) );
  AND U1635 ( .A(n864), .B(n2027), .Z(n2026) );
  XOR U1636 ( .A(n2028), .B(n2029), .Z(n2020) );
  AND U1637 ( .A(n868), .B(n2027), .Z(n2029) );
  XNOR U1638 ( .A(n2028), .B(n2025), .Z(n2027) );
  XOR U1639 ( .A(n2030), .B(n2031), .Z(n2025) );
  AND U1640 ( .A(n871), .B(n2032), .Z(n2031) );
  XOR U1641 ( .A(p_input[1224]), .B(n2030), .Z(n2032) );
  XOR U1642 ( .A(n2033), .B(n2034), .Z(n2030) );
  AND U1643 ( .A(n875), .B(n2035), .Z(n2034) );
  XOR U1644 ( .A(n2036), .B(n2037), .Z(n2028) );
  AND U1645 ( .A(n879), .B(n2035), .Z(n2037) );
  XNOR U1646 ( .A(n2036), .B(n2033), .Z(n2035) );
  XOR U1647 ( .A(n2038), .B(n2039), .Z(n2033) );
  AND U1648 ( .A(n882), .B(n2040), .Z(n2039) );
  XOR U1649 ( .A(p_input[1240]), .B(n2038), .Z(n2040) );
  XOR U1650 ( .A(n2041), .B(n2042), .Z(n2038) );
  AND U1651 ( .A(n886), .B(n2043), .Z(n2042) );
  XOR U1652 ( .A(n2044), .B(n2045), .Z(n2036) );
  AND U1653 ( .A(n890), .B(n2043), .Z(n2045) );
  XNOR U1654 ( .A(n2044), .B(n2041), .Z(n2043) );
  XOR U1655 ( .A(n2046), .B(n2047), .Z(n2041) );
  AND U1656 ( .A(n893), .B(n2048), .Z(n2047) );
  XOR U1657 ( .A(p_input[1256]), .B(n2046), .Z(n2048) );
  XOR U1658 ( .A(n2049), .B(n2050), .Z(n2046) );
  AND U1659 ( .A(n897), .B(n2051), .Z(n2050) );
  XOR U1660 ( .A(n2052), .B(n2053), .Z(n2044) );
  AND U1661 ( .A(n901), .B(n2051), .Z(n2053) );
  XNOR U1662 ( .A(n2052), .B(n2049), .Z(n2051) );
  XOR U1663 ( .A(n2054), .B(n2055), .Z(n2049) );
  AND U1664 ( .A(n904), .B(n2056), .Z(n2055) );
  XOR U1665 ( .A(p_input[1272]), .B(n2054), .Z(n2056) );
  XOR U1666 ( .A(n2057), .B(n2058), .Z(n2054) );
  AND U1667 ( .A(n908), .B(n2059), .Z(n2058) );
  XOR U1668 ( .A(n2060), .B(n2061), .Z(n2052) );
  AND U1669 ( .A(n912), .B(n2059), .Z(n2061) );
  XNOR U1670 ( .A(n2060), .B(n2057), .Z(n2059) );
  XOR U1671 ( .A(n2062), .B(n2063), .Z(n2057) );
  AND U1672 ( .A(n915), .B(n2064), .Z(n2063) );
  XOR U1673 ( .A(p_input[1288]), .B(n2062), .Z(n2064) );
  XOR U1674 ( .A(n2065), .B(n2066), .Z(n2062) );
  AND U1675 ( .A(n919), .B(n2067), .Z(n2066) );
  XOR U1676 ( .A(n2068), .B(n2069), .Z(n2060) );
  AND U1677 ( .A(n923), .B(n2067), .Z(n2069) );
  XNOR U1678 ( .A(n2068), .B(n2065), .Z(n2067) );
  XOR U1679 ( .A(n2070), .B(n2071), .Z(n2065) );
  AND U1680 ( .A(n926), .B(n2072), .Z(n2071) );
  XOR U1681 ( .A(p_input[1304]), .B(n2070), .Z(n2072) );
  XOR U1682 ( .A(n2073), .B(n2074), .Z(n2070) );
  AND U1683 ( .A(n930), .B(n2075), .Z(n2074) );
  XOR U1684 ( .A(n2076), .B(n2077), .Z(n2068) );
  AND U1685 ( .A(n934), .B(n2075), .Z(n2077) );
  XNOR U1686 ( .A(n2076), .B(n2073), .Z(n2075) );
  XOR U1687 ( .A(n2078), .B(n2079), .Z(n2073) );
  AND U1688 ( .A(n937), .B(n2080), .Z(n2079) );
  XOR U1689 ( .A(p_input[1320]), .B(n2078), .Z(n2080) );
  XOR U1690 ( .A(n2081), .B(n2082), .Z(n2078) );
  AND U1691 ( .A(n941), .B(n2083), .Z(n2082) );
  XOR U1692 ( .A(n2084), .B(n2085), .Z(n2076) );
  AND U1693 ( .A(n945), .B(n2083), .Z(n2085) );
  XNOR U1694 ( .A(n2084), .B(n2081), .Z(n2083) );
  XOR U1695 ( .A(n2086), .B(n2087), .Z(n2081) );
  AND U1696 ( .A(n948), .B(n2088), .Z(n2087) );
  XOR U1697 ( .A(p_input[1336]), .B(n2086), .Z(n2088) );
  XOR U1698 ( .A(n2089), .B(n2090), .Z(n2086) );
  AND U1699 ( .A(n952), .B(n2091), .Z(n2090) );
  XOR U1700 ( .A(n2092), .B(n2093), .Z(n2084) );
  AND U1701 ( .A(n956), .B(n2091), .Z(n2093) );
  XNOR U1702 ( .A(n2092), .B(n2089), .Z(n2091) );
  XOR U1703 ( .A(n2094), .B(n2095), .Z(n2089) );
  AND U1704 ( .A(n959), .B(n2096), .Z(n2095) );
  XOR U1705 ( .A(p_input[1352]), .B(n2094), .Z(n2096) );
  XOR U1706 ( .A(n2097), .B(n2098), .Z(n2094) );
  AND U1707 ( .A(n963), .B(n2099), .Z(n2098) );
  XOR U1708 ( .A(n2100), .B(n2101), .Z(n2092) );
  AND U1709 ( .A(n967), .B(n2099), .Z(n2101) );
  XNOR U1710 ( .A(n2100), .B(n2097), .Z(n2099) );
  XOR U1711 ( .A(n2102), .B(n2103), .Z(n2097) );
  AND U1712 ( .A(n970), .B(n2104), .Z(n2103) );
  XOR U1713 ( .A(p_input[1368]), .B(n2102), .Z(n2104) );
  XOR U1714 ( .A(n2105), .B(n2106), .Z(n2102) );
  AND U1715 ( .A(n974), .B(n2107), .Z(n2106) );
  XOR U1716 ( .A(n2108), .B(n2109), .Z(n2100) );
  AND U1717 ( .A(n978), .B(n2107), .Z(n2109) );
  XNOR U1718 ( .A(n2108), .B(n2105), .Z(n2107) );
  XOR U1719 ( .A(n2110), .B(n2111), .Z(n2105) );
  AND U1720 ( .A(n981), .B(n2112), .Z(n2111) );
  XOR U1721 ( .A(p_input[1384]), .B(n2110), .Z(n2112) );
  XOR U1722 ( .A(n2113), .B(n2114), .Z(n2110) );
  AND U1723 ( .A(n985), .B(n2115), .Z(n2114) );
  XOR U1724 ( .A(n2116), .B(n2117), .Z(n2108) );
  AND U1725 ( .A(n989), .B(n2115), .Z(n2117) );
  XNOR U1726 ( .A(n2116), .B(n2113), .Z(n2115) );
  XOR U1727 ( .A(n2118), .B(n2119), .Z(n2113) );
  AND U1728 ( .A(n992), .B(n2120), .Z(n2119) );
  XOR U1729 ( .A(p_input[1400]), .B(n2118), .Z(n2120) );
  XOR U1730 ( .A(n2121), .B(n2122), .Z(n2118) );
  AND U1731 ( .A(n996), .B(n2123), .Z(n2122) );
  XOR U1732 ( .A(n2124), .B(n2125), .Z(n2116) );
  AND U1733 ( .A(n1000), .B(n2123), .Z(n2125) );
  XNOR U1734 ( .A(n2124), .B(n2121), .Z(n2123) );
  XOR U1735 ( .A(n2126), .B(n2127), .Z(n2121) );
  AND U1736 ( .A(n1003), .B(n2128), .Z(n2127) );
  XOR U1737 ( .A(p_input[1416]), .B(n2126), .Z(n2128) );
  XOR U1738 ( .A(n2129), .B(n2130), .Z(n2126) );
  AND U1739 ( .A(n1007), .B(n2131), .Z(n2130) );
  XOR U1740 ( .A(n2132), .B(n2133), .Z(n2124) );
  AND U1741 ( .A(n1011), .B(n2131), .Z(n2133) );
  XNOR U1742 ( .A(n2132), .B(n2129), .Z(n2131) );
  XOR U1743 ( .A(n2134), .B(n2135), .Z(n2129) );
  AND U1744 ( .A(n1014), .B(n2136), .Z(n2135) );
  XOR U1745 ( .A(p_input[1432]), .B(n2134), .Z(n2136) );
  XOR U1746 ( .A(n2137), .B(n2138), .Z(n2134) );
  AND U1747 ( .A(n1018), .B(n2139), .Z(n2138) );
  XOR U1748 ( .A(n2140), .B(n2141), .Z(n2132) );
  AND U1749 ( .A(n1022), .B(n2139), .Z(n2141) );
  XNOR U1750 ( .A(n2140), .B(n2137), .Z(n2139) );
  XOR U1751 ( .A(n2142), .B(n2143), .Z(n2137) );
  AND U1752 ( .A(n1025), .B(n2144), .Z(n2143) );
  XOR U1753 ( .A(p_input[1448]), .B(n2142), .Z(n2144) );
  XOR U1754 ( .A(n2145), .B(n2146), .Z(n2142) );
  AND U1755 ( .A(n1029), .B(n2147), .Z(n2146) );
  XOR U1756 ( .A(n2148), .B(n2149), .Z(n2140) );
  AND U1757 ( .A(n1033), .B(n2147), .Z(n2149) );
  XNOR U1758 ( .A(n2148), .B(n2145), .Z(n2147) );
  XOR U1759 ( .A(n2150), .B(n2151), .Z(n2145) );
  AND U1760 ( .A(n1036), .B(n2152), .Z(n2151) );
  XOR U1761 ( .A(p_input[1464]), .B(n2150), .Z(n2152) );
  XOR U1762 ( .A(n2153), .B(n2154), .Z(n2150) );
  AND U1763 ( .A(n1040), .B(n2155), .Z(n2154) );
  XOR U1764 ( .A(n2156), .B(n2157), .Z(n2148) );
  AND U1765 ( .A(n1044), .B(n2155), .Z(n2157) );
  XNOR U1766 ( .A(n2156), .B(n2153), .Z(n2155) );
  XOR U1767 ( .A(n2158), .B(n2159), .Z(n2153) );
  AND U1768 ( .A(n1047), .B(n2160), .Z(n2159) );
  XOR U1769 ( .A(p_input[1480]), .B(n2158), .Z(n2160) );
  XOR U1770 ( .A(n2161), .B(n2162), .Z(n2158) );
  AND U1771 ( .A(n1051), .B(n2163), .Z(n2162) );
  XOR U1772 ( .A(n2164), .B(n2165), .Z(n2156) );
  AND U1773 ( .A(n1055), .B(n2163), .Z(n2165) );
  XNOR U1774 ( .A(n2164), .B(n2161), .Z(n2163) );
  XOR U1775 ( .A(n2166), .B(n2167), .Z(n2161) );
  AND U1776 ( .A(n1058), .B(n2168), .Z(n2167) );
  XOR U1777 ( .A(p_input[1496]), .B(n2166), .Z(n2168) );
  XOR U1778 ( .A(n2169), .B(n2170), .Z(n2166) );
  AND U1779 ( .A(n1062), .B(n2171), .Z(n2170) );
  XOR U1780 ( .A(n2172), .B(n2173), .Z(n2164) );
  AND U1781 ( .A(n1066), .B(n2171), .Z(n2173) );
  XNOR U1782 ( .A(n2172), .B(n2169), .Z(n2171) );
  XOR U1783 ( .A(n2174), .B(n2175), .Z(n2169) );
  AND U1784 ( .A(n1069), .B(n2176), .Z(n2175) );
  XOR U1785 ( .A(p_input[1512]), .B(n2174), .Z(n2176) );
  XOR U1786 ( .A(n2177), .B(n2178), .Z(n2174) );
  AND U1787 ( .A(n1073), .B(n2179), .Z(n2178) );
  XOR U1788 ( .A(n2180), .B(n2181), .Z(n2172) );
  AND U1789 ( .A(n1077), .B(n2179), .Z(n2181) );
  XNOR U1790 ( .A(n2180), .B(n2177), .Z(n2179) );
  XOR U1791 ( .A(n2182), .B(n2183), .Z(n2177) );
  AND U1792 ( .A(n1080), .B(n2184), .Z(n2183) );
  XOR U1793 ( .A(p_input[1528]), .B(n2182), .Z(n2184) );
  XOR U1794 ( .A(n2185), .B(n2186), .Z(n2182) );
  AND U1795 ( .A(n1084), .B(n2187), .Z(n2186) );
  XOR U1796 ( .A(n2188), .B(n2189), .Z(n2180) );
  AND U1797 ( .A(n1088), .B(n2187), .Z(n2189) );
  XNOR U1798 ( .A(n2188), .B(n2185), .Z(n2187) );
  XOR U1799 ( .A(n2190), .B(n2191), .Z(n2185) );
  AND U1800 ( .A(n1091), .B(n2192), .Z(n2191) );
  XOR U1801 ( .A(p_input[1544]), .B(n2190), .Z(n2192) );
  XOR U1802 ( .A(n2193), .B(n2194), .Z(n2190) );
  AND U1803 ( .A(n1095), .B(n2195), .Z(n2194) );
  XOR U1804 ( .A(n2196), .B(n2197), .Z(n2188) );
  AND U1805 ( .A(n1099), .B(n2195), .Z(n2197) );
  XNOR U1806 ( .A(n2196), .B(n2193), .Z(n2195) );
  XOR U1807 ( .A(n2198), .B(n2199), .Z(n2193) );
  AND U1808 ( .A(n1102), .B(n2200), .Z(n2199) );
  XOR U1809 ( .A(p_input[1560]), .B(n2198), .Z(n2200) );
  XOR U1810 ( .A(n2201), .B(n2202), .Z(n2198) );
  AND U1811 ( .A(n1106), .B(n2203), .Z(n2202) );
  XOR U1812 ( .A(n2204), .B(n2205), .Z(n2196) );
  AND U1813 ( .A(n1110), .B(n2203), .Z(n2205) );
  XNOR U1814 ( .A(n2204), .B(n2201), .Z(n2203) );
  XOR U1815 ( .A(n2206), .B(n2207), .Z(n2201) );
  AND U1816 ( .A(n1113), .B(n2208), .Z(n2207) );
  XOR U1817 ( .A(p_input[1576]), .B(n2206), .Z(n2208) );
  XOR U1818 ( .A(n2209), .B(n2210), .Z(n2206) );
  AND U1819 ( .A(n1117), .B(n2211), .Z(n2210) );
  XOR U1820 ( .A(n2212), .B(n2213), .Z(n2204) );
  AND U1821 ( .A(n1121), .B(n2211), .Z(n2213) );
  XNOR U1822 ( .A(n2212), .B(n2209), .Z(n2211) );
  XOR U1823 ( .A(n2214), .B(n2215), .Z(n2209) );
  AND U1824 ( .A(n1124), .B(n2216), .Z(n2215) );
  XOR U1825 ( .A(p_input[1592]), .B(n2214), .Z(n2216) );
  XOR U1826 ( .A(n2217), .B(n2218), .Z(n2214) );
  AND U1827 ( .A(n1128), .B(n2219), .Z(n2218) );
  XOR U1828 ( .A(n2220), .B(n2221), .Z(n2212) );
  AND U1829 ( .A(n1132), .B(n2219), .Z(n2221) );
  XNOR U1830 ( .A(n2220), .B(n2217), .Z(n2219) );
  XOR U1831 ( .A(n2222), .B(n2223), .Z(n2217) );
  AND U1832 ( .A(n1135), .B(n2224), .Z(n2223) );
  XOR U1833 ( .A(p_input[1608]), .B(n2222), .Z(n2224) );
  XOR U1834 ( .A(n2225), .B(n2226), .Z(n2222) );
  AND U1835 ( .A(n1139), .B(n2227), .Z(n2226) );
  XOR U1836 ( .A(n2228), .B(n2229), .Z(n2220) );
  AND U1837 ( .A(n1143), .B(n2227), .Z(n2229) );
  XNOR U1838 ( .A(n2228), .B(n2225), .Z(n2227) );
  XOR U1839 ( .A(n2230), .B(n2231), .Z(n2225) );
  AND U1840 ( .A(n1146), .B(n2232), .Z(n2231) );
  XOR U1841 ( .A(p_input[1624]), .B(n2230), .Z(n2232) );
  XOR U1842 ( .A(n2233), .B(n2234), .Z(n2230) );
  AND U1843 ( .A(n1150), .B(n2235), .Z(n2234) );
  XOR U1844 ( .A(n2236), .B(n2237), .Z(n2228) );
  AND U1845 ( .A(n1154), .B(n2235), .Z(n2237) );
  XNOR U1846 ( .A(n2236), .B(n2233), .Z(n2235) );
  XOR U1847 ( .A(n2238), .B(n2239), .Z(n2233) );
  AND U1848 ( .A(n1157), .B(n2240), .Z(n2239) );
  XOR U1849 ( .A(p_input[1640]), .B(n2238), .Z(n2240) );
  XOR U1850 ( .A(n2241), .B(n2242), .Z(n2238) );
  AND U1851 ( .A(n1161), .B(n2243), .Z(n2242) );
  XOR U1852 ( .A(n2244), .B(n2245), .Z(n2236) );
  AND U1853 ( .A(n1165), .B(n2243), .Z(n2245) );
  XNOR U1854 ( .A(n2244), .B(n2241), .Z(n2243) );
  XOR U1855 ( .A(n2246), .B(n2247), .Z(n2241) );
  AND U1856 ( .A(n1168), .B(n2248), .Z(n2247) );
  XOR U1857 ( .A(p_input[1656]), .B(n2246), .Z(n2248) );
  XOR U1858 ( .A(n2249), .B(n2250), .Z(n2246) );
  AND U1859 ( .A(n1172), .B(n2251), .Z(n2250) );
  XOR U1860 ( .A(n2252), .B(n2253), .Z(n2244) );
  AND U1861 ( .A(n1176), .B(n2251), .Z(n2253) );
  XNOR U1862 ( .A(n2252), .B(n2249), .Z(n2251) );
  XOR U1863 ( .A(n2254), .B(n2255), .Z(n2249) );
  AND U1864 ( .A(n1179), .B(n2256), .Z(n2255) );
  XOR U1865 ( .A(p_input[1672]), .B(n2254), .Z(n2256) );
  XOR U1866 ( .A(n2257), .B(n2258), .Z(n2254) );
  AND U1867 ( .A(n1183), .B(n2259), .Z(n2258) );
  XOR U1868 ( .A(n2260), .B(n2261), .Z(n2252) );
  AND U1869 ( .A(n1187), .B(n2259), .Z(n2261) );
  XNOR U1870 ( .A(n2260), .B(n2257), .Z(n2259) );
  XOR U1871 ( .A(n2262), .B(n2263), .Z(n2257) );
  AND U1872 ( .A(n1190), .B(n2264), .Z(n2263) );
  XOR U1873 ( .A(p_input[1688]), .B(n2262), .Z(n2264) );
  XOR U1874 ( .A(n2265), .B(n2266), .Z(n2262) );
  AND U1875 ( .A(n1194), .B(n2267), .Z(n2266) );
  XOR U1876 ( .A(n2268), .B(n2269), .Z(n2260) );
  AND U1877 ( .A(n1198), .B(n2267), .Z(n2269) );
  XNOR U1878 ( .A(n2268), .B(n2265), .Z(n2267) );
  XOR U1879 ( .A(n2270), .B(n2271), .Z(n2265) );
  AND U1880 ( .A(n1201), .B(n2272), .Z(n2271) );
  XOR U1881 ( .A(p_input[1704]), .B(n2270), .Z(n2272) );
  XOR U1882 ( .A(n2273), .B(n2274), .Z(n2270) );
  AND U1883 ( .A(n1205), .B(n2275), .Z(n2274) );
  XOR U1884 ( .A(n2276), .B(n2277), .Z(n2268) );
  AND U1885 ( .A(n1209), .B(n2275), .Z(n2277) );
  XNOR U1886 ( .A(n2276), .B(n2273), .Z(n2275) );
  XOR U1887 ( .A(n2278), .B(n2279), .Z(n2273) );
  AND U1888 ( .A(n1212), .B(n2280), .Z(n2279) );
  XOR U1889 ( .A(p_input[1720]), .B(n2278), .Z(n2280) );
  XOR U1890 ( .A(n2281), .B(n2282), .Z(n2278) );
  AND U1891 ( .A(n1216), .B(n2283), .Z(n2282) );
  XOR U1892 ( .A(n2284), .B(n2285), .Z(n2276) );
  AND U1893 ( .A(n1220), .B(n2283), .Z(n2285) );
  XNOR U1894 ( .A(n2284), .B(n2281), .Z(n2283) );
  XOR U1895 ( .A(n2286), .B(n2287), .Z(n2281) );
  AND U1896 ( .A(n1223), .B(n2288), .Z(n2287) );
  XOR U1897 ( .A(p_input[1736]), .B(n2286), .Z(n2288) );
  XOR U1898 ( .A(n2289), .B(n2290), .Z(n2286) );
  AND U1899 ( .A(n1227), .B(n2291), .Z(n2290) );
  XOR U1900 ( .A(n2292), .B(n2293), .Z(n2284) );
  AND U1901 ( .A(n1231), .B(n2291), .Z(n2293) );
  XNOR U1902 ( .A(n2292), .B(n2289), .Z(n2291) );
  XOR U1903 ( .A(n2294), .B(n2295), .Z(n2289) );
  AND U1904 ( .A(n1234), .B(n2296), .Z(n2295) );
  XOR U1905 ( .A(p_input[1752]), .B(n2294), .Z(n2296) );
  XOR U1906 ( .A(n2297), .B(n2298), .Z(n2294) );
  AND U1907 ( .A(n1238), .B(n2299), .Z(n2298) );
  XOR U1908 ( .A(n2300), .B(n2301), .Z(n2292) );
  AND U1909 ( .A(n1242), .B(n2299), .Z(n2301) );
  XNOR U1910 ( .A(n2300), .B(n2297), .Z(n2299) );
  XOR U1911 ( .A(n2302), .B(n2303), .Z(n2297) );
  AND U1912 ( .A(n1245), .B(n2304), .Z(n2303) );
  XOR U1913 ( .A(p_input[1768]), .B(n2302), .Z(n2304) );
  XOR U1914 ( .A(n2305), .B(n2306), .Z(n2302) );
  AND U1915 ( .A(n1249), .B(n2307), .Z(n2306) );
  XOR U1916 ( .A(n2308), .B(n2309), .Z(n2300) );
  AND U1917 ( .A(n1253), .B(n2307), .Z(n2309) );
  XNOR U1918 ( .A(n2308), .B(n2305), .Z(n2307) );
  XOR U1919 ( .A(n2310), .B(n2311), .Z(n2305) );
  AND U1920 ( .A(n1256), .B(n2312), .Z(n2311) );
  XOR U1921 ( .A(p_input[1784]), .B(n2310), .Z(n2312) );
  XOR U1922 ( .A(n2313), .B(n2314), .Z(n2310) );
  AND U1923 ( .A(n1260), .B(n2315), .Z(n2314) );
  XOR U1924 ( .A(n2316), .B(n2317), .Z(n2308) );
  AND U1925 ( .A(n1264), .B(n2315), .Z(n2317) );
  XNOR U1926 ( .A(n2316), .B(n2313), .Z(n2315) );
  XOR U1927 ( .A(n2318), .B(n2319), .Z(n2313) );
  AND U1928 ( .A(n1267), .B(n2320), .Z(n2319) );
  XOR U1929 ( .A(p_input[1800]), .B(n2318), .Z(n2320) );
  XOR U1930 ( .A(n2321), .B(n2322), .Z(n2318) );
  AND U1931 ( .A(n1271), .B(n2323), .Z(n2322) );
  XOR U1932 ( .A(n2324), .B(n2325), .Z(n2316) );
  AND U1933 ( .A(n1275), .B(n2323), .Z(n2325) );
  XNOR U1934 ( .A(n2324), .B(n2321), .Z(n2323) );
  XOR U1935 ( .A(n2326), .B(n2327), .Z(n2321) );
  AND U1936 ( .A(n1278), .B(n2328), .Z(n2327) );
  XOR U1937 ( .A(p_input[1816]), .B(n2326), .Z(n2328) );
  XOR U1938 ( .A(n2329), .B(n2330), .Z(n2326) );
  AND U1939 ( .A(n1282), .B(n2331), .Z(n2330) );
  XOR U1940 ( .A(n2332), .B(n2333), .Z(n2324) );
  AND U1941 ( .A(n1286), .B(n2331), .Z(n2333) );
  XNOR U1942 ( .A(n2332), .B(n2329), .Z(n2331) );
  XOR U1943 ( .A(n2334), .B(n2335), .Z(n2329) );
  AND U1944 ( .A(n1289), .B(n2336), .Z(n2335) );
  XOR U1945 ( .A(p_input[1832]), .B(n2334), .Z(n2336) );
  XOR U1946 ( .A(n2337), .B(n2338), .Z(n2334) );
  AND U1947 ( .A(n1293), .B(n2339), .Z(n2338) );
  XOR U1948 ( .A(n2340), .B(n2341), .Z(n2332) );
  AND U1949 ( .A(n1297), .B(n2339), .Z(n2341) );
  XNOR U1950 ( .A(n2340), .B(n2337), .Z(n2339) );
  XOR U1951 ( .A(n2342), .B(n2343), .Z(n2337) );
  AND U1952 ( .A(n1300), .B(n2344), .Z(n2343) );
  XOR U1953 ( .A(p_input[1848]), .B(n2342), .Z(n2344) );
  XOR U1954 ( .A(n2345), .B(n2346), .Z(n2342) );
  AND U1955 ( .A(n1304), .B(n2347), .Z(n2346) );
  XOR U1956 ( .A(n2348), .B(n2349), .Z(n2340) );
  AND U1957 ( .A(n1308), .B(n2347), .Z(n2349) );
  XNOR U1958 ( .A(n2348), .B(n2345), .Z(n2347) );
  XOR U1959 ( .A(n2350), .B(n2351), .Z(n2345) );
  AND U1960 ( .A(n1311), .B(n2352), .Z(n2351) );
  XOR U1961 ( .A(p_input[1864]), .B(n2350), .Z(n2352) );
  XOR U1962 ( .A(n2353), .B(n2354), .Z(n2350) );
  AND U1963 ( .A(n1315), .B(n2355), .Z(n2354) );
  XOR U1964 ( .A(n2356), .B(n2357), .Z(n2348) );
  AND U1965 ( .A(n1319), .B(n2355), .Z(n2357) );
  XNOR U1966 ( .A(n2356), .B(n2353), .Z(n2355) );
  XOR U1967 ( .A(n2358), .B(n2359), .Z(n2353) );
  AND U1968 ( .A(n1322), .B(n2360), .Z(n2359) );
  XOR U1969 ( .A(p_input[1880]), .B(n2358), .Z(n2360) );
  XOR U1970 ( .A(n2361), .B(n2362), .Z(n2358) );
  AND U1971 ( .A(n1326), .B(n2363), .Z(n2362) );
  XOR U1972 ( .A(n2364), .B(n2365), .Z(n2356) );
  AND U1973 ( .A(n1330), .B(n2363), .Z(n2365) );
  XNOR U1974 ( .A(n2364), .B(n2361), .Z(n2363) );
  XOR U1975 ( .A(n2366), .B(n2367), .Z(n2361) );
  AND U1976 ( .A(n1333), .B(n2368), .Z(n2367) );
  XOR U1977 ( .A(p_input[1896]), .B(n2366), .Z(n2368) );
  XOR U1978 ( .A(n2369), .B(n2370), .Z(n2366) );
  AND U1979 ( .A(n1337), .B(n2371), .Z(n2370) );
  XOR U1980 ( .A(n2372), .B(n2373), .Z(n2364) );
  AND U1981 ( .A(n1341), .B(n2371), .Z(n2373) );
  XNOR U1982 ( .A(n2372), .B(n2369), .Z(n2371) );
  XOR U1983 ( .A(n2374), .B(n2375), .Z(n2369) );
  AND U1984 ( .A(n1344), .B(n2376), .Z(n2375) );
  XOR U1985 ( .A(p_input[1912]), .B(n2374), .Z(n2376) );
  XOR U1986 ( .A(n2377), .B(n2378), .Z(n2374) );
  AND U1987 ( .A(n1348), .B(n2379), .Z(n2378) );
  XOR U1988 ( .A(n2380), .B(n2381), .Z(n2372) );
  AND U1989 ( .A(n1352), .B(n2379), .Z(n2381) );
  XNOR U1990 ( .A(n2380), .B(n2377), .Z(n2379) );
  XOR U1991 ( .A(n2382), .B(n2383), .Z(n2377) );
  AND U1992 ( .A(n1355), .B(n2384), .Z(n2383) );
  XOR U1993 ( .A(p_input[1928]), .B(n2382), .Z(n2384) );
  XOR U1994 ( .A(n2385), .B(n2386), .Z(n2382) );
  AND U1995 ( .A(n1359), .B(n2387), .Z(n2386) );
  XOR U1996 ( .A(n2388), .B(n2389), .Z(n2380) );
  AND U1997 ( .A(n1363), .B(n2387), .Z(n2389) );
  XNOR U1998 ( .A(n2388), .B(n2385), .Z(n2387) );
  XOR U1999 ( .A(n2390), .B(n2391), .Z(n2385) );
  AND U2000 ( .A(n1366), .B(n2392), .Z(n2391) );
  XOR U2001 ( .A(p_input[1944]), .B(n2390), .Z(n2392) );
  XOR U2002 ( .A(n2393), .B(n2394), .Z(n2390) );
  AND U2003 ( .A(n1370), .B(n2395), .Z(n2394) );
  XOR U2004 ( .A(n2396), .B(n2397), .Z(n2388) );
  AND U2005 ( .A(n1374), .B(n2395), .Z(n2397) );
  XNOR U2006 ( .A(n2396), .B(n2393), .Z(n2395) );
  XOR U2007 ( .A(n2398), .B(n2399), .Z(n2393) );
  AND U2008 ( .A(n1377), .B(n2400), .Z(n2399) );
  XOR U2009 ( .A(p_input[1960]), .B(n2398), .Z(n2400) );
  XOR U2010 ( .A(n2401), .B(n2402), .Z(n2398) );
  AND U2011 ( .A(n1381), .B(n2403), .Z(n2402) );
  XOR U2012 ( .A(n2404), .B(n2405), .Z(n2396) );
  AND U2013 ( .A(n1385), .B(n2403), .Z(n2405) );
  XNOR U2014 ( .A(n2404), .B(n2401), .Z(n2403) );
  XOR U2015 ( .A(n2406), .B(n2407), .Z(n2401) );
  AND U2016 ( .A(n1388), .B(n2408), .Z(n2407) );
  XOR U2017 ( .A(p_input[1976]), .B(n2406), .Z(n2408) );
  XOR U2018 ( .A(n2409), .B(n2410), .Z(n2406) );
  AND U2019 ( .A(n1392), .B(n2411), .Z(n2410) );
  XOR U2020 ( .A(n2412), .B(n2413), .Z(n2404) );
  AND U2021 ( .A(n1396), .B(n2411), .Z(n2413) );
  XNOR U2022 ( .A(n2412), .B(n2409), .Z(n2411) );
  XOR U2023 ( .A(n2414), .B(n2415), .Z(n2409) );
  AND U2024 ( .A(n1399), .B(n2416), .Z(n2415) );
  XOR U2025 ( .A(p_input[1992]), .B(n2414), .Z(n2416) );
  XOR U2026 ( .A(n2417), .B(n2418), .Z(n2414) );
  AND U2027 ( .A(n1403), .B(n2419), .Z(n2418) );
  XOR U2028 ( .A(n2420), .B(n2421), .Z(n2412) );
  AND U2029 ( .A(n1407), .B(n2419), .Z(n2421) );
  XNOR U2030 ( .A(n2420), .B(n2417), .Z(n2419) );
  XOR U2031 ( .A(n2422), .B(n2423), .Z(n2417) );
  AND U2032 ( .A(n1410), .B(n2424), .Z(n2423) );
  XOR U2033 ( .A(p_input[2008]), .B(n2422), .Z(n2424) );
  XNOR U2034 ( .A(n2425), .B(n2426), .Z(n2422) );
  AND U2035 ( .A(n1414), .B(n2427), .Z(n2426) );
  XNOR U2036 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n2428), .Z(n2420) );
  AND U2037 ( .A(n1417), .B(n2427), .Z(n2428) );
  XOR U2038 ( .A(n2429), .B(n2425), .Z(n2427) );
  XOR U2039 ( .A(n5), .B(n2430), .Z(o[23]) );
  AND U2040 ( .A(n30), .B(n2431), .Z(n5) );
  XOR U2041 ( .A(n6), .B(n2430), .Z(n2431) );
  XOR U2042 ( .A(n2432), .B(n2433), .Z(n2430) );
  AND U2043 ( .A(n34), .B(n2434), .Z(n2433) );
  XOR U2044 ( .A(p_input[7]), .B(n2432), .Z(n2434) );
  XOR U2045 ( .A(n2435), .B(n2436), .Z(n2432) );
  AND U2046 ( .A(n38), .B(n2437), .Z(n2436) );
  XOR U2047 ( .A(n2438), .B(n2439), .Z(n6) );
  AND U2048 ( .A(n42), .B(n2437), .Z(n2439) );
  XNOR U2049 ( .A(n2440), .B(n2435), .Z(n2437) );
  XOR U2050 ( .A(n2441), .B(n2442), .Z(n2435) );
  AND U2051 ( .A(n46), .B(n2443), .Z(n2442) );
  XOR U2052 ( .A(p_input[23]), .B(n2441), .Z(n2443) );
  XOR U2053 ( .A(n2444), .B(n2445), .Z(n2441) );
  AND U2054 ( .A(n50), .B(n2446), .Z(n2445) );
  IV U2055 ( .A(n2438), .Z(n2440) );
  XNOR U2056 ( .A(n2447), .B(n2448), .Z(n2438) );
  AND U2057 ( .A(n54), .B(n2446), .Z(n2448) );
  XNOR U2058 ( .A(n2447), .B(n2444), .Z(n2446) );
  XOR U2059 ( .A(n2449), .B(n2450), .Z(n2444) );
  AND U2060 ( .A(n57), .B(n2451), .Z(n2450) );
  XOR U2061 ( .A(p_input[39]), .B(n2449), .Z(n2451) );
  XOR U2062 ( .A(n2452), .B(n2453), .Z(n2449) );
  AND U2063 ( .A(n61), .B(n2454), .Z(n2453) );
  XOR U2064 ( .A(n2455), .B(n2456), .Z(n2447) );
  AND U2065 ( .A(n65), .B(n2454), .Z(n2456) );
  XNOR U2066 ( .A(n2455), .B(n2452), .Z(n2454) );
  XOR U2067 ( .A(n2457), .B(n2458), .Z(n2452) );
  AND U2068 ( .A(n68), .B(n2459), .Z(n2458) );
  XOR U2069 ( .A(p_input[55]), .B(n2457), .Z(n2459) );
  XOR U2070 ( .A(n2460), .B(n2461), .Z(n2457) );
  AND U2071 ( .A(n72), .B(n2462), .Z(n2461) );
  XOR U2072 ( .A(n2463), .B(n2464), .Z(n2455) );
  AND U2073 ( .A(n76), .B(n2462), .Z(n2464) );
  XNOR U2074 ( .A(n2463), .B(n2460), .Z(n2462) );
  XOR U2075 ( .A(n2465), .B(n2466), .Z(n2460) );
  AND U2076 ( .A(n79), .B(n2467), .Z(n2466) );
  XOR U2077 ( .A(p_input[71]), .B(n2465), .Z(n2467) );
  XOR U2078 ( .A(n2468), .B(n2469), .Z(n2465) );
  AND U2079 ( .A(n83), .B(n2470), .Z(n2469) );
  XOR U2080 ( .A(n2471), .B(n2472), .Z(n2463) );
  AND U2081 ( .A(n87), .B(n2470), .Z(n2472) );
  XNOR U2082 ( .A(n2471), .B(n2468), .Z(n2470) );
  XOR U2083 ( .A(n2473), .B(n2474), .Z(n2468) );
  AND U2084 ( .A(n90), .B(n2475), .Z(n2474) );
  XOR U2085 ( .A(p_input[87]), .B(n2473), .Z(n2475) );
  XOR U2086 ( .A(n2476), .B(n2477), .Z(n2473) );
  AND U2087 ( .A(n94), .B(n2478), .Z(n2477) );
  XOR U2088 ( .A(n2479), .B(n2480), .Z(n2471) );
  AND U2089 ( .A(n98), .B(n2478), .Z(n2480) );
  XNOR U2090 ( .A(n2479), .B(n2476), .Z(n2478) );
  XOR U2091 ( .A(n2481), .B(n2482), .Z(n2476) );
  AND U2092 ( .A(n101), .B(n2483), .Z(n2482) );
  XOR U2093 ( .A(p_input[103]), .B(n2481), .Z(n2483) );
  XOR U2094 ( .A(n2484), .B(n2485), .Z(n2481) );
  AND U2095 ( .A(n105), .B(n2486), .Z(n2485) );
  XOR U2096 ( .A(n2487), .B(n2488), .Z(n2479) );
  AND U2097 ( .A(n109), .B(n2486), .Z(n2488) );
  XNOR U2098 ( .A(n2487), .B(n2484), .Z(n2486) );
  XOR U2099 ( .A(n2489), .B(n2490), .Z(n2484) );
  AND U2100 ( .A(n112), .B(n2491), .Z(n2490) );
  XOR U2101 ( .A(p_input[119]), .B(n2489), .Z(n2491) );
  XOR U2102 ( .A(n2492), .B(n2493), .Z(n2489) );
  AND U2103 ( .A(n116), .B(n2494), .Z(n2493) );
  XOR U2104 ( .A(n2495), .B(n2496), .Z(n2487) );
  AND U2105 ( .A(n120), .B(n2494), .Z(n2496) );
  XNOR U2106 ( .A(n2495), .B(n2492), .Z(n2494) );
  XOR U2107 ( .A(n2497), .B(n2498), .Z(n2492) );
  AND U2108 ( .A(n123), .B(n2499), .Z(n2498) );
  XOR U2109 ( .A(p_input[135]), .B(n2497), .Z(n2499) );
  XOR U2110 ( .A(n2500), .B(n2501), .Z(n2497) );
  AND U2111 ( .A(n127), .B(n2502), .Z(n2501) );
  XOR U2112 ( .A(n2503), .B(n2504), .Z(n2495) );
  AND U2113 ( .A(n131), .B(n2502), .Z(n2504) );
  XNOR U2114 ( .A(n2503), .B(n2500), .Z(n2502) );
  XOR U2115 ( .A(n2505), .B(n2506), .Z(n2500) );
  AND U2116 ( .A(n134), .B(n2507), .Z(n2506) );
  XOR U2117 ( .A(p_input[151]), .B(n2505), .Z(n2507) );
  XOR U2118 ( .A(n2508), .B(n2509), .Z(n2505) );
  AND U2119 ( .A(n138), .B(n2510), .Z(n2509) );
  XOR U2120 ( .A(n2511), .B(n2512), .Z(n2503) );
  AND U2121 ( .A(n142), .B(n2510), .Z(n2512) );
  XNOR U2122 ( .A(n2511), .B(n2508), .Z(n2510) );
  XOR U2123 ( .A(n2513), .B(n2514), .Z(n2508) );
  AND U2124 ( .A(n145), .B(n2515), .Z(n2514) );
  XOR U2125 ( .A(p_input[167]), .B(n2513), .Z(n2515) );
  XOR U2126 ( .A(n2516), .B(n2517), .Z(n2513) );
  AND U2127 ( .A(n149), .B(n2518), .Z(n2517) );
  XOR U2128 ( .A(n2519), .B(n2520), .Z(n2511) );
  AND U2129 ( .A(n153), .B(n2518), .Z(n2520) );
  XNOR U2130 ( .A(n2519), .B(n2516), .Z(n2518) );
  XOR U2131 ( .A(n2521), .B(n2522), .Z(n2516) );
  AND U2132 ( .A(n156), .B(n2523), .Z(n2522) );
  XOR U2133 ( .A(p_input[183]), .B(n2521), .Z(n2523) );
  XOR U2134 ( .A(n2524), .B(n2525), .Z(n2521) );
  AND U2135 ( .A(n160), .B(n2526), .Z(n2525) );
  XOR U2136 ( .A(n2527), .B(n2528), .Z(n2519) );
  AND U2137 ( .A(n164), .B(n2526), .Z(n2528) );
  XNOR U2138 ( .A(n2527), .B(n2524), .Z(n2526) );
  XOR U2139 ( .A(n2529), .B(n2530), .Z(n2524) );
  AND U2140 ( .A(n167), .B(n2531), .Z(n2530) );
  XOR U2141 ( .A(p_input[199]), .B(n2529), .Z(n2531) );
  XOR U2142 ( .A(n2532), .B(n2533), .Z(n2529) );
  AND U2143 ( .A(n171), .B(n2534), .Z(n2533) );
  XOR U2144 ( .A(n2535), .B(n2536), .Z(n2527) );
  AND U2145 ( .A(n175), .B(n2534), .Z(n2536) );
  XNOR U2146 ( .A(n2535), .B(n2532), .Z(n2534) );
  XOR U2147 ( .A(n2537), .B(n2538), .Z(n2532) );
  AND U2148 ( .A(n178), .B(n2539), .Z(n2538) );
  XOR U2149 ( .A(p_input[215]), .B(n2537), .Z(n2539) );
  XOR U2150 ( .A(n2540), .B(n2541), .Z(n2537) );
  AND U2151 ( .A(n182), .B(n2542), .Z(n2541) );
  XOR U2152 ( .A(n2543), .B(n2544), .Z(n2535) );
  AND U2153 ( .A(n186), .B(n2542), .Z(n2544) );
  XNOR U2154 ( .A(n2543), .B(n2540), .Z(n2542) );
  XOR U2155 ( .A(n2545), .B(n2546), .Z(n2540) );
  AND U2156 ( .A(n189), .B(n2547), .Z(n2546) );
  XOR U2157 ( .A(p_input[231]), .B(n2545), .Z(n2547) );
  XOR U2158 ( .A(n2548), .B(n2549), .Z(n2545) );
  AND U2159 ( .A(n193), .B(n2550), .Z(n2549) );
  XOR U2160 ( .A(n2551), .B(n2552), .Z(n2543) );
  AND U2161 ( .A(n197), .B(n2550), .Z(n2552) );
  XNOR U2162 ( .A(n2551), .B(n2548), .Z(n2550) );
  XOR U2163 ( .A(n2553), .B(n2554), .Z(n2548) );
  AND U2164 ( .A(n200), .B(n2555), .Z(n2554) );
  XOR U2165 ( .A(p_input[247]), .B(n2553), .Z(n2555) );
  XOR U2166 ( .A(n2556), .B(n2557), .Z(n2553) );
  AND U2167 ( .A(n204), .B(n2558), .Z(n2557) );
  XOR U2168 ( .A(n2559), .B(n2560), .Z(n2551) );
  AND U2169 ( .A(n208), .B(n2558), .Z(n2560) );
  XNOR U2170 ( .A(n2559), .B(n2556), .Z(n2558) );
  XOR U2171 ( .A(n2561), .B(n2562), .Z(n2556) );
  AND U2172 ( .A(n211), .B(n2563), .Z(n2562) );
  XOR U2173 ( .A(p_input[263]), .B(n2561), .Z(n2563) );
  XOR U2174 ( .A(n2564), .B(n2565), .Z(n2561) );
  AND U2175 ( .A(n215), .B(n2566), .Z(n2565) );
  XOR U2176 ( .A(n2567), .B(n2568), .Z(n2559) );
  AND U2177 ( .A(n219), .B(n2566), .Z(n2568) );
  XNOR U2178 ( .A(n2567), .B(n2564), .Z(n2566) );
  XOR U2179 ( .A(n2569), .B(n2570), .Z(n2564) );
  AND U2180 ( .A(n222), .B(n2571), .Z(n2570) );
  XOR U2181 ( .A(p_input[279]), .B(n2569), .Z(n2571) );
  XOR U2182 ( .A(n2572), .B(n2573), .Z(n2569) );
  AND U2183 ( .A(n226), .B(n2574), .Z(n2573) );
  XOR U2184 ( .A(n2575), .B(n2576), .Z(n2567) );
  AND U2185 ( .A(n230), .B(n2574), .Z(n2576) );
  XNOR U2186 ( .A(n2575), .B(n2572), .Z(n2574) );
  XOR U2187 ( .A(n2577), .B(n2578), .Z(n2572) );
  AND U2188 ( .A(n233), .B(n2579), .Z(n2578) );
  XOR U2189 ( .A(p_input[295]), .B(n2577), .Z(n2579) );
  XOR U2190 ( .A(n2580), .B(n2581), .Z(n2577) );
  AND U2191 ( .A(n237), .B(n2582), .Z(n2581) );
  XOR U2192 ( .A(n2583), .B(n2584), .Z(n2575) );
  AND U2193 ( .A(n241), .B(n2582), .Z(n2584) );
  XNOR U2194 ( .A(n2583), .B(n2580), .Z(n2582) );
  XOR U2195 ( .A(n2585), .B(n2586), .Z(n2580) );
  AND U2196 ( .A(n244), .B(n2587), .Z(n2586) );
  XOR U2197 ( .A(p_input[311]), .B(n2585), .Z(n2587) );
  XOR U2198 ( .A(n2588), .B(n2589), .Z(n2585) );
  AND U2199 ( .A(n248), .B(n2590), .Z(n2589) );
  XOR U2200 ( .A(n2591), .B(n2592), .Z(n2583) );
  AND U2201 ( .A(n252), .B(n2590), .Z(n2592) );
  XNOR U2202 ( .A(n2591), .B(n2588), .Z(n2590) );
  XOR U2203 ( .A(n2593), .B(n2594), .Z(n2588) );
  AND U2204 ( .A(n255), .B(n2595), .Z(n2594) );
  XOR U2205 ( .A(p_input[327]), .B(n2593), .Z(n2595) );
  XOR U2206 ( .A(n2596), .B(n2597), .Z(n2593) );
  AND U2207 ( .A(n259), .B(n2598), .Z(n2597) );
  XOR U2208 ( .A(n2599), .B(n2600), .Z(n2591) );
  AND U2209 ( .A(n263), .B(n2598), .Z(n2600) );
  XNOR U2210 ( .A(n2599), .B(n2596), .Z(n2598) );
  XOR U2211 ( .A(n2601), .B(n2602), .Z(n2596) );
  AND U2212 ( .A(n266), .B(n2603), .Z(n2602) );
  XOR U2213 ( .A(p_input[343]), .B(n2601), .Z(n2603) );
  XOR U2214 ( .A(n2604), .B(n2605), .Z(n2601) );
  AND U2215 ( .A(n270), .B(n2606), .Z(n2605) );
  XOR U2216 ( .A(n2607), .B(n2608), .Z(n2599) );
  AND U2217 ( .A(n274), .B(n2606), .Z(n2608) );
  XNOR U2218 ( .A(n2607), .B(n2604), .Z(n2606) );
  XOR U2219 ( .A(n2609), .B(n2610), .Z(n2604) );
  AND U2220 ( .A(n277), .B(n2611), .Z(n2610) );
  XOR U2221 ( .A(p_input[359]), .B(n2609), .Z(n2611) );
  XOR U2222 ( .A(n2612), .B(n2613), .Z(n2609) );
  AND U2223 ( .A(n281), .B(n2614), .Z(n2613) );
  XOR U2224 ( .A(n2615), .B(n2616), .Z(n2607) );
  AND U2225 ( .A(n285), .B(n2614), .Z(n2616) );
  XNOR U2226 ( .A(n2615), .B(n2612), .Z(n2614) );
  XOR U2227 ( .A(n2617), .B(n2618), .Z(n2612) );
  AND U2228 ( .A(n288), .B(n2619), .Z(n2618) );
  XOR U2229 ( .A(p_input[375]), .B(n2617), .Z(n2619) );
  XOR U2230 ( .A(n2620), .B(n2621), .Z(n2617) );
  AND U2231 ( .A(n292), .B(n2622), .Z(n2621) );
  XOR U2232 ( .A(n2623), .B(n2624), .Z(n2615) );
  AND U2233 ( .A(n296), .B(n2622), .Z(n2624) );
  XNOR U2234 ( .A(n2623), .B(n2620), .Z(n2622) );
  XOR U2235 ( .A(n2625), .B(n2626), .Z(n2620) );
  AND U2236 ( .A(n299), .B(n2627), .Z(n2626) );
  XOR U2237 ( .A(p_input[391]), .B(n2625), .Z(n2627) );
  XOR U2238 ( .A(n2628), .B(n2629), .Z(n2625) );
  AND U2239 ( .A(n303), .B(n2630), .Z(n2629) );
  XOR U2240 ( .A(n2631), .B(n2632), .Z(n2623) );
  AND U2241 ( .A(n307), .B(n2630), .Z(n2632) );
  XNOR U2242 ( .A(n2631), .B(n2628), .Z(n2630) );
  XOR U2243 ( .A(n2633), .B(n2634), .Z(n2628) );
  AND U2244 ( .A(n310), .B(n2635), .Z(n2634) );
  XOR U2245 ( .A(p_input[407]), .B(n2633), .Z(n2635) );
  XOR U2246 ( .A(n2636), .B(n2637), .Z(n2633) );
  AND U2247 ( .A(n314), .B(n2638), .Z(n2637) );
  XOR U2248 ( .A(n2639), .B(n2640), .Z(n2631) );
  AND U2249 ( .A(n318), .B(n2638), .Z(n2640) );
  XNOR U2250 ( .A(n2639), .B(n2636), .Z(n2638) );
  XOR U2251 ( .A(n2641), .B(n2642), .Z(n2636) );
  AND U2252 ( .A(n321), .B(n2643), .Z(n2642) );
  XOR U2253 ( .A(p_input[423]), .B(n2641), .Z(n2643) );
  XOR U2254 ( .A(n2644), .B(n2645), .Z(n2641) );
  AND U2255 ( .A(n325), .B(n2646), .Z(n2645) );
  XOR U2256 ( .A(n2647), .B(n2648), .Z(n2639) );
  AND U2257 ( .A(n329), .B(n2646), .Z(n2648) );
  XNOR U2258 ( .A(n2647), .B(n2644), .Z(n2646) );
  XOR U2259 ( .A(n2649), .B(n2650), .Z(n2644) );
  AND U2260 ( .A(n332), .B(n2651), .Z(n2650) );
  XOR U2261 ( .A(p_input[439]), .B(n2649), .Z(n2651) );
  XOR U2262 ( .A(n2652), .B(n2653), .Z(n2649) );
  AND U2263 ( .A(n336), .B(n2654), .Z(n2653) );
  XOR U2264 ( .A(n2655), .B(n2656), .Z(n2647) );
  AND U2265 ( .A(n340), .B(n2654), .Z(n2656) );
  XNOR U2266 ( .A(n2655), .B(n2652), .Z(n2654) );
  XOR U2267 ( .A(n2657), .B(n2658), .Z(n2652) );
  AND U2268 ( .A(n343), .B(n2659), .Z(n2658) );
  XOR U2269 ( .A(p_input[455]), .B(n2657), .Z(n2659) );
  XOR U2270 ( .A(n2660), .B(n2661), .Z(n2657) );
  AND U2271 ( .A(n347), .B(n2662), .Z(n2661) );
  XOR U2272 ( .A(n2663), .B(n2664), .Z(n2655) );
  AND U2273 ( .A(n351), .B(n2662), .Z(n2664) );
  XNOR U2274 ( .A(n2663), .B(n2660), .Z(n2662) );
  XOR U2275 ( .A(n2665), .B(n2666), .Z(n2660) );
  AND U2276 ( .A(n354), .B(n2667), .Z(n2666) );
  XOR U2277 ( .A(p_input[471]), .B(n2665), .Z(n2667) );
  XOR U2278 ( .A(n2668), .B(n2669), .Z(n2665) );
  AND U2279 ( .A(n358), .B(n2670), .Z(n2669) );
  XOR U2280 ( .A(n2671), .B(n2672), .Z(n2663) );
  AND U2281 ( .A(n362), .B(n2670), .Z(n2672) );
  XNOR U2282 ( .A(n2671), .B(n2668), .Z(n2670) );
  XOR U2283 ( .A(n2673), .B(n2674), .Z(n2668) );
  AND U2284 ( .A(n365), .B(n2675), .Z(n2674) );
  XOR U2285 ( .A(p_input[487]), .B(n2673), .Z(n2675) );
  XOR U2286 ( .A(n2676), .B(n2677), .Z(n2673) );
  AND U2287 ( .A(n369), .B(n2678), .Z(n2677) );
  XOR U2288 ( .A(n2679), .B(n2680), .Z(n2671) );
  AND U2289 ( .A(n373), .B(n2678), .Z(n2680) );
  XNOR U2290 ( .A(n2679), .B(n2676), .Z(n2678) );
  XOR U2291 ( .A(n2681), .B(n2682), .Z(n2676) );
  AND U2292 ( .A(n376), .B(n2683), .Z(n2682) );
  XOR U2293 ( .A(p_input[503]), .B(n2681), .Z(n2683) );
  XOR U2294 ( .A(n2684), .B(n2685), .Z(n2681) );
  AND U2295 ( .A(n380), .B(n2686), .Z(n2685) );
  XOR U2296 ( .A(n2687), .B(n2688), .Z(n2679) );
  AND U2297 ( .A(n384), .B(n2686), .Z(n2688) );
  XNOR U2298 ( .A(n2687), .B(n2684), .Z(n2686) );
  XOR U2299 ( .A(n2689), .B(n2690), .Z(n2684) );
  AND U2300 ( .A(n387), .B(n2691), .Z(n2690) );
  XOR U2301 ( .A(p_input[519]), .B(n2689), .Z(n2691) );
  XOR U2302 ( .A(n2692), .B(n2693), .Z(n2689) );
  AND U2303 ( .A(n391), .B(n2694), .Z(n2693) );
  XOR U2304 ( .A(n2695), .B(n2696), .Z(n2687) );
  AND U2305 ( .A(n395), .B(n2694), .Z(n2696) );
  XNOR U2306 ( .A(n2695), .B(n2692), .Z(n2694) );
  XOR U2307 ( .A(n2697), .B(n2698), .Z(n2692) );
  AND U2308 ( .A(n398), .B(n2699), .Z(n2698) );
  XOR U2309 ( .A(p_input[535]), .B(n2697), .Z(n2699) );
  XOR U2310 ( .A(n2700), .B(n2701), .Z(n2697) );
  AND U2311 ( .A(n402), .B(n2702), .Z(n2701) );
  XOR U2312 ( .A(n2703), .B(n2704), .Z(n2695) );
  AND U2313 ( .A(n406), .B(n2702), .Z(n2704) );
  XNOR U2314 ( .A(n2703), .B(n2700), .Z(n2702) );
  XOR U2315 ( .A(n2705), .B(n2706), .Z(n2700) );
  AND U2316 ( .A(n409), .B(n2707), .Z(n2706) );
  XOR U2317 ( .A(p_input[551]), .B(n2705), .Z(n2707) );
  XOR U2318 ( .A(n2708), .B(n2709), .Z(n2705) );
  AND U2319 ( .A(n413), .B(n2710), .Z(n2709) );
  XOR U2320 ( .A(n2711), .B(n2712), .Z(n2703) );
  AND U2321 ( .A(n417), .B(n2710), .Z(n2712) );
  XNOR U2322 ( .A(n2711), .B(n2708), .Z(n2710) );
  XOR U2323 ( .A(n2713), .B(n2714), .Z(n2708) );
  AND U2324 ( .A(n420), .B(n2715), .Z(n2714) );
  XOR U2325 ( .A(p_input[567]), .B(n2713), .Z(n2715) );
  XOR U2326 ( .A(n2716), .B(n2717), .Z(n2713) );
  AND U2327 ( .A(n424), .B(n2718), .Z(n2717) );
  XOR U2328 ( .A(n2719), .B(n2720), .Z(n2711) );
  AND U2329 ( .A(n428), .B(n2718), .Z(n2720) );
  XNOR U2330 ( .A(n2719), .B(n2716), .Z(n2718) );
  XOR U2331 ( .A(n2721), .B(n2722), .Z(n2716) );
  AND U2332 ( .A(n431), .B(n2723), .Z(n2722) );
  XOR U2333 ( .A(p_input[583]), .B(n2721), .Z(n2723) );
  XOR U2334 ( .A(n2724), .B(n2725), .Z(n2721) );
  AND U2335 ( .A(n435), .B(n2726), .Z(n2725) );
  XOR U2336 ( .A(n2727), .B(n2728), .Z(n2719) );
  AND U2337 ( .A(n439), .B(n2726), .Z(n2728) );
  XNOR U2338 ( .A(n2727), .B(n2724), .Z(n2726) );
  XOR U2339 ( .A(n2729), .B(n2730), .Z(n2724) );
  AND U2340 ( .A(n442), .B(n2731), .Z(n2730) );
  XOR U2341 ( .A(p_input[599]), .B(n2729), .Z(n2731) );
  XOR U2342 ( .A(n2732), .B(n2733), .Z(n2729) );
  AND U2343 ( .A(n446), .B(n2734), .Z(n2733) );
  XOR U2344 ( .A(n2735), .B(n2736), .Z(n2727) );
  AND U2345 ( .A(n450), .B(n2734), .Z(n2736) );
  XNOR U2346 ( .A(n2735), .B(n2732), .Z(n2734) );
  XOR U2347 ( .A(n2737), .B(n2738), .Z(n2732) );
  AND U2348 ( .A(n453), .B(n2739), .Z(n2738) );
  XOR U2349 ( .A(p_input[615]), .B(n2737), .Z(n2739) );
  XOR U2350 ( .A(n2740), .B(n2741), .Z(n2737) );
  AND U2351 ( .A(n457), .B(n2742), .Z(n2741) );
  XOR U2352 ( .A(n2743), .B(n2744), .Z(n2735) );
  AND U2353 ( .A(n461), .B(n2742), .Z(n2744) );
  XNOR U2354 ( .A(n2743), .B(n2740), .Z(n2742) );
  XOR U2355 ( .A(n2745), .B(n2746), .Z(n2740) );
  AND U2356 ( .A(n464), .B(n2747), .Z(n2746) );
  XOR U2357 ( .A(p_input[631]), .B(n2745), .Z(n2747) );
  XOR U2358 ( .A(n2748), .B(n2749), .Z(n2745) );
  AND U2359 ( .A(n468), .B(n2750), .Z(n2749) );
  XOR U2360 ( .A(n2751), .B(n2752), .Z(n2743) );
  AND U2361 ( .A(n472), .B(n2750), .Z(n2752) );
  XNOR U2362 ( .A(n2751), .B(n2748), .Z(n2750) );
  XOR U2363 ( .A(n2753), .B(n2754), .Z(n2748) );
  AND U2364 ( .A(n475), .B(n2755), .Z(n2754) );
  XOR U2365 ( .A(p_input[647]), .B(n2753), .Z(n2755) );
  XOR U2366 ( .A(n2756), .B(n2757), .Z(n2753) );
  AND U2367 ( .A(n479), .B(n2758), .Z(n2757) );
  XOR U2368 ( .A(n2759), .B(n2760), .Z(n2751) );
  AND U2369 ( .A(n483), .B(n2758), .Z(n2760) );
  XNOR U2370 ( .A(n2759), .B(n2756), .Z(n2758) );
  XOR U2371 ( .A(n2761), .B(n2762), .Z(n2756) );
  AND U2372 ( .A(n486), .B(n2763), .Z(n2762) );
  XOR U2373 ( .A(p_input[663]), .B(n2761), .Z(n2763) );
  XOR U2374 ( .A(n2764), .B(n2765), .Z(n2761) );
  AND U2375 ( .A(n490), .B(n2766), .Z(n2765) );
  XOR U2376 ( .A(n2767), .B(n2768), .Z(n2759) );
  AND U2377 ( .A(n494), .B(n2766), .Z(n2768) );
  XNOR U2378 ( .A(n2767), .B(n2764), .Z(n2766) );
  XOR U2379 ( .A(n2769), .B(n2770), .Z(n2764) );
  AND U2380 ( .A(n497), .B(n2771), .Z(n2770) );
  XOR U2381 ( .A(p_input[679]), .B(n2769), .Z(n2771) );
  XOR U2382 ( .A(n2772), .B(n2773), .Z(n2769) );
  AND U2383 ( .A(n501), .B(n2774), .Z(n2773) );
  XOR U2384 ( .A(n2775), .B(n2776), .Z(n2767) );
  AND U2385 ( .A(n505), .B(n2774), .Z(n2776) );
  XNOR U2386 ( .A(n2775), .B(n2772), .Z(n2774) );
  XOR U2387 ( .A(n2777), .B(n2778), .Z(n2772) );
  AND U2388 ( .A(n508), .B(n2779), .Z(n2778) );
  XOR U2389 ( .A(p_input[695]), .B(n2777), .Z(n2779) );
  XOR U2390 ( .A(n2780), .B(n2781), .Z(n2777) );
  AND U2391 ( .A(n512), .B(n2782), .Z(n2781) );
  XOR U2392 ( .A(n2783), .B(n2784), .Z(n2775) );
  AND U2393 ( .A(n516), .B(n2782), .Z(n2784) );
  XNOR U2394 ( .A(n2783), .B(n2780), .Z(n2782) );
  XOR U2395 ( .A(n2785), .B(n2786), .Z(n2780) );
  AND U2396 ( .A(n519), .B(n2787), .Z(n2786) );
  XOR U2397 ( .A(p_input[711]), .B(n2785), .Z(n2787) );
  XOR U2398 ( .A(n2788), .B(n2789), .Z(n2785) );
  AND U2399 ( .A(n523), .B(n2790), .Z(n2789) );
  XOR U2400 ( .A(n2791), .B(n2792), .Z(n2783) );
  AND U2401 ( .A(n527), .B(n2790), .Z(n2792) );
  XNOR U2402 ( .A(n2791), .B(n2788), .Z(n2790) );
  XOR U2403 ( .A(n2793), .B(n2794), .Z(n2788) );
  AND U2404 ( .A(n530), .B(n2795), .Z(n2794) );
  XOR U2405 ( .A(p_input[727]), .B(n2793), .Z(n2795) );
  XOR U2406 ( .A(n2796), .B(n2797), .Z(n2793) );
  AND U2407 ( .A(n534), .B(n2798), .Z(n2797) );
  XOR U2408 ( .A(n2799), .B(n2800), .Z(n2791) );
  AND U2409 ( .A(n538), .B(n2798), .Z(n2800) );
  XNOR U2410 ( .A(n2799), .B(n2796), .Z(n2798) );
  XOR U2411 ( .A(n2801), .B(n2802), .Z(n2796) );
  AND U2412 ( .A(n541), .B(n2803), .Z(n2802) );
  XOR U2413 ( .A(p_input[743]), .B(n2801), .Z(n2803) );
  XOR U2414 ( .A(n2804), .B(n2805), .Z(n2801) );
  AND U2415 ( .A(n545), .B(n2806), .Z(n2805) );
  XOR U2416 ( .A(n2807), .B(n2808), .Z(n2799) );
  AND U2417 ( .A(n549), .B(n2806), .Z(n2808) );
  XNOR U2418 ( .A(n2807), .B(n2804), .Z(n2806) );
  XOR U2419 ( .A(n2809), .B(n2810), .Z(n2804) );
  AND U2420 ( .A(n552), .B(n2811), .Z(n2810) );
  XOR U2421 ( .A(p_input[759]), .B(n2809), .Z(n2811) );
  XOR U2422 ( .A(n2812), .B(n2813), .Z(n2809) );
  AND U2423 ( .A(n556), .B(n2814), .Z(n2813) );
  XOR U2424 ( .A(n2815), .B(n2816), .Z(n2807) );
  AND U2425 ( .A(n560), .B(n2814), .Z(n2816) );
  XNOR U2426 ( .A(n2815), .B(n2812), .Z(n2814) );
  XOR U2427 ( .A(n2817), .B(n2818), .Z(n2812) );
  AND U2428 ( .A(n563), .B(n2819), .Z(n2818) );
  XOR U2429 ( .A(p_input[775]), .B(n2817), .Z(n2819) );
  XOR U2430 ( .A(n2820), .B(n2821), .Z(n2817) );
  AND U2431 ( .A(n567), .B(n2822), .Z(n2821) );
  XOR U2432 ( .A(n2823), .B(n2824), .Z(n2815) );
  AND U2433 ( .A(n571), .B(n2822), .Z(n2824) );
  XNOR U2434 ( .A(n2823), .B(n2820), .Z(n2822) );
  XOR U2435 ( .A(n2825), .B(n2826), .Z(n2820) );
  AND U2436 ( .A(n574), .B(n2827), .Z(n2826) );
  XOR U2437 ( .A(p_input[791]), .B(n2825), .Z(n2827) );
  XOR U2438 ( .A(n2828), .B(n2829), .Z(n2825) );
  AND U2439 ( .A(n578), .B(n2830), .Z(n2829) );
  XOR U2440 ( .A(n2831), .B(n2832), .Z(n2823) );
  AND U2441 ( .A(n582), .B(n2830), .Z(n2832) );
  XNOR U2442 ( .A(n2831), .B(n2828), .Z(n2830) );
  XOR U2443 ( .A(n2833), .B(n2834), .Z(n2828) );
  AND U2444 ( .A(n585), .B(n2835), .Z(n2834) );
  XOR U2445 ( .A(p_input[807]), .B(n2833), .Z(n2835) );
  XOR U2446 ( .A(n2836), .B(n2837), .Z(n2833) );
  AND U2447 ( .A(n589), .B(n2838), .Z(n2837) );
  XOR U2448 ( .A(n2839), .B(n2840), .Z(n2831) );
  AND U2449 ( .A(n593), .B(n2838), .Z(n2840) );
  XNOR U2450 ( .A(n2839), .B(n2836), .Z(n2838) );
  XOR U2451 ( .A(n2841), .B(n2842), .Z(n2836) );
  AND U2452 ( .A(n596), .B(n2843), .Z(n2842) );
  XOR U2453 ( .A(p_input[823]), .B(n2841), .Z(n2843) );
  XOR U2454 ( .A(n2844), .B(n2845), .Z(n2841) );
  AND U2455 ( .A(n600), .B(n2846), .Z(n2845) );
  XOR U2456 ( .A(n2847), .B(n2848), .Z(n2839) );
  AND U2457 ( .A(n604), .B(n2846), .Z(n2848) );
  XNOR U2458 ( .A(n2847), .B(n2844), .Z(n2846) );
  XOR U2459 ( .A(n2849), .B(n2850), .Z(n2844) );
  AND U2460 ( .A(n607), .B(n2851), .Z(n2850) );
  XOR U2461 ( .A(p_input[839]), .B(n2849), .Z(n2851) );
  XOR U2462 ( .A(n2852), .B(n2853), .Z(n2849) );
  AND U2463 ( .A(n611), .B(n2854), .Z(n2853) );
  XOR U2464 ( .A(n2855), .B(n2856), .Z(n2847) );
  AND U2465 ( .A(n615), .B(n2854), .Z(n2856) );
  XNOR U2466 ( .A(n2855), .B(n2852), .Z(n2854) );
  XOR U2467 ( .A(n2857), .B(n2858), .Z(n2852) );
  AND U2468 ( .A(n618), .B(n2859), .Z(n2858) );
  XOR U2469 ( .A(p_input[855]), .B(n2857), .Z(n2859) );
  XOR U2470 ( .A(n2860), .B(n2861), .Z(n2857) );
  AND U2471 ( .A(n622), .B(n2862), .Z(n2861) );
  XOR U2472 ( .A(n2863), .B(n2864), .Z(n2855) );
  AND U2473 ( .A(n626), .B(n2862), .Z(n2864) );
  XNOR U2474 ( .A(n2863), .B(n2860), .Z(n2862) );
  XOR U2475 ( .A(n2865), .B(n2866), .Z(n2860) );
  AND U2476 ( .A(n629), .B(n2867), .Z(n2866) );
  XOR U2477 ( .A(p_input[871]), .B(n2865), .Z(n2867) );
  XOR U2478 ( .A(n2868), .B(n2869), .Z(n2865) );
  AND U2479 ( .A(n633), .B(n2870), .Z(n2869) );
  XOR U2480 ( .A(n2871), .B(n2872), .Z(n2863) );
  AND U2481 ( .A(n637), .B(n2870), .Z(n2872) );
  XNOR U2482 ( .A(n2871), .B(n2868), .Z(n2870) );
  XOR U2483 ( .A(n2873), .B(n2874), .Z(n2868) );
  AND U2484 ( .A(n640), .B(n2875), .Z(n2874) );
  XOR U2485 ( .A(p_input[887]), .B(n2873), .Z(n2875) );
  XOR U2486 ( .A(n2876), .B(n2877), .Z(n2873) );
  AND U2487 ( .A(n644), .B(n2878), .Z(n2877) );
  XOR U2488 ( .A(n2879), .B(n2880), .Z(n2871) );
  AND U2489 ( .A(n648), .B(n2878), .Z(n2880) );
  XNOR U2490 ( .A(n2879), .B(n2876), .Z(n2878) );
  XOR U2491 ( .A(n2881), .B(n2882), .Z(n2876) );
  AND U2492 ( .A(n651), .B(n2883), .Z(n2882) );
  XOR U2493 ( .A(p_input[903]), .B(n2881), .Z(n2883) );
  XOR U2494 ( .A(n2884), .B(n2885), .Z(n2881) );
  AND U2495 ( .A(n655), .B(n2886), .Z(n2885) );
  XOR U2496 ( .A(n2887), .B(n2888), .Z(n2879) );
  AND U2497 ( .A(n659), .B(n2886), .Z(n2888) );
  XNOR U2498 ( .A(n2887), .B(n2884), .Z(n2886) );
  XOR U2499 ( .A(n2889), .B(n2890), .Z(n2884) );
  AND U2500 ( .A(n662), .B(n2891), .Z(n2890) );
  XOR U2501 ( .A(p_input[919]), .B(n2889), .Z(n2891) );
  XOR U2502 ( .A(n2892), .B(n2893), .Z(n2889) );
  AND U2503 ( .A(n666), .B(n2894), .Z(n2893) );
  XOR U2504 ( .A(n2895), .B(n2896), .Z(n2887) );
  AND U2505 ( .A(n670), .B(n2894), .Z(n2896) );
  XNOR U2506 ( .A(n2895), .B(n2892), .Z(n2894) );
  XOR U2507 ( .A(n2897), .B(n2898), .Z(n2892) );
  AND U2508 ( .A(n673), .B(n2899), .Z(n2898) );
  XOR U2509 ( .A(p_input[935]), .B(n2897), .Z(n2899) );
  XOR U2510 ( .A(n2900), .B(n2901), .Z(n2897) );
  AND U2511 ( .A(n677), .B(n2902), .Z(n2901) );
  XOR U2512 ( .A(n2903), .B(n2904), .Z(n2895) );
  AND U2513 ( .A(n681), .B(n2902), .Z(n2904) );
  XNOR U2514 ( .A(n2903), .B(n2900), .Z(n2902) );
  XOR U2515 ( .A(n2905), .B(n2906), .Z(n2900) );
  AND U2516 ( .A(n684), .B(n2907), .Z(n2906) );
  XOR U2517 ( .A(p_input[951]), .B(n2905), .Z(n2907) );
  XOR U2518 ( .A(n2908), .B(n2909), .Z(n2905) );
  AND U2519 ( .A(n688), .B(n2910), .Z(n2909) );
  XOR U2520 ( .A(n2911), .B(n2912), .Z(n2903) );
  AND U2521 ( .A(n692), .B(n2910), .Z(n2912) );
  XNOR U2522 ( .A(n2911), .B(n2908), .Z(n2910) );
  XOR U2523 ( .A(n2913), .B(n2914), .Z(n2908) );
  AND U2524 ( .A(n695), .B(n2915), .Z(n2914) );
  XOR U2525 ( .A(p_input[967]), .B(n2913), .Z(n2915) );
  XOR U2526 ( .A(n2916), .B(n2917), .Z(n2913) );
  AND U2527 ( .A(n699), .B(n2918), .Z(n2917) );
  XOR U2528 ( .A(n2919), .B(n2920), .Z(n2911) );
  AND U2529 ( .A(n703), .B(n2918), .Z(n2920) );
  XNOR U2530 ( .A(n2919), .B(n2916), .Z(n2918) );
  XOR U2531 ( .A(n2921), .B(n2922), .Z(n2916) );
  AND U2532 ( .A(n706), .B(n2923), .Z(n2922) );
  XOR U2533 ( .A(p_input[983]), .B(n2921), .Z(n2923) );
  XOR U2534 ( .A(n2924), .B(n2925), .Z(n2921) );
  AND U2535 ( .A(n710), .B(n2926), .Z(n2925) );
  XOR U2536 ( .A(n2927), .B(n2928), .Z(n2919) );
  AND U2537 ( .A(n714), .B(n2926), .Z(n2928) );
  XNOR U2538 ( .A(n2927), .B(n2924), .Z(n2926) );
  XOR U2539 ( .A(n2929), .B(n2930), .Z(n2924) );
  AND U2540 ( .A(n717), .B(n2931), .Z(n2930) );
  XOR U2541 ( .A(p_input[999]), .B(n2929), .Z(n2931) );
  XOR U2542 ( .A(n2932), .B(n2933), .Z(n2929) );
  AND U2543 ( .A(n721), .B(n2934), .Z(n2933) );
  XOR U2544 ( .A(n2935), .B(n2936), .Z(n2927) );
  AND U2545 ( .A(n725), .B(n2934), .Z(n2936) );
  XNOR U2546 ( .A(n2935), .B(n2932), .Z(n2934) );
  XOR U2547 ( .A(n2937), .B(n2938), .Z(n2932) );
  AND U2548 ( .A(n728), .B(n2939), .Z(n2938) );
  XOR U2549 ( .A(p_input[1015]), .B(n2937), .Z(n2939) );
  XOR U2550 ( .A(n2940), .B(n2941), .Z(n2937) );
  AND U2551 ( .A(n732), .B(n2942), .Z(n2941) );
  XOR U2552 ( .A(n2943), .B(n2944), .Z(n2935) );
  AND U2553 ( .A(n736), .B(n2942), .Z(n2944) );
  XNOR U2554 ( .A(n2943), .B(n2940), .Z(n2942) );
  XOR U2555 ( .A(n2945), .B(n2946), .Z(n2940) );
  AND U2556 ( .A(n739), .B(n2947), .Z(n2946) );
  XOR U2557 ( .A(p_input[1031]), .B(n2945), .Z(n2947) );
  XOR U2558 ( .A(n2948), .B(n2949), .Z(n2945) );
  AND U2559 ( .A(n743), .B(n2950), .Z(n2949) );
  XOR U2560 ( .A(n2951), .B(n2952), .Z(n2943) );
  AND U2561 ( .A(n747), .B(n2950), .Z(n2952) );
  XNOR U2562 ( .A(n2951), .B(n2948), .Z(n2950) );
  XOR U2563 ( .A(n2953), .B(n2954), .Z(n2948) );
  AND U2564 ( .A(n750), .B(n2955), .Z(n2954) );
  XOR U2565 ( .A(p_input[1047]), .B(n2953), .Z(n2955) );
  XOR U2566 ( .A(n2956), .B(n2957), .Z(n2953) );
  AND U2567 ( .A(n754), .B(n2958), .Z(n2957) );
  XOR U2568 ( .A(n2959), .B(n2960), .Z(n2951) );
  AND U2569 ( .A(n758), .B(n2958), .Z(n2960) );
  XNOR U2570 ( .A(n2959), .B(n2956), .Z(n2958) );
  XOR U2571 ( .A(n2961), .B(n2962), .Z(n2956) );
  AND U2572 ( .A(n761), .B(n2963), .Z(n2962) );
  XOR U2573 ( .A(p_input[1063]), .B(n2961), .Z(n2963) );
  XOR U2574 ( .A(n2964), .B(n2965), .Z(n2961) );
  AND U2575 ( .A(n765), .B(n2966), .Z(n2965) );
  XOR U2576 ( .A(n2967), .B(n2968), .Z(n2959) );
  AND U2577 ( .A(n769), .B(n2966), .Z(n2968) );
  XNOR U2578 ( .A(n2967), .B(n2964), .Z(n2966) );
  XOR U2579 ( .A(n2969), .B(n2970), .Z(n2964) );
  AND U2580 ( .A(n772), .B(n2971), .Z(n2970) );
  XOR U2581 ( .A(p_input[1079]), .B(n2969), .Z(n2971) );
  XOR U2582 ( .A(n2972), .B(n2973), .Z(n2969) );
  AND U2583 ( .A(n776), .B(n2974), .Z(n2973) );
  XOR U2584 ( .A(n2975), .B(n2976), .Z(n2967) );
  AND U2585 ( .A(n780), .B(n2974), .Z(n2976) );
  XNOR U2586 ( .A(n2975), .B(n2972), .Z(n2974) );
  XOR U2587 ( .A(n2977), .B(n2978), .Z(n2972) );
  AND U2588 ( .A(n783), .B(n2979), .Z(n2978) );
  XOR U2589 ( .A(p_input[1095]), .B(n2977), .Z(n2979) );
  XOR U2590 ( .A(n2980), .B(n2981), .Z(n2977) );
  AND U2591 ( .A(n787), .B(n2982), .Z(n2981) );
  XOR U2592 ( .A(n2983), .B(n2984), .Z(n2975) );
  AND U2593 ( .A(n791), .B(n2982), .Z(n2984) );
  XNOR U2594 ( .A(n2983), .B(n2980), .Z(n2982) );
  XOR U2595 ( .A(n2985), .B(n2986), .Z(n2980) );
  AND U2596 ( .A(n794), .B(n2987), .Z(n2986) );
  XOR U2597 ( .A(p_input[1111]), .B(n2985), .Z(n2987) );
  XOR U2598 ( .A(n2988), .B(n2989), .Z(n2985) );
  AND U2599 ( .A(n798), .B(n2990), .Z(n2989) );
  XOR U2600 ( .A(n2991), .B(n2992), .Z(n2983) );
  AND U2601 ( .A(n802), .B(n2990), .Z(n2992) );
  XNOR U2602 ( .A(n2991), .B(n2988), .Z(n2990) );
  XOR U2603 ( .A(n2993), .B(n2994), .Z(n2988) );
  AND U2604 ( .A(n805), .B(n2995), .Z(n2994) );
  XOR U2605 ( .A(p_input[1127]), .B(n2993), .Z(n2995) );
  XOR U2606 ( .A(n2996), .B(n2997), .Z(n2993) );
  AND U2607 ( .A(n809), .B(n2998), .Z(n2997) );
  XOR U2608 ( .A(n2999), .B(n3000), .Z(n2991) );
  AND U2609 ( .A(n813), .B(n2998), .Z(n3000) );
  XNOR U2610 ( .A(n2999), .B(n2996), .Z(n2998) );
  XOR U2611 ( .A(n3001), .B(n3002), .Z(n2996) );
  AND U2612 ( .A(n816), .B(n3003), .Z(n3002) );
  XOR U2613 ( .A(p_input[1143]), .B(n3001), .Z(n3003) );
  XOR U2614 ( .A(n3004), .B(n3005), .Z(n3001) );
  AND U2615 ( .A(n820), .B(n3006), .Z(n3005) );
  XOR U2616 ( .A(n3007), .B(n3008), .Z(n2999) );
  AND U2617 ( .A(n824), .B(n3006), .Z(n3008) );
  XNOR U2618 ( .A(n3007), .B(n3004), .Z(n3006) );
  XOR U2619 ( .A(n3009), .B(n3010), .Z(n3004) );
  AND U2620 ( .A(n827), .B(n3011), .Z(n3010) );
  XOR U2621 ( .A(p_input[1159]), .B(n3009), .Z(n3011) );
  XOR U2622 ( .A(n3012), .B(n3013), .Z(n3009) );
  AND U2623 ( .A(n831), .B(n3014), .Z(n3013) );
  XOR U2624 ( .A(n3015), .B(n3016), .Z(n3007) );
  AND U2625 ( .A(n835), .B(n3014), .Z(n3016) );
  XNOR U2626 ( .A(n3015), .B(n3012), .Z(n3014) );
  XOR U2627 ( .A(n3017), .B(n3018), .Z(n3012) );
  AND U2628 ( .A(n838), .B(n3019), .Z(n3018) );
  XOR U2629 ( .A(p_input[1175]), .B(n3017), .Z(n3019) );
  XOR U2630 ( .A(n3020), .B(n3021), .Z(n3017) );
  AND U2631 ( .A(n842), .B(n3022), .Z(n3021) );
  XOR U2632 ( .A(n3023), .B(n3024), .Z(n3015) );
  AND U2633 ( .A(n846), .B(n3022), .Z(n3024) );
  XNOR U2634 ( .A(n3023), .B(n3020), .Z(n3022) );
  XOR U2635 ( .A(n3025), .B(n3026), .Z(n3020) );
  AND U2636 ( .A(n849), .B(n3027), .Z(n3026) );
  XOR U2637 ( .A(p_input[1191]), .B(n3025), .Z(n3027) );
  XOR U2638 ( .A(n3028), .B(n3029), .Z(n3025) );
  AND U2639 ( .A(n853), .B(n3030), .Z(n3029) );
  XOR U2640 ( .A(n3031), .B(n3032), .Z(n3023) );
  AND U2641 ( .A(n857), .B(n3030), .Z(n3032) );
  XNOR U2642 ( .A(n3031), .B(n3028), .Z(n3030) );
  XOR U2643 ( .A(n3033), .B(n3034), .Z(n3028) );
  AND U2644 ( .A(n860), .B(n3035), .Z(n3034) );
  XOR U2645 ( .A(p_input[1207]), .B(n3033), .Z(n3035) );
  XOR U2646 ( .A(n3036), .B(n3037), .Z(n3033) );
  AND U2647 ( .A(n864), .B(n3038), .Z(n3037) );
  XOR U2648 ( .A(n3039), .B(n3040), .Z(n3031) );
  AND U2649 ( .A(n868), .B(n3038), .Z(n3040) );
  XNOR U2650 ( .A(n3039), .B(n3036), .Z(n3038) );
  XOR U2651 ( .A(n3041), .B(n3042), .Z(n3036) );
  AND U2652 ( .A(n871), .B(n3043), .Z(n3042) );
  XOR U2653 ( .A(p_input[1223]), .B(n3041), .Z(n3043) );
  XOR U2654 ( .A(n3044), .B(n3045), .Z(n3041) );
  AND U2655 ( .A(n875), .B(n3046), .Z(n3045) );
  XOR U2656 ( .A(n3047), .B(n3048), .Z(n3039) );
  AND U2657 ( .A(n879), .B(n3046), .Z(n3048) );
  XNOR U2658 ( .A(n3047), .B(n3044), .Z(n3046) );
  XOR U2659 ( .A(n3049), .B(n3050), .Z(n3044) );
  AND U2660 ( .A(n882), .B(n3051), .Z(n3050) );
  XOR U2661 ( .A(p_input[1239]), .B(n3049), .Z(n3051) );
  XOR U2662 ( .A(n3052), .B(n3053), .Z(n3049) );
  AND U2663 ( .A(n886), .B(n3054), .Z(n3053) );
  XOR U2664 ( .A(n3055), .B(n3056), .Z(n3047) );
  AND U2665 ( .A(n890), .B(n3054), .Z(n3056) );
  XNOR U2666 ( .A(n3055), .B(n3052), .Z(n3054) );
  XOR U2667 ( .A(n3057), .B(n3058), .Z(n3052) );
  AND U2668 ( .A(n893), .B(n3059), .Z(n3058) );
  XOR U2669 ( .A(p_input[1255]), .B(n3057), .Z(n3059) );
  XOR U2670 ( .A(n3060), .B(n3061), .Z(n3057) );
  AND U2671 ( .A(n897), .B(n3062), .Z(n3061) );
  XOR U2672 ( .A(n3063), .B(n3064), .Z(n3055) );
  AND U2673 ( .A(n901), .B(n3062), .Z(n3064) );
  XNOR U2674 ( .A(n3063), .B(n3060), .Z(n3062) );
  XOR U2675 ( .A(n3065), .B(n3066), .Z(n3060) );
  AND U2676 ( .A(n904), .B(n3067), .Z(n3066) );
  XOR U2677 ( .A(p_input[1271]), .B(n3065), .Z(n3067) );
  XOR U2678 ( .A(n3068), .B(n3069), .Z(n3065) );
  AND U2679 ( .A(n908), .B(n3070), .Z(n3069) );
  XOR U2680 ( .A(n3071), .B(n3072), .Z(n3063) );
  AND U2681 ( .A(n912), .B(n3070), .Z(n3072) );
  XNOR U2682 ( .A(n3071), .B(n3068), .Z(n3070) );
  XOR U2683 ( .A(n3073), .B(n3074), .Z(n3068) );
  AND U2684 ( .A(n915), .B(n3075), .Z(n3074) );
  XOR U2685 ( .A(p_input[1287]), .B(n3073), .Z(n3075) );
  XOR U2686 ( .A(n3076), .B(n3077), .Z(n3073) );
  AND U2687 ( .A(n919), .B(n3078), .Z(n3077) );
  XOR U2688 ( .A(n3079), .B(n3080), .Z(n3071) );
  AND U2689 ( .A(n923), .B(n3078), .Z(n3080) );
  XNOR U2690 ( .A(n3079), .B(n3076), .Z(n3078) );
  XOR U2691 ( .A(n3081), .B(n3082), .Z(n3076) );
  AND U2692 ( .A(n926), .B(n3083), .Z(n3082) );
  XOR U2693 ( .A(p_input[1303]), .B(n3081), .Z(n3083) );
  XOR U2694 ( .A(n3084), .B(n3085), .Z(n3081) );
  AND U2695 ( .A(n930), .B(n3086), .Z(n3085) );
  XOR U2696 ( .A(n3087), .B(n3088), .Z(n3079) );
  AND U2697 ( .A(n934), .B(n3086), .Z(n3088) );
  XNOR U2698 ( .A(n3087), .B(n3084), .Z(n3086) );
  XOR U2699 ( .A(n3089), .B(n3090), .Z(n3084) );
  AND U2700 ( .A(n937), .B(n3091), .Z(n3090) );
  XOR U2701 ( .A(p_input[1319]), .B(n3089), .Z(n3091) );
  XOR U2702 ( .A(n3092), .B(n3093), .Z(n3089) );
  AND U2703 ( .A(n941), .B(n3094), .Z(n3093) );
  XOR U2704 ( .A(n3095), .B(n3096), .Z(n3087) );
  AND U2705 ( .A(n945), .B(n3094), .Z(n3096) );
  XNOR U2706 ( .A(n3095), .B(n3092), .Z(n3094) );
  XOR U2707 ( .A(n3097), .B(n3098), .Z(n3092) );
  AND U2708 ( .A(n948), .B(n3099), .Z(n3098) );
  XOR U2709 ( .A(p_input[1335]), .B(n3097), .Z(n3099) );
  XOR U2710 ( .A(n3100), .B(n3101), .Z(n3097) );
  AND U2711 ( .A(n952), .B(n3102), .Z(n3101) );
  XOR U2712 ( .A(n3103), .B(n3104), .Z(n3095) );
  AND U2713 ( .A(n956), .B(n3102), .Z(n3104) );
  XNOR U2714 ( .A(n3103), .B(n3100), .Z(n3102) );
  XOR U2715 ( .A(n3105), .B(n3106), .Z(n3100) );
  AND U2716 ( .A(n959), .B(n3107), .Z(n3106) );
  XOR U2717 ( .A(p_input[1351]), .B(n3105), .Z(n3107) );
  XOR U2718 ( .A(n3108), .B(n3109), .Z(n3105) );
  AND U2719 ( .A(n963), .B(n3110), .Z(n3109) );
  XOR U2720 ( .A(n3111), .B(n3112), .Z(n3103) );
  AND U2721 ( .A(n967), .B(n3110), .Z(n3112) );
  XNOR U2722 ( .A(n3111), .B(n3108), .Z(n3110) );
  XOR U2723 ( .A(n3113), .B(n3114), .Z(n3108) );
  AND U2724 ( .A(n970), .B(n3115), .Z(n3114) );
  XOR U2725 ( .A(p_input[1367]), .B(n3113), .Z(n3115) );
  XOR U2726 ( .A(n3116), .B(n3117), .Z(n3113) );
  AND U2727 ( .A(n974), .B(n3118), .Z(n3117) );
  XOR U2728 ( .A(n3119), .B(n3120), .Z(n3111) );
  AND U2729 ( .A(n978), .B(n3118), .Z(n3120) );
  XNOR U2730 ( .A(n3119), .B(n3116), .Z(n3118) );
  XOR U2731 ( .A(n3121), .B(n3122), .Z(n3116) );
  AND U2732 ( .A(n981), .B(n3123), .Z(n3122) );
  XOR U2733 ( .A(p_input[1383]), .B(n3121), .Z(n3123) );
  XOR U2734 ( .A(n3124), .B(n3125), .Z(n3121) );
  AND U2735 ( .A(n985), .B(n3126), .Z(n3125) );
  XOR U2736 ( .A(n3127), .B(n3128), .Z(n3119) );
  AND U2737 ( .A(n989), .B(n3126), .Z(n3128) );
  XNOR U2738 ( .A(n3127), .B(n3124), .Z(n3126) );
  XOR U2739 ( .A(n3129), .B(n3130), .Z(n3124) );
  AND U2740 ( .A(n992), .B(n3131), .Z(n3130) );
  XOR U2741 ( .A(p_input[1399]), .B(n3129), .Z(n3131) );
  XOR U2742 ( .A(n3132), .B(n3133), .Z(n3129) );
  AND U2743 ( .A(n996), .B(n3134), .Z(n3133) );
  XOR U2744 ( .A(n3135), .B(n3136), .Z(n3127) );
  AND U2745 ( .A(n1000), .B(n3134), .Z(n3136) );
  XNOR U2746 ( .A(n3135), .B(n3132), .Z(n3134) );
  XOR U2747 ( .A(n3137), .B(n3138), .Z(n3132) );
  AND U2748 ( .A(n1003), .B(n3139), .Z(n3138) );
  XOR U2749 ( .A(p_input[1415]), .B(n3137), .Z(n3139) );
  XOR U2750 ( .A(n3140), .B(n3141), .Z(n3137) );
  AND U2751 ( .A(n1007), .B(n3142), .Z(n3141) );
  XOR U2752 ( .A(n3143), .B(n3144), .Z(n3135) );
  AND U2753 ( .A(n1011), .B(n3142), .Z(n3144) );
  XNOR U2754 ( .A(n3143), .B(n3140), .Z(n3142) );
  XOR U2755 ( .A(n3145), .B(n3146), .Z(n3140) );
  AND U2756 ( .A(n1014), .B(n3147), .Z(n3146) );
  XOR U2757 ( .A(p_input[1431]), .B(n3145), .Z(n3147) );
  XOR U2758 ( .A(n3148), .B(n3149), .Z(n3145) );
  AND U2759 ( .A(n1018), .B(n3150), .Z(n3149) );
  XOR U2760 ( .A(n3151), .B(n3152), .Z(n3143) );
  AND U2761 ( .A(n1022), .B(n3150), .Z(n3152) );
  XNOR U2762 ( .A(n3151), .B(n3148), .Z(n3150) );
  XOR U2763 ( .A(n3153), .B(n3154), .Z(n3148) );
  AND U2764 ( .A(n1025), .B(n3155), .Z(n3154) );
  XOR U2765 ( .A(p_input[1447]), .B(n3153), .Z(n3155) );
  XOR U2766 ( .A(n3156), .B(n3157), .Z(n3153) );
  AND U2767 ( .A(n1029), .B(n3158), .Z(n3157) );
  XOR U2768 ( .A(n3159), .B(n3160), .Z(n3151) );
  AND U2769 ( .A(n1033), .B(n3158), .Z(n3160) );
  XNOR U2770 ( .A(n3159), .B(n3156), .Z(n3158) );
  XOR U2771 ( .A(n3161), .B(n3162), .Z(n3156) );
  AND U2772 ( .A(n1036), .B(n3163), .Z(n3162) );
  XOR U2773 ( .A(p_input[1463]), .B(n3161), .Z(n3163) );
  XOR U2774 ( .A(n3164), .B(n3165), .Z(n3161) );
  AND U2775 ( .A(n1040), .B(n3166), .Z(n3165) );
  XOR U2776 ( .A(n3167), .B(n3168), .Z(n3159) );
  AND U2777 ( .A(n1044), .B(n3166), .Z(n3168) );
  XNOR U2778 ( .A(n3167), .B(n3164), .Z(n3166) );
  XOR U2779 ( .A(n3169), .B(n3170), .Z(n3164) );
  AND U2780 ( .A(n1047), .B(n3171), .Z(n3170) );
  XOR U2781 ( .A(p_input[1479]), .B(n3169), .Z(n3171) );
  XOR U2782 ( .A(n3172), .B(n3173), .Z(n3169) );
  AND U2783 ( .A(n1051), .B(n3174), .Z(n3173) );
  XOR U2784 ( .A(n3175), .B(n3176), .Z(n3167) );
  AND U2785 ( .A(n1055), .B(n3174), .Z(n3176) );
  XNOR U2786 ( .A(n3175), .B(n3172), .Z(n3174) );
  XOR U2787 ( .A(n3177), .B(n3178), .Z(n3172) );
  AND U2788 ( .A(n1058), .B(n3179), .Z(n3178) );
  XOR U2789 ( .A(p_input[1495]), .B(n3177), .Z(n3179) );
  XOR U2790 ( .A(n3180), .B(n3181), .Z(n3177) );
  AND U2791 ( .A(n1062), .B(n3182), .Z(n3181) );
  XOR U2792 ( .A(n3183), .B(n3184), .Z(n3175) );
  AND U2793 ( .A(n1066), .B(n3182), .Z(n3184) );
  XNOR U2794 ( .A(n3183), .B(n3180), .Z(n3182) );
  XOR U2795 ( .A(n3185), .B(n3186), .Z(n3180) );
  AND U2796 ( .A(n1069), .B(n3187), .Z(n3186) );
  XOR U2797 ( .A(p_input[1511]), .B(n3185), .Z(n3187) );
  XOR U2798 ( .A(n3188), .B(n3189), .Z(n3185) );
  AND U2799 ( .A(n1073), .B(n3190), .Z(n3189) );
  XOR U2800 ( .A(n3191), .B(n3192), .Z(n3183) );
  AND U2801 ( .A(n1077), .B(n3190), .Z(n3192) );
  XNOR U2802 ( .A(n3191), .B(n3188), .Z(n3190) );
  XOR U2803 ( .A(n3193), .B(n3194), .Z(n3188) );
  AND U2804 ( .A(n1080), .B(n3195), .Z(n3194) );
  XOR U2805 ( .A(p_input[1527]), .B(n3193), .Z(n3195) );
  XOR U2806 ( .A(n3196), .B(n3197), .Z(n3193) );
  AND U2807 ( .A(n1084), .B(n3198), .Z(n3197) );
  XOR U2808 ( .A(n3199), .B(n3200), .Z(n3191) );
  AND U2809 ( .A(n1088), .B(n3198), .Z(n3200) );
  XNOR U2810 ( .A(n3199), .B(n3196), .Z(n3198) );
  XOR U2811 ( .A(n3201), .B(n3202), .Z(n3196) );
  AND U2812 ( .A(n1091), .B(n3203), .Z(n3202) );
  XOR U2813 ( .A(p_input[1543]), .B(n3201), .Z(n3203) );
  XOR U2814 ( .A(n3204), .B(n3205), .Z(n3201) );
  AND U2815 ( .A(n1095), .B(n3206), .Z(n3205) );
  XOR U2816 ( .A(n3207), .B(n3208), .Z(n3199) );
  AND U2817 ( .A(n1099), .B(n3206), .Z(n3208) );
  XNOR U2818 ( .A(n3207), .B(n3204), .Z(n3206) );
  XOR U2819 ( .A(n3209), .B(n3210), .Z(n3204) );
  AND U2820 ( .A(n1102), .B(n3211), .Z(n3210) );
  XOR U2821 ( .A(p_input[1559]), .B(n3209), .Z(n3211) );
  XOR U2822 ( .A(n3212), .B(n3213), .Z(n3209) );
  AND U2823 ( .A(n1106), .B(n3214), .Z(n3213) );
  XOR U2824 ( .A(n3215), .B(n3216), .Z(n3207) );
  AND U2825 ( .A(n1110), .B(n3214), .Z(n3216) );
  XNOR U2826 ( .A(n3215), .B(n3212), .Z(n3214) );
  XOR U2827 ( .A(n3217), .B(n3218), .Z(n3212) );
  AND U2828 ( .A(n1113), .B(n3219), .Z(n3218) );
  XOR U2829 ( .A(p_input[1575]), .B(n3217), .Z(n3219) );
  XOR U2830 ( .A(n3220), .B(n3221), .Z(n3217) );
  AND U2831 ( .A(n1117), .B(n3222), .Z(n3221) );
  XOR U2832 ( .A(n3223), .B(n3224), .Z(n3215) );
  AND U2833 ( .A(n1121), .B(n3222), .Z(n3224) );
  XNOR U2834 ( .A(n3223), .B(n3220), .Z(n3222) );
  XOR U2835 ( .A(n3225), .B(n3226), .Z(n3220) );
  AND U2836 ( .A(n1124), .B(n3227), .Z(n3226) );
  XOR U2837 ( .A(p_input[1591]), .B(n3225), .Z(n3227) );
  XOR U2838 ( .A(n3228), .B(n3229), .Z(n3225) );
  AND U2839 ( .A(n1128), .B(n3230), .Z(n3229) );
  XOR U2840 ( .A(n3231), .B(n3232), .Z(n3223) );
  AND U2841 ( .A(n1132), .B(n3230), .Z(n3232) );
  XNOR U2842 ( .A(n3231), .B(n3228), .Z(n3230) );
  XOR U2843 ( .A(n3233), .B(n3234), .Z(n3228) );
  AND U2844 ( .A(n1135), .B(n3235), .Z(n3234) );
  XOR U2845 ( .A(p_input[1607]), .B(n3233), .Z(n3235) );
  XOR U2846 ( .A(n3236), .B(n3237), .Z(n3233) );
  AND U2847 ( .A(n1139), .B(n3238), .Z(n3237) );
  XOR U2848 ( .A(n3239), .B(n3240), .Z(n3231) );
  AND U2849 ( .A(n1143), .B(n3238), .Z(n3240) );
  XNOR U2850 ( .A(n3239), .B(n3236), .Z(n3238) );
  XOR U2851 ( .A(n3241), .B(n3242), .Z(n3236) );
  AND U2852 ( .A(n1146), .B(n3243), .Z(n3242) );
  XOR U2853 ( .A(p_input[1623]), .B(n3241), .Z(n3243) );
  XOR U2854 ( .A(n3244), .B(n3245), .Z(n3241) );
  AND U2855 ( .A(n1150), .B(n3246), .Z(n3245) );
  XOR U2856 ( .A(n3247), .B(n3248), .Z(n3239) );
  AND U2857 ( .A(n1154), .B(n3246), .Z(n3248) );
  XNOR U2858 ( .A(n3247), .B(n3244), .Z(n3246) );
  XOR U2859 ( .A(n3249), .B(n3250), .Z(n3244) );
  AND U2860 ( .A(n1157), .B(n3251), .Z(n3250) );
  XOR U2861 ( .A(p_input[1639]), .B(n3249), .Z(n3251) );
  XOR U2862 ( .A(n3252), .B(n3253), .Z(n3249) );
  AND U2863 ( .A(n1161), .B(n3254), .Z(n3253) );
  XOR U2864 ( .A(n3255), .B(n3256), .Z(n3247) );
  AND U2865 ( .A(n1165), .B(n3254), .Z(n3256) );
  XNOR U2866 ( .A(n3255), .B(n3252), .Z(n3254) );
  XOR U2867 ( .A(n3257), .B(n3258), .Z(n3252) );
  AND U2868 ( .A(n1168), .B(n3259), .Z(n3258) );
  XOR U2869 ( .A(p_input[1655]), .B(n3257), .Z(n3259) );
  XOR U2870 ( .A(n3260), .B(n3261), .Z(n3257) );
  AND U2871 ( .A(n1172), .B(n3262), .Z(n3261) );
  XOR U2872 ( .A(n3263), .B(n3264), .Z(n3255) );
  AND U2873 ( .A(n1176), .B(n3262), .Z(n3264) );
  XNOR U2874 ( .A(n3263), .B(n3260), .Z(n3262) );
  XOR U2875 ( .A(n3265), .B(n3266), .Z(n3260) );
  AND U2876 ( .A(n1179), .B(n3267), .Z(n3266) );
  XOR U2877 ( .A(p_input[1671]), .B(n3265), .Z(n3267) );
  XOR U2878 ( .A(n3268), .B(n3269), .Z(n3265) );
  AND U2879 ( .A(n1183), .B(n3270), .Z(n3269) );
  XOR U2880 ( .A(n3271), .B(n3272), .Z(n3263) );
  AND U2881 ( .A(n1187), .B(n3270), .Z(n3272) );
  XNOR U2882 ( .A(n3271), .B(n3268), .Z(n3270) );
  XOR U2883 ( .A(n3273), .B(n3274), .Z(n3268) );
  AND U2884 ( .A(n1190), .B(n3275), .Z(n3274) );
  XOR U2885 ( .A(p_input[1687]), .B(n3273), .Z(n3275) );
  XOR U2886 ( .A(n3276), .B(n3277), .Z(n3273) );
  AND U2887 ( .A(n1194), .B(n3278), .Z(n3277) );
  XOR U2888 ( .A(n3279), .B(n3280), .Z(n3271) );
  AND U2889 ( .A(n1198), .B(n3278), .Z(n3280) );
  XNOR U2890 ( .A(n3279), .B(n3276), .Z(n3278) );
  XOR U2891 ( .A(n3281), .B(n3282), .Z(n3276) );
  AND U2892 ( .A(n1201), .B(n3283), .Z(n3282) );
  XOR U2893 ( .A(p_input[1703]), .B(n3281), .Z(n3283) );
  XOR U2894 ( .A(n3284), .B(n3285), .Z(n3281) );
  AND U2895 ( .A(n1205), .B(n3286), .Z(n3285) );
  XOR U2896 ( .A(n3287), .B(n3288), .Z(n3279) );
  AND U2897 ( .A(n1209), .B(n3286), .Z(n3288) );
  XNOR U2898 ( .A(n3287), .B(n3284), .Z(n3286) );
  XOR U2899 ( .A(n3289), .B(n3290), .Z(n3284) );
  AND U2900 ( .A(n1212), .B(n3291), .Z(n3290) );
  XOR U2901 ( .A(p_input[1719]), .B(n3289), .Z(n3291) );
  XOR U2902 ( .A(n3292), .B(n3293), .Z(n3289) );
  AND U2903 ( .A(n1216), .B(n3294), .Z(n3293) );
  XOR U2904 ( .A(n3295), .B(n3296), .Z(n3287) );
  AND U2905 ( .A(n1220), .B(n3294), .Z(n3296) );
  XNOR U2906 ( .A(n3295), .B(n3292), .Z(n3294) );
  XOR U2907 ( .A(n3297), .B(n3298), .Z(n3292) );
  AND U2908 ( .A(n1223), .B(n3299), .Z(n3298) );
  XOR U2909 ( .A(p_input[1735]), .B(n3297), .Z(n3299) );
  XOR U2910 ( .A(n3300), .B(n3301), .Z(n3297) );
  AND U2911 ( .A(n1227), .B(n3302), .Z(n3301) );
  XOR U2912 ( .A(n3303), .B(n3304), .Z(n3295) );
  AND U2913 ( .A(n1231), .B(n3302), .Z(n3304) );
  XNOR U2914 ( .A(n3303), .B(n3300), .Z(n3302) );
  XOR U2915 ( .A(n3305), .B(n3306), .Z(n3300) );
  AND U2916 ( .A(n1234), .B(n3307), .Z(n3306) );
  XOR U2917 ( .A(p_input[1751]), .B(n3305), .Z(n3307) );
  XOR U2918 ( .A(n3308), .B(n3309), .Z(n3305) );
  AND U2919 ( .A(n1238), .B(n3310), .Z(n3309) );
  XOR U2920 ( .A(n3311), .B(n3312), .Z(n3303) );
  AND U2921 ( .A(n1242), .B(n3310), .Z(n3312) );
  XNOR U2922 ( .A(n3311), .B(n3308), .Z(n3310) );
  XOR U2923 ( .A(n3313), .B(n3314), .Z(n3308) );
  AND U2924 ( .A(n1245), .B(n3315), .Z(n3314) );
  XOR U2925 ( .A(p_input[1767]), .B(n3313), .Z(n3315) );
  XOR U2926 ( .A(n3316), .B(n3317), .Z(n3313) );
  AND U2927 ( .A(n1249), .B(n3318), .Z(n3317) );
  XOR U2928 ( .A(n3319), .B(n3320), .Z(n3311) );
  AND U2929 ( .A(n1253), .B(n3318), .Z(n3320) );
  XNOR U2930 ( .A(n3319), .B(n3316), .Z(n3318) );
  XOR U2931 ( .A(n3321), .B(n3322), .Z(n3316) );
  AND U2932 ( .A(n1256), .B(n3323), .Z(n3322) );
  XOR U2933 ( .A(p_input[1783]), .B(n3321), .Z(n3323) );
  XOR U2934 ( .A(n3324), .B(n3325), .Z(n3321) );
  AND U2935 ( .A(n1260), .B(n3326), .Z(n3325) );
  XOR U2936 ( .A(n3327), .B(n3328), .Z(n3319) );
  AND U2937 ( .A(n1264), .B(n3326), .Z(n3328) );
  XNOR U2938 ( .A(n3327), .B(n3324), .Z(n3326) );
  XOR U2939 ( .A(n3329), .B(n3330), .Z(n3324) );
  AND U2940 ( .A(n1267), .B(n3331), .Z(n3330) );
  XOR U2941 ( .A(p_input[1799]), .B(n3329), .Z(n3331) );
  XOR U2942 ( .A(n3332), .B(n3333), .Z(n3329) );
  AND U2943 ( .A(n1271), .B(n3334), .Z(n3333) );
  XOR U2944 ( .A(n3335), .B(n3336), .Z(n3327) );
  AND U2945 ( .A(n1275), .B(n3334), .Z(n3336) );
  XNOR U2946 ( .A(n3335), .B(n3332), .Z(n3334) );
  XOR U2947 ( .A(n3337), .B(n3338), .Z(n3332) );
  AND U2948 ( .A(n1278), .B(n3339), .Z(n3338) );
  XOR U2949 ( .A(p_input[1815]), .B(n3337), .Z(n3339) );
  XOR U2950 ( .A(n3340), .B(n3341), .Z(n3337) );
  AND U2951 ( .A(n1282), .B(n3342), .Z(n3341) );
  XOR U2952 ( .A(n3343), .B(n3344), .Z(n3335) );
  AND U2953 ( .A(n1286), .B(n3342), .Z(n3344) );
  XNOR U2954 ( .A(n3343), .B(n3340), .Z(n3342) );
  XOR U2955 ( .A(n3345), .B(n3346), .Z(n3340) );
  AND U2956 ( .A(n1289), .B(n3347), .Z(n3346) );
  XOR U2957 ( .A(p_input[1831]), .B(n3345), .Z(n3347) );
  XOR U2958 ( .A(n3348), .B(n3349), .Z(n3345) );
  AND U2959 ( .A(n1293), .B(n3350), .Z(n3349) );
  XOR U2960 ( .A(n3351), .B(n3352), .Z(n3343) );
  AND U2961 ( .A(n1297), .B(n3350), .Z(n3352) );
  XNOR U2962 ( .A(n3351), .B(n3348), .Z(n3350) );
  XOR U2963 ( .A(n3353), .B(n3354), .Z(n3348) );
  AND U2964 ( .A(n1300), .B(n3355), .Z(n3354) );
  XOR U2965 ( .A(p_input[1847]), .B(n3353), .Z(n3355) );
  XOR U2966 ( .A(n3356), .B(n3357), .Z(n3353) );
  AND U2967 ( .A(n1304), .B(n3358), .Z(n3357) );
  XOR U2968 ( .A(n3359), .B(n3360), .Z(n3351) );
  AND U2969 ( .A(n1308), .B(n3358), .Z(n3360) );
  XNOR U2970 ( .A(n3359), .B(n3356), .Z(n3358) );
  XOR U2971 ( .A(n3361), .B(n3362), .Z(n3356) );
  AND U2972 ( .A(n1311), .B(n3363), .Z(n3362) );
  XOR U2973 ( .A(p_input[1863]), .B(n3361), .Z(n3363) );
  XOR U2974 ( .A(n3364), .B(n3365), .Z(n3361) );
  AND U2975 ( .A(n1315), .B(n3366), .Z(n3365) );
  XOR U2976 ( .A(n3367), .B(n3368), .Z(n3359) );
  AND U2977 ( .A(n1319), .B(n3366), .Z(n3368) );
  XNOR U2978 ( .A(n3367), .B(n3364), .Z(n3366) );
  XOR U2979 ( .A(n3369), .B(n3370), .Z(n3364) );
  AND U2980 ( .A(n1322), .B(n3371), .Z(n3370) );
  XOR U2981 ( .A(p_input[1879]), .B(n3369), .Z(n3371) );
  XOR U2982 ( .A(n3372), .B(n3373), .Z(n3369) );
  AND U2983 ( .A(n1326), .B(n3374), .Z(n3373) );
  XOR U2984 ( .A(n3375), .B(n3376), .Z(n3367) );
  AND U2985 ( .A(n1330), .B(n3374), .Z(n3376) );
  XNOR U2986 ( .A(n3375), .B(n3372), .Z(n3374) );
  XOR U2987 ( .A(n3377), .B(n3378), .Z(n3372) );
  AND U2988 ( .A(n1333), .B(n3379), .Z(n3378) );
  XOR U2989 ( .A(p_input[1895]), .B(n3377), .Z(n3379) );
  XOR U2990 ( .A(n3380), .B(n3381), .Z(n3377) );
  AND U2991 ( .A(n1337), .B(n3382), .Z(n3381) );
  XOR U2992 ( .A(n3383), .B(n3384), .Z(n3375) );
  AND U2993 ( .A(n1341), .B(n3382), .Z(n3384) );
  XNOR U2994 ( .A(n3383), .B(n3380), .Z(n3382) );
  XOR U2995 ( .A(n3385), .B(n3386), .Z(n3380) );
  AND U2996 ( .A(n1344), .B(n3387), .Z(n3386) );
  XOR U2997 ( .A(p_input[1911]), .B(n3385), .Z(n3387) );
  XOR U2998 ( .A(n3388), .B(n3389), .Z(n3385) );
  AND U2999 ( .A(n1348), .B(n3390), .Z(n3389) );
  XOR U3000 ( .A(n3391), .B(n3392), .Z(n3383) );
  AND U3001 ( .A(n1352), .B(n3390), .Z(n3392) );
  XNOR U3002 ( .A(n3391), .B(n3388), .Z(n3390) );
  XOR U3003 ( .A(n3393), .B(n3394), .Z(n3388) );
  AND U3004 ( .A(n1355), .B(n3395), .Z(n3394) );
  XOR U3005 ( .A(p_input[1927]), .B(n3393), .Z(n3395) );
  XOR U3006 ( .A(n3396), .B(n3397), .Z(n3393) );
  AND U3007 ( .A(n1359), .B(n3398), .Z(n3397) );
  XOR U3008 ( .A(n3399), .B(n3400), .Z(n3391) );
  AND U3009 ( .A(n1363), .B(n3398), .Z(n3400) );
  XNOR U3010 ( .A(n3399), .B(n3396), .Z(n3398) );
  XOR U3011 ( .A(n3401), .B(n3402), .Z(n3396) );
  AND U3012 ( .A(n1366), .B(n3403), .Z(n3402) );
  XOR U3013 ( .A(p_input[1943]), .B(n3401), .Z(n3403) );
  XOR U3014 ( .A(n3404), .B(n3405), .Z(n3401) );
  AND U3015 ( .A(n1370), .B(n3406), .Z(n3405) );
  XOR U3016 ( .A(n3407), .B(n3408), .Z(n3399) );
  AND U3017 ( .A(n1374), .B(n3406), .Z(n3408) );
  XNOR U3018 ( .A(n3407), .B(n3404), .Z(n3406) );
  XOR U3019 ( .A(n3409), .B(n3410), .Z(n3404) );
  AND U3020 ( .A(n1377), .B(n3411), .Z(n3410) );
  XOR U3021 ( .A(p_input[1959]), .B(n3409), .Z(n3411) );
  XOR U3022 ( .A(n3412), .B(n3413), .Z(n3409) );
  AND U3023 ( .A(n1381), .B(n3414), .Z(n3413) );
  XOR U3024 ( .A(n3415), .B(n3416), .Z(n3407) );
  AND U3025 ( .A(n1385), .B(n3414), .Z(n3416) );
  XNOR U3026 ( .A(n3415), .B(n3412), .Z(n3414) );
  XOR U3027 ( .A(n3417), .B(n3418), .Z(n3412) );
  AND U3028 ( .A(n1388), .B(n3419), .Z(n3418) );
  XOR U3029 ( .A(p_input[1975]), .B(n3417), .Z(n3419) );
  XOR U3030 ( .A(n3420), .B(n3421), .Z(n3417) );
  AND U3031 ( .A(n1392), .B(n3422), .Z(n3421) );
  XOR U3032 ( .A(n3423), .B(n3424), .Z(n3415) );
  AND U3033 ( .A(n1396), .B(n3422), .Z(n3424) );
  XNOR U3034 ( .A(n3423), .B(n3420), .Z(n3422) );
  XOR U3035 ( .A(n3425), .B(n3426), .Z(n3420) );
  AND U3036 ( .A(n1399), .B(n3427), .Z(n3426) );
  XOR U3037 ( .A(p_input[1991]), .B(n3425), .Z(n3427) );
  XOR U3038 ( .A(n3428), .B(n3429), .Z(n3425) );
  AND U3039 ( .A(n1403), .B(n3430), .Z(n3429) );
  XOR U3040 ( .A(n3431), .B(n3432), .Z(n3423) );
  AND U3041 ( .A(n1407), .B(n3430), .Z(n3432) );
  XNOR U3042 ( .A(n3431), .B(n3428), .Z(n3430) );
  XOR U3043 ( .A(n3433), .B(n3434), .Z(n3428) );
  AND U3044 ( .A(n1410), .B(n3435), .Z(n3434) );
  XOR U3045 ( .A(p_input[2007]), .B(n3433), .Z(n3435) );
  XNOR U3046 ( .A(n3436), .B(n3437), .Z(n3433) );
  AND U3047 ( .A(n1414), .B(n3438), .Z(n3437) );
  XNOR U3048 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n3439), .Z(n3431) );
  AND U3049 ( .A(n1417), .B(n3438), .Z(n3439) );
  XOR U3050 ( .A(n3440), .B(n3436), .Z(n3438) );
  IV U3051 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .Z(n3436) );
  IV U3052 ( .A(\knn_comb_/min_val_out[0][7] ), .Z(n3440) );
  XOR U3053 ( .A(n7), .B(n3441), .Z(o[22]) );
  AND U3054 ( .A(n30), .B(n3442), .Z(n7) );
  XOR U3055 ( .A(n8), .B(n3441), .Z(n3442) );
  XOR U3056 ( .A(n3443), .B(n3444), .Z(n3441) );
  AND U3057 ( .A(n34), .B(n3445), .Z(n3444) );
  XOR U3058 ( .A(p_input[6]), .B(n3443), .Z(n3445) );
  XOR U3059 ( .A(n3446), .B(n3447), .Z(n3443) );
  AND U3060 ( .A(n38), .B(n3448), .Z(n3447) );
  XOR U3061 ( .A(n3449), .B(n3450), .Z(n8) );
  AND U3062 ( .A(n42), .B(n3448), .Z(n3450) );
  XNOR U3063 ( .A(n3451), .B(n3446), .Z(n3448) );
  XOR U3064 ( .A(n3452), .B(n3453), .Z(n3446) );
  AND U3065 ( .A(n46), .B(n3454), .Z(n3453) );
  XOR U3066 ( .A(p_input[22]), .B(n3452), .Z(n3454) );
  XOR U3067 ( .A(n3455), .B(n3456), .Z(n3452) );
  AND U3068 ( .A(n50), .B(n3457), .Z(n3456) );
  IV U3069 ( .A(n3449), .Z(n3451) );
  XNOR U3070 ( .A(n3458), .B(n3459), .Z(n3449) );
  AND U3071 ( .A(n54), .B(n3457), .Z(n3459) );
  XNOR U3072 ( .A(n3458), .B(n3455), .Z(n3457) );
  XOR U3073 ( .A(n3460), .B(n3461), .Z(n3455) );
  AND U3074 ( .A(n57), .B(n3462), .Z(n3461) );
  XOR U3075 ( .A(p_input[38]), .B(n3460), .Z(n3462) );
  XOR U3076 ( .A(n3463), .B(n3464), .Z(n3460) );
  AND U3077 ( .A(n61), .B(n3465), .Z(n3464) );
  XOR U3078 ( .A(n3466), .B(n3467), .Z(n3458) );
  AND U3079 ( .A(n65), .B(n3465), .Z(n3467) );
  XNOR U3080 ( .A(n3466), .B(n3463), .Z(n3465) );
  XOR U3081 ( .A(n3468), .B(n3469), .Z(n3463) );
  AND U3082 ( .A(n68), .B(n3470), .Z(n3469) );
  XOR U3083 ( .A(p_input[54]), .B(n3468), .Z(n3470) );
  XOR U3084 ( .A(n3471), .B(n3472), .Z(n3468) );
  AND U3085 ( .A(n72), .B(n3473), .Z(n3472) );
  XOR U3086 ( .A(n3474), .B(n3475), .Z(n3466) );
  AND U3087 ( .A(n76), .B(n3473), .Z(n3475) );
  XNOR U3088 ( .A(n3474), .B(n3471), .Z(n3473) );
  XOR U3089 ( .A(n3476), .B(n3477), .Z(n3471) );
  AND U3090 ( .A(n79), .B(n3478), .Z(n3477) );
  XOR U3091 ( .A(p_input[70]), .B(n3476), .Z(n3478) );
  XOR U3092 ( .A(n3479), .B(n3480), .Z(n3476) );
  AND U3093 ( .A(n83), .B(n3481), .Z(n3480) );
  XOR U3094 ( .A(n3482), .B(n3483), .Z(n3474) );
  AND U3095 ( .A(n87), .B(n3481), .Z(n3483) );
  XNOR U3096 ( .A(n3482), .B(n3479), .Z(n3481) );
  XOR U3097 ( .A(n3484), .B(n3485), .Z(n3479) );
  AND U3098 ( .A(n90), .B(n3486), .Z(n3485) );
  XOR U3099 ( .A(p_input[86]), .B(n3484), .Z(n3486) );
  XOR U3100 ( .A(n3487), .B(n3488), .Z(n3484) );
  AND U3101 ( .A(n94), .B(n3489), .Z(n3488) );
  XOR U3102 ( .A(n3490), .B(n3491), .Z(n3482) );
  AND U3103 ( .A(n98), .B(n3489), .Z(n3491) );
  XNOR U3104 ( .A(n3490), .B(n3487), .Z(n3489) );
  XOR U3105 ( .A(n3492), .B(n3493), .Z(n3487) );
  AND U3106 ( .A(n101), .B(n3494), .Z(n3493) );
  XOR U3107 ( .A(p_input[102]), .B(n3492), .Z(n3494) );
  XOR U3108 ( .A(n3495), .B(n3496), .Z(n3492) );
  AND U3109 ( .A(n105), .B(n3497), .Z(n3496) );
  XOR U3110 ( .A(n3498), .B(n3499), .Z(n3490) );
  AND U3111 ( .A(n109), .B(n3497), .Z(n3499) );
  XNOR U3112 ( .A(n3498), .B(n3495), .Z(n3497) );
  XOR U3113 ( .A(n3500), .B(n3501), .Z(n3495) );
  AND U3114 ( .A(n112), .B(n3502), .Z(n3501) );
  XOR U3115 ( .A(p_input[118]), .B(n3500), .Z(n3502) );
  XOR U3116 ( .A(n3503), .B(n3504), .Z(n3500) );
  AND U3117 ( .A(n116), .B(n3505), .Z(n3504) );
  XOR U3118 ( .A(n3506), .B(n3507), .Z(n3498) );
  AND U3119 ( .A(n120), .B(n3505), .Z(n3507) );
  XNOR U3120 ( .A(n3506), .B(n3503), .Z(n3505) );
  XOR U3121 ( .A(n3508), .B(n3509), .Z(n3503) );
  AND U3122 ( .A(n123), .B(n3510), .Z(n3509) );
  XOR U3123 ( .A(p_input[134]), .B(n3508), .Z(n3510) );
  XOR U3124 ( .A(n3511), .B(n3512), .Z(n3508) );
  AND U3125 ( .A(n127), .B(n3513), .Z(n3512) );
  XOR U3126 ( .A(n3514), .B(n3515), .Z(n3506) );
  AND U3127 ( .A(n131), .B(n3513), .Z(n3515) );
  XNOR U3128 ( .A(n3514), .B(n3511), .Z(n3513) );
  XOR U3129 ( .A(n3516), .B(n3517), .Z(n3511) );
  AND U3130 ( .A(n134), .B(n3518), .Z(n3517) );
  XOR U3131 ( .A(p_input[150]), .B(n3516), .Z(n3518) );
  XOR U3132 ( .A(n3519), .B(n3520), .Z(n3516) );
  AND U3133 ( .A(n138), .B(n3521), .Z(n3520) );
  XOR U3134 ( .A(n3522), .B(n3523), .Z(n3514) );
  AND U3135 ( .A(n142), .B(n3521), .Z(n3523) );
  XNOR U3136 ( .A(n3522), .B(n3519), .Z(n3521) );
  XOR U3137 ( .A(n3524), .B(n3525), .Z(n3519) );
  AND U3138 ( .A(n145), .B(n3526), .Z(n3525) );
  XOR U3139 ( .A(p_input[166]), .B(n3524), .Z(n3526) );
  XOR U3140 ( .A(n3527), .B(n3528), .Z(n3524) );
  AND U3141 ( .A(n149), .B(n3529), .Z(n3528) );
  XOR U3142 ( .A(n3530), .B(n3531), .Z(n3522) );
  AND U3143 ( .A(n153), .B(n3529), .Z(n3531) );
  XNOR U3144 ( .A(n3530), .B(n3527), .Z(n3529) );
  XOR U3145 ( .A(n3532), .B(n3533), .Z(n3527) );
  AND U3146 ( .A(n156), .B(n3534), .Z(n3533) );
  XOR U3147 ( .A(p_input[182]), .B(n3532), .Z(n3534) );
  XOR U3148 ( .A(n3535), .B(n3536), .Z(n3532) );
  AND U3149 ( .A(n160), .B(n3537), .Z(n3536) );
  XOR U3150 ( .A(n3538), .B(n3539), .Z(n3530) );
  AND U3151 ( .A(n164), .B(n3537), .Z(n3539) );
  XNOR U3152 ( .A(n3538), .B(n3535), .Z(n3537) );
  XOR U3153 ( .A(n3540), .B(n3541), .Z(n3535) );
  AND U3154 ( .A(n167), .B(n3542), .Z(n3541) );
  XOR U3155 ( .A(p_input[198]), .B(n3540), .Z(n3542) );
  XOR U3156 ( .A(n3543), .B(n3544), .Z(n3540) );
  AND U3157 ( .A(n171), .B(n3545), .Z(n3544) );
  XOR U3158 ( .A(n3546), .B(n3547), .Z(n3538) );
  AND U3159 ( .A(n175), .B(n3545), .Z(n3547) );
  XNOR U3160 ( .A(n3546), .B(n3543), .Z(n3545) );
  XOR U3161 ( .A(n3548), .B(n3549), .Z(n3543) );
  AND U3162 ( .A(n178), .B(n3550), .Z(n3549) );
  XOR U3163 ( .A(p_input[214]), .B(n3548), .Z(n3550) );
  XOR U3164 ( .A(n3551), .B(n3552), .Z(n3548) );
  AND U3165 ( .A(n182), .B(n3553), .Z(n3552) );
  XOR U3166 ( .A(n3554), .B(n3555), .Z(n3546) );
  AND U3167 ( .A(n186), .B(n3553), .Z(n3555) );
  XNOR U3168 ( .A(n3554), .B(n3551), .Z(n3553) );
  XOR U3169 ( .A(n3556), .B(n3557), .Z(n3551) );
  AND U3170 ( .A(n189), .B(n3558), .Z(n3557) );
  XOR U3171 ( .A(p_input[230]), .B(n3556), .Z(n3558) );
  XOR U3172 ( .A(n3559), .B(n3560), .Z(n3556) );
  AND U3173 ( .A(n193), .B(n3561), .Z(n3560) );
  XOR U3174 ( .A(n3562), .B(n3563), .Z(n3554) );
  AND U3175 ( .A(n197), .B(n3561), .Z(n3563) );
  XNOR U3176 ( .A(n3562), .B(n3559), .Z(n3561) );
  XOR U3177 ( .A(n3564), .B(n3565), .Z(n3559) );
  AND U3178 ( .A(n200), .B(n3566), .Z(n3565) );
  XOR U3179 ( .A(p_input[246]), .B(n3564), .Z(n3566) );
  XOR U3180 ( .A(n3567), .B(n3568), .Z(n3564) );
  AND U3181 ( .A(n204), .B(n3569), .Z(n3568) );
  XOR U3182 ( .A(n3570), .B(n3571), .Z(n3562) );
  AND U3183 ( .A(n208), .B(n3569), .Z(n3571) );
  XNOR U3184 ( .A(n3570), .B(n3567), .Z(n3569) );
  XOR U3185 ( .A(n3572), .B(n3573), .Z(n3567) );
  AND U3186 ( .A(n211), .B(n3574), .Z(n3573) );
  XOR U3187 ( .A(p_input[262]), .B(n3572), .Z(n3574) );
  XOR U3188 ( .A(n3575), .B(n3576), .Z(n3572) );
  AND U3189 ( .A(n215), .B(n3577), .Z(n3576) );
  XOR U3190 ( .A(n3578), .B(n3579), .Z(n3570) );
  AND U3191 ( .A(n219), .B(n3577), .Z(n3579) );
  XNOR U3192 ( .A(n3578), .B(n3575), .Z(n3577) );
  XOR U3193 ( .A(n3580), .B(n3581), .Z(n3575) );
  AND U3194 ( .A(n222), .B(n3582), .Z(n3581) );
  XOR U3195 ( .A(p_input[278]), .B(n3580), .Z(n3582) );
  XOR U3196 ( .A(n3583), .B(n3584), .Z(n3580) );
  AND U3197 ( .A(n226), .B(n3585), .Z(n3584) );
  XOR U3198 ( .A(n3586), .B(n3587), .Z(n3578) );
  AND U3199 ( .A(n230), .B(n3585), .Z(n3587) );
  XNOR U3200 ( .A(n3586), .B(n3583), .Z(n3585) );
  XOR U3201 ( .A(n3588), .B(n3589), .Z(n3583) );
  AND U3202 ( .A(n233), .B(n3590), .Z(n3589) );
  XOR U3203 ( .A(p_input[294]), .B(n3588), .Z(n3590) );
  XOR U3204 ( .A(n3591), .B(n3592), .Z(n3588) );
  AND U3205 ( .A(n237), .B(n3593), .Z(n3592) );
  XOR U3206 ( .A(n3594), .B(n3595), .Z(n3586) );
  AND U3207 ( .A(n241), .B(n3593), .Z(n3595) );
  XNOR U3208 ( .A(n3594), .B(n3591), .Z(n3593) );
  XOR U3209 ( .A(n3596), .B(n3597), .Z(n3591) );
  AND U3210 ( .A(n244), .B(n3598), .Z(n3597) );
  XOR U3211 ( .A(p_input[310]), .B(n3596), .Z(n3598) );
  XOR U3212 ( .A(n3599), .B(n3600), .Z(n3596) );
  AND U3213 ( .A(n248), .B(n3601), .Z(n3600) );
  XOR U3214 ( .A(n3602), .B(n3603), .Z(n3594) );
  AND U3215 ( .A(n252), .B(n3601), .Z(n3603) );
  XNOR U3216 ( .A(n3602), .B(n3599), .Z(n3601) );
  XOR U3217 ( .A(n3604), .B(n3605), .Z(n3599) );
  AND U3218 ( .A(n255), .B(n3606), .Z(n3605) );
  XOR U3219 ( .A(p_input[326]), .B(n3604), .Z(n3606) );
  XOR U3220 ( .A(n3607), .B(n3608), .Z(n3604) );
  AND U3221 ( .A(n259), .B(n3609), .Z(n3608) );
  XOR U3222 ( .A(n3610), .B(n3611), .Z(n3602) );
  AND U3223 ( .A(n263), .B(n3609), .Z(n3611) );
  XNOR U3224 ( .A(n3610), .B(n3607), .Z(n3609) );
  XOR U3225 ( .A(n3612), .B(n3613), .Z(n3607) );
  AND U3226 ( .A(n266), .B(n3614), .Z(n3613) );
  XOR U3227 ( .A(p_input[342]), .B(n3612), .Z(n3614) );
  XOR U3228 ( .A(n3615), .B(n3616), .Z(n3612) );
  AND U3229 ( .A(n270), .B(n3617), .Z(n3616) );
  XOR U3230 ( .A(n3618), .B(n3619), .Z(n3610) );
  AND U3231 ( .A(n274), .B(n3617), .Z(n3619) );
  XNOR U3232 ( .A(n3618), .B(n3615), .Z(n3617) );
  XOR U3233 ( .A(n3620), .B(n3621), .Z(n3615) );
  AND U3234 ( .A(n277), .B(n3622), .Z(n3621) );
  XOR U3235 ( .A(p_input[358]), .B(n3620), .Z(n3622) );
  XOR U3236 ( .A(n3623), .B(n3624), .Z(n3620) );
  AND U3237 ( .A(n281), .B(n3625), .Z(n3624) );
  XOR U3238 ( .A(n3626), .B(n3627), .Z(n3618) );
  AND U3239 ( .A(n285), .B(n3625), .Z(n3627) );
  XNOR U3240 ( .A(n3626), .B(n3623), .Z(n3625) );
  XOR U3241 ( .A(n3628), .B(n3629), .Z(n3623) );
  AND U3242 ( .A(n288), .B(n3630), .Z(n3629) );
  XOR U3243 ( .A(p_input[374]), .B(n3628), .Z(n3630) );
  XOR U3244 ( .A(n3631), .B(n3632), .Z(n3628) );
  AND U3245 ( .A(n292), .B(n3633), .Z(n3632) );
  XOR U3246 ( .A(n3634), .B(n3635), .Z(n3626) );
  AND U3247 ( .A(n296), .B(n3633), .Z(n3635) );
  XNOR U3248 ( .A(n3634), .B(n3631), .Z(n3633) );
  XOR U3249 ( .A(n3636), .B(n3637), .Z(n3631) );
  AND U3250 ( .A(n299), .B(n3638), .Z(n3637) );
  XOR U3251 ( .A(p_input[390]), .B(n3636), .Z(n3638) );
  XOR U3252 ( .A(n3639), .B(n3640), .Z(n3636) );
  AND U3253 ( .A(n303), .B(n3641), .Z(n3640) );
  XOR U3254 ( .A(n3642), .B(n3643), .Z(n3634) );
  AND U3255 ( .A(n307), .B(n3641), .Z(n3643) );
  XNOR U3256 ( .A(n3642), .B(n3639), .Z(n3641) );
  XOR U3257 ( .A(n3644), .B(n3645), .Z(n3639) );
  AND U3258 ( .A(n310), .B(n3646), .Z(n3645) );
  XOR U3259 ( .A(p_input[406]), .B(n3644), .Z(n3646) );
  XOR U3260 ( .A(n3647), .B(n3648), .Z(n3644) );
  AND U3261 ( .A(n314), .B(n3649), .Z(n3648) );
  XOR U3262 ( .A(n3650), .B(n3651), .Z(n3642) );
  AND U3263 ( .A(n318), .B(n3649), .Z(n3651) );
  XNOR U3264 ( .A(n3650), .B(n3647), .Z(n3649) );
  XOR U3265 ( .A(n3652), .B(n3653), .Z(n3647) );
  AND U3266 ( .A(n321), .B(n3654), .Z(n3653) );
  XOR U3267 ( .A(p_input[422]), .B(n3652), .Z(n3654) );
  XOR U3268 ( .A(n3655), .B(n3656), .Z(n3652) );
  AND U3269 ( .A(n325), .B(n3657), .Z(n3656) );
  XOR U3270 ( .A(n3658), .B(n3659), .Z(n3650) );
  AND U3271 ( .A(n329), .B(n3657), .Z(n3659) );
  XNOR U3272 ( .A(n3658), .B(n3655), .Z(n3657) );
  XOR U3273 ( .A(n3660), .B(n3661), .Z(n3655) );
  AND U3274 ( .A(n332), .B(n3662), .Z(n3661) );
  XOR U3275 ( .A(p_input[438]), .B(n3660), .Z(n3662) );
  XOR U3276 ( .A(n3663), .B(n3664), .Z(n3660) );
  AND U3277 ( .A(n336), .B(n3665), .Z(n3664) );
  XOR U3278 ( .A(n3666), .B(n3667), .Z(n3658) );
  AND U3279 ( .A(n340), .B(n3665), .Z(n3667) );
  XNOR U3280 ( .A(n3666), .B(n3663), .Z(n3665) );
  XOR U3281 ( .A(n3668), .B(n3669), .Z(n3663) );
  AND U3282 ( .A(n343), .B(n3670), .Z(n3669) );
  XOR U3283 ( .A(p_input[454]), .B(n3668), .Z(n3670) );
  XOR U3284 ( .A(n3671), .B(n3672), .Z(n3668) );
  AND U3285 ( .A(n347), .B(n3673), .Z(n3672) );
  XOR U3286 ( .A(n3674), .B(n3675), .Z(n3666) );
  AND U3287 ( .A(n351), .B(n3673), .Z(n3675) );
  XNOR U3288 ( .A(n3674), .B(n3671), .Z(n3673) );
  XOR U3289 ( .A(n3676), .B(n3677), .Z(n3671) );
  AND U3290 ( .A(n354), .B(n3678), .Z(n3677) );
  XOR U3291 ( .A(p_input[470]), .B(n3676), .Z(n3678) );
  XOR U3292 ( .A(n3679), .B(n3680), .Z(n3676) );
  AND U3293 ( .A(n358), .B(n3681), .Z(n3680) );
  XOR U3294 ( .A(n3682), .B(n3683), .Z(n3674) );
  AND U3295 ( .A(n362), .B(n3681), .Z(n3683) );
  XNOR U3296 ( .A(n3682), .B(n3679), .Z(n3681) );
  XOR U3297 ( .A(n3684), .B(n3685), .Z(n3679) );
  AND U3298 ( .A(n365), .B(n3686), .Z(n3685) );
  XOR U3299 ( .A(p_input[486]), .B(n3684), .Z(n3686) );
  XOR U3300 ( .A(n3687), .B(n3688), .Z(n3684) );
  AND U3301 ( .A(n369), .B(n3689), .Z(n3688) );
  XOR U3302 ( .A(n3690), .B(n3691), .Z(n3682) );
  AND U3303 ( .A(n373), .B(n3689), .Z(n3691) );
  XNOR U3304 ( .A(n3690), .B(n3687), .Z(n3689) );
  XOR U3305 ( .A(n3692), .B(n3693), .Z(n3687) );
  AND U3306 ( .A(n376), .B(n3694), .Z(n3693) );
  XOR U3307 ( .A(p_input[502]), .B(n3692), .Z(n3694) );
  XOR U3308 ( .A(n3695), .B(n3696), .Z(n3692) );
  AND U3309 ( .A(n380), .B(n3697), .Z(n3696) );
  XOR U3310 ( .A(n3698), .B(n3699), .Z(n3690) );
  AND U3311 ( .A(n384), .B(n3697), .Z(n3699) );
  XNOR U3312 ( .A(n3698), .B(n3695), .Z(n3697) );
  XOR U3313 ( .A(n3700), .B(n3701), .Z(n3695) );
  AND U3314 ( .A(n387), .B(n3702), .Z(n3701) );
  XOR U3315 ( .A(p_input[518]), .B(n3700), .Z(n3702) );
  XOR U3316 ( .A(n3703), .B(n3704), .Z(n3700) );
  AND U3317 ( .A(n391), .B(n3705), .Z(n3704) );
  XOR U3318 ( .A(n3706), .B(n3707), .Z(n3698) );
  AND U3319 ( .A(n395), .B(n3705), .Z(n3707) );
  XNOR U3320 ( .A(n3706), .B(n3703), .Z(n3705) );
  XOR U3321 ( .A(n3708), .B(n3709), .Z(n3703) );
  AND U3322 ( .A(n398), .B(n3710), .Z(n3709) );
  XOR U3323 ( .A(p_input[534]), .B(n3708), .Z(n3710) );
  XOR U3324 ( .A(n3711), .B(n3712), .Z(n3708) );
  AND U3325 ( .A(n402), .B(n3713), .Z(n3712) );
  XOR U3326 ( .A(n3714), .B(n3715), .Z(n3706) );
  AND U3327 ( .A(n406), .B(n3713), .Z(n3715) );
  XNOR U3328 ( .A(n3714), .B(n3711), .Z(n3713) );
  XOR U3329 ( .A(n3716), .B(n3717), .Z(n3711) );
  AND U3330 ( .A(n409), .B(n3718), .Z(n3717) );
  XOR U3331 ( .A(p_input[550]), .B(n3716), .Z(n3718) );
  XOR U3332 ( .A(n3719), .B(n3720), .Z(n3716) );
  AND U3333 ( .A(n413), .B(n3721), .Z(n3720) );
  XOR U3334 ( .A(n3722), .B(n3723), .Z(n3714) );
  AND U3335 ( .A(n417), .B(n3721), .Z(n3723) );
  XNOR U3336 ( .A(n3722), .B(n3719), .Z(n3721) );
  XOR U3337 ( .A(n3724), .B(n3725), .Z(n3719) );
  AND U3338 ( .A(n420), .B(n3726), .Z(n3725) );
  XOR U3339 ( .A(p_input[566]), .B(n3724), .Z(n3726) );
  XOR U3340 ( .A(n3727), .B(n3728), .Z(n3724) );
  AND U3341 ( .A(n424), .B(n3729), .Z(n3728) );
  XOR U3342 ( .A(n3730), .B(n3731), .Z(n3722) );
  AND U3343 ( .A(n428), .B(n3729), .Z(n3731) );
  XNOR U3344 ( .A(n3730), .B(n3727), .Z(n3729) );
  XOR U3345 ( .A(n3732), .B(n3733), .Z(n3727) );
  AND U3346 ( .A(n431), .B(n3734), .Z(n3733) );
  XOR U3347 ( .A(p_input[582]), .B(n3732), .Z(n3734) );
  XOR U3348 ( .A(n3735), .B(n3736), .Z(n3732) );
  AND U3349 ( .A(n435), .B(n3737), .Z(n3736) );
  XOR U3350 ( .A(n3738), .B(n3739), .Z(n3730) );
  AND U3351 ( .A(n439), .B(n3737), .Z(n3739) );
  XNOR U3352 ( .A(n3738), .B(n3735), .Z(n3737) );
  XOR U3353 ( .A(n3740), .B(n3741), .Z(n3735) );
  AND U3354 ( .A(n442), .B(n3742), .Z(n3741) );
  XOR U3355 ( .A(p_input[598]), .B(n3740), .Z(n3742) );
  XOR U3356 ( .A(n3743), .B(n3744), .Z(n3740) );
  AND U3357 ( .A(n446), .B(n3745), .Z(n3744) );
  XOR U3358 ( .A(n3746), .B(n3747), .Z(n3738) );
  AND U3359 ( .A(n450), .B(n3745), .Z(n3747) );
  XNOR U3360 ( .A(n3746), .B(n3743), .Z(n3745) );
  XOR U3361 ( .A(n3748), .B(n3749), .Z(n3743) );
  AND U3362 ( .A(n453), .B(n3750), .Z(n3749) );
  XOR U3363 ( .A(p_input[614]), .B(n3748), .Z(n3750) );
  XOR U3364 ( .A(n3751), .B(n3752), .Z(n3748) );
  AND U3365 ( .A(n457), .B(n3753), .Z(n3752) );
  XOR U3366 ( .A(n3754), .B(n3755), .Z(n3746) );
  AND U3367 ( .A(n461), .B(n3753), .Z(n3755) );
  XNOR U3368 ( .A(n3754), .B(n3751), .Z(n3753) );
  XOR U3369 ( .A(n3756), .B(n3757), .Z(n3751) );
  AND U3370 ( .A(n464), .B(n3758), .Z(n3757) );
  XOR U3371 ( .A(p_input[630]), .B(n3756), .Z(n3758) );
  XOR U3372 ( .A(n3759), .B(n3760), .Z(n3756) );
  AND U3373 ( .A(n468), .B(n3761), .Z(n3760) );
  XOR U3374 ( .A(n3762), .B(n3763), .Z(n3754) );
  AND U3375 ( .A(n472), .B(n3761), .Z(n3763) );
  XNOR U3376 ( .A(n3762), .B(n3759), .Z(n3761) );
  XOR U3377 ( .A(n3764), .B(n3765), .Z(n3759) );
  AND U3378 ( .A(n475), .B(n3766), .Z(n3765) );
  XOR U3379 ( .A(p_input[646]), .B(n3764), .Z(n3766) );
  XOR U3380 ( .A(n3767), .B(n3768), .Z(n3764) );
  AND U3381 ( .A(n479), .B(n3769), .Z(n3768) );
  XOR U3382 ( .A(n3770), .B(n3771), .Z(n3762) );
  AND U3383 ( .A(n483), .B(n3769), .Z(n3771) );
  XNOR U3384 ( .A(n3770), .B(n3767), .Z(n3769) );
  XOR U3385 ( .A(n3772), .B(n3773), .Z(n3767) );
  AND U3386 ( .A(n486), .B(n3774), .Z(n3773) );
  XOR U3387 ( .A(p_input[662]), .B(n3772), .Z(n3774) );
  XOR U3388 ( .A(n3775), .B(n3776), .Z(n3772) );
  AND U3389 ( .A(n490), .B(n3777), .Z(n3776) );
  XOR U3390 ( .A(n3778), .B(n3779), .Z(n3770) );
  AND U3391 ( .A(n494), .B(n3777), .Z(n3779) );
  XNOR U3392 ( .A(n3778), .B(n3775), .Z(n3777) );
  XOR U3393 ( .A(n3780), .B(n3781), .Z(n3775) );
  AND U3394 ( .A(n497), .B(n3782), .Z(n3781) );
  XOR U3395 ( .A(p_input[678]), .B(n3780), .Z(n3782) );
  XOR U3396 ( .A(n3783), .B(n3784), .Z(n3780) );
  AND U3397 ( .A(n501), .B(n3785), .Z(n3784) );
  XOR U3398 ( .A(n3786), .B(n3787), .Z(n3778) );
  AND U3399 ( .A(n505), .B(n3785), .Z(n3787) );
  XNOR U3400 ( .A(n3786), .B(n3783), .Z(n3785) );
  XOR U3401 ( .A(n3788), .B(n3789), .Z(n3783) );
  AND U3402 ( .A(n508), .B(n3790), .Z(n3789) );
  XOR U3403 ( .A(p_input[694]), .B(n3788), .Z(n3790) );
  XOR U3404 ( .A(n3791), .B(n3792), .Z(n3788) );
  AND U3405 ( .A(n512), .B(n3793), .Z(n3792) );
  XOR U3406 ( .A(n3794), .B(n3795), .Z(n3786) );
  AND U3407 ( .A(n516), .B(n3793), .Z(n3795) );
  XNOR U3408 ( .A(n3794), .B(n3791), .Z(n3793) );
  XOR U3409 ( .A(n3796), .B(n3797), .Z(n3791) );
  AND U3410 ( .A(n519), .B(n3798), .Z(n3797) );
  XOR U3411 ( .A(p_input[710]), .B(n3796), .Z(n3798) );
  XOR U3412 ( .A(n3799), .B(n3800), .Z(n3796) );
  AND U3413 ( .A(n523), .B(n3801), .Z(n3800) );
  XOR U3414 ( .A(n3802), .B(n3803), .Z(n3794) );
  AND U3415 ( .A(n527), .B(n3801), .Z(n3803) );
  XNOR U3416 ( .A(n3802), .B(n3799), .Z(n3801) );
  XOR U3417 ( .A(n3804), .B(n3805), .Z(n3799) );
  AND U3418 ( .A(n530), .B(n3806), .Z(n3805) );
  XOR U3419 ( .A(p_input[726]), .B(n3804), .Z(n3806) );
  XOR U3420 ( .A(n3807), .B(n3808), .Z(n3804) );
  AND U3421 ( .A(n534), .B(n3809), .Z(n3808) );
  XOR U3422 ( .A(n3810), .B(n3811), .Z(n3802) );
  AND U3423 ( .A(n538), .B(n3809), .Z(n3811) );
  XNOR U3424 ( .A(n3810), .B(n3807), .Z(n3809) );
  XOR U3425 ( .A(n3812), .B(n3813), .Z(n3807) );
  AND U3426 ( .A(n541), .B(n3814), .Z(n3813) );
  XOR U3427 ( .A(p_input[742]), .B(n3812), .Z(n3814) );
  XOR U3428 ( .A(n3815), .B(n3816), .Z(n3812) );
  AND U3429 ( .A(n545), .B(n3817), .Z(n3816) );
  XOR U3430 ( .A(n3818), .B(n3819), .Z(n3810) );
  AND U3431 ( .A(n549), .B(n3817), .Z(n3819) );
  XNOR U3432 ( .A(n3818), .B(n3815), .Z(n3817) );
  XOR U3433 ( .A(n3820), .B(n3821), .Z(n3815) );
  AND U3434 ( .A(n552), .B(n3822), .Z(n3821) );
  XOR U3435 ( .A(p_input[758]), .B(n3820), .Z(n3822) );
  XOR U3436 ( .A(n3823), .B(n3824), .Z(n3820) );
  AND U3437 ( .A(n556), .B(n3825), .Z(n3824) );
  XOR U3438 ( .A(n3826), .B(n3827), .Z(n3818) );
  AND U3439 ( .A(n560), .B(n3825), .Z(n3827) );
  XNOR U3440 ( .A(n3826), .B(n3823), .Z(n3825) );
  XOR U3441 ( .A(n3828), .B(n3829), .Z(n3823) );
  AND U3442 ( .A(n563), .B(n3830), .Z(n3829) );
  XOR U3443 ( .A(p_input[774]), .B(n3828), .Z(n3830) );
  XOR U3444 ( .A(n3831), .B(n3832), .Z(n3828) );
  AND U3445 ( .A(n567), .B(n3833), .Z(n3832) );
  XOR U3446 ( .A(n3834), .B(n3835), .Z(n3826) );
  AND U3447 ( .A(n571), .B(n3833), .Z(n3835) );
  XNOR U3448 ( .A(n3834), .B(n3831), .Z(n3833) );
  XOR U3449 ( .A(n3836), .B(n3837), .Z(n3831) );
  AND U3450 ( .A(n574), .B(n3838), .Z(n3837) );
  XOR U3451 ( .A(p_input[790]), .B(n3836), .Z(n3838) );
  XOR U3452 ( .A(n3839), .B(n3840), .Z(n3836) );
  AND U3453 ( .A(n578), .B(n3841), .Z(n3840) );
  XOR U3454 ( .A(n3842), .B(n3843), .Z(n3834) );
  AND U3455 ( .A(n582), .B(n3841), .Z(n3843) );
  XNOR U3456 ( .A(n3842), .B(n3839), .Z(n3841) );
  XOR U3457 ( .A(n3844), .B(n3845), .Z(n3839) );
  AND U3458 ( .A(n585), .B(n3846), .Z(n3845) );
  XOR U3459 ( .A(p_input[806]), .B(n3844), .Z(n3846) );
  XOR U3460 ( .A(n3847), .B(n3848), .Z(n3844) );
  AND U3461 ( .A(n589), .B(n3849), .Z(n3848) );
  XOR U3462 ( .A(n3850), .B(n3851), .Z(n3842) );
  AND U3463 ( .A(n593), .B(n3849), .Z(n3851) );
  XNOR U3464 ( .A(n3850), .B(n3847), .Z(n3849) );
  XOR U3465 ( .A(n3852), .B(n3853), .Z(n3847) );
  AND U3466 ( .A(n596), .B(n3854), .Z(n3853) );
  XOR U3467 ( .A(p_input[822]), .B(n3852), .Z(n3854) );
  XOR U3468 ( .A(n3855), .B(n3856), .Z(n3852) );
  AND U3469 ( .A(n600), .B(n3857), .Z(n3856) );
  XOR U3470 ( .A(n3858), .B(n3859), .Z(n3850) );
  AND U3471 ( .A(n604), .B(n3857), .Z(n3859) );
  XNOR U3472 ( .A(n3858), .B(n3855), .Z(n3857) );
  XOR U3473 ( .A(n3860), .B(n3861), .Z(n3855) );
  AND U3474 ( .A(n607), .B(n3862), .Z(n3861) );
  XOR U3475 ( .A(p_input[838]), .B(n3860), .Z(n3862) );
  XOR U3476 ( .A(n3863), .B(n3864), .Z(n3860) );
  AND U3477 ( .A(n611), .B(n3865), .Z(n3864) );
  XOR U3478 ( .A(n3866), .B(n3867), .Z(n3858) );
  AND U3479 ( .A(n615), .B(n3865), .Z(n3867) );
  XNOR U3480 ( .A(n3866), .B(n3863), .Z(n3865) );
  XOR U3481 ( .A(n3868), .B(n3869), .Z(n3863) );
  AND U3482 ( .A(n618), .B(n3870), .Z(n3869) );
  XOR U3483 ( .A(p_input[854]), .B(n3868), .Z(n3870) );
  XOR U3484 ( .A(n3871), .B(n3872), .Z(n3868) );
  AND U3485 ( .A(n622), .B(n3873), .Z(n3872) );
  XOR U3486 ( .A(n3874), .B(n3875), .Z(n3866) );
  AND U3487 ( .A(n626), .B(n3873), .Z(n3875) );
  XNOR U3488 ( .A(n3874), .B(n3871), .Z(n3873) );
  XOR U3489 ( .A(n3876), .B(n3877), .Z(n3871) );
  AND U3490 ( .A(n629), .B(n3878), .Z(n3877) );
  XOR U3491 ( .A(p_input[870]), .B(n3876), .Z(n3878) );
  XOR U3492 ( .A(n3879), .B(n3880), .Z(n3876) );
  AND U3493 ( .A(n633), .B(n3881), .Z(n3880) );
  XOR U3494 ( .A(n3882), .B(n3883), .Z(n3874) );
  AND U3495 ( .A(n637), .B(n3881), .Z(n3883) );
  XNOR U3496 ( .A(n3882), .B(n3879), .Z(n3881) );
  XOR U3497 ( .A(n3884), .B(n3885), .Z(n3879) );
  AND U3498 ( .A(n640), .B(n3886), .Z(n3885) );
  XOR U3499 ( .A(p_input[886]), .B(n3884), .Z(n3886) );
  XOR U3500 ( .A(n3887), .B(n3888), .Z(n3884) );
  AND U3501 ( .A(n644), .B(n3889), .Z(n3888) );
  XOR U3502 ( .A(n3890), .B(n3891), .Z(n3882) );
  AND U3503 ( .A(n648), .B(n3889), .Z(n3891) );
  XNOR U3504 ( .A(n3890), .B(n3887), .Z(n3889) );
  XOR U3505 ( .A(n3892), .B(n3893), .Z(n3887) );
  AND U3506 ( .A(n651), .B(n3894), .Z(n3893) );
  XOR U3507 ( .A(p_input[902]), .B(n3892), .Z(n3894) );
  XOR U3508 ( .A(n3895), .B(n3896), .Z(n3892) );
  AND U3509 ( .A(n655), .B(n3897), .Z(n3896) );
  XOR U3510 ( .A(n3898), .B(n3899), .Z(n3890) );
  AND U3511 ( .A(n659), .B(n3897), .Z(n3899) );
  XNOR U3512 ( .A(n3898), .B(n3895), .Z(n3897) );
  XOR U3513 ( .A(n3900), .B(n3901), .Z(n3895) );
  AND U3514 ( .A(n662), .B(n3902), .Z(n3901) );
  XOR U3515 ( .A(p_input[918]), .B(n3900), .Z(n3902) );
  XOR U3516 ( .A(n3903), .B(n3904), .Z(n3900) );
  AND U3517 ( .A(n666), .B(n3905), .Z(n3904) );
  XOR U3518 ( .A(n3906), .B(n3907), .Z(n3898) );
  AND U3519 ( .A(n670), .B(n3905), .Z(n3907) );
  XNOR U3520 ( .A(n3906), .B(n3903), .Z(n3905) );
  XOR U3521 ( .A(n3908), .B(n3909), .Z(n3903) );
  AND U3522 ( .A(n673), .B(n3910), .Z(n3909) );
  XOR U3523 ( .A(p_input[934]), .B(n3908), .Z(n3910) );
  XOR U3524 ( .A(n3911), .B(n3912), .Z(n3908) );
  AND U3525 ( .A(n677), .B(n3913), .Z(n3912) );
  XOR U3526 ( .A(n3914), .B(n3915), .Z(n3906) );
  AND U3527 ( .A(n681), .B(n3913), .Z(n3915) );
  XNOR U3528 ( .A(n3914), .B(n3911), .Z(n3913) );
  XOR U3529 ( .A(n3916), .B(n3917), .Z(n3911) );
  AND U3530 ( .A(n684), .B(n3918), .Z(n3917) );
  XOR U3531 ( .A(p_input[950]), .B(n3916), .Z(n3918) );
  XOR U3532 ( .A(n3919), .B(n3920), .Z(n3916) );
  AND U3533 ( .A(n688), .B(n3921), .Z(n3920) );
  XOR U3534 ( .A(n3922), .B(n3923), .Z(n3914) );
  AND U3535 ( .A(n692), .B(n3921), .Z(n3923) );
  XNOR U3536 ( .A(n3922), .B(n3919), .Z(n3921) );
  XOR U3537 ( .A(n3924), .B(n3925), .Z(n3919) );
  AND U3538 ( .A(n695), .B(n3926), .Z(n3925) );
  XOR U3539 ( .A(p_input[966]), .B(n3924), .Z(n3926) );
  XOR U3540 ( .A(n3927), .B(n3928), .Z(n3924) );
  AND U3541 ( .A(n699), .B(n3929), .Z(n3928) );
  XOR U3542 ( .A(n3930), .B(n3931), .Z(n3922) );
  AND U3543 ( .A(n703), .B(n3929), .Z(n3931) );
  XNOR U3544 ( .A(n3930), .B(n3927), .Z(n3929) );
  XOR U3545 ( .A(n3932), .B(n3933), .Z(n3927) );
  AND U3546 ( .A(n706), .B(n3934), .Z(n3933) );
  XOR U3547 ( .A(p_input[982]), .B(n3932), .Z(n3934) );
  XOR U3548 ( .A(n3935), .B(n3936), .Z(n3932) );
  AND U3549 ( .A(n710), .B(n3937), .Z(n3936) );
  XOR U3550 ( .A(n3938), .B(n3939), .Z(n3930) );
  AND U3551 ( .A(n714), .B(n3937), .Z(n3939) );
  XNOR U3552 ( .A(n3938), .B(n3935), .Z(n3937) );
  XOR U3553 ( .A(n3940), .B(n3941), .Z(n3935) );
  AND U3554 ( .A(n717), .B(n3942), .Z(n3941) );
  XOR U3555 ( .A(p_input[998]), .B(n3940), .Z(n3942) );
  XOR U3556 ( .A(n3943), .B(n3944), .Z(n3940) );
  AND U3557 ( .A(n721), .B(n3945), .Z(n3944) );
  XOR U3558 ( .A(n3946), .B(n3947), .Z(n3938) );
  AND U3559 ( .A(n725), .B(n3945), .Z(n3947) );
  XNOR U3560 ( .A(n3946), .B(n3943), .Z(n3945) );
  XOR U3561 ( .A(n3948), .B(n3949), .Z(n3943) );
  AND U3562 ( .A(n728), .B(n3950), .Z(n3949) );
  XOR U3563 ( .A(p_input[1014]), .B(n3948), .Z(n3950) );
  XOR U3564 ( .A(n3951), .B(n3952), .Z(n3948) );
  AND U3565 ( .A(n732), .B(n3953), .Z(n3952) );
  XOR U3566 ( .A(n3954), .B(n3955), .Z(n3946) );
  AND U3567 ( .A(n736), .B(n3953), .Z(n3955) );
  XNOR U3568 ( .A(n3954), .B(n3951), .Z(n3953) );
  XOR U3569 ( .A(n3956), .B(n3957), .Z(n3951) );
  AND U3570 ( .A(n739), .B(n3958), .Z(n3957) );
  XOR U3571 ( .A(p_input[1030]), .B(n3956), .Z(n3958) );
  XOR U3572 ( .A(n3959), .B(n3960), .Z(n3956) );
  AND U3573 ( .A(n743), .B(n3961), .Z(n3960) );
  XOR U3574 ( .A(n3962), .B(n3963), .Z(n3954) );
  AND U3575 ( .A(n747), .B(n3961), .Z(n3963) );
  XNOR U3576 ( .A(n3962), .B(n3959), .Z(n3961) );
  XOR U3577 ( .A(n3964), .B(n3965), .Z(n3959) );
  AND U3578 ( .A(n750), .B(n3966), .Z(n3965) );
  XOR U3579 ( .A(p_input[1046]), .B(n3964), .Z(n3966) );
  XOR U3580 ( .A(n3967), .B(n3968), .Z(n3964) );
  AND U3581 ( .A(n754), .B(n3969), .Z(n3968) );
  XOR U3582 ( .A(n3970), .B(n3971), .Z(n3962) );
  AND U3583 ( .A(n758), .B(n3969), .Z(n3971) );
  XNOR U3584 ( .A(n3970), .B(n3967), .Z(n3969) );
  XOR U3585 ( .A(n3972), .B(n3973), .Z(n3967) );
  AND U3586 ( .A(n761), .B(n3974), .Z(n3973) );
  XOR U3587 ( .A(p_input[1062]), .B(n3972), .Z(n3974) );
  XOR U3588 ( .A(n3975), .B(n3976), .Z(n3972) );
  AND U3589 ( .A(n765), .B(n3977), .Z(n3976) );
  XOR U3590 ( .A(n3978), .B(n3979), .Z(n3970) );
  AND U3591 ( .A(n769), .B(n3977), .Z(n3979) );
  XNOR U3592 ( .A(n3978), .B(n3975), .Z(n3977) );
  XOR U3593 ( .A(n3980), .B(n3981), .Z(n3975) );
  AND U3594 ( .A(n772), .B(n3982), .Z(n3981) );
  XOR U3595 ( .A(p_input[1078]), .B(n3980), .Z(n3982) );
  XOR U3596 ( .A(n3983), .B(n3984), .Z(n3980) );
  AND U3597 ( .A(n776), .B(n3985), .Z(n3984) );
  XOR U3598 ( .A(n3986), .B(n3987), .Z(n3978) );
  AND U3599 ( .A(n780), .B(n3985), .Z(n3987) );
  XNOR U3600 ( .A(n3986), .B(n3983), .Z(n3985) );
  XOR U3601 ( .A(n3988), .B(n3989), .Z(n3983) );
  AND U3602 ( .A(n783), .B(n3990), .Z(n3989) );
  XOR U3603 ( .A(p_input[1094]), .B(n3988), .Z(n3990) );
  XOR U3604 ( .A(n3991), .B(n3992), .Z(n3988) );
  AND U3605 ( .A(n787), .B(n3993), .Z(n3992) );
  XOR U3606 ( .A(n3994), .B(n3995), .Z(n3986) );
  AND U3607 ( .A(n791), .B(n3993), .Z(n3995) );
  XNOR U3608 ( .A(n3994), .B(n3991), .Z(n3993) );
  XOR U3609 ( .A(n3996), .B(n3997), .Z(n3991) );
  AND U3610 ( .A(n794), .B(n3998), .Z(n3997) );
  XOR U3611 ( .A(p_input[1110]), .B(n3996), .Z(n3998) );
  XOR U3612 ( .A(n3999), .B(n4000), .Z(n3996) );
  AND U3613 ( .A(n798), .B(n4001), .Z(n4000) );
  XOR U3614 ( .A(n4002), .B(n4003), .Z(n3994) );
  AND U3615 ( .A(n802), .B(n4001), .Z(n4003) );
  XNOR U3616 ( .A(n4002), .B(n3999), .Z(n4001) );
  XOR U3617 ( .A(n4004), .B(n4005), .Z(n3999) );
  AND U3618 ( .A(n805), .B(n4006), .Z(n4005) );
  XOR U3619 ( .A(p_input[1126]), .B(n4004), .Z(n4006) );
  XOR U3620 ( .A(n4007), .B(n4008), .Z(n4004) );
  AND U3621 ( .A(n809), .B(n4009), .Z(n4008) );
  XOR U3622 ( .A(n4010), .B(n4011), .Z(n4002) );
  AND U3623 ( .A(n813), .B(n4009), .Z(n4011) );
  XNOR U3624 ( .A(n4010), .B(n4007), .Z(n4009) );
  XOR U3625 ( .A(n4012), .B(n4013), .Z(n4007) );
  AND U3626 ( .A(n816), .B(n4014), .Z(n4013) );
  XOR U3627 ( .A(p_input[1142]), .B(n4012), .Z(n4014) );
  XOR U3628 ( .A(n4015), .B(n4016), .Z(n4012) );
  AND U3629 ( .A(n820), .B(n4017), .Z(n4016) );
  XOR U3630 ( .A(n4018), .B(n4019), .Z(n4010) );
  AND U3631 ( .A(n824), .B(n4017), .Z(n4019) );
  XNOR U3632 ( .A(n4018), .B(n4015), .Z(n4017) );
  XOR U3633 ( .A(n4020), .B(n4021), .Z(n4015) );
  AND U3634 ( .A(n827), .B(n4022), .Z(n4021) );
  XOR U3635 ( .A(p_input[1158]), .B(n4020), .Z(n4022) );
  XOR U3636 ( .A(n4023), .B(n4024), .Z(n4020) );
  AND U3637 ( .A(n831), .B(n4025), .Z(n4024) );
  XOR U3638 ( .A(n4026), .B(n4027), .Z(n4018) );
  AND U3639 ( .A(n835), .B(n4025), .Z(n4027) );
  XNOR U3640 ( .A(n4026), .B(n4023), .Z(n4025) );
  XOR U3641 ( .A(n4028), .B(n4029), .Z(n4023) );
  AND U3642 ( .A(n838), .B(n4030), .Z(n4029) );
  XOR U3643 ( .A(p_input[1174]), .B(n4028), .Z(n4030) );
  XOR U3644 ( .A(n4031), .B(n4032), .Z(n4028) );
  AND U3645 ( .A(n842), .B(n4033), .Z(n4032) );
  XOR U3646 ( .A(n4034), .B(n4035), .Z(n4026) );
  AND U3647 ( .A(n846), .B(n4033), .Z(n4035) );
  XNOR U3648 ( .A(n4034), .B(n4031), .Z(n4033) );
  XOR U3649 ( .A(n4036), .B(n4037), .Z(n4031) );
  AND U3650 ( .A(n849), .B(n4038), .Z(n4037) );
  XOR U3651 ( .A(p_input[1190]), .B(n4036), .Z(n4038) );
  XOR U3652 ( .A(n4039), .B(n4040), .Z(n4036) );
  AND U3653 ( .A(n853), .B(n4041), .Z(n4040) );
  XOR U3654 ( .A(n4042), .B(n4043), .Z(n4034) );
  AND U3655 ( .A(n857), .B(n4041), .Z(n4043) );
  XNOR U3656 ( .A(n4042), .B(n4039), .Z(n4041) );
  XOR U3657 ( .A(n4044), .B(n4045), .Z(n4039) );
  AND U3658 ( .A(n860), .B(n4046), .Z(n4045) );
  XOR U3659 ( .A(p_input[1206]), .B(n4044), .Z(n4046) );
  XOR U3660 ( .A(n4047), .B(n4048), .Z(n4044) );
  AND U3661 ( .A(n864), .B(n4049), .Z(n4048) );
  XOR U3662 ( .A(n4050), .B(n4051), .Z(n4042) );
  AND U3663 ( .A(n868), .B(n4049), .Z(n4051) );
  XNOR U3664 ( .A(n4050), .B(n4047), .Z(n4049) );
  XOR U3665 ( .A(n4052), .B(n4053), .Z(n4047) );
  AND U3666 ( .A(n871), .B(n4054), .Z(n4053) );
  XOR U3667 ( .A(p_input[1222]), .B(n4052), .Z(n4054) );
  XOR U3668 ( .A(n4055), .B(n4056), .Z(n4052) );
  AND U3669 ( .A(n875), .B(n4057), .Z(n4056) );
  XOR U3670 ( .A(n4058), .B(n4059), .Z(n4050) );
  AND U3671 ( .A(n879), .B(n4057), .Z(n4059) );
  XNOR U3672 ( .A(n4058), .B(n4055), .Z(n4057) );
  XOR U3673 ( .A(n4060), .B(n4061), .Z(n4055) );
  AND U3674 ( .A(n882), .B(n4062), .Z(n4061) );
  XOR U3675 ( .A(p_input[1238]), .B(n4060), .Z(n4062) );
  XOR U3676 ( .A(n4063), .B(n4064), .Z(n4060) );
  AND U3677 ( .A(n886), .B(n4065), .Z(n4064) );
  XOR U3678 ( .A(n4066), .B(n4067), .Z(n4058) );
  AND U3679 ( .A(n890), .B(n4065), .Z(n4067) );
  XNOR U3680 ( .A(n4066), .B(n4063), .Z(n4065) );
  XOR U3681 ( .A(n4068), .B(n4069), .Z(n4063) );
  AND U3682 ( .A(n893), .B(n4070), .Z(n4069) );
  XOR U3683 ( .A(p_input[1254]), .B(n4068), .Z(n4070) );
  XOR U3684 ( .A(n4071), .B(n4072), .Z(n4068) );
  AND U3685 ( .A(n897), .B(n4073), .Z(n4072) );
  XOR U3686 ( .A(n4074), .B(n4075), .Z(n4066) );
  AND U3687 ( .A(n901), .B(n4073), .Z(n4075) );
  XNOR U3688 ( .A(n4074), .B(n4071), .Z(n4073) );
  XOR U3689 ( .A(n4076), .B(n4077), .Z(n4071) );
  AND U3690 ( .A(n904), .B(n4078), .Z(n4077) );
  XOR U3691 ( .A(p_input[1270]), .B(n4076), .Z(n4078) );
  XOR U3692 ( .A(n4079), .B(n4080), .Z(n4076) );
  AND U3693 ( .A(n908), .B(n4081), .Z(n4080) );
  XOR U3694 ( .A(n4082), .B(n4083), .Z(n4074) );
  AND U3695 ( .A(n912), .B(n4081), .Z(n4083) );
  XNOR U3696 ( .A(n4082), .B(n4079), .Z(n4081) );
  XOR U3697 ( .A(n4084), .B(n4085), .Z(n4079) );
  AND U3698 ( .A(n915), .B(n4086), .Z(n4085) );
  XOR U3699 ( .A(p_input[1286]), .B(n4084), .Z(n4086) );
  XOR U3700 ( .A(n4087), .B(n4088), .Z(n4084) );
  AND U3701 ( .A(n919), .B(n4089), .Z(n4088) );
  XOR U3702 ( .A(n4090), .B(n4091), .Z(n4082) );
  AND U3703 ( .A(n923), .B(n4089), .Z(n4091) );
  XNOR U3704 ( .A(n4090), .B(n4087), .Z(n4089) );
  XOR U3705 ( .A(n4092), .B(n4093), .Z(n4087) );
  AND U3706 ( .A(n926), .B(n4094), .Z(n4093) );
  XOR U3707 ( .A(p_input[1302]), .B(n4092), .Z(n4094) );
  XOR U3708 ( .A(n4095), .B(n4096), .Z(n4092) );
  AND U3709 ( .A(n930), .B(n4097), .Z(n4096) );
  XOR U3710 ( .A(n4098), .B(n4099), .Z(n4090) );
  AND U3711 ( .A(n934), .B(n4097), .Z(n4099) );
  XNOR U3712 ( .A(n4098), .B(n4095), .Z(n4097) );
  XOR U3713 ( .A(n4100), .B(n4101), .Z(n4095) );
  AND U3714 ( .A(n937), .B(n4102), .Z(n4101) );
  XOR U3715 ( .A(p_input[1318]), .B(n4100), .Z(n4102) );
  XOR U3716 ( .A(n4103), .B(n4104), .Z(n4100) );
  AND U3717 ( .A(n941), .B(n4105), .Z(n4104) );
  XOR U3718 ( .A(n4106), .B(n4107), .Z(n4098) );
  AND U3719 ( .A(n945), .B(n4105), .Z(n4107) );
  XNOR U3720 ( .A(n4106), .B(n4103), .Z(n4105) );
  XOR U3721 ( .A(n4108), .B(n4109), .Z(n4103) );
  AND U3722 ( .A(n948), .B(n4110), .Z(n4109) );
  XOR U3723 ( .A(p_input[1334]), .B(n4108), .Z(n4110) );
  XOR U3724 ( .A(n4111), .B(n4112), .Z(n4108) );
  AND U3725 ( .A(n952), .B(n4113), .Z(n4112) );
  XOR U3726 ( .A(n4114), .B(n4115), .Z(n4106) );
  AND U3727 ( .A(n956), .B(n4113), .Z(n4115) );
  XNOR U3728 ( .A(n4114), .B(n4111), .Z(n4113) );
  XOR U3729 ( .A(n4116), .B(n4117), .Z(n4111) );
  AND U3730 ( .A(n959), .B(n4118), .Z(n4117) );
  XOR U3731 ( .A(p_input[1350]), .B(n4116), .Z(n4118) );
  XOR U3732 ( .A(n4119), .B(n4120), .Z(n4116) );
  AND U3733 ( .A(n963), .B(n4121), .Z(n4120) );
  XOR U3734 ( .A(n4122), .B(n4123), .Z(n4114) );
  AND U3735 ( .A(n967), .B(n4121), .Z(n4123) );
  XNOR U3736 ( .A(n4122), .B(n4119), .Z(n4121) );
  XOR U3737 ( .A(n4124), .B(n4125), .Z(n4119) );
  AND U3738 ( .A(n970), .B(n4126), .Z(n4125) );
  XOR U3739 ( .A(p_input[1366]), .B(n4124), .Z(n4126) );
  XOR U3740 ( .A(n4127), .B(n4128), .Z(n4124) );
  AND U3741 ( .A(n974), .B(n4129), .Z(n4128) );
  XOR U3742 ( .A(n4130), .B(n4131), .Z(n4122) );
  AND U3743 ( .A(n978), .B(n4129), .Z(n4131) );
  XNOR U3744 ( .A(n4130), .B(n4127), .Z(n4129) );
  XOR U3745 ( .A(n4132), .B(n4133), .Z(n4127) );
  AND U3746 ( .A(n981), .B(n4134), .Z(n4133) );
  XOR U3747 ( .A(p_input[1382]), .B(n4132), .Z(n4134) );
  XOR U3748 ( .A(n4135), .B(n4136), .Z(n4132) );
  AND U3749 ( .A(n985), .B(n4137), .Z(n4136) );
  XOR U3750 ( .A(n4138), .B(n4139), .Z(n4130) );
  AND U3751 ( .A(n989), .B(n4137), .Z(n4139) );
  XNOR U3752 ( .A(n4138), .B(n4135), .Z(n4137) );
  XOR U3753 ( .A(n4140), .B(n4141), .Z(n4135) );
  AND U3754 ( .A(n992), .B(n4142), .Z(n4141) );
  XOR U3755 ( .A(p_input[1398]), .B(n4140), .Z(n4142) );
  XOR U3756 ( .A(n4143), .B(n4144), .Z(n4140) );
  AND U3757 ( .A(n996), .B(n4145), .Z(n4144) );
  XOR U3758 ( .A(n4146), .B(n4147), .Z(n4138) );
  AND U3759 ( .A(n1000), .B(n4145), .Z(n4147) );
  XNOR U3760 ( .A(n4146), .B(n4143), .Z(n4145) );
  XOR U3761 ( .A(n4148), .B(n4149), .Z(n4143) );
  AND U3762 ( .A(n1003), .B(n4150), .Z(n4149) );
  XOR U3763 ( .A(p_input[1414]), .B(n4148), .Z(n4150) );
  XOR U3764 ( .A(n4151), .B(n4152), .Z(n4148) );
  AND U3765 ( .A(n1007), .B(n4153), .Z(n4152) );
  XOR U3766 ( .A(n4154), .B(n4155), .Z(n4146) );
  AND U3767 ( .A(n1011), .B(n4153), .Z(n4155) );
  XNOR U3768 ( .A(n4154), .B(n4151), .Z(n4153) );
  XOR U3769 ( .A(n4156), .B(n4157), .Z(n4151) );
  AND U3770 ( .A(n1014), .B(n4158), .Z(n4157) );
  XOR U3771 ( .A(p_input[1430]), .B(n4156), .Z(n4158) );
  XOR U3772 ( .A(n4159), .B(n4160), .Z(n4156) );
  AND U3773 ( .A(n1018), .B(n4161), .Z(n4160) );
  XOR U3774 ( .A(n4162), .B(n4163), .Z(n4154) );
  AND U3775 ( .A(n1022), .B(n4161), .Z(n4163) );
  XNOR U3776 ( .A(n4162), .B(n4159), .Z(n4161) );
  XOR U3777 ( .A(n4164), .B(n4165), .Z(n4159) );
  AND U3778 ( .A(n1025), .B(n4166), .Z(n4165) );
  XOR U3779 ( .A(p_input[1446]), .B(n4164), .Z(n4166) );
  XOR U3780 ( .A(n4167), .B(n4168), .Z(n4164) );
  AND U3781 ( .A(n1029), .B(n4169), .Z(n4168) );
  XOR U3782 ( .A(n4170), .B(n4171), .Z(n4162) );
  AND U3783 ( .A(n1033), .B(n4169), .Z(n4171) );
  XNOR U3784 ( .A(n4170), .B(n4167), .Z(n4169) );
  XOR U3785 ( .A(n4172), .B(n4173), .Z(n4167) );
  AND U3786 ( .A(n1036), .B(n4174), .Z(n4173) );
  XOR U3787 ( .A(p_input[1462]), .B(n4172), .Z(n4174) );
  XOR U3788 ( .A(n4175), .B(n4176), .Z(n4172) );
  AND U3789 ( .A(n1040), .B(n4177), .Z(n4176) );
  XOR U3790 ( .A(n4178), .B(n4179), .Z(n4170) );
  AND U3791 ( .A(n1044), .B(n4177), .Z(n4179) );
  XNOR U3792 ( .A(n4178), .B(n4175), .Z(n4177) );
  XOR U3793 ( .A(n4180), .B(n4181), .Z(n4175) );
  AND U3794 ( .A(n1047), .B(n4182), .Z(n4181) );
  XOR U3795 ( .A(p_input[1478]), .B(n4180), .Z(n4182) );
  XOR U3796 ( .A(n4183), .B(n4184), .Z(n4180) );
  AND U3797 ( .A(n1051), .B(n4185), .Z(n4184) );
  XOR U3798 ( .A(n4186), .B(n4187), .Z(n4178) );
  AND U3799 ( .A(n1055), .B(n4185), .Z(n4187) );
  XNOR U3800 ( .A(n4186), .B(n4183), .Z(n4185) );
  XOR U3801 ( .A(n4188), .B(n4189), .Z(n4183) );
  AND U3802 ( .A(n1058), .B(n4190), .Z(n4189) );
  XOR U3803 ( .A(p_input[1494]), .B(n4188), .Z(n4190) );
  XOR U3804 ( .A(n4191), .B(n4192), .Z(n4188) );
  AND U3805 ( .A(n1062), .B(n4193), .Z(n4192) );
  XOR U3806 ( .A(n4194), .B(n4195), .Z(n4186) );
  AND U3807 ( .A(n1066), .B(n4193), .Z(n4195) );
  XNOR U3808 ( .A(n4194), .B(n4191), .Z(n4193) );
  XOR U3809 ( .A(n4196), .B(n4197), .Z(n4191) );
  AND U3810 ( .A(n1069), .B(n4198), .Z(n4197) );
  XOR U3811 ( .A(p_input[1510]), .B(n4196), .Z(n4198) );
  XOR U3812 ( .A(n4199), .B(n4200), .Z(n4196) );
  AND U3813 ( .A(n1073), .B(n4201), .Z(n4200) );
  XOR U3814 ( .A(n4202), .B(n4203), .Z(n4194) );
  AND U3815 ( .A(n1077), .B(n4201), .Z(n4203) );
  XNOR U3816 ( .A(n4202), .B(n4199), .Z(n4201) );
  XOR U3817 ( .A(n4204), .B(n4205), .Z(n4199) );
  AND U3818 ( .A(n1080), .B(n4206), .Z(n4205) );
  XOR U3819 ( .A(p_input[1526]), .B(n4204), .Z(n4206) );
  XOR U3820 ( .A(n4207), .B(n4208), .Z(n4204) );
  AND U3821 ( .A(n1084), .B(n4209), .Z(n4208) );
  XOR U3822 ( .A(n4210), .B(n4211), .Z(n4202) );
  AND U3823 ( .A(n1088), .B(n4209), .Z(n4211) );
  XNOR U3824 ( .A(n4210), .B(n4207), .Z(n4209) );
  XOR U3825 ( .A(n4212), .B(n4213), .Z(n4207) );
  AND U3826 ( .A(n1091), .B(n4214), .Z(n4213) );
  XOR U3827 ( .A(p_input[1542]), .B(n4212), .Z(n4214) );
  XOR U3828 ( .A(n4215), .B(n4216), .Z(n4212) );
  AND U3829 ( .A(n1095), .B(n4217), .Z(n4216) );
  XOR U3830 ( .A(n4218), .B(n4219), .Z(n4210) );
  AND U3831 ( .A(n1099), .B(n4217), .Z(n4219) );
  XNOR U3832 ( .A(n4218), .B(n4215), .Z(n4217) );
  XOR U3833 ( .A(n4220), .B(n4221), .Z(n4215) );
  AND U3834 ( .A(n1102), .B(n4222), .Z(n4221) );
  XOR U3835 ( .A(p_input[1558]), .B(n4220), .Z(n4222) );
  XOR U3836 ( .A(n4223), .B(n4224), .Z(n4220) );
  AND U3837 ( .A(n1106), .B(n4225), .Z(n4224) );
  XOR U3838 ( .A(n4226), .B(n4227), .Z(n4218) );
  AND U3839 ( .A(n1110), .B(n4225), .Z(n4227) );
  XNOR U3840 ( .A(n4226), .B(n4223), .Z(n4225) );
  XOR U3841 ( .A(n4228), .B(n4229), .Z(n4223) );
  AND U3842 ( .A(n1113), .B(n4230), .Z(n4229) );
  XOR U3843 ( .A(p_input[1574]), .B(n4228), .Z(n4230) );
  XOR U3844 ( .A(n4231), .B(n4232), .Z(n4228) );
  AND U3845 ( .A(n1117), .B(n4233), .Z(n4232) );
  XOR U3846 ( .A(n4234), .B(n4235), .Z(n4226) );
  AND U3847 ( .A(n1121), .B(n4233), .Z(n4235) );
  XNOR U3848 ( .A(n4234), .B(n4231), .Z(n4233) );
  XOR U3849 ( .A(n4236), .B(n4237), .Z(n4231) );
  AND U3850 ( .A(n1124), .B(n4238), .Z(n4237) );
  XOR U3851 ( .A(p_input[1590]), .B(n4236), .Z(n4238) );
  XOR U3852 ( .A(n4239), .B(n4240), .Z(n4236) );
  AND U3853 ( .A(n1128), .B(n4241), .Z(n4240) );
  XOR U3854 ( .A(n4242), .B(n4243), .Z(n4234) );
  AND U3855 ( .A(n1132), .B(n4241), .Z(n4243) );
  XNOR U3856 ( .A(n4242), .B(n4239), .Z(n4241) );
  XOR U3857 ( .A(n4244), .B(n4245), .Z(n4239) );
  AND U3858 ( .A(n1135), .B(n4246), .Z(n4245) );
  XOR U3859 ( .A(p_input[1606]), .B(n4244), .Z(n4246) );
  XOR U3860 ( .A(n4247), .B(n4248), .Z(n4244) );
  AND U3861 ( .A(n1139), .B(n4249), .Z(n4248) );
  XOR U3862 ( .A(n4250), .B(n4251), .Z(n4242) );
  AND U3863 ( .A(n1143), .B(n4249), .Z(n4251) );
  XNOR U3864 ( .A(n4250), .B(n4247), .Z(n4249) );
  XOR U3865 ( .A(n4252), .B(n4253), .Z(n4247) );
  AND U3866 ( .A(n1146), .B(n4254), .Z(n4253) );
  XOR U3867 ( .A(p_input[1622]), .B(n4252), .Z(n4254) );
  XOR U3868 ( .A(n4255), .B(n4256), .Z(n4252) );
  AND U3869 ( .A(n1150), .B(n4257), .Z(n4256) );
  XOR U3870 ( .A(n4258), .B(n4259), .Z(n4250) );
  AND U3871 ( .A(n1154), .B(n4257), .Z(n4259) );
  XNOR U3872 ( .A(n4258), .B(n4255), .Z(n4257) );
  XOR U3873 ( .A(n4260), .B(n4261), .Z(n4255) );
  AND U3874 ( .A(n1157), .B(n4262), .Z(n4261) );
  XOR U3875 ( .A(p_input[1638]), .B(n4260), .Z(n4262) );
  XOR U3876 ( .A(n4263), .B(n4264), .Z(n4260) );
  AND U3877 ( .A(n1161), .B(n4265), .Z(n4264) );
  XOR U3878 ( .A(n4266), .B(n4267), .Z(n4258) );
  AND U3879 ( .A(n1165), .B(n4265), .Z(n4267) );
  XNOR U3880 ( .A(n4266), .B(n4263), .Z(n4265) );
  XOR U3881 ( .A(n4268), .B(n4269), .Z(n4263) );
  AND U3882 ( .A(n1168), .B(n4270), .Z(n4269) );
  XOR U3883 ( .A(p_input[1654]), .B(n4268), .Z(n4270) );
  XOR U3884 ( .A(n4271), .B(n4272), .Z(n4268) );
  AND U3885 ( .A(n1172), .B(n4273), .Z(n4272) );
  XOR U3886 ( .A(n4274), .B(n4275), .Z(n4266) );
  AND U3887 ( .A(n1176), .B(n4273), .Z(n4275) );
  XNOR U3888 ( .A(n4274), .B(n4271), .Z(n4273) );
  XOR U3889 ( .A(n4276), .B(n4277), .Z(n4271) );
  AND U3890 ( .A(n1179), .B(n4278), .Z(n4277) );
  XOR U3891 ( .A(p_input[1670]), .B(n4276), .Z(n4278) );
  XOR U3892 ( .A(n4279), .B(n4280), .Z(n4276) );
  AND U3893 ( .A(n1183), .B(n4281), .Z(n4280) );
  XOR U3894 ( .A(n4282), .B(n4283), .Z(n4274) );
  AND U3895 ( .A(n1187), .B(n4281), .Z(n4283) );
  XNOR U3896 ( .A(n4282), .B(n4279), .Z(n4281) );
  XOR U3897 ( .A(n4284), .B(n4285), .Z(n4279) );
  AND U3898 ( .A(n1190), .B(n4286), .Z(n4285) );
  XOR U3899 ( .A(p_input[1686]), .B(n4284), .Z(n4286) );
  XOR U3900 ( .A(n4287), .B(n4288), .Z(n4284) );
  AND U3901 ( .A(n1194), .B(n4289), .Z(n4288) );
  XOR U3902 ( .A(n4290), .B(n4291), .Z(n4282) );
  AND U3903 ( .A(n1198), .B(n4289), .Z(n4291) );
  XNOR U3904 ( .A(n4290), .B(n4287), .Z(n4289) );
  XOR U3905 ( .A(n4292), .B(n4293), .Z(n4287) );
  AND U3906 ( .A(n1201), .B(n4294), .Z(n4293) );
  XOR U3907 ( .A(p_input[1702]), .B(n4292), .Z(n4294) );
  XOR U3908 ( .A(n4295), .B(n4296), .Z(n4292) );
  AND U3909 ( .A(n1205), .B(n4297), .Z(n4296) );
  XOR U3910 ( .A(n4298), .B(n4299), .Z(n4290) );
  AND U3911 ( .A(n1209), .B(n4297), .Z(n4299) );
  XNOR U3912 ( .A(n4298), .B(n4295), .Z(n4297) );
  XOR U3913 ( .A(n4300), .B(n4301), .Z(n4295) );
  AND U3914 ( .A(n1212), .B(n4302), .Z(n4301) );
  XOR U3915 ( .A(p_input[1718]), .B(n4300), .Z(n4302) );
  XOR U3916 ( .A(n4303), .B(n4304), .Z(n4300) );
  AND U3917 ( .A(n1216), .B(n4305), .Z(n4304) );
  XOR U3918 ( .A(n4306), .B(n4307), .Z(n4298) );
  AND U3919 ( .A(n1220), .B(n4305), .Z(n4307) );
  XNOR U3920 ( .A(n4306), .B(n4303), .Z(n4305) );
  XOR U3921 ( .A(n4308), .B(n4309), .Z(n4303) );
  AND U3922 ( .A(n1223), .B(n4310), .Z(n4309) );
  XOR U3923 ( .A(p_input[1734]), .B(n4308), .Z(n4310) );
  XOR U3924 ( .A(n4311), .B(n4312), .Z(n4308) );
  AND U3925 ( .A(n1227), .B(n4313), .Z(n4312) );
  XOR U3926 ( .A(n4314), .B(n4315), .Z(n4306) );
  AND U3927 ( .A(n1231), .B(n4313), .Z(n4315) );
  XNOR U3928 ( .A(n4314), .B(n4311), .Z(n4313) );
  XOR U3929 ( .A(n4316), .B(n4317), .Z(n4311) );
  AND U3930 ( .A(n1234), .B(n4318), .Z(n4317) );
  XOR U3931 ( .A(p_input[1750]), .B(n4316), .Z(n4318) );
  XOR U3932 ( .A(n4319), .B(n4320), .Z(n4316) );
  AND U3933 ( .A(n1238), .B(n4321), .Z(n4320) );
  XOR U3934 ( .A(n4322), .B(n4323), .Z(n4314) );
  AND U3935 ( .A(n1242), .B(n4321), .Z(n4323) );
  XNOR U3936 ( .A(n4322), .B(n4319), .Z(n4321) );
  XOR U3937 ( .A(n4324), .B(n4325), .Z(n4319) );
  AND U3938 ( .A(n1245), .B(n4326), .Z(n4325) );
  XOR U3939 ( .A(p_input[1766]), .B(n4324), .Z(n4326) );
  XOR U3940 ( .A(n4327), .B(n4328), .Z(n4324) );
  AND U3941 ( .A(n1249), .B(n4329), .Z(n4328) );
  XOR U3942 ( .A(n4330), .B(n4331), .Z(n4322) );
  AND U3943 ( .A(n1253), .B(n4329), .Z(n4331) );
  XNOR U3944 ( .A(n4330), .B(n4327), .Z(n4329) );
  XOR U3945 ( .A(n4332), .B(n4333), .Z(n4327) );
  AND U3946 ( .A(n1256), .B(n4334), .Z(n4333) );
  XOR U3947 ( .A(p_input[1782]), .B(n4332), .Z(n4334) );
  XOR U3948 ( .A(n4335), .B(n4336), .Z(n4332) );
  AND U3949 ( .A(n1260), .B(n4337), .Z(n4336) );
  XOR U3950 ( .A(n4338), .B(n4339), .Z(n4330) );
  AND U3951 ( .A(n1264), .B(n4337), .Z(n4339) );
  XNOR U3952 ( .A(n4338), .B(n4335), .Z(n4337) );
  XOR U3953 ( .A(n4340), .B(n4341), .Z(n4335) );
  AND U3954 ( .A(n1267), .B(n4342), .Z(n4341) );
  XOR U3955 ( .A(p_input[1798]), .B(n4340), .Z(n4342) );
  XOR U3956 ( .A(n4343), .B(n4344), .Z(n4340) );
  AND U3957 ( .A(n1271), .B(n4345), .Z(n4344) );
  XOR U3958 ( .A(n4346), .B(n4347), .Z(n4338) );
  AND U3959 ( .A(n1275), .B(n4345), .Z(n4347) );
  XNOR U3960 ( .A(n4346), .B(n4343), .Z(n4345) );
  XOR U3961 ( .A(n4348), .B(n4349), .Z(n4343) );
  AND U3962 ( .A(n1278), .B(n4350), .Z(n4349) );
  XOR U3963 ( .A(p_input[1814]), .B(n4348), .Z(n4350) );
  XOR U3964 ( .A(n4351), .B(n4352), .Z(n4348) );
  AND U3965 ( .A(n1282), .B(n4353), .Z(n4352) );
  XOR U3966 ( .A(n4354), .B(n4355), .Z(n4346) );
  AND U3967 ( .A(n1286), .B(n4353), .Z(n4355) );
  XNOR U3968 ( .A(n4354), .B(n4351), .Z(n4353) );
  XOR U3969 ( .A(n4356), .B(n4357), .Z(n4351) );
  AND U3970 ( .A(n1289), .B(n4358), .Z(n4357) );
  XOR U3971 ( .A(p_input[1830]), .B(n4356), .Z(n4358) );
  XOR U3972 ( .A(n4359), .B(n4360), .Z(n4356) );
  AND U3973 ( .A(n1293), .B(n4361), .Z(n4360) );
  XOR U3974 ( .A(n4362), .B(n4363), .Z(n4354) );
  AND U3975 ( .A(n1297), .B(n4361), .Z(n4363) );
  XNOR U3976 ( .A(n4362), .B(n4359), .Z(n4361) );
  XOR U3977 ( .A(n4364), .B(n4365), .Z(n4359) );
  AND U3978 ( .A(n1300), .B(n4366), .Z(n4365) );
  XOR U3979 ( .A(p_input[1846]), .B(n4364), .Z(n4366) );
  XOR U3980 ( .A(n4367), .B(n4368), .Z(n4364) );
  AND U3981 ( .A(n1304), .B(n4369), .Z(n4368) );
  XOR U3982 ( .A(n4370), .B(n4371), .Z(n4362) );
  AND U3983 ( .A(n1308), .B(n4369), .Z(n4371) );
  XNOR U3984 ( .A(n4370), .B(n4367), .Z(n4369) );
  XOR U3985 ( .A(n4372), .B(n4373), .Z(n4367) );
  AND U3986 ( .A(n1311), .B(n4374), .Z(n4373) );
  XOR U3987 ( .A(p_input[1862]), .B(n4372), .Z(n4374) );
  XOR U3988 ( .A(n4375), .B(n4376), .Z(n4372) );
  AND U3989 ( .A(n1315), .B(n4377), .Z(n4376) );
  XOR U3990 ( .A(n4378), .B(n4379), .Z(n4370) );
  AND U3991 ( .A(n1319), .B(n4377), .Z(n4379) );
  XNOR U3992 ( .A(n4378), .B(n4375), .Z(n4377) );
  XOR U3993 ( .A(n4380), .B(n4381), .Z(n4375) );
  AND U3994 ( .A(n1322), .B(n4382), .Z(n4381) );
  XOR U3995 ( .A(p_input[1878]), .B(n4380), .Z(n4382) );
  XOR U3996 ( .A(n4383), .B(n4384), .Z(n4380) );
  AND U3997 ( .A(n1326), .B(n4385), .Z(n4384) );
  XOR U3998 ( .A(n4386), .B(n4387), .Z(n4378) );
  AND U3999 ( .A(n1330), .B(n4385), .Z(n4387) );
  XNOR U4000 ( .A(n4386), .B(n4383), .Z(n4385) );
  XOR U4001 ( .A(n4388), .B(n4389), .Z(n4383) );
  AND U4002 ( .A(n1333), .B(n4390), .Z(n4389) );
  XOR U4003 ( .A(p_input[1894]), .B(n4388), .Z(n4390) );
  XOR U4004 ( .A(n4391), .B(n4392), .Z(n4388) );
  AND U4005 ( .A(n1337), .B(n4393), .Z(n4392) );
  XOR U4006 ( .A(n4394), .B(n4395), .Z(n4386) );
  AND U4007 ( .A(n1341), .B(n4393), .Z(n4395) );
  XNOR U4008 ( .A(n4394), .B(n4391), .Z(n4393) );
  XOR U4009 ( .A(n4396), .B(n4397), .Z(n4391) );
  AND U4010 ( .A(n1344), .B(n4398), .Z(n4397) );
  XOR U4011 ( .A(p_input[1910]), .B(n4396), .Z(n4398) );
  XOR U4012 ( .A(n4399), .B(n4400), .Z(n4396) );
  AND U4013 ( .A(n1348), .B(n4401), .Z(n4400) );
  XOR U4014 ( .A(n4402), .B(n4403), .Z(n4394) );
  AND U4015 ( .A(n1352), .B(n4401), .Z(n4403) );
  XNOR U4016 ( .A(n4402), .B(n4399), .Z(n4401) );
  XOR U4017 ( .A(n4404), .B(n4405), .Z(n4399) );
  AND U4018 ( .A(n1355), .B(n4406), .Z(n4405) );
  XOR U4019 ( .A(p_input[1926]), .B(n4404), .Z(n4406) );
  XOR U4020 ( .A(n4407), .B(n4408), .Z(n4404) );
  AND U4021 ( .A(n1359), .B(n4409), .Z(n4408) );
  XOR U4022 ( .A(n4410), .B(n4411), .Z(n4402) );
  AND U4023 ( .A(n1363), .B(n4409), .Z(n4411) );
  XNOR U4024 ( .A(n4410), .B(n4407), .Z(n4409) );
  XOR U4025 ( .A(n4412), .B(n4413), .Z(n4407) );
  AND U4026 ( .A(n1366), .B(n4414), .Z(n4413) );
  XOR U4027 ( .A(p_input[1942]), .B(n4412), .Z(n4414) );
  XOR U4028 ( .A(n4415), .B(n4416), .Z(n4412) );
  AND U4029 ( .A(n1370), .B(n4417), .Z(n4416) );
  XOR U4030 ( .A(n4418), .B(n4419), .Z(n4410) );
  AND U4031 ( .A(n1374), .B(n4417), .Z(n4419) );
  XNOR U4032 ( .A(n4418), .B(n4415), .Z(n4417) );
  XOR U4033 ( .A(n4420), .B(n4421), .Z(n4415) );
  AND U4034 ( .A(n1377), .B(n4422), .Z(n4421) );
  XOR U4035 ( .A(p_input[1958]), .B(n4420), .Z(n4422) );
  XOR U4036 ( .A(n4423), .B(n4424), .Z(n4420) );
  AND U4037 ( .A(n1381), .B(n4425), .Z(n4424) );
  XOR U4038 ( .A(n4426), .B(n4427), .Z(n4418) );
  AND U4039 ( .A(n1385), .B(n4425), .Z(n4427) );
  XNOR U4040 ( .A(n4426), .B(n4423), .Z(n4425) );
  XOR U4041 ( .A(n4428), .B(n4429), .Z(n4423) );
  AND U4042 ( .A(n1388), .B(n4430), .Z(n4429) );
  XOR U4043 ( .A(p_input[1974]), .B(n4428), .Z(n4430) );
  XOR U4044 ( .A(n4431), .B(n4432), .Z(n4428) );
  AND U4045 ( .A(n1392), .B(n4433), .Z(n4432) );
  XOR U4046 ( .A(n4434), .B(n4435), .Z(n4426) );
  AND U4047 ( .A(n1396), .B(n4433), .Z(n4435) );
  XNOR U4048 ( .A(n4434), .B(n4431), .Z(n4433) );
  XOR U4049 ( .A(n4436), .B(n4437), .Z(n4431) );
  AND U4050 ( .A(n1399), .B(n4438), .Z(n4437) );
  XOR U4051 ( .A(p_input[1990]), .B(n4436), .Z(n4438) );
  XOR U4052 ( .A(n4439), .B(n4440), .Z(n4436) );
  AND U4053 ( .A(n1403), .B(n4441), .Z(n4440) );
  XOR U4054 ( .A(n4442), .B(n4443), .Z(n4434) );
  AND U4055 ( .A(n1407), .B(n4441), .Z(n4443) );
  XNOR U4056 ( .A(n4442), .B(n4439), .Z(n4441) );
  XOR U4057 ( .A(n4444), .B(n4445), .Z(n4439) );
  AND U4058 ( .A(n1410), .B(n4446), .Z(n4445) );
  XOR U4059 ( .A(p_input[2006]), .B(n4444), .Z(n4446) );
  XNOR U4060 ( .A(n4447), .B(n4448), .Z(n4444) );
  AND U4061 ( .A(n1414), .B(n4449), .Z(n4448) );
  XNOR U4062 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n4450), .Z(n4442) );
  AND U4063 ( .A(n1417), .B(n4449), .Z(n4450) );
  XOR U4064 ( .A(n4451), .B(n4447), .Z(n4449) );
  XOR U4065 ( .A(n9), .B(n4452), .Z(o[21]) );
  AND U4066 ( .A(n30), .B(n4453), .Z(n9) );
  XOR U4067 ( .A(n10), .B(n4452), .Z(n4453) );
  XOR U4068 ( .A(n4454), .B(n4455), .Z(n4452) );
  AND U4069 ( .A(n34), .B(n4456), .Z(n4455) );
  XOR U4070 ( .A(p_input[5]), .B(n4454), .Z(n4456) );
  XOR U4071 ( .A(n4457), .B(n4458), .Z(n4454) );
  AND U4072 ( .A(n38), .B(n4459), .Z(n4458) );
  XOR U4073 ( .A(n4460), .B(n4461), .Z(n10) );
  AND U4074 ( .A(n42), .B(n4459), .Z(n4461) );
  XNOR U4075 ( .A(n4462), .B(n4457), .Z(n4459) );
  XOR U4076 ( .A(n4463), .B(n4464), .Z(n4457) );
  AND U4077 ( .A(n46), .B(n4465), .Z(n4464) );
  XOR U4078 ( .A(p_input[21]), .B(n4463), .Z(n4465) );
  XOR U4079 ( .A(n4466), .B(n4467), .Z(n4463) );
  AND U4080 ( .A(n50), .B(n4468), .Z(n4467) );
  IV U4081 ( .A(n4460), .Z(n4462) );
  XNOR U4082 ( .A(n4469), .B(n4470), .Z(n4460) );
  AND U4083 ( .A(n54), .B(n4468), .Z(n4470) );
  XNOR U4084 ( .A(n4469), .B(n4466), .Z(n4468) );
  XOR U4085 ( .A(n4471), .B(n4472), .Z(n4466) );
  AND U4086 ( .A(n57), .B(n4473), .Z(n4472) );
  XOR U4087 ( .A(p_input[37]), .B(n4471), .Z(n4473) );
  XOR U4088 ( .A(n4474), .B(n4475), .Z(n4471) );
  AND U4089 ( .A(n61), .B(n4476), .Z(n4475) );
  XOR U4090 ( .A(n4477), .B(n4478), .Z(n4469) );
  AND U4091 ( .A(n65), .B(n4476), .Z(n4478) );
  XNOR U4092 ( .A(n4477), .B(n4474), .Z(n4476) );
  XOR U4093 ( .A(n4479), .B(n4480), .Z(n4474) );
  AND U4094 ( .A(n68), .B(n4481), .Z(n4480) );
  XOR U4095 ( .A(p_input[53]), .B(n4479), .Z(n4481) );
  XOR U4096 ( .A(n4482), .B(n4483), .Z(n4479) );
  AND U4097 ( .A(n72), .B(n4484), .Z(n4483) );
  XOR U4098 ( .A(n4485), .B(n4486), .Z(n4477) );
  AND U4099 ( .A(n76), .B(n4484), .Z(n4486) );
  XNOR U4100 ( .A(n4485), .B(n4482), .Z(n4484) );
  XOR U4101 ( .A(n4487), .B(n4488), .Z(n4482) );
  AND U4102 ( .A(n79), .B(n4489), .Z(n4488) );
  XOR U4103 ( .A(p_input[69]), .B(n4487), .Z(n4489) );
  XOR U4104 ( .A(n4490), .B(n4491), .Z(n4487) );
  AND U4105 ( .A(n83), .B(n4492), .Z(n4491) );
  XOR U4106 ( .A(n4493), .B(n4494), .Z(n4485) );
  AND U4107 ( .A(n87), .B(n4492), .Z(n4494) );
  XNOR U4108 ( .A(n4493), .B(n4490), .Z(n4492) );
  XOR U4109 ( .A(n4495), .B(n4496), .Z(n4490) );
  AND U4110 ( .A(n90), .B(n4497), .Z(n4496) );
  XOR U4111 ( .A(p_input[85]), .B(n4495), .Z(n4497) );
  XOR U4112 ( .A(n4498), .B(n4499), .Z(n4495) );
  AND U4113 ( .A(n94), .B(n4500), .Z(n4499) );
  XOR U4114 ( .A(n4501), .B(n4502), .Z(n4493) );
  AND U4115 ( .A(n98), .B(n4500), .Z(n4502) );
  XNOR U4116 ( .A(n4501), .B(n4498), .Z(n4500) );
  XOR U4117 ( .A(n4503), .B(n4504), .Z(n4498) );
  AND U4118 ( .A(n101), .B(n4505), .Z(n4504) );
  XOR U4119 ( .A(p_input[101]), .B(n4503), .Z(n4505) );
  XOR U4120 ( .A(n4506), .B(n4507), .Z(n4503) );
  AND U4121 ( .A(n105), .B(n4508), .Z(n4507) );
  XOR U4122 ( .A(n4509), .B(n4510), .Z(n4501) );
  AND U4123 ( .A(n109), .B(n4508), .Z(n4510) );
  XNOR U4124 ( .A(n4509), .B(n4506), .Z(n4508) );
  XOR U4125 ( .A(n4511), .B(n4512), .Z(n4506) );
  AND U4126 ( .A(n112), .B(n4513), .Z(n4512) );
  XOR U4127 ( .A(p_input[117]), .B(n4511), .Z(n4513) );
  XOR U4128 ( .A(n4514), .B(n4515), .Z(n4511) );
  AND U4129 ( .A(n116), .B(n4516), .Z(n4515) );
  XOR U4130 ( .A(n4517), .B(n4518), .Z(n4509) );
  AND U4131 ( .A(n120), .B(n4516), .Z(n4518) );
  XNOR U4132 ( .A(n4517), .B(n4514), .Z(n4516) );
  XOR U4133 ( .A(n4519), .B(n4520), .Z(n4514) );
  AND U4134 ( .A(n123), .B(n4521), .Z(n4520) );
  XOR U4135 ( .A(p_input[133]), .B(n4519), .Z(n4521) );
  XOR U4136 ( .A(n4522), .B(n4523), .Z(n4519) );
  AND U4137 ( .A(n127), .B(n4524), .Z(n4523) );
  XOR U4138 ( .A(n4525), .B(n4526), .Z(n4517) );
  AND U4139 ( .A(n131), .B(n4524), .Z(n4526) );
  XNOR U4140 ( .A(n4525), .B(n4522), .Z(n4524) );
  XOR U4141 ( .A(n4527), .B(n4528), .Z(n4522) );
  AND U4142 ( .A(n134), .B(n4529), .Z(n4528) );
  XOR U4143 ( .A(p_input[149]), .B(n4527), .Z(n4529) );
  XOR U4144 ( .A(n4530), .B(n4531), .Z(n4527) );
  AND U4145 ( .A(n138), .B(n4532), .Z(n4531) );
  XOR U4146 ( .A(n4533), .B(n4534), .Z(n4525) );
  AND U4147 ( .A(n142), .B(n4532), .Z(n4534) );
  XNOR U4148 ( .A(n4533), .B(n4530), .Z(n4532) );
  XOR U4149 ( .A(n4535), .B(n4536), .Z(n4530) );
  AND U4150 ( .A(n145), .B(n4537), .Z(n4536) );
  XOR U4151 ( .A(p_input[165]), .B(n4535), .Z(n4537) );
  XOR U4152 ( .A(n4538), .B(n4539), .Z(n4535) );
  AND U4153 ( .A(n149), .B(n4540), .Z(n4539) );
  XOR U4154 ( .A(n4541), .B(n4542), .Z(n4533) );
  AND U4155 ( .A(n153), .B(n4540), .Z(n4542) );
  XNOR U4156 ( .A(n4541), .B(n4538), .Z(n4540) );
  XOR U4157 ( .A(n4543), .B(n4544), .Z(n4538) );
  AND U4158 ( .A(n156), .B(n4545), .Z(n4544) );
  XOR U4159 ( .A(p_input[181]), .B(n4543), .Z(n4545) );
  XOR U4160 ( .A(n4546), .B(n4547), .Z(n4543) );
  AND U4161 ( .A(n160), .B(n4548), .Z(n4547) );
  XOR U4162 ( .A(n4549), .B(n4550), .Z(n4541) );
  AND U4163 ( .A(n164), .B(n4548), .Z(n4550) );
  XNOR U4164 ( .A(n4549), .B(n4546), .Z(n4548) );
  XOR U4165 ( .A(n4551), .B(n4552), .Z(n4546) );
  AND U4166 ( .A(n167), .B(n4553), .Z(n4552) );
  XOR U4167 ( .A(p_input[197]), .B(n4551), .Z(n4553) );
  XOR U4168 ( .A(n4554), .B(n4555), .Z(n4551) );
  AND U4169 ( .A(n171), .B(n4556), .Z(n4555) );
  XOR U4170 ( .A(n4557), .B(n4558), .Z(n4549) );
  AND U4171 ( .A(n175), .B(n4556), .Z(n4558) );
  XNOR U4172 ( .A(n4557), .B(n4554), .Z(n4556) );
  XOR U4173 ( .A(n4559), .B(n4560), .Z(n4554) );
  AND U4174 ( .A(n178), .B(n4561), .Z(n4560) );
  XOR U4175 ( .A(p_input[213]), .B(n4559), .Z(n4561) );
  XOR U4176 ( .A(n4562), .B(n4563), .Z(n4559) );
  AND U4177 ( .A(n182), .B(n4564), .Z(n4563) );
  XOR U4178 ( .A(n4565), .B(n4566), .Z(n4557) );
  AND U4179 ( .A(n186), .B(n4564), .Z(n4566) );
  XNOR U4180 ( .A(n4565), .B(n4562), .Z(n4564) );
  XOR U4181 ( .A(n4567), .B(n4568), .Z(n4562) );
  AND U4182 ( .A(n189), .B(n4569), .Z(n4568) );
  XOR U4183 ( .A(p_input[229]), .B(n4567), .Z(n4569) );
  XOR U4184 ( .A(n4570), .B(n4571), .Z(n4567) );
  AND U4185 ( .A(n193), .B(n4572), .Z(n4571) );
  XOR U4186 ( .A(n4573), .B(n4574), .Z(n4565) );
  AND U4187 ( .A(n197), .B(n4572), .Z(n4574) );
  XNOR U4188 ( .A(n4573), .B(n4570), .Z(n4572) );
  XOR U4189 ( .A(n4575), .B(n4576), .Z(n4570) );
  AND U4190 ( .A(n200), .B(n4577), .Z(n4576) );
  XOR U4191 ( .A(p_input[245]), .B(n4575), .Z(n4577) );
  XOR U4192 ( .A(n4578), .B(n4579), .Z(n4575) );
  AND U4193 ( .A(n204), .B(n4580), .Z(n4579) );
  XOR U4194 ( .A(n4581), .B(n4582), .Z(n4573) );
  AND U4195 ( .A(n208), .B(n4580), .Z(n4582) );
  XNOR U4196 ( .A(n4581), .B(n4578), .Z(n4580) );
  XOR U4197 ( .A(n4583), .B(n4584), .Z(n4578) );
  AND U4198 ( .A(n211), .B(n4585), .Z(n4584) );
  XOR U4199 ( .A(p_input[261]), .B(n4583), .Z(n4585) );
  XOR U4200 ( .A(n4586), .B(n4587), .Z(n4583) );
  AND U4201 ( .A(n215), .B(n4588), .Z(n4587) );
  XOR U4202 ( .A(n4589), .B(n4590), .Z(n4581) );
  AND U4203 ( .A(n219), .B(n4588), .Z(n4590) );
  XNOR U4204 ( .A(n4589), .B(n4586), .Z(n4588) );
  XOR U4205 ( .A(n4591), .B(n4592), .Z(n4586) );
  AND U4206 ( .A(n222), .B(n4593), .Z(n4592) );
  XOR U4207 ( .A(p_input[277]), .B(n4591), .Z(n4593) );
  XOR U4208 ( .A(n4594), .B(n4595), .Z(n4591) );
  AND U4209 ( .A(n226), .B(n4596), .Z(n4595) );
  XOR U4210 ( .A(n4597), .B(n4598), .Z(n4589) );
  AND U4211 ( .A(n230), .B(n4596), .Z(n4598) );
  XNOR U4212 ( .A(n4597), .B(n4594), .Z(n4596) );
  XOR U4213 ( .A(n4599), .B(n4600), .Z(n4594) );
  AND U4214 ( .A(n233), .B(n4601), .Z(n4600) );
  XOR U4215 ( .A(p_input[293]), .B(n4599), .Z(n4601) );
  XOR U4216 ( .A(n4602), .B(n4603), .Z(n4599) );
  AND U4217 ( .A(n237), .B(n4604), .Z(n4603) );
  XOR U4218 ( .A(n4605), .B(n4606), .Z(n4597) );
  AND U4219 ( .A(n241), .B(n4604), .Z(n4606) );
  XNOR U4220 ( .A(n4605), .B(n4602), .Z(n4604) );
  XOR U4221 ( .A(n4607), .B(n4608), .Z(n4602) );
  AND U4222 ( .A(n244), .B(n4609), .Z(n4608) );
  XOR U4223 ( .A(p_input[309]), .B(n4607), .Z(n4609) );
  XOR U4224 ( .A(n4610), .B(n4611), .Z(n4607) );
  AND U4225 ( .A(n248), .B(n4612), .Z(n4611) );
  XOR U4226 ( .A(n4613), .B(n4614), .Z(n4605) );
  AND U4227 ( .A(n252), .B(n4612), .Z(n4614) );
  XNOR U4228 ( .A(n4613), .B(n4610), .Z(n4612) );
  XOR U4229 ( .A(n4615), .B(n4616), .Z(n4610) );
  AND U4230 ( .A(n255), .B(n4617), .Z(n4616) );
  XOR U4231 ( .A(p_input[325]), .B(n4615), .Z(n4617) );
  XOR U4232 ( .A(n4618), .B(n4619), .Z(n4615) );
  AND U4233 ( .A(n259), .B(n4620), .Z(n4619) );
  XOR U4234 ( .A(n4621), .B(n4622), .Z(n4613) );
  AND U4235 ( .A(n263), .B(n4620), .Z(n4622) );
  XNOR U4236 ( .A(n4621), .B(n4618), .Z(n4620) );
  XOR U4237 ( .A(n4623), .B(n4624), .Z(n4618) );
  AND U4238 ( .A(n266), .B(n4625), .Z(n4624) );
  XOR U4239 ( .A(p_input[341]), .B(n4623), .Z(n4625) );
  XOR U4240 ( .A(n4626), .B(n4627), .Z(n4623) );
  AND U4241 ( .A(n270), .B(n4628), .Z(n4627) );
  XOR U4242 ( .A(n4629), .B(n4630), .Z(n4621) );
  AND U4243 ( .A(n274), .B(n4628), .Z(n4630) );
  XNOR U4244 ( .A(n4629), .B(n4626), .Z(n4628) );
  XOR U4245 ( .A(n4631), .B(n4632), .Z(n4626) );
  AND U4246 ( .A(n277), .B(n4633), .Z(n4632) );
  XOR U4247 ( .A(p_input[357]), .B(n4631), .Z(n4633) );
  XOR U4248 ( .A(n4634), .B(n4635), .Z(n4631) );
  AND U4249 ( .A(n281), .B(n4636), .Z(n4635) );
  XOR U4250 ( .A(n4637), .B(n4638), .Z(n4629) );
  AND U4251 ( .A(n285), .B(n4636), .Z(n4638) );
  XNOR U4252 ( .A(n4637), .B(n4634), .Z(n4636) );
  XOR U4253 ( .A(n4639), .B(n4640), .Z(n4634) );
  AND U4254 ( .A(n288), .B(n4641), .Z(n4640) );
  XOR U4255 ( .A(p_input[373]), .B(n4639), .Z(n4641) );
  XOR U4256 ( .A(n4642), .B(n4643), .Z(n4639) );
  AND U4257 ( .A(n292), .B(n4644), .Z(n4643) );
  XOR U4258 ( .A(n4645), .B(n4646), .Z(n4637) );
  AND U4259 ( .A(n296), .B(n4644), .Z(n4646) );
  XNOR U4260 ( .A(n4645), .B(n4642), .Z(n4644) );
  XOR U4261 ( .A(n4647), .B(n4648), .Z(n4642) );
  AND U4262 ( .A(n299), .B(n4649), .Z(n4648) );
  XOR U4263 ( .A(p_input[389]), .B(n4647), .Z(n4649) );
  XOR U4264 ( .A(n4650), .B(n4651), .Z(n4647) );
  AND U4265 ( .A(n303), .B(n4652), .Z(n4651) );
  XOR U4266 ( .A(n4653), .B(n4654), .Z(n4645) );
  AND U4267 ( .A(n307), .B(n4652), .Z(n4654) );
  XNOR U4268 ( .A(n4653), .B(n4650), .Z(n4652) );
  XOR U4269 ( .A(n4655), .B(n4656), .Z(n4650) );
  AND U4270 ( .A(n310), .B(n4657), .Z(n4656) );
  XOR U4271 ( .A(p_input[405]), .B(n4655), .Z(n4657) );
  XOR U4272 ( .A(n4658), .B(n4659), .Z(n4655) );
  AND U4273 ( .A(n314), .B(n4660), .Z(n4659) );
  XOR U4274 ( .A(n4661), .B(n4662), .Z(n4653) );
  AND U4275 ( .A(n318), .B(n4660), .Z(n4662) );
  XNOR U4276 ( .A(n4661), .B(n4658), .Z(n4660) );
  XOR U4277 ( .A(n4663), .B(n4664), .Z(n4658) );
  AND U4278 ( .A(n321), .B(n4665), .Z(n4664) );
  XOR U4279 ( .A(p_input[421]), .B(n4663), .Z(n4665) );
  XOR U4280 ( .A(n4666), .B(n4667), .Z(n4663) );
  AND U4281 ( .A(n325), .B(n4668), .Z(n4667) );
  XOR U4282 ( .A(n4669), .B(n4670), .Z(n4661) );
  AND U4283 ( .A(n329), .B(n4668), .Z(n4670) );
  XNOR U4284 ( .A(n4669), .B(n4666), .Z(n4668) );
  XOR U4285 ( .A(n4671), .B(n4672), .Z(n4666) );
  AND U4286 ( .A(n332), .B(n4673), .Z(n4672) );
  XOR U4287 ( .A(p_input[437]), .B(n4671), .Z(n4673) );
  XOR U4288 ( .A(n4674), .B(n4675), .Z(n4671) );
  AND U4289 ( .A(n336), .B(n4676), .Z(n4675) );
  XOR U4290 ( .A(n4677), .B(n4678), .Z(n4669) );
  AND U4291 ( .A(n340), .B(n4676), .Z(n4678) );
  XNOR U4292 ( .A(n4677), .B(n4674), .Z(n4676) );
  XOR U4293 ( .A(n4679), .B(n4680), .Z(n4674) );
  AND U4294 ( .A(n343), .B(n4681), .Z(n4680) );
  XOR U4295 ( .A(p_input[453]), .B(n4679), .Z(n4681) );
  XOR U4296 ( .A(n4682), .B(n4683), .Z(n4679) );
  AND U4297 ( .A(n347), .B(n4684), .Z(n4683) );
  XOR U4298 ( .A(n4685), .B(n4686), .Z(n4677) );
  AND U4299 ( .A(n351), .B(n4684), .Z(n4686) );
  XNOR U4300 ( .A(n4685), .B(n4682), .Z(n4684) );
  XOR U4301 ( .A(n4687), .B(n4688), .Z(n4682) );
  AND U4302 ( .A(n354), .B(n4689), .Z(n4688) );
  XOR U4303 ( .A(p_input[469]), .B(n4687), .Z(n4689) );
  XOR U4304 ( .A(n4690), .B(n4691), .Z(n4687) );
  AND U4305 ( .A(n358), .B(n4692), .Z(n4691) );
  XOR U4306 ( .A(n4693), .B(n4694), .Z(n4685) );
  AND U4307 ( .A(n362), .B(n4692), .Z(n4694) );
  XNOR U4308 ( .A(n4693), .B(n4690), .Z(n4692) );
  XOR U4309 ( .A(n4695), .B(n4696), .Z(n4690) );
  AND U4310 ( .A(n365), .B(n4697), .Z(n4696) );
  XOR U4311 ( .A(p_input[485]), .B(n4695), .Z(n4697) );
  XOR U4312 ( .A(n4698), .B(n4699), .Z(n4695) );
  AND U4313 ( .A(n369), .B(n4700), .Z(n4699) );
  XOR U4314 ( .A(n4701), .B(n4702), .Z(n4693) );
  AND U4315 ( .A(n373), .B(n4700), .Z(n4702) );
  XNOR U4316 ( .A(n4701), .B(n4698), .Z(n4700) );
  XOR U4317 ( .A(n4703), .B(n4704), .Z(n4698) );
  AND U4318 ( .A(n376), .B(n4705), .Z(n4704) );
  XOR U4319 ( .A(p_input[501]), .B(n4703), .Z(n4705) );
  XOR U4320 ( .A(n4706), .B(n4707), .Z(n4703) );
  AND U4321 ( .A(n380), .B(n4708), .Z(n4707) );
  XOR U4322 ( .A(n4709), .B(n4710), .Z(n4701) );
  AND U4323 ( .A(n384), .B(n4708), .Z(n4710) );
  XNOR U4324 ( .A(n4709), .B(n4706), .Z(n4708) );
  XOR U4325 ( .A(n4711), .B(n4712), .Z(n4706) );
  AND U4326 ( .A(n387), .B(n4713), .Z(n4712) );
  XOR U4327 ( .A(p_input[517]), .B(n4711), .Z(n4713) );
  XOR U4328 ( .A(n4714), .B(n4715), .Z(n4711) );
  AND U4329 ( .A(n391), .B(n4716), .Z(n4715) );
  XOR U4330 ( .A(n4717), .B(n4718), .Z(n4709) );
  AND U4331 ( .A(n395), .B(n4716), .Z(n4718) );
  XNOR U4332 ( .A(n4717), .B(n4714), .Z(n4716) );
  XOR U4333 ( .A(n4719), .B(n4720), .Z(n4714) );
  AND U4334 ( .A(n398), .B(n4721), .Z(n4720) );
  XOR U4335 ( .A(p_input[533]), .B(n4719), .Z(n4721) );
  XOR U4336 ( .A(n4722), .B(n4723), .Z(n4719) );
  AND U4337 ( .A(n402), .B(n4724), .Z(n4723) );
  XOR U4338 ( .A(n4725), .B(n4726), .Z(n4717) );
  AND U4339 ( .A(n406), .B(n4724), .Z(n4726) );
  XNOR U4340 ( .A(n4725), .B(n4722), .Z(n4724) );
  XOR U4341 ( .A(n4727), .B(n4728), .Z(n4722) );
  AND U4342 ( .A(n409), .B(n4729), .Z(n4728) );
  XOR U4343 ( .A(p_input[549]), .B(n4727), .Z(n4729) );
  XOR U4344 ( .A(n4730), .B(n4731), .Z(n4727) );
  AND U4345 ( .A(n413), .B(n4732), .Z(n4731) );
  XOR U4346 ( .A(n4733), .B(n4734), .Z(n4725) );
  AND U4347 ( .A(n417), .B(n4732), .Z(n4734) );
  XNOR U4348 ( .A(n4733), .B(n4730), .Z(n4732) );
  XOR U4349 ( .A(n4735), .B(n4736), .Z(n4730) );
  AND U4350 ( .A(n420), .B(n4737), .Z(n4736) );
  XOR U4351 ( .A(p_input[565]), .B(n4735), .Z(n4737) );
  XOR U4352 ( .A(n4738), .B(n4739), .Z(n4735) );
  AND U4353 ( .A(n424), .B(n4740), .Z(n4739) );
  XOR U4354 ( .A(n4741), .B(n4742), .Z(n4733) );
  AND U4355 ( .A(n428), .B(n4740), .Z(n4742) );
  XNOR U4356 ( .A(n4741), .B(n4738), .Z(n4740) );
  XOR U4357 ( .A(n4743), .B(n4744), .Z(n4738) );
  AND U4358 ( .A(n431), .B(n4745), .Z(n4744) );
  XOR U4359 ( .A(p_input[581]), .B(n4743), .Z(n4745) );
  XOR U4360 ( .A(n4746), .B(n4747), .Z(n4743) );
  AND U4361 ( .A(n435), .B(n4748), .Z(n4747) );
  XOR U4362 ( .A(n4749), .B(n4750), .Z(n4741) );
  AND U4363 ( .A(n439), .B(n4748), .Z(n4750) );
  XNOR U4364 ( .A(n4749), .B(n4746), .Z(n4748) );
  XOR U4365 ( .A(n4751), .B(n4752), .Z(n4746) );
  AND U4366 ( .A(n442), .B(n4753), .Z(n4752) );
  XOR U4367 ( .A(p_input[597]), .B(n4751), .Z(n4753) );
  XOR U4368 ( .A(n4754), .B(n4755), .Z(n4751) );
  AND U4369 ( .A(n446), .B(n4756), .Z(n4755) );
  XOR U4370 ( .A(n4757), .B(n4758), .Z(n4749) );
  AND U4371 ( .A(n450), .B(n4756), .Z(n4758) );
  XNOR U4372 ( .A(n4757), .B(n4754), .Z(n4756) );
  XOR U4373 ( .A(n4759), .B(n4760), .Z(n4754) );
  AND U4374 ( .A(n453), .B(n4761), .Z(n4760) );
  XOR U4375 ( .A(p_input[613]), .B(n4759), .Z(n4761) );
  XOR U4376 ( .A(n4762), .B(n4763), .Z(n4759) );
  AND U4377 ( .A(n457), .B(n4764), .Z(n4763) );
  XOR U4378 ( .A(n4765), .B(n4766), .Z(n4757) );
  AND U4379 ( .A(n461), .B(n4764), .Z(n4766) );
  XNOR U4380 ( .A(n4765), .B(n4762), .Z(n4764) );
  XOR U4381 ( .A(n4767), .B(n4768), .Z(n4762) );
  AND U4382 ( .A(n464), .B(n4769), .Z(n4768) );
  XOR U4383 ( .A(p_input[629]), .B(n4767), .Z(n4769) );
  XOR U4384 ( .A(n4770), .B(n4771), .Z(n4767) );
  AND U4385 ( .A(n468), .B(n4772), .Z(n4771) );
  XOR U4386 ( .A(n4773), .B(n4774), .Z(n4765) );
  AND U4387 ( .A(n472), .B(n4772), .Z(n4774) );
  XNOR U4388 ( .A(n4773), .B(n4770), .Z(n4772) );
  XOR U4389 ( .A(n4775), .B(n4776), .Z(n4770) );
  AND U4390 ( .A(n475), .B(n4777), .Z(n4776) );
  XOR U4391 ( .A(p_input[645]), .B(n4775), .Z(n4777) );
  XOR U4392 ( .A(n4778), .B(n4779), .Z(n4775) );
  AND U4393 ( .A(n479), .B(n4780), .Z(n4779) );
  XOR U4394 ( .A(n4781), .B(n4782), .Z(n4773) );
  AND U4395 ( .A(n483), .B(n4780), .Z(n4782) );
  XNOR U4396 ( .A(n4781), .B(n4778), .Z(n4780) );
  XOR U4397 ( .A(n4783), .B(n4784), .Z(n4778) );
  AND U4398 ( .A(n486), .B(n4785), .Z(n4784) );
  XOR U4399 ( .A(p_input[661]), .B(n4783), .Z(n4785) );
  XOR U4400 ( .A(n4786), .B(n4787), .Z(n4783) );
  AND U4401 ( .A(n490), .B(n4788), .Z(n4787) );
  XOR U4402 ( .A(n4789), .B(n4790), .Z(n4781) );
  AND U4403 ( .A(n494), .B(n4788), .Z(n4790) );
  XNOR U4404 ( .A(n4789), .B(n4786), .Z(n4788) );
  XOR U4405 ( .A(n4791), .B(n4792), .Z(n4786) );
  AND U4406 ( .A(n497), .B(n4793), .Z(n4792) );
  XOR U4407 ( .A(p_input[677]), .B(n4791), .Z(n4793) );
  XOR U4408 ( .A(n4794), .B(n4795), .Z(n4791) );
  AND U4409 ( .A(n501), .B(n4796), .Z(n4795) );
  XOR U4410 ( .A(n4797), .B(n4798), .Z(n4789) );
  AND U4411 ( .A(n505), .B(n4796), .Z(n4798) );
  XNOR U4412 ( .A(n4797), .B(n4794), .Z(n4796) );
  XOR U4413 ( .A(n4799), .B(n4800), .Z(n4794) );
  AND U4414 ( .A(n508), .B(n4801), .Z(n4800) );
  XOR U4415 ( .A(p_input[693]), .B(n4799), .Z(n4801) );
  XOR U4416 ( .A(n4802), .B(n4803), .Z(n4799) );
  AND U4417 ( .A(n512), .B(n4804), .Z(n4803) );
  XOR U4418 ( .A(n4805), .B(n4806), .Z(n4797) );
  AND U4419 ( .A(n516), .B(n4804), .Z(n4806) );
  XNOR U4420 ( .A(n4805), .B(n4802), .Z(n4804) );
  XOR U4421 ( .A(n4807), .B(n4808), .Z(n4802) );
  AND U4422 ( .A(n519), .B(n4809), .Z(n4808) );
  XOR U4423 ( .A(p_input[709]), .B(n4807), .Z(n4809) );
  XOR U4424 ( .A(n4810), .B(n4811), .Z(n4807) );
  AND U4425 ( .A(n523), .B(n4812), .Z(n4811) );
  XOR U4426 ( .A(n4813), .B(n4814), .Z(n4805) );
  AND U4427 ( .A(n527), .B(n4812), .Z(n4814) );
  XNOR U4428 ( .A(n4813), .B(n4810), .Z(n4812) );
  XOR U4429 ( .A(n4815), .B(n4816), .Z(n4810) );
  AND U4430 ( .A(n530), .B(n4817), .Z(n4816) );
  XOR U4431 ( .A(p_input[725]), .B(n4815), .Z(n4817) );
  XOR U4432 ( .A(n4818), .B(n4819), .Z(n4815) );
  AND U4433 ( .A(n534), .B(n4820), .Z(n4819) );
  XOR U4434 ( .A(n4821), .B(n4822), .Z(n4813) );
  AND U4435 ( .A(n538), .B(n4820), .Z(n4822) );
  XNOR U4436 ( .A(n4821), .B(n4818), .Z(n4820) );
  XOR U4437 ( .A(n4823), .B(n4824), .Z(n4818) );
  AND U4438 ( .A(n541), .B(n4825), .Z(n4824) );
  XOR U4439 ( .A(p_input[741]), .B(n4823), .Z(n4825) );
  XOR U4440 ( .A(n4826), .B(n4827), .Z(n4823) );
  AND U4441 ( .A(n545), .B(n4828), .Z(n4827) );
  XOR U4442 ( .A(n4829), .B(n4830), .Z(n4821) );
  AND U4443 ( .A(n549), .B(n4828), .Z(n4830) );
  XNOR U4444 ( .A(n4829), .B(n4826), .Z(n4828) );
  XOR U4445 ( .A(n4831), .B(n4832), .Z(n4826) );
  AND U4446 ( .A(n552), .B(n4833), .Z(n4832) );
  XOR U4447 ( .A(p_input[757]), .B(n4831), .Z(n4833) );
  XOR U4448 ( .A(n4834), .B(n4835), .Z(n4831) );
  AND U4449 ( .A(n556), .B(n4836), .Z(n4835) );
  XOR U4450 ( .A(n4837), .B(n4838), .Z(n4829) );
  AND U4451 ( .A(n560), .B(n4836), .Z(n4838) );
  XNOR U4452 ( .A(n4837), .B(n4834), .Z(n4836) );
  XOR U4453 ( .A(n4839), .B(n4840), .Z(n4834) );
  AND U4454 ( .A(n563), .B(n4841), .Z(n4840) );
  XOR U4455 ( .A(p_input[773]), .B(n4839), .Z(n4841) );
  XOR U4456 ( .A(n4842), .B(n4843), .Z(n4839) );
  AND U4457 ( .A(n567), .B(n4844), .Z(n4843) );
  XOR U4458 ( .A(n4845), .B(n4846), .Z(n4837) );
  AND U4459 ( .A(n571), .B(n4844), .Z(n4846) );
  XNOR U4460 ( .A(n4845), .B(n4842), .Z(n4844) );
  XOR U4461 ( .A(n4847), .B(n4848), .Z(n4842) );
  AND U4462 ( .A(n574), .B(n4849), .Z(n4848) );
  XOR U4463 ( .A(p_input[789]), .B(n4847), .Z(n4849) );
  XOR U4464 ( .A(n4850), .B(n4851), .Z(n4847) );
  AND U4465 ( .A(n578), .B(n4852), .Z(n4851) );
  XOR U4466 ( .A(n4853), .B(n4854), .Z(n4845) );
  AND U4467 ( .A(n582), .B(n4852), .Z(n4854) );
  XNOR U4468 ( .A(n4853), .B(n4850), .Z(n4852) );
  XOR U4469 ( .A(n4855), .B(n4856), .Z(n4850) );
  AND U4470 ( .A(n585), .B(n4857), .Z(n4856) );
  XOR U4471 ( .A(p_input[805]), .B(n4855), .Z(n4857) );
  XOR U4472 ( .A(n4858), .B(n4859), .Z(n4855) );
  AND U4473 ( .A(n589), .B(n4860), .Z(n4859) );
  XOR U4474 ( .A(n4861), .B(n4862), .Z(n4853) );
  AND U4475 ( .A(n593), .B(n4860), .Z(n4862) );
  XNOR U4476 ( .A(n4861), .B(n4858), .Z(n4860) );
  XOR U4477 ( .A(n4863), .B(n4864), .Z(n4858) );
  AND U4478 ( .A(n596), .B(n4865), .Z(n4864) );
  XOR U4479 ( .A(p_input[821]), .B(n4863), .Z(n4865) );
  XOR U4480 ( .A(n4866), .B(n4867), .Z(n4863) );
  AND U4481 ( .A(n600), .B(n4868), .Z(n4867) );
  XOR U4482 ( .A(n4869), .B(n4870), .Z(n4861) );
  AND U4483 ( .A(n604), .B(n4868), .Z(n4870) );
  XNOR U4484 ( .A(n4869), .B(n4866), .Z(n4868) );
  XOR U4485 ( .A(n4871), .B(n4872), .Z(n4866) );
  AND U4486 ( .A(n607), .B(n4873), .Z(n4872) );
  XOR U4487 ( .A(p_input[837]), .B(n4871), .Z(n4873) );
  XOR U4488 ( .A(n4874), .B(n4875), .Z(n4871) );
  AND U4489 ( .A(n611), .B(n4876), .Z(n4875) );
  XOR U4490 ( .A(n4877), .B(n4878), .Z(n4869) );
  AND U4491 ( .A(n615), .B(n4876), .Z(n4878) );
  XNOR U4492 ( .A(n4877), .B(n4874), .Z(n4876) );
  XOR U4493 ( .A(n4879), .B(n4880), .Z(n4874) );
  AND U4494 ( .A(n618), .B(n4881), .Z(n4880) );
  XOR U4495 ( .A(p_input[853]), .B(n4879), .Z(n4881) );
  XOR U4496 ( .A(n4882), .B(n4883), .Z(n4879) );
  AND U4497 ( .A(n622), .B(n4884), .Z(n4883) );
  XOR U4498 ( .A(n4885), .B(n4886), .Z(n4877) );
  AND U4499 ( .A(n626), .B(n4884), .Z(n4886) );
  XNOR U4500 ( .A(n4885), .B(n4882), .Z(n4884) );
  XOR U4501 ( .A(n4887), .B(n4888), .Z(n4882) );
  AND U4502 ( .A(n629), .B(n4889), .Z(n4888) );
  XOR U4503 ( .A(p_input[869]), .B(n4887), .Z(n4889) );
  XOR U4504 ( .A(n4890), .B(n4891), .Z(n4887) );
  AND U4505 ( .A(n633), .B(n4892), .Z(n4891) );
  XOR U4506 ( .A(n4893), .B(n4894), .Z(n4885) );
  AND U4507 ( .A(n637), .B(n4892), .Z(n4894) );
  XNOR U4508 ( .A(n4893), .B(n4890), .Z(n4892) );
  XOR U4509 ( .A(n4895), .B(n4896), .Z(n4890) );
  AND U4510 ( .A(n640), .B(n4897), .Z(n4896) );
  XOR U4511 ( .A(p_input[885]), .B(n4895), .Z(n4897) );
  XOR U4512 ( .A(n4898), .B(n4899), .Z(n4895) );
  AND U4513 ( .A(n644), .B(n4900), .Z(n4899) );
  XOR U4514 ( .A(n4901), .B(n4902), .Z(n4893) );
  AND U4515 ( .A(n648), .B(n4900), .Z(n4902) );
  XNOR U4516 ( .A(n4901), .B(n4898), .Z(n4900) );
  XOR U4517 ( .A(n4903), .B(n4904), .Z(n4898) );
  AND U4518 ( .A(n651), .B(n4905), .Z(n4904) );
  XOR U4519 ( .A(p_input[901]), .B(n4903), .Z(n4905) );
  XOR U4520 ( .A(n4906), .B(n4907), .Z(n4903) );
  AND U4521 ( .A(n655), .B(n4908), .Z(n4907) );
  XOR U4522 ( .A(n4909), .B(n4910), .Z(n4901) );
  AND U4523 ( .A(n659), .B(n4908), .Z(n4910) );
  XNOR U4524 ( .A(n4909), .B(n4906), .Z(n4908) );
  XOR U4525 ( .A(n4911), .B(n4912), .Z(n4906) );
  AND U4526 ( .A(n662), .B(n4913), .Z(n4912) );
  XOR U4527 ( .A(p_input[917]), .B(n4911), .Z(n4913) );
  XOR U4528 ( .A(n4914), .B(n4915), .Z(n4911) );
  AND U4529 ( .A(n666), .B(n4916), .Z(n4915) );
  XOR U4530 ( .A(n4917), .B(n4918), .Z(n4909) );
  AND U4531 ( .A(n670), .B(n4916), .Z(n4918) );
  XNOR U4532 ( .A(n4917), .B(n4914), .Z(n4916) );
  XOR U4533 ( .A(n4919), .B(n4920), .Z(n4914) );
  AND U4534 ( .A(n673), .B(n4921), .Z(n4920) );
  XOR U4535 ( .A(p_input[933]), .B(n4919), .Z(n4921) );
  XOR U4536 ( .A(n4922), .B(n4923), .Z(n4919) );
  AND U4537 ( .A(n677), .B(n4924), .Z(n4923) );
  XOR U4538 ( .A(n4925), .B(n4926), .Z(n4917) );
  AND U4539 ( .A(n681), .B(n4924), .Z(n4926) );
  XNOR U4540 ( .A(n4925), .B(n4922), .Z(n4924) );
  XOR U4541 ( .A(n4927), .B(n4928), .Z(n4922) );
  AND U4542 ( .A(n684), .B(n4929), .Z(n4928) );
  XOR U4543 ( .A(p_input[949]), .B(n4927), .Z(n4929) );
  XOR U4544 ( .A(n4930), .B(n4931), .Z(n4927) );
  AND U4545 ( .A(n688), .B(n4932), .Z(n4931) );
  XOR U4546 ( .A(n4933), .B(n4934), .Z(n4925) );
  AND U4547 ( .A(n692), .B(n4932), .Z(n4934) );
  XNOR U4548 ( .A(n4933), .B(n4930), .Z(n4932) );
  XOR U4549 ( .A(n4935), .B(n4936), .Z(n4930) );
  AND U4550 ( .A(n695), .B(n4937), .Z(n4936) );
  XOR U4551 ( .A(p_input[965]), .B(n4935), .Z(n4937) );
  XOR U4552 ( .A(n4938), .B(n4939), .Z(n4935) );
  AND U4553 ( .A(n699), .B(n4940), .Z(n4939) );
  XOR U4554 ( .A(n4941), .B(n4942), .Z(n4933) );
  AND U4555 ( .A(n703), .B(n4940), .Z(n4942) );
  XNOR U4556 ( .A(n4941), .B(n4938), .Z(n4940) );
  XOR U4557 ( .A(n4943), .B(n4944), .Z(n4938) );
  AND U4558 ( .A(n706), .B(n4945), .Z(n4944) );
  XOR U4559 ( .A(p_input[981]), .B(n4943), .Z(n4945) );
  XOR U4560 ( .A(n4946), .B(n4947), .Z(n4943) );
  AND U4561 ( .A(n710), .B(n4948), .Z(n4947) );
  XOR U4562 ( .A(n4949), .B(n4950), .Z(n4941) );
  AND U4563 ( .A(n714), .B(n4948), .Z(n4950) );
  XNOR U4564 ( .A(n4949), .B(n4946), .Z(n4948) );
  XOR U4565 ( .A(n4951), .B(n4952), .Z(n4946) );
  AND U4566 ( .A(n717), .B(n4953), .Z(n4952) );
  XOR U4567 ( .A(p_input[997]), .B(n4951), .Z(n4953) );
  XOR U4568 ( .A(n4954), .B(n4955), .Z(n4951) );
  AND U4569 ( .A(n721), .B(n4956), .Z(n4955) );
  XOR U4570 ( .A(n4957), .B(n4958), .Z(n4949) );
  AND U4571 ( .A(n725), .B(n4956), .Z(n4958) );
  XNOR U4572 ( .A(n4957), .B(n4954), .Z(n4956) );
  XOR U4573 ( .A(n4959), .B(n4960), .Z(n4954) );
  AND U4574 ( .A(n728), .B(n4961), .Z(n4960) );
  XOR U4575 ( .A(p_input[1013]), .B(n4959), .Z(n4961) );
  XOR U4576 ( .A(n4962), .B(n4963), .Z(n4959) );
  AND U4577 ( .A(n732), .B(n4964), .Z(n4963) );
  XOR U4578 ( .A(n4965), .B(n4966), .Z(n4957) );
  AND U4579 ( .A(n736), .B(n4964), .Z(n4966) );
  XNOR U4580 ( .A(n4965), .B(n4962), .Z(n4964) );
  XOR U4581 ( .A(n4967), .B(n4968), .Z(n4962) );
  AND U4582 ( .A(n739), .B(n4969), .Z(n4968) );
  XOR U4583 ( .A(p_input[1029]), .B(n4967), .Z(n4969) );
  XOR U4584 ( .A(n4970), .B(n4971), .Z(n4967) );
  AND U4585 ( .A(n743), .B(n4972), .Z(n4971) );
  XOR U4586 ( .A(n4973), .B(n4974), .Z(n4965) );
  AND U4587 ( .A(n747), .B(n4972), .Z(n4974) );
  XNOR U4588 ( .A(n4973), .B(n4970), .Z(n4972) );
  XOR U4589 ( .A(n4975), .B(n4976), .Z(n4970) );
  AND U4590 ( .A(n750), .B(n4977), .Z(n4976) );
  XOR U4591 ( .A(p_input[1045]), .B(n4975), .Z(n4977) );
  XOR U4592 ( .A(n4978), .B(n4979), .Z(n4975) );
  AND U4593 ( .A(n754), .B(n4980), .Z(n4979) );
  XOR U4594 ( .A(n4981), .B(n4982), .Z(n4973) );
  AND U4595 ( .A(n758), .B(n4980), .Z(n4982) );
  XNOR U4596 ( .A(n4981), .B(n4978), .Z(n4980) );
  XOR U4597 ( .A(n4983), .B(n4984), .Z(n4978) );
  AND U4598 ( .A(n761), .B(n4985), .Z(n4984) );
  XOR U4599 ( .A(p_input[1061]), .B(n4983), .Z(n4985) );
  XOR U4600 ( .A(n4986), .B(n4987), .Z(n4983) );
  AND U4601 ( .A(n765), .B(n4988), .Z(n4987) );
  XOR U4602 ( .A(n4989), .B(n4990), .Z(n4981) );
  AND U4603 ( .A(n769), .B(n4988), .Z(n4990) );
  XNOR U4604 ( .A(n4989), .B(n4986), .Z(n4988) );
  XOR U4605 ( .A(n4991), .B(n4992), .Z(n4986) );
  AND U4606 ( .A(n772), .B(n4993), .Z(n4992) );
  XOR U4607 ( .A(p_input[1077]), .B(n4991), .Z(n4993) );
  XOR U4608 ( .A(n4994), .B(n4995), .Z(n4991) );
  AND U4609 ( .A(n776), .B(n4996), .Z(n4995) );
  XOR U4610 ( .A(n4997), .B(n4998), .Z(n4989) );
  AND U4611 ( .A(n780), .B(n4996), .Z(n4998) );
  XNOR U4612 ( .A(n4997), .B(n4994), .Z(n4996) );
  XOR U4613 ( .A(n4999), .B(n5000), .Z(n4994) );
  AND U4614 ( .A(n783), .B(n5001), .Z(n5000) );
  XOR U4615 ( .A(p_input[1093]), .B(n4999), .Z(n5001) );
  XOR U4616 ( .A(n5002), .B(n5003), .Z(n4999) );
  AND U4617 ( .A(n787), .B(n5004), .Z(n5003) );
  XOR U4618 ( .A(n5005), .B(n5006), .Z(n4997) );
  AND U4619 ( .A(n791), .B(n5004), .Z(n5006) );
  XNOR U4620 ( .A(n5005), .B(n5002), .Z(n5004) );
  XOR U4621 ( .A(n5007), .B(n5008), .Z(n5002) );
  AND U4622 ( .A(n794), .B(n5009), .Z(n5008) );
  XOR U4623 ( .A(p_input[1109]), .B(n5007), .Z(n5009) );
  XOR U4624 ( .A(n5010), .B(n5011), .Z(n5007) );
  AND U4625 ( .A(n798), .B(n5012), .Z(n5011) );
  XOR U4626 ( .A(n5013), .B(n5014), .Z(n5005) );
  AND U4627 ( .A(n802), .B(n5012), .Z(n5014) );
  XNOR U4628 ( .A(n5013), .B(n5010), .Z(n5012) );
  XOR U4629 ( .A(n5015), .B(n5016), .Z(n5010) );
  AND U4630 ( .A(n805), .B(n5017), .Z(n5016) );
  XOR U4631 ( .A(p_input[1125]), .B(n5015), .Z(n5017) );
  XOR U4632 ( .A(n5018), .B(n5019), .Z(n5015) );
  AND U4633 ( .A(n809), .B(n5020), .Z(n5019) );
  XOR U4634 ( .A(n5021), .B(n5022), .Z(n5013) );
  AND U4635 ( .A(n813), .B(n5020), .Z(n5022) );
  XNOR U4636 ( .A(n5021), .B(n5018), .Z(n5020) );
  XOR U4637 ( .A(n5023), .B(n5024), .Z(n5018) );
  AND U4638 ( .A(n816), .B(n5025), .Z(n5024) );
  XOR U4639 ( .A(p_input[1141]), .B(n5023), .Z(n5025) );
  XOR U4640 ( .A(n5026), .B(n5027), .Z(n5023) );
  AND U4641 ( .A(n820), .B(n5028), .Z(n5027) );
  XOR U4642 ( .A(n5029), .B(n5030), .Z(n5021) );
  AND U4643 ( .A(n824), .B(n5028), .Z(n5030) );
  XNOR U4644 ( .A(n5029), .B(n5026), .Z(n5028) );
  XOR U4645 ( .A(n5031), .B(n5032), .Z(n5026) );
  AND U4646 ( .A(n827), .B(n5033), .Z(n5032) );
  XOR U4647 ( .A(p_input[1157]), .B(n5031), .Z(n5033) );
  XOR U4648 ( .A(n5034), .B(n5035), .Z(n5031) );
  AND U4649 ( .A(n831), .B(n5036), .Z(n5035) );
  XOR U4650 ( .A(n5037), .B(n5038), .Z(n5029) );
  AND U4651 ( .A(n835), .B(n5036), .Z(n5038) );
  XNOR U4652 ( .A(n5037), .B(n5034), .Z(n5036) );
  XOR U4653 ( .A(n5039), .B(n5040), .Z(n5034) );
  AND U4654 ( .A(n838), .B(n5041), .Z(n5040) );
  XOR U4655 ( .A(p_input[1173]), .B(n5039), .Z(n5041) );
  XOR U4656 ( .A(n5042), .B(n5043), .Z(n5039) );
  AND U4657 ( .A(n842), .B(n5044), .Z(n5043) );
  XOR U4658 ( .A(n5045), .B(n5046), .Z(n5037) );
  AND U4659 ( .A(n846), .B(n5044), .Z(n5046) );
  XNOR U4660 ( .A(n5045), .B(n5042), .Z(n5044) );
  XOR U4661 ( .A(n5047), .B(n5048), .Z(n5042) );
  AND U4662 ( .A(n849), .B(n5049), .Z(n5048) );
  XOR U4663 ( .A(p_input[1189]), .B(n5047), .Z(n5049) );
  XOR U4664 ( .A(n5050), .B(n5051), .Z(n5047) );
  AND U4665 ( .A(n853), .B(n5052), .Z(n5051) );
  XOR U4666 ( .A(n5053), .B(n5054), .Z(n5045) );
  AND U4667 ( .A(n857), .B(n5052), .Z(n5054) );
  XNOR U4668 ( .A(n5053), .B(n5050), .Z(n5052) );
  XOR U4669 ( .A(n5055), .B(n5056), .Z(n5050) );
  AND U4670 ( .A(n860), .B(n5057), .Z(n5056) );
  XOR U4671 ( .A(p_input[1205]), .B(n5055), .Z(n5057) );
  XOR U4672 ( .A(n5058), .B(n5059), .Z(n5055) );
  AND U4673 ( .A(n864), .B(n5060), .Z(n5059) );
  XOR U4674 ( .A(n5061), .B(n5062), .Z(n5053) );
  AND U4675 ( .A(n868), .B(n5060), .Z(n5062) );
  XNOR U4676 ( .A(n5061), .B(n5058), .Z(n5060) );
  XOR U4677 ( .A(n5063), .B(n5064), .Z(n5058) );
  AND U4678 ( .A(n871), .B(n5065), .Z(n5064) );
  XOR U4679 ( .A(p_input[1221]), .B(n5063), .Z(n5065) );
  XOR U4680 ( .A(n5066), .B(n5067), .Z(n5063) );
  AND U4681 ( .A(n875), .B(n5068), .Z(n5067) );
  XOR U4682 ( .A(n5069), .B(n5070), .Z(n5061) );
  AND U4683 ( .A(n879), .B(n5068), .Z(n5070) );
  XNOR U4684 ( .A(n5069), .B(n5066), .Z(n5068) );
  XOR U4685 ( .A(n5071), .B(n5072), .Z(n5066) );
  AND U4686 ( .A(n882), .B(n5073), .Z(n5072) );
  XOR U4687 ( .A(p_input[1237]), .B(n5071), .Z(n5073) );
  XOR U4688 ( .A(n5074), .B(n5075), .Z(n5071) );
  AND U4689 ( .A(n886), .B(n5076), .Z(n5075) );
  XOR U4690 ( .A(n5077), .B(n5078), .Z(n5069) );
  AND U4691 ( .A(n890), .B(n5076), .Z(n5078) );
  XNOR U4692 ( .A(n5077), .B(n5074), .Z(n5076) );
  XOR U4693 ( .A(n5079), .B(n5080), .Z(n5074) );
  AND U4694 ( .A(n893), .B(n5081), .Z(n5080) );
  XOR U4695 ( .A(p_input[1253]), .B(n5079), .Z(n5081) );
  XOR U4696 ( .A(n5082), .B(n5083), .Z(n5079) );
  AND U4697 ( .A(n897), .B(n5084), .Z(n5083) );
  XOR U4698 ( .A(n5085), .B(n5086), .Z(n5077) );
  AND U4699 ( .A(n901), .B(n5084), .Z(n5086) );
  XNOR U4700 ( .A(n5085), .B(n5082), .Z(n5084) );
  XOR U4701 ( .A(n5087), .B(n5088), .Z(n5082) );
  AND U4702 ( .A(n904), .B(n5089), .Z(n5088) );
  XOR U4703 ( .A(p_input[1269]), .B(n5087), .Z(n5089) );
  XOR U4704 ( .A(n5090), .B(n5091), .Z(n5087) );
  AND U4705 ( .A(n908), .B(n5092), .Z(n5091) );
  XOR U4706 ( .A(n5093), .B(n5094), .Z(n5085) );
  AND U4707 ( .A(n912), .B(n5092), .Z(n5094) );
  XNOR U4708 ( .A(n5093), .B(n5090), .Z(n5092) );
  XOR U4709 ( .A(n5095), .B(n5096), .Z(n5090) );
  AND U4710 ( .A(n915), .B(n5097), .Z(n5096) );
  XOR U4711 ( .A(p_input[1285]), .B(n5095), .Z(n5097) );
  XOR U4712 ( .A(n5098), .B(n5099), .Z(n5095) );
  AND U4713 ( .A(n919), .B(n5100), .Z(n5099) );
  XOR U4714 ( .A(n5101), .B(n5102), .Z(n5093) );
  AND U4715 ( .A(n923), .B(n5100), .Z(n5102) );
  XNOR U4716 ( .A(n5101), .B(n5098), .Z(n5100) );
  XOR U4717 ( .A(n5103), .B(n5104), .Z(n5098) );
  AND U4718 ( .A(n926), .B(n5105), .Z(n5104) );
  XOR U4719 ( .A(p_input[1301]), .B(n5103), .Z(n5105) );
  XOR U4720 ( .A(n5106), .B(n5107), .Z(n5103) );
  AND U4721 ( .A(n930), .B(n5108), .Z(n5107) );
  XOR U4722 ( .A(n5109), .B(n5110), .Z(n5101) );
  AND U4723 ( .A(n934), .B(n5108), .Z(n5110) );
  XNOR U4724 ( .A(n5109), .B(n5106), .Z(n5108) );
  XOR U4725 ( .A(n5111), .B(n5112), .Z(n5106) );
  AND U4726 ( .A(n937), .B(n5113), .Z(n5112) );
  XOR U4727 ( .A(p_input[1317]), .B(n5111), .Z(n5113) );
  XOR U4728 ( .A(n5114), .B(n5115), .Z(n5111) );
  AND U4729 ( .A(n941), .B(n5116), .Z(n5115) );
  XOR U4730 ( .A(n5117), .B(n5118), .Z(n5109) );
  AND U4731 ( .A(n945), .B(n5116), .Z(n5118) );
  XNOR U4732 ( .A(n5117), .B(n5114), .Z(n5116) );
  XOR U4733 ( .A(n5119), .B(n5120), .Z(n5114) );
  AND U4734 ( .A(n948), .B(n5121), .Z(n5120) );
  XOR U4735 ( .A(p_input[1333]), .B(n5119), .Z(n5121) );
  XOR U4736 ( .A(n5122), .B(n5123), .Z(n5119) );
  AND U4737 ( .A(n952), .B(n5124), .Z(n5123) );
  XOR U4738 ( .A(n5125), .B(n5126), .Z(n5117) );
  AND U4739 ( .A(n956), .B(n5124), .Z(n5126) );
  XNOR U4740 ( .A(n5125), .B(n5122), .Z(n5124) );
  XOR U4741 ( .A(n5127), .B(n5128), .Z(n5122) );
  AND U4742 ( .A(n959), .B(n5129), .Z(n5128) );
  XOR U4743 ( .A(p_input[1349]), .B(n5127), .Z(n5129) );
  XOR U4744 ( .A(n5130), .B(n5131), .Z(n5127) );
  AND U4745 ( .A(n963), .B(n5132), .Z(n5131) );
  XOR U4746 ( .A(n5133), .B(n5134), .Z(n5125) );
  AND U4747 ( .A(n967), .B(n5132), .Z(n5134) );
  XNOR U4748 ( .A(n5133), .B(n5130), .Z(n5132) );
  XOR U4749 ( .A(n5135), .B(n5136), .Z(n5130) );
  AND U4750 ( .A(n970), .B(n5137), .Z(n5136) );
  XOR U4751 ( .A(p_input[1365]), .B(n5135), .Z(n5137) );
  XOR U4752 ( .A(n5138), .B(n5139), .Z(n5135) );
  AND U4753 ( .A(n974), .B(n5140), .Z(n5139) );
  XOR U4754 ( .A(n5141), .B(n5142), .Z(n5133) );
  AND U4755 ( .A(n978), .B(n5140), .Z(n5142) );
  XNOR U4756 ( .A(n5141), .B(n5138), .Z(n5140) );
  XOR U4757 ( .A(n5143), .B(n5144), .Z(n5138) );
  AND U4758 ( .A(n981), .B(n5145), .Z(n5144) );
  XOR U4759 ( .A(p_input[1381]), .B(n5143), .Z(n5145) );
  XOR U4760 ( .A(n5146), .B(n5147), .Z(n5143) );
  AND U4761 ( .A(n985), .B(n5148), .Z(n5147) );
  XOR U4762 ( .A(n5149), .B(n5150), .Z(n5141) );
  AND U4763 ( .A(n989), .B(n5148), .Z(n5150) );
  XNOR U4764 ( .A(n5149), .B(n5146), .Z(n5148) );
  XOR U4765 ( .A(n5151), .B(n5152), .Z(n5146) );
  AND U4766 ( .A(n992), .B(n5153), .Z(n5152) );
  XOR U4767 ( .A(p_input[1397]), .B(n5151), .Z(n5153) );
  XOR U4768 ( .A(n5154), .B(n5155), .Z(n5151) );
  AND U4769 ( .A(n996), .B(n5156), .Z(n5155) );
  XOR U4770 ( .A(n5157), .B(n5158), .Z(n5149) );
  AND U4771 ( .A(n1000), .B(n5156), .Z(n5158) );
  XNOR U4772 ( .A(n5157), .B(n5154), .Z(n5156) );
  XOR U4773 ( .A(n5159), .B(n5160), .Z(n5154) );
  AND U4774 ( .A(n1003), .B(n5161), .Z(n5160) );
  XOR U4775 ( .A(p_input[1413]), .B(n5159), .Z(n5161) );
  XOR U4776 ( .A(n5162), .B(n5163), .Z(n5159) );
  AND U4777 ( .A(n1007), .B(n5164), .Z(n5163) );
  XOR U4778 ( .A(n5165), .B(n5166), .Z(n5157) );
  AND U4779 ( .A(n1011), .B(n5164), .Z(n5166) );
  XNOR U4780 ( .A(n5165), .B(n5162), .Z(n5164) );
  XOR U4781 ( .A(n5167), .B(n5168), .Z(n5162) );
  AND U4782 ( .A(n1014), .B(n5169), .Z(n5168) );
  XOR U4783 ( .A(p_input[1429]), .B(n5167), .Z(n5169) );
  XOR U4784 ( .A(n5170), .B(n5171), .Z(n5167) );
  AND U4785 ( .A(n1018), .B(n5172), .Z(n5171) );
  XOR U4786 ( .A(n5173), .B(n5174), .Z(n5165) );
  AND U4787 ( .A(n1022), .B(n5172), .Z(n5174) );
  XNOR U4788 ( .A(n5173), .B(n5170), .Z(n5172) );
  XOR U4789 ( .A(n5175), .B(n5176), .Z(n5170) );
  AND U4790 ( .A(n1025), .B(n5177), .Z(n5176) );
  XOR U4791 ( .A(p_input[1445]), .B(n5175), .Z(n5177) );
  XOR U4792 ( .A(n5178), .B(n5179), .Z(n5175) );
  AND U4793 ( .A(n1029), .B(n5180), .Z(n5179) );
  XOR U4794 ( .A(n5181), .B(n5182), .Z(n5173) );
  AND U4795 ( .A(n1033), .B(n5180), .Z(n5182) );
  XNOR U4796 ( .A(n5181), .B(n5178), .Z(n5180) );
  XOR U4797 ( .A(n5183), .B(n5184), .Z(n5178) );
  AND U4798 ( .A(n1036), .B(n5185), .Z(n5184) );
  XOR U4799 ( .A(p_input[1461]), .B(n5183), .Z(n5185) );
  XOR U4800 ( .A(n5186), .B(n5187), .Z(n5183) );
  AND U4801 ( .A(n1040), .B(n5188), .Z(n5187) );
  XOR U4802 ( .A(n5189), .B(n5190), .Z(n5181) );
  AND U4803 ( .A(n1044), .B(n5188), .Z(n5190) );
  XNOR U4804 ( .A(n5189), .B(n5186), .Z(n5188) );
  XOR U4805 ( .A(n5191), .B(n5192), .Z(n5186) );
  AND U4806 ( .A(n1047), .B(n5193), .Z(n5192) );
  XOR U4807 ( .A(p_input[1477]), .B(n5191), .Z(n5193) );
  XOR U4808 ( .A(n5194), .B(n5195), .Z(n5191) );
  AND U4809 ( .A(n1051), .B(n5196), .Z(n5195) );
  XOR U4810 ( .A(n5197), .B(n5198), .Z(n5189) );
  AND U4811 ( .A(n1055), .B(n5196), .Z(n5198) );
  XNOR U4812 ( .A(n5197), .B(n5194), .Z(n5196) );
  XOR U4813 ( .A(n5199), .B(n5200), .Z(n5194) );
  AND U4814 ( .A(n1058), .B(n5201), .Z(n5200) );
  XOR U4815 ( .A(p_input[1493]), .B(n5199), .Z(n5201) );
  XOR U4816 ( .A(n5202), .B(n5203), .Z(n5199) );
  AND U4817 ( .A(n1062), .B(n5204), .Z(n5203) );
  XOR U4818 ( .A(n5205), .B(n5206), .Z(n5197) );
  AND U4819 ( .A(n1066), .B(n5204), .Z(n5206) );
  XNOR U4820 ( .A(n5205), .B(n5202), .Z(n5204) );
  XOR U4821 ( .A(n5207), .B(n5208), .Z(n5202) );
  AND U4822 ( .A(n1069), .B(n5209), .Z(n5208) );
  XOR U4823 ( .A(p_input[1509]), .B(n5207), .Z(n5209) );
  XOR U4824 ( .A(n5210), .B(n5211), .Z(n5207) );
  AND U4825 ( .A(n1073), .B(n5212), .Z(n5211) );
  XOR U4826 ( .A(n5213), .B(n5214), .Z(n5205) );
  AND U4827 ( .A(n1077), .B(n5212), .Z(n5214) );
  XNOR U4828 ( .A(n5213), .B(n5210), .Z(n5212) );
  XOR U4829 ( .A(n5215), .B(n5216), .Z(n5210) );
  AND U4830 ( .A(n1080), .B(n5217), .Z(n5216) );
  XOR U4831 ( .A(p_input[1525]), .B(n5215), .Z(n5217) );
  XOR U4832 ( .A(n5218), .B(n5219), .Z(n5215) );
  AND U4833 ( .A(n1084), .B(n5220), .Z(n5219) );
  XOR U4834 ( .A(n5221), .B(n5222), .Z(n5213) );
  AND U4835 ( .A(n1088), .B(n5220), .Z(n5222) );
  XNOR U4836 ( .A(n5221), .B(n5218), .Z(n5220) );
  XOR U4837 ( .A(n5223), .B(n5224), .Z(n5218) );
  AND U4838 ( .A(n1091), .B(n5225), .Z(n5224) );
  XOR U4839 ( .A(p_input[1541]), .B(n5223), .Z(n5225) );
  XOR U4840 ( .A(n5226), .B(n5227), .Z(n5223) );
  AND U4841 ( .A(n1095), .B(n5228), .Z(n5227) );
  XOR U4842 ( .A(n5229), .B(n5230), .Z(n5221) );
  AND U4843 ( .A(n1099), .B(n5228), .Z(n5230) );
  XNOR U4844 ( .A(n5229), .B(n5226), .Z(n5228) );
  XOR U4845 ( .A(n5231), .B(n5232), .Z(n5226) );
  AND U4846 ( .A(n1102), .B(n5233), .Z(n5232) );
  XOR U4847 ( .A(p_input[1557]), .B(n5231), .Z(n5233) );
  XOR U4848 ( .A(n5234), .B(n5235), .Z(n5231) );
  AND U4849 ( .A(n1106), .B(n5236), .Z(n5235) );
  XOR U4850 ( .A(n5237), .B(n5238), .Z(n5229) );
  AND U4851 ( .A(n1110), .B(n5236), .Z(n5238) );
  XNOR U4852 ( .A(n5237), .B(n5234), .Z(n5236) );
  XOR U4853 ( .A(n5239), .B(n5240), .Z(n5234) );
  AND U4854 ( .A(n1113), .B(n5241), .Z(n5240) );
  XOR U4855 ( .A(p_input[1573]), .B(n5239), .Z(n5241) );
  XOR U4856 ( .A(n5242), .B(n5243), .Z(n5239) );
  AND U4857 ( .A(n1117), .B(n5244), .Z(n5243) );
  XOR U4858 ( .A(n5245), .B(n5246), .Z(n5237) );
  AND U4859 ( .A(n1121), .B(n5244), .Z(n5246) );
  XNOR U4860 ( .A(n5245), .B(n5242), .Z(n5244) );
  XOR U4861 ( .A(n5247), .B(n5248), .Z(n5242) );
  AND U4862 ( .A(n1124), .B(n5249), .Z(n5248) );
  XOR U4863 ( .A(p_input[1589]), .B(n5247), .Z(n5249) );
  XOR U4864 ( .A(n5250), .B(n5251), .Z(n5247) );
  AND U4865 ( .A(n1128), .B(n5252), .Z(n5251) );
  XOR U4866 ( .A(n5253), .B(n5254), .Z(n5245) );
  AND U4867 ( .A(n1132), .B(n5252), .Z(n5254) );
  XNOR U4868 ( .A(n5253), .B(n5250), .Z(n5252) );
  XOR U4869 ( .A(n5255), .B(n5256), .Z(n5250) );
  AND U4870 ( .A(n1135), .B(n5257), .Z(n5256) );
  XOR U4871 ( .A(p_input[1605]), .B(n5255), .Z(n5257) );
  XOR U4872 ( .A(n5258), .B(n5259), .Z(n5255) );
  AND U4873 ( .A(n1139), .B(n5260), .Z(n5259) );
  XOR U4874 ( .A(n5261), .B(n5262), .Z(n5253) );
  AND U4875 ( .A(n1143), .B(n5260), .Z(n5262) );
  XNOR U4876 ( .A(n5261), .B(n5258), .Z(n5260) );
  XOR U4877 ( .A(n5263), .B(n5264), .Z(n5258) );
  AND U4878 ( .A(n1146), .B(n5265), .Z(n5264) );
  XOR U4879 ( .A(p_input[1621]), .B(n5263), .Z(n5265) );
  XOR U4880 ( .A(n5266), .B(n5267), .Z(n5263) );
  AND U4881 ( .A(n1150), .B(n5268), .Z(n5267) );
  XOR U4882 ( .A(n5269), .B(n5270), .Z(n5261) );
  AND U4883 ( .A(n1154), .B(n5268), .Z(n5270) );
  XNOR U4884 ( .A(n5269), .B(n5266), .Z(n5268) );
  XOR U4885 ( .A(n5271), .B(n5272), .Z(n5266) );
  AND U4886 ( .A(n1157), .B(n5273), .Z(n5272) );
  XOR U4887 ( .A(p_input[1637]), .B(n5271), .Z(n5273) );
  XOR U4888 ( .A(n5274), .B(n5275), .Z(n5271) );
  AND U4889 ( .A(n1161), .B(n5276), .Z(n5275) );
  XOR U4890 ( .A(n5277), .B(n5278), .Z(n5269) );
  AND U4891 ( .A(n1165), .B(n5276), .Z(n5278) );
  XNOR U4892 ( .A(n5277), .B(n5274), .Z(n5276) );
  XOR U4893 ( .A(n5279), .B(n5280), .Z(n5274) );
  AND U4894 ( .A(n1168), .B(n5281), .Z(n5280) );
  XOR U4895 ( .A(p_input[1653]), .B(n5279), .Z(n5281) );
  XOR U4896 ( .A(n5282), .B(n5283), .Z(n5279) );
  AND U4897 ( .A(n1172), .B(n5284), .Z(n5283) );
  XOR U4898 ( .A(n5285), .B(n5286), .Z(n5277) );
  AND U4899 ( .A(n1176), .B(n5284), .Z(n5286) );
  XNOR U4900 ( .A(n5285), .B(n5282), .Z(n5284) );
  XOR U4901 ( .A(n5287), .B(n5288), .Z(n5282) );
  AND U4902 ( .A(n1179), .B(n5289), .Z(n5288) );
  XOR U4903 ( .A(p_input[1669]), .B(n5287), .Z(n5289) );
  XOR U4904 ( .A(n5290), .B(n5291), .Z(n5287) );
  AND U4905 ( .A(n1183), .B(n5292), .Z(n5291) );
  XOR U4906 ( .A(n5293), .B(n5294), .Z(n5285) );
  AND U4907 ( .A(n1187), .B(n5292), .Z(n5294) );
  XNOR U4908 ( .A(n5293), .B(n5290), .Z(n5292) );
  XOR U4909 ( .A(n5295), .B(n5296), .Z(n5290) );
  AND U4910 ( .A(n1190), .B(n5297), .Z(n5296) );
  XOR U4911 ( .A(p_input[1685]), .B(n5295), .Z(n5297) );
  XOR U4912 ( .A(n5298), .B(n5299), .Z(n5295) );
  AND U4913 ( .A(n1194), .B(n5300), .Z(n5299) );
  XOR U4914 ( .A(n5301), .B(n5302), .Z(n5293) );
  AND U4915 ( .A(n1198), .B(n5300), .Z(n5302) );
  XNOR U4916 ( .A(n5301), .B(n5298), .Z(n5300) );
  XOR U4917 ( .A(n5303), .B(n5304), .Z(n5298) );
  AND U4918 ( .A(n1201), .B(n5305), .Z(n5304) );
  XOR U4919 ( .A(p_input[1701]), .B(n5303), .Z(n5305) );
  XOR U4920 ( .A(n5306), .B(n5307), .Z(n5303) );
  AND U4921 ( .A(n1205), .B(n5308), .Z(n5307) );
  XOR U4922 ( .A(n5309), .B(n5310), .Z(n5301) );
  AND U4923 ( .A(n1209), .B(n5308), .Z(n5310) );
  XNOR U4924 ( .A(n5309), .B(n5306), .Z(n5308) );
  XOR U4925 ( .A(n5311), .B(n5312), .Z(n5306) );
  AND U4926 ( .A(n1212), .B(n5313), .Z(n5312) );
  XOR U4927 ( .A(p_input[1717]), .B(n5311), .Z(n5313) );
  XOR U4928 ( .A(n5314), .B(n5315), .Z(n5311) );
  AND U4929 ( .A(n1216), .B(n5316), .Z(n5315) );
  XOR U4930 ( .A(n5317), .B(n5318), .Z(n5309) );
  AND U4931 ( .A(n1220), .B(n5316), .Z(n5318) );
  XNOR U4932 ( .A(n5317), .B(n5314), .Z(n5316) );
  XOR U4933 ( .A(n5319), .B(n5320), .Z(n5314) );
  AND U4934 ( .A(n1223), .B(n5321), .Z(n5320) );
  XOR U4935 ( .A(p_input[1733]), .B(n5319), .Z(n5321) );
  XOR U4936 ( .A(n5322), .B(n5323), .Z(n5319) );
  AND U4937 ( .A(n1227), .B(n5324), .Z(n5323) );
  XOR U4938 ( .A(n5325), .B(n5326), .Z(n5317) );
  AND U4939 ( .A(n1231), .B(n5324), .Z(n5326) );
  XNOR U4940 ( .A(n5325), .B(n5322), .Z(n5324) );
  XOR U4941 ( .A(n5327), .B(n5328), .Z(n5322) );
  AND U4942 ( .A(n1234), .B(n5329), .Z(n5328) );
  XOR U4943 ( .A(p_input[1749]), .B(n5327), .Z(n5329) );
  XOR U4944 ( .A(n5330), .B(n5331), .Z(n5327) );
  AND U4945 ( .A(n1238), .B(n5332), .Z(n5331) );
  XOR U4946 ( .A(n5333), .B(n5334), .Z(n5325) );
  AND U4947 ( .A(n1242), .B(n5332), .Z(n5334) );
  XNOR U4948 ( .A(n5333), .B(n5330), .Z(n5332) );
  XOR U4949 ( .A(n5335), .B(n5336), .Z(n5330) );
  AND U4950 ( .A(n1245), .B(n5337), .Z(n5336) );
  XOR U4951 ( .A(p_input[1765]), .B(n5335), .Z(n5337) );
  XOR U4952 ( .A(n5338), .B(n5339), .Z(n5335) );
  AND U4953 ( .A(n1249), .B(n5340), .Z(n5339) );
  XOR U4954 ( .A(n5341), .B(n5342), .Z(n5333) );
  AND U4955 ( .A(n1253), .B(n5340), .Z(n5342) );
  XNOR U4956 ( .A(n5341), .B(n5338), .Z(n5340) );
  XOR U4957 ( .A(n5343), .B(n5344), .Z(n5338) );
  AND U4958 ( .A(n1256), .B(n5345), .Z(n5344) );
  XOR U4959 ( .A(p_input[1781]), .B(n5343), .Z(n5345) );
  XOR U4960 ( .A(n5346), .B(n5347), .Z(n5343) );
  AND U4961 ( .A(n1260), .B(n5348), .Z(n5347) );
  XOR U4962 ( .A(n5349), .B(n5350), .Z(n5341) );
  AND U4963 ( .A(n1264), .B(n5348), .Z(n5350) );
  XNOR U4964 ( .A(n5349), .B(n5346), .Z(n5348) );
  XOR U4965 ( .A(n5351), .B(n5352), .Z(n5346) );
  AND U4966 ( .A(n1267), .B(n5353), .Z(n5352) );
  XOR U4967 ( .A(p_input[1797]), .B(n5351), .Z(n5353) );
  XOR U4968 ( .A(n5354), .B(n5355), .Z(n5351) );
  AND U4969 ( .A(n1271), .B(n5356), .Z(n5355) );
  XOR U4970 ( .A(n5357), .B(n5358), .Z(n5349) );
  AND U4971 ( .A(n1275), .B(n5356), .Z(n5358) );
  XNOR U4972 ( .A(n5357), .B(n5354), .Z(n5356) );
  XOR U4973 ( .A(n5359), .B(n5360), .Z(n5354) );
  AND U4974 ( .A(n1278), .B(n5361), .Z(n5360) );
  XOR U4975 ( .A(p_input[1813]), .B(n5359), .Z(n5361) );
  XOR U4976 ( .A(n5362), .B(n5363), .Z(n5359) );
  AND U4977 ( .A(n1282), .B(n5364), .Z(n5363) );
  XOR U4978 ( .A(n5365), .B(n5366), .Z(n5357) );
  AND U4979 ( .A(n1286), .B(n5364), .Z(n5366) );
  XNOR U4980 ( .A(n5365), .B(n5362), .Z(n5364) );
  XOR U4981 ( .A(n5367), .B(n5368), .Z(n5362) );
  AND U4982 ( .A(n1289), .B(n5369), .Z(n5368) );
  XOR U4983 ( .A(p_input[1829]), .B(n5367), .Z(n5369) );
  XOR U4984 ( .A(n5370), .B(n5371), .Z(n5367) );
  AND U4985 ( .A(n1293), .B(n5372), .Z(n5371) );
  XOR U4986 ( .A(n5373), .B(n5374), .Z(n5365) );
  AND U4987 ( .A(n1297), .B(n5372), .Z(n5374) );
  XNOR U4988 ( .A(n5373), .B(n5370), .Z(n5372) );
  XOR U4989 ( .A(n5375), .B(n5376), .Z(n5370) );
  AND U4990 ( .A(n1300), .B(n5377), .Z(n5376) );
  XOR U4991 ( .A(p_input[1845]), .B(n5375), .Z(n5377) );
  XOR U4992 ( .A(n5378), .B(n5379), .Z(n5375) );
  AND U4993 ( .A(n1304), .B(n5380), .Z(n5379) );
  XOR U4994 ( .A(n5381), .B(n5382), .Z(n5373) );
  AND U4995 ( .A(n1308), .B(n5380), .Z(n5382) );
  XNOR U4996 ( .A(n5381), .B(n5378), .Z(n5380) );
  XOR U4997 ( .A(n5383), .B(n5384), .Z(n5378) );
  AND U4998 ( .A(n1311), .B(n5385), .Z(n5384) );
  XOR U4999 ( .A(p_input[1861]), .B(n5383), .Z(n5385) );
  XOR U5000 ( .A(n5386), .B(n5387), .Z(n5383) );
  AND U5001 ( .A(n1315), .B(n5388), .Z(n5387) );
  XOR U5002 ( .A(n5389), .B(n5390), .Z(n5381) );
  AND U5003 ( .A(n1319), .B(n5388), .Z(n5390) );
  XNOR U5004 ( .A(n5389), .B(n5386), .Z(n5388) );
  XOR U5005 ( .A(n5391), .B(n5392), .Z(n5386) );
  AND U5006 ( .A(n1322), .B(n5393), .Z(n5392) );
  XOR U5007 ( .A(p_input[1877]), .B(n5391), .Z(n5393) );
  XOR U5008 ( .A(n5394), .B(n5395), .Z(n5391) );
  AND U5009 ( .A(n1326), .B(n5396), .Z(n5395) );
  XOR U5010 ( .A(n5397), .B(n5398), .Z(n5389) );
  AND U5011 ( .A(n1330), .B(n5396), .Z(n5398) );
  XNOR U5012 ( .A(n5397), .B(n5394), .Z(n5396) );
  XOR U5013 ( .A(n5399), .B(n5400), .Z(n5394) );
  AND U5014 ( .A(n1333), .B(n5401), .Z(n5400) );
  XOR U5015 ( .A(p_input[1893]), .B(n5399), .Z(n5401) );
  XOR U5016 ( .A(n5402), .B(n5403), .Z(n5399) );
  AND U5017 ( .A(n1337), .B(n5404), .Z(n5403) );
  XOR U5018 ( .A(n5405), .B(n5406), .Z(n5397) );
  AND U5019 ( .A(n1341), .B(n5404), .Z(n5406) );
  XNOR U5020 ( .A(n5405), .B(n5402), .Z(n5404) );
  XOR U5021 ( .A(n5407), .B(n5408), .Z(n5402) );
  AND U5022 ( .A(n1344), .B(n5409), .Z(n5408) );
  XOR U5023 ( .A(p_input[1909]), .B(n5407), .Z(n5409) );
  XOR U5024 ( .A(n5410), .B(n5411), .Z(n5407) );
  AND U5025 ( .A(n1348), .B(n5412), .Z(n5411) );
  XOR U5026 ( .A(n5413), .B(n5414), .Z(n5405) );
  AND U5027 ( .A(n1352), .B(n5412), .Z(n5414) );
  XNOR U5028 ( .A(n5413), .B(n5410), .Z(n5412) );
  XOR U5029 ( .A(n5415), .B(n5416), .Z(n5410) );
  AND U5030 ( .A(n1355), .B(n5417), .Z(n5416) );
  XOR U5031 ( .A(p_input[1925]), .B(n5415), .Z(n5417) );
  XOR U5032 ( .A(n5418), .B(n5419), .Z(n5415) );
  AND U5033 ( .A(n1359), .B(n5420), .Z(n5419) );
  XOR U5034 ( .A(n5421), .B(n5422), .Z(n5413) );
  AND U5035 ( .A(n1363), .B(n5420), .Z(n5422) );
  XNOR U5036 ( .A(n5421), .B(n5418), .Z(n5420) );
  XOR U5037 ( .A(n5423), .B(n5424), .Z(n5418) );
  AND U5038 ( .A(n1366), .B(n5425), .Z(n5424) );
  XOR U5039 ( .A(p_input[1941]), .B(n5423), .Z(n5425) );
  XOR U5040 ( .A(n5426), .B(n5427), .Z(n5423) );
  AND U5041 ( .A(n1370), .B(n5428), .Z(n5427) );
  XOR U5042 ( .A(n5429), .B(n5430), .Z(n5421) );
  AND U5043 ( .A(n1374), .B(n5428), .Z(n5430) );
  XNOR U5044 ( .A(n5429), .B(n5426), .Z(n5428) );
  XOR U5045 ( .A(n5431), .B(n5432), .Z(n5426) );
  AND U5046 ( .A(n1377), .B(n5433), .Z(n5432) );
  XOR U5047 ( .A(p_input[1957]), .B(n5431), .Z(n5433) );
  XOR U5048 ( .A(n5434), .B(n5435), .Z(n5431) );
  AND U5049 ( .A(n1381), .B(n5436), .Z(n5435) );
  XOR U5050 ( .A(n5437), .B(n5438), .Z(n5429) );
  AND U5051 ( .A(n1385), .B(n5436), .Z(n5438) );
  XNOR U5052 ( .A(n5437), .B(n5434), .Z(n5436) );
  XOR U5053 ( .A(n5439), .B(n5440), .Z(n5434) );
  AND U5054 ( .A(n1388), .B(n5441), .Z(n5440) );
  XOR U5055 ( .A(p_input[1973]), .B(n5439), .Z(n5441) );
  XOR U5056 ( .A(n5442), .B(n5443), .Z(n5439) );
  AND U5057 ( .A(n1392), .B(n5444), .Z(n5443) );
  XOR U5058 ( .A(n5445), .B(n5446), .Z(n5437) );
  AND U5059 ( .A(n1396), .B(n5444), .Z(n5446) );
  XNOR U5060 ( .A(n5445), .B(n5442), .Z(n5444) );
  XOR U5061 ( .A(n5447), .B(n5448), .Z(n5442) );
  AND U5062 ( .A(n1399), .B(n5449), .Z(n5448) );
  XOR U5063 ( .A(p_input[1989]), .B(n5447), .Z(n5449) );
  XOR U5064 ( .A(n5450), .B(n5451), .Z(n5447) );
  AND U5065 ( .A(n1403), .B(n5452), .Z(n5451) );
  XOR U5066 ( .A(n5453), .B(n5454), .Z(n5445) );
  AND U5067 ( .A(n1407), .B(n5452), .Z(n5454) );
  XNOR U5068 ( .A(n5453), .B(n5450), .Z(n5452) );
  XOR U5069 ( .A(n5455), .B(n5456), .Z(n5450) );
  AND U5070 ( .A(n1410), .B(n5457), .Z(n5456) );
  XOR U5071 ( .A(p_input[2005]), .B(n5455), .Z(n5457) );
  XNOR U5072 ( .A(n5458), .B(n5459), .Z(n5455) );
  AND U5073 ( .A(n1414), .B(n5460), .Z(n5459) );
  XNOR U5074 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n5461), .Z(n5453) );
  AND U5075 ( .A(n1417), .B(n5460), .Z(n5461) );
  XOR U5076 ( .A(n5462), .B(n5458), .Z(n5460) );
  XOR U5077 ( .A(n11), .B(n5463), .Z(o[20]) );
  AND U5078 ( .A(n30), .B(n5464), .Z(n11) );
  XOR U5079 ( .A(n12), .B(n5463), .Z(n5464) );
  XOR U5080 ( .A(n5465), .B(n5466), .Z(n5463) );
  AND U5081 ( .A(n34), .B(n5467), .Z(n5466) );
  XOR U5082 ( .A(p_input[4]), .B(n5465), .Z(n5467) );
  XOR U5083 ( .A(n5468), .B(n5469), .Z(n5465) );
  AND U5084 ( .A(n38), .B(n5470), .Z(n5469) );
  XOR U5085 ( .A(n5471), .B(n5472), .Z(n12) );
  AND U5086 ( .A(n42), .B(n5470), .Z(n5472) );
  XNOR U5087 ( .A(n5473), .B(n5468), .Z(n5470) );
  XOR U5088 ( .A(n5474), .B(n5475), .Z(n5468) );
  AND U5089 ( .A(n46), .B(n5476), .Z(n5475) );
  XOR U5090 ( .A(p_input[20]), .B(n5474), .Z(n5476) );
  XOR U5091 ( .A(n5477), .B(n5478), .Z(n5474) );
  AND U5092 ( .A(n50), .B(n5479), .Z(n5478) );
  IV U5093 ( .A(n5471), .Z(n5473) );
  XNOR U5094 ( .A(n5480), .B(n5481), .Z(n5471) );
  AND U5095 ( .A(n54), .B(n5479), .Z(n5481) );
  XNOR U5096 ( .A(n5480), .B(n5477), .Z(n5479) );
  XOR U5097 ( .A(n5482), .B(n5483), .Z(n5477) );
  AND U5098 ( .A(n57), .B(n5484), .Z(n5483) );
  XOR U5099 ( .A(p_input[36]), .B(n5482), .Z(n5484) );
  XOR U5100 ( .A(n5485), .B(n5486), .Z(n5482) );
  AND U5101 ( .A(n61), .B(n5487), .Z(n5486) );
  XOR U5102 ( .A(n5488), .B(n5489), .Z(n5480) );
  AND U5103 ( .A(n65), .B(n5487), .Z(n5489) );
  XNOR U5104 ( .A(n5488), .B(n5485), .Z(n5487) );
  XOR U5105 ( .A(n5490), .B(n5491), .Z(n5485) );
  AND U5106 ( .A(n68), .B(n5492), .Z(n5491) );
  XOR U5107 ( .A(p_input[52]), .B(n5490), .Z(n5492) );
  XOR U5108 ( .A(n5493), .B(n5494), .Z(n5490) );
  AND U5109 ( .A(n72), .B(n5495), .Z(n5494) );
  XOR U5110 ( .A(n5496), .B(n5497), .Z(n5488) );
  AND U5111 ( .A(n76), .B(n5495), .Z(n5497) );
  XNOR U5112 ( .A(n5496), .B(n5493), .Z(n5495) );
  XOR U5113 ( .A(n5498), .B(n5499), .Z(n5493) );
  AND U5114 ( .A(n79), .B(n5500), .Z(n5499) );
  XOR U5115 ( .A(p_input[68]), .B(n5498), .Z(n5500) );
  XOR U5116 ( .A(n5501), .B(n5502), .Z(n5498) );
  AND U5117 ( .A(n83), .B(n5503), .Z(n5502) );
  XOR U5118 ( .A(n5504), .B(n5505), .Z(n5496) );
  AND U5119 ( .A(n87), .B(n5503), .Z(n5505) );
  XNOR U5120 ( .A(n5504), .B(n5501), .Z(n5503) );
  XOR U5121 ( .A(n5506), .B(n5507), .Z(n5501) );
  AND U5122 ( .A(n90), .B(n5508), .Z(n5507) );
  XOR U5123 ( .A(p_input[84]), .B(n5506), .Z(n5508) );
  XOR U5124 ( .A(n5509), .B(n5510), .Z(n5506) );
  AND U5125 ( .A(n94), .B(n5511), .Z(n5510) );
  XOR U5126 ( .A(n5512), .B(n5513), .Z(n5504) );
  AND U5127 ( .A(n98), .B(n5511), .Z(n5513) );
  XNOR U5128 ( .A(n5512), .B(n5509), .Z(n5511) );
  XOR U5129 ( .A(n5514), .B(n5515), .Z(n5509) );
  AND U5130 ( .A(n101), .B(n5516), .Z(n5515) );
  XOR U5131 ( .A(p_input[100]), .B(n5514), .Z(n5516) );
  XOR U5132 ( .A(n5517), .B(n5518), .Z(n5514) );
  AND U5133 ( .A(n105), .B(n5519), .Z(n5518) );
  XOR U5134 ( .A(n5520), .B(n5521), .Z(n5512) );
  AND U5135 ( .A(n109), .B(n5519), .Z(n5521) );
  XNOR U5136 ( .A(n5520), .B(n5517), .Z(n5519) );
  XOR U5137 ( .A(n5522), .B(n5523), .Z(n5517) );
  AND U5138 ( .A(n112), .B(n5524), .Z(n5523) );
  XOR U5139 ( .A(p_input[116]), .B(n5522), .Z(n5524) );
  XOR U5140 ( .A(n5525), .B(n5526), .Z(n5522) );
  AND U5141 ( .A(n116), .B(n5527), .Z(n5526) );
  XOR U5142 ( .A(n5528), .B(n5529), .Z(n5520) );
  AND U5143 ( .A(n120), .B(n5527), .Z(n5529) );
  XNOR U5144 ( .A(n5528), .B(n5525), .Z(n5527) );
  XOR U5145 ( .A(n5530), .B(n5531), .Z(n5525) );
  AND U5146 ( .A(n123), .B(n5532), .Z(n5531) );
  XOR U5147 ( .A(p_input[132]), .B(n5530), .Z(n5532) );
  XOR U5148 ( .A(n5533), .B(n5534), .Z(n5530) );
  AND U5149 ( .A(n127), .B(n5535), .Z(n5534) );
  XOR U5150 ( .A(n5536), .B(n5537), .Z(n5528) );
  AND U5151 ( .A(n131), .B(n5535), .Z(n5537) );
  XNOR U5152 ( .A(n5536), .B(n5533), .Z(n5535) );
  XOR U5153 ( .A(n5538), .B(n5539), .Z(n5533) );
  AND U5154 ( .A(n134), .B(n5540), .Z(n5539) );
  XOR U5155 ( .A(p_input[148]), .B(n5538), .Z(n5540) );
  XOR U5156 ( .A(n5541), .B(n5542), .Z(n5538) );
  AND U5157 ( .A(n138), .B(n5543), .Z(n5542) );
  XOR U5158 ( .A(n5544), .B(n5545), .Z(n5536) );
  AND U5159 ( .A(n142), .B(n5543), .Z(n5545) );
  XNOR U5160 ( .A(n5544), .B(n5541), .Z(n5543) );
  XOR U5161 ( .A(n5546), .B(n5547), .Z(n5541) );
  AND U5162 ( .A(n145), .B(n5548), .Z(n5547) );
  XOR U5163 ( .A(p_input[164]), .B(n5546), .Z(n5548) );
  XOR U5164 ( .A(n5549), .B(n5550), .Z(n5546) );
  AND U5165 ( .A(n149), .B(n5551), .Z(n5550) );
  XOR U5166 ( .A(n5552), .B(n5553), .Z(n5544) );
  AND U5167 ( .A(n153), .B(n5551), .Z(n5553) );
  XNOR U5168 ( .A(n5552), .B(n5549), .Z(n5551) );
  XOR U5169 ( .A(n5554), .B(n5555), .Z(n5549) );
  AND U5170 ( .A(n156), .B(n5556), .Z(n5555) );
  XOR U5171 ( .A(p_input[180]), .B(n5554), .Z(n5556) );
  XOR U5172 ( .A(n5557), .B(n5558), .Z(n5554) );
  AND U5173 ( .A(n160), .B(n5559), .Z(n5558) );
  XOR U5174 ( .A(n5560), .B(n5561), .Z(n5552) );
  AND U5175 ( .A(n164), .B(n5559), .Z(n5561) );
  XNOR U5176 ( .A(n5560), .B(n5557), .Z(n5559) );
  XOR U5177 ( .A(n5562), .B(n5563), .Z(n5557) );
  AND U5178 ( .A(n167), .B(n5564), .Z(n5563) );
  XOR U5179 ( .A(p_input[196]), .B(n5562), .Z(n5564) );
  XOR U5180 ( .A(n5565), .B(n5566), .Z(n5562) );
  AND U5181 ( .A(n171), .B(n5567), .Z(n5566) );
  XOR U5182 ( .A(n5568), .B(n5569), .Z(n5560) );
  AND U5183 ( .A(n175), .B(n5567), .Z(n5569) );
  XNOR U5184 ( .A(n5568), .B(n5565), .Z(n5567) );
  XOR U5185 ( .A(n5570), .B(n5571), .Z(n5565) );
  AND U5186 ( .A(n178), .B(n5572), .Z(n5571) );
  XOR U5187 ( .A(p_input[212]), .B(n5570), .Z(n5572) );
  XOR U5188 ( .A(n5573), .B(n5574), .Z(n5570) );
  AND U5189 ( .A(n182), .B(n5575), .Z(n5574) );
  XOR U5190 ( .A(n5576), .B(n5577), .Z(n5568) );
  AND U5191 ( .A(n186), .B(n5575), .Z(n5577) );
  XNOR U5192 ( .A(n5576), .B(n5573), .Z(n5575) );
  XOR U5193 ( .A(n5578), .B(n5579), .Z(n5573) );
  AND U5194 ( .A(n189), .B(n5580), .Z(n5579) );
  XOR U5195 ( .A(p_input[228]), .B(n5578), .Z(n5580) );
  XOR U5196 ( .A(n5581), .B(n5582), .Z(n5578) );
  AND U5197 ( .A(n193), .B(n5583), .Z(n5582) );
  XOR U5198 ( .A(n5584), .B(n5585), .Z(n5576) );
  AND U5199 ( .A(n197), .B(n5583), .Z(n5585) );
  XNOR U5200 ( .A(n5584), .B(n5581), .Z(n5583) );
  XOR U5201 ( .A(n5586), .B(n5587), .Z(n5581) );
  AND U5202 ( .A(n200), .B(n5588), .Z(n5587) );
  XOR U5203 ( .A(p_input[244]), .B(n5586), .Z(n5588) );
  XOR U5204 ( .A(n5589), .B(n5590), .Z(n5586) );
  AND U5205 ( .A(n204), .B(n5591), .Z(n5590) );
  XOR U5206 ( .A(n5592), .B(n5593), .Z(n5584) );
  AND U5207 ( .A(n208), .B(n5591), .Z(n5593) );
  XNOR U5208 ( .A(n5592), .B(n5589), .Z(n5591) );
  XOR U5209 ( .A(n5594), .B(n5595), .Z(n5589) );
  AND U5210 ( .A(n211), .B(n5596), .Z(n5595) );
  XOR U5211 ( .A(p_input[260]), .B(n5594), .Z(n5596) );
  XOR U5212 ( .A(n5597), .B(n5598), .Z(n5594) );
  AND U5213 ( .A(n215), .B(n5599), .Z(n5598) );
  XOR U5214 ( .A(n5600), .B(n5601), .Z(n5592) );
  AND U5215 ( .A(n219), .B(n5599), .Z(n5601) );
  XNOR U5216 ( .A(n5600), .B(n5597), .Z(n5599) );
  XOR U5217 ( .A(n5602), .B(n5603), .Z(n5597) );
  AND U5218 ( .A(n222), .B(n5604), .Z(n5603) );
  XOR U5219 ( .A(p_input[276]), .B(n5602), .Z(n5604) );
  XOR U5220 ( .A(n5605), .B(n5606), .Z(n5602) );
  AND U5221 ( .A(n226), .B(n5607), .Z(n5606) );
  XOR U5222 ( .A(n5608), .B(n5609), .Z(n5600) );
  AND U5223 ( .A(n230), .B(n5607), .Z(n5609) );
  XNOR U5224 ( .A(n5608), .B(n5605), .Z(n5607) );
  XOR U5225 ( .A(n5610), .B(n5611), .Z(n5605) );
  AND U5226 ( .A(n233), .B(n5612), .Z(n5611) );
  XOR U5227 ( .A(p_input[292]), .B(n5610), .Z(n5612) );
  XOR U5228 ( .A(n5613), .B(n5614), .Z(n5610) );
  AND U5229 ( .A(n237), .B(n5615), .Z(n5614) );
  XOR U5230 ( .A(n5616), .B(n5617), .Z(n5608) );
  AND U5231 ( .A(n241), .B(n5615), .Z(n5617) );
  XNOR U5232 ( .A(n5616), .B(n5613), .Z(n5615) );
  XOR U5233 ( .A(n5618), .B(n5619), .Z(n5613) );
  AND U5234 ( .A(n244), .B(n5620), .Z(n5619) );
  XOR U5235 ( .A(p_input[308]), .B(n5618), .Z(n5620) );
  XOR U5236 ( .A(n5621), .B(n5622), .Z(n5618) );
  AND U5237 ( .A(n248), .B(n5623), .Z(n5622) );
  XOR U5238 ( .A(n5624), .B(n5625), .Z(n5616) );
  AND U5239 ( .A(n252), .B(n5623), .Z(n5625) );
  XNOR U5240 ( .A(n5624), .B(n5621), .Z(n5623) );
  XOR U5241 ( .A(n5626), .B(n5627), .Z(n5621) );
  AND U5242 ( .A(n255), .B(n5628), .Z(n5627) );
  XOR U5243 ( .A(p_input[324]), .B(n5626), .Z(n5628) );
  XOR U5244 ( .A(n5629), .B(n5630), .Z(n5626) );
  AND U5245 ( .A(n259), .B(n5631), .Z(n5630) );
  XOR U5246 ( .A(n5632), .B(n5633), .Z(n5624) );
  AND U5247 ( .A(n263), .B(n5631), .Z(n5633) );
  XNOR U5248 ( .A(n5632), .B(n5629), .Z(n5631) );
  XOR U5249 ( .A(n5634), .B(n5635), .Z(n5629) );
  AND U5250 ( .A(n266), .B(n5636), .Z(n5635) );
  XOR U5251 ( .A(p_input[340]), .B(n5634), .Z(n5636) );
  XOR U5252 ( .A(n5637), .B(n5638), .Z(n5634) );
  AND U5253 ( .A(n270), .B(n5639), .Z(n5638) );
  XOR U5254 ( .A(n5640), .B(n5641), .Z(n5632) );
  AND U5255 ( .A(n274), .B(n5639), .Z(n5641) );
  XNOR U5256 ( .A(n5640), .B(n5637), .Z(n5639) );
  XOR U5257 ( .A(n5642), .B(n5643), .Z(n5637) );
  AND U5258 ( .A(n277), .B(n5644), .Z(n5643) );
  XOR U5259 ( .A(p_input[356]), .B(n5642), .Z(n5644) );
  XOR U5260 ( .A(n5645), .B(n5646), .Z(n5642) );
  AND U5261 ( .A(n281), .B(n5647), .Z(n5646) );
  XOR U5262 ( .A(n5648), .B(n5649), .Z(n5640) );
  AND U5263 ( .A(n285), .B(n5647), .Z(n5649) );
  XNOR U5264 ( .A(n5648), .B(n5645), .Z(n5647) );
  XOR U5265 ( .A(n5650), .B(n5651), .Z(n5645) );
  AND U5266 ( .A(n288), .B(n5652), .Z(n5651) );
  XOR U5267 ( .A(p_input[372]), .B(n5650), .Z(n5652) );
  XOR U5268 ( .A(n5653), .B(n5654), .Z(n5650) );
  AND U5269 ( .A(n292), .B(n5655), .Z(n5654) );
  XOR U5270 ( .A(n5656), .B(n5657), .Z(n5648) );
  AND U5271 ( .A(n296), .B(n5655), .Z(n5657) );
  XNOR U5272 ( .A(n5656), .B(n5653), .Z(n5655) );
  XOR U5273 ( .A(n5658), .B(n5659), .Z(n5653) );
  AND U5274 ( .A(n299), .B(n5660), .Z(n5659) );
  XOR U5275 ( .A(p_input[388]), .B(n5658), .Z(n5660) );
  XOR U5276 ( .A(n5661), .B(n5662), .Z(n5658) );
  AND U5277 ( .A(n303), .B(n5663), .Z(n5662) );
  XOR U5278 ( .A(n5664), .B(n5665), .Z(n5656) );
  AND U5279 ( .A(n307), .B(n5663), .Z(n5665) );
  XNOR U5280 ( .A(n5664), .B(n5661), .Z(n5663) );
  XOR U5281 ( .A(n5666), .B(n5667), .Z(n5661) );
  AND U5282 ( .A(n310), .B(n5668), .Z(n5667) );
  XOR U5283 ( .A(p_input[404]), .B(n5666), .Z(n5668) );
  XOR U5284 ( .A(n5669), .B(n5670), .Z(n5666) );
  AND U5285 ( .A(n314), .B(n5671), .Z(n5670) );
  XOR U5286 ( .A(n5672), .B(n5673), .Z(n5664) );
  AND U5287 ( .A(n318), .B(n5671), .Z(n5673) );
  XNOR U5288 ( .A(n5672), .B(n5669), .Z(n5671) );
  XOR U5289 ( .A(n5674), .B(n5675), .Z(n5669) );
  AND U5290 ( .A(n321), .B(n5676), .Z(n5675) );
  XOR U5291 ( .A(p_input[420]), .B(n5674), .Z(n5676) );
  XOR U5292 ( .A(n5677), .B(n5678), .Z(n5674) );
  AND U5293 ( .A(n325), .B(n5679), .Z(n5678) );
  XOR U5294 ( .A(n5680), .B(n5681), .Z(n5672) );
  AND U5295 ( .A(n329), .B(n5679), .Z(n5681) );
  XNOR U5296 ( .A(n5680), .B(n5677), .Z(n5679) );
  XOR U5297 ( .A(n5682), .B(n5683), .Z(n5677) );
  AND U5298 ( .A(n332), .B(n5684), .Z(n5683) );
  XOR U5299 ( .A(p_input[436]), .B(n5682), .Z(n5684) );
  XOR U5300 ( .A(n5685), .B(n5686), .Z(n5682) );
  AND U5301 ( .A(n336), .B(n5687), .Z(n5686) );
  XOR U5302 ( .A(n5688), .B(n5689), .Z(n5680) );
  AND U5303 ( .A(n340), .B(n5687), .Z(n5689) );
  XNOR U5304 ( .A(n5688), .B(n5685), .Z(n5687) );
  XOR U5305 ( .A(n5690), .B(n5691), .Z(n5685) );
  AND U5306 ( .A(n343), .B(n5692), .Z(n5691) );
  XOR U5307 ( .A(p_input[452]), .B(n5690), .Z(n5692) );
  XOR U5308 ( .A(n5693), .B(n5694), .Z(n5690) );
  AND U5309 ( .A(n347), .B(n5695), .Z(n5694) );
  XOR U5310 ( .A(n5696), .B(n5697), .Z(n5688) );
  AND U5311 ( .A(n351), .B(n5695), .Z(n5697) );
  XNOR U5312 ( .A(n5696), .B(n5693), .Z(n5695) );
  XOR U5313 ( .A(n5698), .B(n5699), .Z(n5693) );
  AND U5314 ( .A(n354), .B(n5700), .Z(n5699) );
  XOR U5315 ( .A(p_input[468]), .B(n5698), .Z(n5700) );
  XOR U5316 ( .A(n5701), .B(n5702), .Z(n5698) );
  AND U5317 ( .A(n358), .B(n5703), .Z(n5702) );
  XOR U5318 ( .A(n5704), .B(n5705), .Z(n5696) );
  AND U5319 ( .A(n362), .B(n5703), .Z(n5705) );
  XNOR U5320 ( .A(n5704), .B(n5701), .Z(n5703) );
  XOR U5321 ( .A(n5706), .B(n5707), .Z(n5701) );
  AND U5322 ( .A(n365), .B(n5708), .Z(n5707) );
  XOR U5323 ( .A(p_input[484]), .B(n5706), .Z(n5708) );
  XOR U5324 ( .A(n5709), .B(n5710), .Z(n5706) );
  AND U5325 ( .A(n369), .B(n5711), .Z(n5710) );
  XOR U5326 ( .A(n5712), .B(n5713), .Z(n5704) );
  AND U5327 ( .A(n373), .B(n5711), .Z(n5713) );
  XNOR U5328 ( .A(n5712), .B(n5709), .Z(n5711) );
  XOR U5329 ( .A(n5714), .B(n5715), .Z(n5709) );
  AND U5330 ( .A(n376), .B(n5716), .Z(n5715) );
  XOR U5331 ( .A(p_input[500]), .B(n5714), .Z(n5716) );
  XOR U5332 ( .A(n5717), .B(n5718), .Z(n5714) );
  AND U5333 ( .A(n380), .B(n5719), .Z(n5718) );
  XOR U5334 ( .A(n5720), .B(n5721), .Z(n5712) );
  AND U5335 ( .A(n384), .B(n5719), .Z(n5721) );
  XNOR U5336 ( .A(n5720), .B(n5717), .Z(n5719) );
  XOR U5337 ( .A(n5722), .B(n5723), .Z(n5717) );
  AND U5338 ( .A(n387), .B(n5724), .Z(n5723) );
  XOR U5339 ( .A(p_input[516]), .B(n5722), .Z(n5724) );
  XOR U5340 ( .A(n5725), .B(n5726), .Z(n5722) );
  AND U5341 ( .A(n391), .B(n5727), .Z(n5726) );
  XOR U5342 ( .A(n5728), .B(n5729), .Z(n5720) );
  AND U5343 ( .A(n395), .B(n5727), .Z(n5729) );
  XNOR U5344 ( .A(n5728), .B(n5725), .Z(n5727) );
  XOR U5345 ( .A(n5730), .B(n5731), .Z(n5725) );
  AND U5346 ( .A(n398), .B(n5732), .Z(n5731) );
  XOR U5347 ( .A(p_input[532]), .B(n5730), .Z(n5732) );
  XOR U5348 ( .A(n5733), .B(n5734), .Z(n5730) );
  AND U5349 ( .A(n402), .B(n5735), .Z(n5734) );
  XOR U5350 ( .A(n5736), .B(n5737), .Z(n5728) );
  AND U5351 ( .A(n406), .B(n5735), .Z(n5737) );
  XNOR U5352 ( .A(n5736), .B(n5733), .Z(n5735) );
  XOR U5353 ( .A(n5738), .B(n5739), .Z(n5733) );
  AND U5354 ( .A(n409), .B(n5740), .Z(n5739) );
  XOR U5355 ( .A(p_input[548]), .B(n5738), .Z(n5740) );
  XOR U5356 ( .A(n5741), .B(n5742), .Z(n5738) );
  AND U5357 ( .A(n413), .B(n5743), .Z(n5742) );
  XOR U5358 ( .A(n5744), .B(n5745), .Z(n5736) );
  AND U5359 ( .A(n417), .B(n5743), .Z(n5745) );
  XNOR U5360 ( .A(n5744), .B(n5741), .Z(n5743) );
  XOR U5361 ( .A(n5746), .B(n5747), .Z(n5741) );
  AND U5362 ( .A(n420), .B(n5748), .Z(n5747) );
  XOR U5363 ( .A(p_input[564]), .B(n5746), .Z(n5748) );
  XOR U5364 ( .A(n5749), .B(n5750), .Z(n5746) );
  AND U5365 ( .A(n424), .B(n5751), .Z(n5750) );
  XOR U5366 ( .A(n5752), .B(n5753), .Z(n5744) );
  AND U5367 ( .A(n428), .B(n5751), .Z(n5753) );
  XNOR U5368 ( .A(n5752), .B(n5749), .Z(n5751) );
  XOR U5369 ( .A(n5754), .B(n5755), .Z(n5749) );
  AND U5370 ( .A(n431), .B(n5756), .Z(n5755) );
  XOR U5371 ( .A(p_input[580]), .B(n5754), .Z(n5756) );
  XOR U5372 ( .A(n5757), .B(n5758), .Z(n5754) );
  AND U5373 ( .A(n435), .B(n5759), .Z(n5758) );
  XOR U5374 ( .A(n5760), .B(n5761), .Z(n5752) );
  AND U5375 ( .A(n439), .B(n5759), .Z(n5761) );
  XNOR U5376 ( .A(n5760), .B(n5757), .Z(n5759) );
  XOR U5377 ( .A(n5762), .B(n5763), .Z(n5757) );
  AND U5378 ( .A(n442), .B(n5764), .Z(n5763) );
  XOR U5379 ( .A(p_input[596]), .B(n5762), .Z(n5764) );
  XOR U5380 ( .A(n5765), .B(n5766), .Z(n5762) );
  AND U5381 ( .A(n446), .B(n5767), .Z(n5766) );
  XOR U5382 ( .A(n5768), .B(n5769), .Z(n5760) );
  AND U5383 ( .A(n450), .B(n5767), .Z(n5769) );
  XNOR U5384 ( .A(n5768), .B(n5765), .Z(n5767) );
  XOR U5385 ( .A(n5770), .B(n5771), .Z(n5765) );
  AND U5386 ( .A(n453), .B(n5772), .Z(n5771) );
  XOR U5387 ( .A(p_input[612]), .B(n5770), .Z(n5772) );
  XOR U5388 ( .A(n5773), .B(n5774), .Z(n5770) );
  AND U5389 ( .A(n457), .B(n5775), .Z(n5774) );
  XOR U5390 ( .A(n5776), .B(n5777), .Z(n5768) );
  AND U5391 ( .A(n461), .B(n5775), .Z(n5777) );
  XNOR U5392 ( .A(n5776), .B(n5773), .Z(n5775) );
  XOR U5393 ( .A(n5778), .B(n5779), .Z(n5773) );
  AND U5394 ( .A(n464), .B(n5780), .Z(n5779) );
  XOR U5395 ( .A(p_input[628]), .B(n5778), .Z(n5780) );
  XOR U5396 ( .A(n5781), .B(n5782), .Z(n5778) );
  AND U5397 ( .A(n468), .B(n5783), .Z(n5782) );
  XOR U5398 ( .A(n5784), .B(n5785), .Z(n5776) );
  AND U5399 ( .A(n472), .B(n5783), .Z(n5785) );
  XNOR U5400 ( .A(n5784), .B(n5781), .Z(n5783) );
  XOR U5401 ( .A(n5786), .B(n5787), .Z(n5781) );
  AND U5402 ( .A(n475), .B(n5788), .Z(n5787) );
  XOR U5403 ( .A(p_input[644]), .B(n5786), .Z(n5788) );
  XOR U5404 ( .A(n5789), .B(n5790), .Z(n5786) );
  AND U5405 ( .A(n479), .B(n5791), .Z(n5790) );
  XOR U5406 ( .A(n5792), .B(n5793), .Z(n5784) );
  AND U5407 ( .A(n483), .B(n5791), .Z(n5793) );
  XNOR U5408 ( .A(n5792), .B(n5789), .Z(n5791) );
  XOR U5409 ( .A(n5794), .B(n5795), .Z(n5789) );
  AND U5410 ( .A(n486), .B(n5796), .Z(n5795) );
  XOR U5411 ( .A(p_input[660]), .B(n5794), .Z(n5796) );
  XOR U5412 ( .A(n5797), .B(n5798), .Z(n5794) );
  AND U5413 ( .A(n490), .B(n5799), .Z(n5798) );
  XOR U5414 ( .A(n5800), .B(n5801), .Z(n5792) );
  AND U5415 ( .A(n494), .B(n5799), .Z(n5801) );
  XNOR U5416 ( .A(n5800), .B(n5797), .Z(n5799) );
  XOR U5417 ( .A(n5802), .B(n5803), .Z(n5797) );
  AND U5418 ( .A(n497), .B(n5804), .Z(n5803) );
  XOR U5419 ( .A(p_input[676]), .B(n5802), .Z(n5804) );
  XOR U5420 ( .A(n5805), .B(n5806), .Z(n5802) );
  AND U5421 ( .A(n501), .B(n5807), .Z(n5806) );
  XOR U5422 ( .A(n5808), .B(n5809), .Z(n5800) );
  AND U5423 ( .A(n505), .B(n5807), .Z(n5809) );
  XNOR U5424 ( .A(n5808), .B(n5805), .Z(n5807) );
  XOR U5425 ( .A(n5810), .B(n5811), .Z(n5805) );
  AND U5426 ( .A(n508), .B(n5812), .Z(n5811) );
  XOR U5427 ( .A(p_input[692]), .B(n5810), .Z(n5812) );
  XOR U5428 ( .A(n5813), .B(n5814), .Z(n5810) );
  AND U5429 ( .A(n512), .B(n5815), .Z(n5814) );
  XOR U5430 ( .A(n5816), .B(n5817), .Z(n5808) );
  AND U5431 ( .A(n516), .B(n5815), .Z(n5817) );
  XNOR U5432 ( .A(n5816), .B(n5813), .Z(n5815) );
  XOR U5433 ( .A(n5818), .B(n5819), .Z(n5813) );
  AND U5434 ( .A(n519), .B(n5820), .Z(n5819) );
  XOR U5435 ( .A(p_input[708]), .B(n5818), .Z(n5820) );
  XOR U5436 ( .A(n5821), .B(n5822), .Z(n5818) );
  AND U5437 ( .A(n523), .B(n5823), .Z(n5822) );
  XOR U5438 ( .A(n5824), .B(n5825), .Z(n5816) );
  AND U5439 ( .A(n527), .B(n5823), .Z(n5825) );
  XNOR U5440 ( .A(n5824), .B(n5821), .Z(n5823) );
  XOR U5441 ( .A(n5826), .B(n5827), .Z(n5821) );
  AND U5442 ( .A(n530), .B(n5828), .Z(n5827) );
  XOR U5443 ( .A(p_input[724]), .B(n5826), .Z(n5828) );
  XOR U5444 ( .A(n5829), .B(n5830), .Z(n5826) );
  AND U5445 ( .A(n534), .B(n5831), .Z(n5830) );
  XOR U5446 ( .A(n5832), .B(n5833), .Z(n5824) );
  AND U5447 ( .A(n538), .B(n5831), .Z(n5833) );
  XNOR U5448 ( .A(n5832), .B(n5829), .Z(n5831) );
  XOR U5449 ( .A(n5834), .B(n5835), .Z(n5829) );
  AND U5450 ( .A(n541), .B(n5836), .Z(n5835) );
  XOR U5451 ( .A(p_input[740]), .B(n5834), .Z(n5836) );
  XOR U5452 ( .A(n5837), .B(n5838), .Z(n5834) );
  AND U5453 ( .A(n545), .B(n5839), .Z(n5838) );
  XOR U5454 ( .A(n5840), .B(n5841), .Z(n5832) );
  AND U5455 ( .A(n549), .B(n5839), .Z(n5841) );
  XNOR U5456 ( .A(n5840), .B(n5837), .Z(n5839) );
  XOR U5457 ( .A(n5842), .B(n5843), .Z(n5837) );
  AND U5458 ( .A(n552), .B(n5844), .Z(n5843) );
  XOR U5459 ( .A(p_input[756]), .B(n5842), .Z(n5844) );
  XOR U5460 ( .A(n5845), .B(n5846), .Z(n5842) );
  AND U5461 ( .A(n556), .B(n5847), .Z(n5846) );
  XOR U5462 ( .A(n5848), .B(n5849), .Z(n5840) );
  AND U5463 ( .A(n560), .B(n5847), .Z(n5849) );
  XNOR U5464 ( .A(n5848), .B(n5845), .Z(n5847) );
  XOR U5465 ( .A(n5850), .B(n5851), .Z(n5845) );
  AND U5466 ( .A(n563), .B(n5852), .Z(n5851) );
  XOR U5467 ( .A(p_input[772]), .B(n5850), .Z(n5852) );
  XOR U5468 ( .A(n5853), .B(n5854), .Z(n5850) );
  AND U5469 ( .A(n567), .B(n5855), .Z(n5854) );
  XOR U5470 ( .A(n5856), .B(n5857), .Z(n5848) );
  AND U5471 ( .A(n571), .B(n5855), .Z(n5857) );
  XNOR U5472 ( .A(n5856), .B(n5853), .Z(n5855) );
  XOR U5473 ( .A(n5858), .B(n5859), .Z(n5853) );
  AND U5474 ( .A(n574), .B(n5860), .Z(n5859) );
  XOR U5475 ( .A(p_input[788]), .B(n5858), .Z(n5860) );
  XOR U5476 ( .A(n5861), .B(n5862), .Z(n5858) );
  AND U5477 ( .A(n578), .B(n5863), .Z(n5862) );
  XOR U5478 ( .A(n5864), .B(n5865), .Z(n5856) );
  AND U5479 ( .A(n582), .B(n5863), .Z(n5865) );
  XNOR U5480 ( .A(n5864), .B(n5861), .Z(n5863) );
  XOR U5481 ( .A(n5866), .B(n5867), .Z(n5861) );
  AND U5482 ( .A(n585), .B(n5868), .Z(n5867) );
  XOR U5483 ( .A(p_input[804]), .B(n5866), .Z(n5868) );
  XOR U5484 ( .A(n5869), .B(n5870), .Z(n5866) );
  AND U5485 ( .A(n589), .B(n5871), .Z(n5870) );
  XOR U5486 ( .A(n5872), .B(n5873), .Z(n5864) );
  AND U5487 ( .A(n593), .B(n5871), .Z(n5873) );
  XNOR U5488 ( .A(n5872), .B(n5869), .Z(n5871) );
  XOR U5489 ( .A(n5874), .B(n5875), .Z(n5869) );
  AND U5490 ( .A(n596), .B(n5876), .Z(n5875) );
  XOR U5491 ( .A(p_input[820]), .B(n5874), .Z(n5876) );
  XOR U5492 ( .A(n5877), .B(n5878), .Z(n5874) );
  AND U5493 ( .A(n600), .B(n5879), .Z(n5878) );
  XOR U5494 ( .A(n5880), .B(n5881), .Z(n5872) );
  AND U5495 ( .A(n604), .B(n5879), .Z(n5881) );
  XNOR U5496 ( .A(n5880), .B(n5877), .Z(n5879) );
  XOR U5497 ( .A(n5882), .B(n5883), .Z(n5877) );
  AND U5498 ( .A(n607), .B(n5884), .Z(n5883) );
  XOR U5499 ( .A(p_input[836]), .B(n5882), .Z(n5884) );
  XOR U5500 ( .A(n5885), .B(n5886), .Z(n5882) );
  AND U5501 ( .A(n611), .B(n5887), .Z(n5886) );
  XOR U5502 ( .A(n5888), .B(n5889), .Z(n5880) );
  AND U5503 ( .A(n615), .B(n5887), .Z(n5889) );
  XNOR U5504 ( .A(n5888), .B(n5885), .Z(n5887) );
  XOR U5505 ( .A(n5890), .B(n5891), .Z(n5885) );
  AND U5506 ( .A(n618), .B(n5892), .Z(n5891) );
  XOR U5507 ( .A(p_input[852]), .B(n5890), .Z(n5892) );
  XOR U5508 ( .A(n5893), .B(n5894), .Z(n5890) );
  AND U5509 ( .A(n622), .B(n5895), .Z(n5894) );
  XOR U5510 ( .A(n5896), .B(n5897), .Z(n5888) );
  AND U5511 ( .A(n626), .B(n5895), .Z(n5897) );
  XNOR U5512 ( .A(n5896), .B(n5893), .Z(n5895) );
  XOR U5513 ( .A(n5898), .B(n5899), .Z(n5893) );
  AND U5514 ( .A(n629), .B(n5900), .Z(n5899) );
  XOR U5515 ( .A(p_input[868]), .B(n5898), .Z(n5900) );
  XOR U5516 ( .A(n5901), .B(n5902), .Z(n5898) );
  AND U5517 ( .A(n633), .B(n5903), .Z(n5902) );
  XOR U5518 ( .A(n5904), .B(n5905), .Z(n5896) );
  AND U5519 ( .A(n637), .B(n5903), .Z(n5905) );
  XNOR U5520 ( .A(n5904), .B(n5901), .Z(n5903) );
  XOR U5521 ( .A(n5906), .B(n5907), .Z(n5901) );
  AND U5522 ( .A(n640), .B(n5908), .Z(n5907) );
  XOR U5523 ( .A(p_input[884]), .B(n5906), .Z(n5908) );
  XOR U5524 ( .A(n5909), .B(n5910), .Z(n5906) );
  AND U5525 ( .A(n644), .B(n5911), .Z(n5910) );
  XOR U5526 ( .A(n5912), .B(n5913), .Z(n5904) );
  AND U5527 ( .A(n648), .B(n5911), .Z(n5913) );
  XNOR U5528 ( .A(n5912), .B(n5909), .Z(n5911) );
  XOR U5529 ( .A(n5914), .B(n5915), .Z(n5909) );
  AND U5530 ( .A(n651), .B(n5916), .Z(n5915) );
  XOR U5531 ( .A(p_input[900]), .B(n5914), .Z(n5916) );
  XOR U5532 ( .A(n5917), .B(n5918), .Z(n5914) );
  AND U5533 ( .A(n655), .B(n5919), .Z(n5918) );
  XOR U5534 ( .A(n5920), .B(n5921), .Z(n5912) );
  AND U5535 ( .A(n659), .B(n5919), .Z(n5921) );
  XNOR U5536 ( .A(n5920), .B(n5917), .Z(n5919) );
  XOR U5537 ( .A(n5922), .B(n5923), .Z(n5917) );
  AND U5538 ( .A(n662), .B(n5924), .Z(n5923) );
  XOR U5539 ( .A(p_input[916]), .B(n5922), .Z(n5924) );
  XOR U5540 ( .A(n5925), .B(n5926), .Z(n5922) );
  AND U5541 ( .A(n666), .B(n5927), .Z(n5926) );
  XOR U5542 ( .A(n5928), .B(n5929), .Z(n5920) );
  AND U5543 ( .A(n670), .B(n5927), .Z(n5929) );
  XNOR U5544 ( .A(n5928), .B(n5925), .Z(n5927) );
  XOR U5545 ( .A(n5930), .B(n5931), .Z(n5925) );
  AND U5546 ( .A(n673), .B(n5932), .Z(n5931) );
  XOR U5547 ( .A(p_input[932]), .B(n5930), .Z(n5932) );
  XOR U5548 ( .A(n5933), .B(n5934), .Z(n5930) );
  AND U5549 ( .A(n677), .B(n5935), .Z(n5934) );
  XOR U5550 ( .A(n5936), .B(n5937), .Z(n5928) );
  AND U5551 ( .A(n681), .B(n5935), .Z(n5937) );
  XNOR U5552 ( .A(n5936), .B(n5933), .Z(n5935) );
  XOR U5553 ( .A(n5938), .B(n5939), .Z(n5933) );
  AND U5554 ( .A(n684), .B(n5940), .Z(n5939) );
  XOR U5555 ( .A(p_input[948]), .B(n5938), .Z(n5940) );
  XOR U5556 ( .A(n5941), .B(n5942), .Z(n5938) );
  AND U5557 ( .A(n688), .B(n5943), .Z(n5942) );
  XOR U5558 ( .A(n5944), .B(n5945), .Z(n5936) );
  AND U5559 ( .A(n692), .B(n5943), .Z(n5945) );
  XNOR U5560 ( .A(n5944), .B(n5941), .Z(n5943) );
  XOR U5561 ( .A(n5946), .B(n5947), .Z(n5941) );
  AND U5562 ( .A(n695), .B(n5948), .Z(n5947) );
  XOR U5563 ( .A(p_input[964]), .B(n5946), .Z(n5948) );
  XOR U5564 ( .A(n5949), .B(n5950), .Z(n5946) );
  AND U5565 ( .A(n699), .B(n5951), .Z(n5950) );
  XOR U5566 ( .A(n5952), .B(n5953), .Z(n5944) );
  AND U5567 ( .A(n703), .B(n5951), .Z(n5953) );
  XNOR U5568 ( .A(n5952), .B(n5949), .Z(n5951) );
  XOR U5569 ( .A(n5954), .B(n5955), .Z(n5949) );
  AND U5570 ( .A(n706), .B(n5956), .Z(n5955) );
  XOR U5571 ( .A(p_input[980]), .B(n5954), .Z(n5956) );
  XOR U5572 ( .A(n5957), .B(n5958), .Z(n5954) );
  AND U5573 ( .A(n710), .B(n5959), .Z(n5958) );
  XOR U5574 ( .A(n5960), .B(n5961), .Z(n5952) );
  AND U5575 ( .A(n714), .B(n5959), .Z(n5961) );
  XNOR U5576 ( .A(n5960), .B(n5957), .Z(n5959) );
  XOR U5577 ( .A(n5962), .B(n5963), .Z(n5957) );
  AND U5578 ( .A(n717), .B(n5964), .Z(n5963) );
  XOR U5579 ( .A(p_input[996]), .B(n5962), .Z(n5964) );
  XOR U5580 ( .A(n5965), .B(n5966), .Z(n5962) );
  AND U5581 ( .A(n721), .B(n5967), .Z(n5966) );
  XOR U5582 ( .A(n5968), .B(n5969), .Z(n5960) );
  AND U5583 ( .A(n725), .B(n5967), .Z(n5969) );
  XNOR U5584 ( .A(n5968), .B(n5965), .Z(n5967) );
  XOR U5585 ( .A(n5970), .B(n5971), .Z(n5965) );
  AND U5586 ( .A(n728), .B(n5972), .Z(n5971) );
  XOR U5587 ( .A(p_input[1012]), .B(n5970), .Z(n5972) );
  XOR U5588 ( .A(n5973), .B(n5974), .Z(n5970) );
  AND U5589 ( .A(n732), .B(n5975), .Z(n5974) );
  XOR U5590 ( .A(n5976), .B(n5977), .Z(n5968) );
  AND U5591 ( .A(n736), .B(n5975), .Z(n5977) );
  XNOR U5592 ( .A(n5976), .B(n5973), .Z(n5975) );
  XOR U5593 ( .A(n5978), .B(n5979), .Z(n5973) );
  AND U5594 ( .A(n739), .B(n5980), .Z(n5979) );
  XOR U5595 ( .A(p_input[1028]), .B(n5978), .Z(n5980) );
  XOR U5596 ( .A(n5981), .B(n5982), .Z(n5978) );
  AND U5597 ( .A(n743), .B(n5983), .Z(n5982) );
  XOR U5598 ( .A(n5984), .B(n5985), .Z(n5976) );
  AND U5599 ( .A(n747), .B(n5983), .Z(n5985) );
  XNOR U5600 ( .A(n5984), .B(n5981), .Z(n5983) );
  XOR U5601 ( .A(n5986), .B(n5987), .Z(n5981) );
  AND U5602 ( .A(n750), .B(n5988), .Z(n5987) );
  XOR U5603 ( .A(p_input[1044]), .B(n5986), .Z(n5988) );
  XOR U5604 ( .A(n5989), .B(n5990), .Z(n5986) );
  AND U5605 ( .A(n754), .B(n5991), .Z(n5990) );
  XOR U5606 ( .A(n5992), .B(n5993), .Z(n5984) );
  AND U5607 ( .A(n758), .B(n5991), .Z(n5993) );
  XNOR U5608 ( .A(n5992), .B(n5989), .Z(n5991) );
  XOR U5609 ( .A(n5994), .B(n5995), .Z(n5989) );
  AND U5610 ( .A(n761), .B(n5996), .Z(n5995) );
  XOR U5611 ( .A(p_input[1060]), .B(n5994), .Z(n5996) );
  XOR U5612 ( .A(n5997), .B(n5998), .Z(n5994) );
  AND U5613 ( .A(n765), .B(n5999), .Z(n5998) );
  XOR U5614 ( .A(n6000), .B(n6001), .Z(n5992) );
  AND U5615 ( .A(n769), .B(n5999), .Z(n6001) );
  XNOR U5616 ( .A(n6000), .B(n5997), .Z(n5999) );
  XOR U5617 ( .A(n6002), .B(n6003), .Z(n5997) );
  AND U5618 ( .A(n772), .B(n6004), .Z(n6003) );
  XOR U5619 ( .A(p_input[1076]), .B(n6002), .Z(n6004) );
  XOR U5620 ( .A(n6005), .B(n6006), .Z(n6002) );
  AND U5621 ( .A(n776), .B(n6007), .Z(n6006) );
  XOR U5622 ( .A(n6008), .B(n6009), .Z(n6000) );
  AND U5623 ( .A(n780), .B(n6007), .Z(n6009) );
  XNOR U5624 ( .A(n6008), .B(n6005), .Z(n6007) );
  XOR U5625 ( .A(n6010), .B(n6011), .Z(n6005) );
  AND U5626 ( .A(n783), .B(n6012), .Z(n6011) );
  XOR U5627 ( .A(p_input[1092]), .B(n6010), .Z(n6012) );
  XOR U5628 ( .A(n6013), .B(n6014), .Z(n6010) );
  AND U5629 ( .A(n787), .B(n6015), .Z(n6014) );
  XOR U5630 ( .A(n6016), .B(n6017), .Z(n6008) );
  AND U5631 ( .A(n791), .B(n6015), .Z(n6017) );
  XNOR U5632 ( .A(n6016), .B(n6013), .Z(n6015) );
  XOR U5633 ( .A(n6018), .B(n6019), .Z(n6013) );
  AND U5634 ( .A(n794), .B(n6020), .Z(n6019) );
  XOR U5635 ( .A(p_input[1108]), .B(n6018), .Z(n6020) );
  XOR U5636 ( .A(n6021), .B(n6022), .Z(n6018) );
  AND U5637 ( .A(n798), .B(n6023), .Z(n6022) );
  XOR U5638 ( .A(n6024), .B(n6025), .Z(n6016) );
  AND U5639 ( .A(n802), .B(n6023), .Z(n6025) );
  XNOR U5640 ( .A(n6024), .B(n6021), .Z(n6023) );
  XOR U5641 ( .A(n6026), .B(n6027), .Z(n6021) );
  AND U5642 ( .A(n805), .B(n6028), .Z(n6027) );
  XOR U5643 ( .A(p_input[1124]), .B(n6026), .Z(n6028) );
  XOR U5644 ( .A(n6029), .B(n6030), .Z(n6026) );
  AND U5645 ( .A(n809), .B(n6031), .Z(n6030) );
  XOR U5646 ( .A(n6032), .B(n6033), .Z(n6024) );
  AND U5647 ( .A(n813), .B(n6031), .Z(n6033) );
  XNOR U5648 ( .A(n6032), .B(n6029), .Z(n6031) );
  XOR U5649 ( .A(n6034), .B(n6035), .Z(n6029) );
  AND U5650 ( .A(n816), .B(n6036), .Z(n6035) );
  XOR U5651 ( .A(p_input[1140]), .B(n6034), .Z(n6036) );
  XOR U5652 ( .A(n6037), .B(n6038), .Z(n6034) );
  AND U5653 ( .A(n820), .B(n6039), .Z(n6038) );
  XOR U5654 ( .A(n6040), .B(n6041), .Z(n6032) );
  AND U5655 ( .A(n824), .B(n6039), .Z(n6041) );
  XNOR U5656 ( .A(n6040), .B(n6037), .Z(n6039) );
  XOR U5657 ( .A(n6042), .B(n6043), .Z(n6037) );
  AND U5658 ( .A(n827), .B(n6044), .Z(n6043) );
  XOR U5659 ( .A(p_input[1156]), .B(n6042), .Z(n6044) );
  XOR U5660 ( .A(n6045), .B(n6046), .Z(n6042) );
  AND U5661 ( .A(n831), .B(n6047), .Z(n6046) );
  XOR U5662 ( .A(n6048), .B(n6049), .Z(n6040) );
  AND U5663 ( .A(n835), .B(n6047), .Z(n6049) );
  XNOR U5664 ( .A(n6048), .B(n6045), .Z(n6047) );
  XOR U5665 ( .A(n6050), .B(n6051), .Z(n6045) );
  AND U5666 ( .A(n838), .B(n6052), .Z(n6051) );
  XOR U5667 ( .A(p_input[1172]), .B(n6050), .Z(n6052) );
  XOR U5668 ( .A(n6053), .B(n6054), .Z(n6050) );
  AND U5669 ( .A(n842), .B(n6055), .Z(n6054) );
  XOR U5670 ( .A(n6056), .B(n6057), .Z(n6048) );
  AND U5671 ( .A(n846), .B(n6055), .Z(n6057) );
  XNOR U5672 ( .A(n6056), .B(n6053), .Z(n6055) );
  XOR U5673 ( .A(n6058), .B(n6059), .Z(n6053) );
  AND U5674 ( .A(n849), .B(n6060), .Z(n6059) );
  XOR U5675 ( .A(p_input[1188]), .B(n6058), .Z(n6060) );
  XOR U5676 ( .A(n6061), .B(n6062), .Z(n6058) );
  AND U5677 ( .A(n853), .B(n6063), .Z(n6062) );
  XOR U5678 ( .A(n6064), .B(n6065), .Z(n6056) );
  AND U5679 ( .A(n857), .B(n6063), .Z(n6065) );
  XNOR U5680 ( .A(n6064), .B(n6061), .Z(n6063) );
  XOR U5681 ( .A(n6066), .B(n6067), .Z(n6061) );
  AND U5682 ( .A(n860), .B(n6068), .Z(n6067) );
  XOR U5683 ( .A(p_input[1204]), .B(n6066), .Z(n6068) );
  XOR U5684 ( .A(n6069), .B(n6070), .Z(n6066) );
  AND U5685 ( .A(n864), .B(n6071), .Z(n6070) );
  XOR U5686 ( .A(n6072), .B(n6073), .Z(n6064) );
  AND U5687 ( .A(n868), .B(n6071), .Z(n6073) );
  XNOR U5688 ( .A(n6072), .B(n6069), .Z(n6071) );
  XOR U5689 ( .A(n6074), .B(n6075), .Z(n6069) );
  AND U5690 ( .A(n871), .B(n6076), .Z(n6075) );
  XOR U5691 ( .A(p_input[1220]), .B(n6074), .Z(n6076) );
  XOR U5692 ( .A(n6077), .B(n6078), .Z(n6074) );
  AND U5693 ( .A(n875), .B(n6079), .Z(n6078) );
  XOR U5694 ( .A(n6080), .B(n6081), .Z(n6072) );
  AND U5695 ( .A(n879), .B(n6079), .Z(n6081) );
  XNOR U5696 ( .A(n6080), .B(n6077), .Z(n6079) );
  XOR U5697 ( .A(n6082), .B(n6083), .Z(n6077) );
  AND U5698 ( .A(n882), .B(n6084), .Z(n6083) );
  XOR U5699 ( .A(p_input[1236]), .B(n6082), .Z(n6084) );
  XOR U5700 ( .A(n6085), .B(n6086), .Z(n6082) );
  AND U5701 ( .A(n886), .B(n6087), .Z(n6086) );
  XOR U5702 ( .A(n6088), .B(n6089), .Z(n6080) );
  AND U5703 ( .A(n890), .B(n6087), .Z(n6089) );
  XNOR U5704 ( .A(n6088), .B(n6085), .Z(n6087) );
  XOR U5705 ( .A(n6090), .B(n6091), .Z(n6085) );
  AND U5706 ( .A(n893), .B(n6092), .Z(n6091) );
  XOR U5707 ( .A(p_input[1252]), .B(n6090), .Z(n6092) );
  XOR U5708 ( .A(n6093), .B(n6094), .Z(n6090) );
  AND U5709 ( .A(n897), .B(n6095), .Z(n6094) );
  XOR U5710 ( .A(n6096), .B(n6097), .Z(n6088) );
  AND U5711 ( .A(n901), .B(n6095), .Z(n6097) );
  XNOR U5712 ( .A(n6096), .B(n6093), .Z(n6095) );
  XOR U5713 ( .A(n6098), .B(n6099), .Z(n6093) );
  AND U5714 ( .A(n904), .B(n6100), .Z(n6099) );
  XOR U5715 ( .A(p_input[1268]), .B(n6098), .Z(n6100) );
  XOR U5716 ( .A(n6101), .B(n6102), .Z(n6098) );
  AND U5717 ( .A(n908), .B(n6103), .Z(n6102) );
  XOR U5718 ( .A(n6104), .B(n6105), .Z(n6096) );
  AND U5719 ( .A(n912), .B(n6103), .Z(n6105) );
  XNOR U5720 ( .A(n6104), .B(n6101), .Z(n6103) );
  XOR U5721 ( .A(n6106), .B(n6107), .Z(n6101) );
  AND U5722 ( .A(n915), .B(n6108), .Z(n6107) );
  XOR U5723 ( .A(p_input[1284]), .B(n6106), .Z(n6108) );
  XOR U5724 ( .A(n6109), .B(n6110), .Z(n6106) );
  AND U5725 ( .A(n919), .B(n6111), .Z(n6110) );
  XOR U5726 ( .A(n6112), .B(n6113), .Z(n6104) );
  AND U5727 ( .A(n923), .B(n6111), .Z(n6113) );
  XNOR U5728 ( .A(n6112), .B(n6109), .Z(n6111) );
  XOR U5729 ( .A(n6114), .B(n6115), .Z(n6109) );
  AND U5730 ( .A(n926), .B(n6116), .Z(n6115) );
  XOR U5731 ( .A(p_input[1300]), .B(n6114), .Z(n6116) );
  XOR U5732 ( .A(n6117), .B(n6118), .Z(n6114) );
  AND U5733 ( .A(n930), .B(n6119), .Z(n6118) );
  XOR U5734 ( .A(n6120), .B(n6121), .Z(n6112) );
  AND U5735 ( .A(n934), .B(n6119), .Z(n6121) );
  XNOR U5736 ( .A(n6120), .B(n6117), .Z(n6119) );
  XOR U5737 ( .A(n6122), .B(n6123), .Z(n6117) );
  AND U5738 ( .A(n937), .B(n6124), .Z(n6123) );
  XOR U5739 ( .A(p_input[1316]), .B(n6122), .Z(n6124) );
  XOR U5740 ( .A(n6125), .B(n6126), .Z(n6122) );
  AND U5741 ( .A(n941), .B(n6127), .Z(n6126) );
  XOR U5742 ( .A(n6128), .B(n6129), .Z(n6120) );
  AND U5743 ( .A(n945), .B(n6127), .Z(n6129) );
  XNOR U5744 ( .A(n6128), .B(n6125), .Z(n6127) );
  XOR U5745 ( .A(n6130), .B(n6131), .Z(n6125) );
  AND U5746 ( .A(n948), .B(n6132), .Z(n6131) );
  XOR U5747 ( .A(p_input[1332]), .B(n6130), .Z(n6132) );
  XOR U5748 ( .A(n6133), .B(n6134), .Z(n6130) );
  AND U5749 ( .A(n952), .B(n6135), .Z(n6134) );
  XOR U5750 ( .A(n6136), .B(n6137), .Z(n6128) );
  AND U5751 ( .A(n956), .B(n6135), .Z(n6137) );
  XNOR U5752 ( .A(n6136), .B(n6133), .Z(n6135) );
  XOR U5753 ( .A(n6138), .B(n6139), .Z(n6133) );
  AND U5754 ( .A(n959), .B(n6140), .Z(n6139) );
  XOR U5755 ( .A(p_input[1348]), .B(n6138), .Z(n6140) );
  XOR U5756 ( .A(n6141), .B(n6142), .Z(n6138) );
  AND U5757 ( .A(n963), .B(n6143), .Z(n6142) );
  XOR U5758 ( .A(n6144), .B(n6145), .Z(n6136) );
  AND U5759 ( .A(n967), .B(n6143), .Z(n6145) );
  XNOR U5760 ( .A(n6144), .B(n6141), .Z(n6143) );
  XOR U5761 ( .A(n6146), .B(n6147), .Z(n6141) );
  AND U5762 ( .A(n970), .B(n6148), .Z(n6147) );
  XOR U5763 ( .A(p_input[1364]), .B(n6146), .Z(n6148) );
  XOR U5764 ( .A(n6149), .B(n6150), .Z(n6146) );
  AND U5765 ( .A(n974), .B(n6151), .Z(n6150) );
  XOR U5766 ( .A(n6152), .B(n6153), .Z(n6144) );
  AND U5767 ( .A(n978), .B(n6151), .Z(n6153) );
  XNOR U5768 ( .A(n6152), .B(n6149), .Z(n6151) );
  XOR U5769 ( .A(n6154), .B(n6155), .Z(n6149) );
  AND U5770 ( .A(n981), .B(n6156), .Z(n6155) );
  XOR U5771 ( .A(p_input[1380]), .B(n6154), .Z(n6156) );
  XOR U5772 ( .A(n6157), .B(n6158), .Z(n6154) );
  AND U5773 ( .A(n985), .B(n6159), .Z(n6158) );
  XOR U5774 ( .A(n6160), .B(n6161), .Z(n6152) );
  AND U5775 ( .A(n989), .B(n6159), .Z(n6161) );
  XNOR U5776 ( .A(n6160), .B(n6157), .Z(n6159) );
  XOR U5777 ( .A(n6162), .B(n6163), .Z(n6157) );
  AND U5778 ( .A(n992), .B(n6164), .Z(n6163) );
  XOR U5779 ( .A(p_input[1396]), .B(n6162), .Z(n6164) );
  XOR U5780 ( .A(n6165), .B(n6166), .Z(n6162) );
  AND U5781 ( .A(n996), .B(n6167), .Z(n6166) );
  XOR U5782 ( .A(n6168), .B(n6169), .Z(n6160) );
  AND U5783 ( .A(n1000), .B(n6167), .Z(n6169) );
  XNOR U5784 ( .A(n6168), .B(n6165), .Z(n6167) );
  XOR U5785 ( .A(n6170), .B(n6171), .Z(n6165) );
  AND U5786 ( .A(n1003), .B(n6172), .Z(n6171) );
  XOR U5787 ( .A(p_input[1412]), .B(n6170), .Z(n6172) );
  XOR U5788 ( .A(n6173), .B(n6174), .Z(n6170) );
  AND U5789 ( .A(n1007), .B(n6175), .Z(n6174) );
  XOR U5790 ( .A(n6176), .B(n6177), .Z(n6168) );
  AND U5791 ( .A(n1011), .B(n6175), .Z(n6177) );
  XNOR U5792 ( .A(n6176), .B(n6173), .Z(n6175) );
  XOR U5793 ( .A(n6178), .B(n6179), .Z(n6173) );
  AND U5794 ( .A(n1014), .B(n6180), .Z(n6179) );
  XOR U5795 ( .A(p_input[1428]), .B(n6178), .Z(n6180) );
  XOR U5796 ( .A(n6181), .B(n6182), .Z(n6178) );
  AND U5797 ( .A(n1018), .B(n6183), .Z(n6182) );
  XOR U5798 ( .A(n6184), .B(n6185), .Z(n6176) );
  AND U5799 ( .A(n1022), .B(n6183), .Z(n6185) );
  XNOR U5800 ( .A(n6184), .B(n6181), .Z(n6183) );
  XOR U5801 ( .A(n6186), .B(n6187), .Z(n6181) );
  AND U5802 ( .A(n1025), .B(n6188), .Z(n6187) );
  XOR U5803 ( .A(p_input[1444]), .B(n6186), .Z(n6188) );
  XOR U5804 ( .A(n6189), .B(n6190), .Z(n6186) );
  AND U5805 ( .A(n1029), .B(n6191), .Z(n6190) );
  XOR U5806 ( .A(n6192), .B(n6193), .Z(n6184) );
  AND U5807 ( .A(n1033), .B(n6191), .Z(n6193) );
  XNOR U5808 ( .A(n6192), .B(n6189), .Z(n6191) );
  XOR U5809 ( .A(n6194), .B(n6195), .Z(n6189) );
  AND U5810 ( .A(n1036), .B(n6196), .Z(n6195) );
  XOR U5811 ( .A(p_input[1460]), .B(n6194), .Z(n6196) );
  XOR U5812 ( .A(n6197), .B(n6198), .Z(n6194) );
  AND U5813 ( .A(n1040), .B(n6199), .Z(n6198) );
  XOR U5814 ( .A(n6200), .B(n6201), .Z(n6192) );
  AND U5815 ( .A(n1044), .B(n6199), .Z(n6201) );
  XNOR U5816 ( .A(n6200), .B(n6197), .Z(n6199) );
  XOR U5817 ( .A(n6202), .B(n6203), .Z(n6197) );
  AND U5818 ( .A(n1047), .B(n6204), .Z(n6203) );
  XOR U5819 ( .A(p_input[1476]), .B(n6202), .Z(n6204) );
  XOR U5820 ( .A(n6205), .B(n6206), .Z(n6202) );
  AND U5821 ( .A(n1051), .B(n6207), .Z(n6206) );
  XOR U5822 ( .A(n6208), .B(n6209), .Z(n6200) );
  AND U5823 ( .A(n1055), .B(n6207), .Z(n6209) );
  XNOR U5824 ( .A(n6208), .B(n6205), .Z(n6207) );
  XOR U5825 ( .A(n6210), .B(n6211), .Z(n6205) );
  AND U5826 ( .A(n1058), .B(n6212), .Z(n6211) );
  XOR U5827 ( .A(p_input[1492]), .B(n6210), .Z(n6212) );
  XOR U5828 ( .A(n6213), .B(n6214), .Z(n6210) );
  AND U5829 ( .A(n1062), .B(n6215), .Z(n6214) );
  XOR U5830 ( .A(n6216), .B(n6217), .Z(n6208) );
  AND U5831 ( .A(n1066), .B(n6215), .Z(n6217) );
  XNOR U5832 ( .A(n6216), .B(n6213), .Z(n6215) );
  XOR U5833 ( .A(n6218), .B(n6219), .Z(n6213) );
  AND U5834 ( .A(n1069), .B(n6220), .Z(n6219) );
  XOR U5835 ( .A(p_input[1508]), .B(n6218), .Z(n6220) );
  XOR U5836 ( .A(n6221), .B(n6222), .Z(n6218) );
  AND U5837 ( .A(n1073), .B(n6223), .Z(n6222) );
  XOR U5838 ( .A(n6224), .B(n6225), .Z(n6216) );
  AND U5839 ( .A(n1077), .B(n6223), .Z(n6225) );
  XNOR U5840 ( .A(n6224), .B(n6221), .Z(n6223) );
  XOR U5841 ( .A(n6226), .B(n6227), .Z(n6221) );
  AND U5842 ( .A(n1080), .B(n6228), .Z(n6227) );
  XOR U5843 ( .A(p_input[1524]), .B(n6226), .Z(n6228) );
  XOR U5844 ( .A(n6229), .B(n6230), .Z(n6226) );
  AND U5845 ( .A(n1084), .B(n6231), .Z(n6230) );
  XOR U5846 ( .A(n6232), .B(n6233), .Z(n6224) );
  AND U5847 ( .A(n1088), .B(n6231), .Z(n6233) );
  XNOR U5848 ( .A(n6232), .B(n6229), .Z(n6231) );
  XOR U5849 ( .A(n6234), .B(n6235), .Z(n6229) );
  AND U5850 ( .A(n1091), .B(n6236), .Z(n6235) );
  XOR U5851 ( .A(p_input[1540]), .B(n6234), .Z(n6236) );
  XOR U5852 ( .A(n6237), .B(n6238), .Z(n6234) );
  AND U5853 ( .A(n1095), .B(n6239), .Z(n6238) );
  XOR U5854 ( .A(n6240), .B(n6241), .Z(n6232) );
  AND U5855 ( .A(n1099), .B(n6239), .Z(n6241) );
  XNOR U5856 ( .A(n6240), .B(n6237), .Z(n6239) );
  XOR U5857 ( .A(n6242), .B(n6243), .Z(n6237) );
  AND U5858 ( .A(n1102), .B(n6244), .Z(n6243) );
  XOR U5859 ( .A(p_input[1556]), .B(n6242), .Z(n6244) );
  XOR U5860 ( .A(n6245), .B(n6246), .Z(n6242) );
  AND U5861 ( .A(n1106), .B(n6247), .Z(n6246) );
  XOR U5862 ( .A(n6248), .B(n6249), .Z(n6240) );
  AND U5863 ( .A(n1110), .B(n6247), .Z(n6249) );
  XNOR U5864 ( .A(n6248), .B(n6245), .Z(n6247) );
  XOR U5865 ( .A(n6250), .B(n6251), .Z(n6245) );
  AND U5866 ( .A(n1113), .B(n6252), .Z(n6251) );
  XOR U5867 ( .A(p_input[1572]), .B(n6250), .Z(n6252) );
  XOR U5868 ( .A(n6253), .B(n6254), .Z(n6250) );
  AND U5869 ( .A(n1117), .B(n6255), .Z(n6254) );
  XOR U5870 ( .A(n6256), .B(n6257), .Z(n6248) );
  AND U5871 ( .A(n1121), .B(n6255), .Z(n6257) );
  XNOR U5872 ( .A(n6256), .B(n6253), .Z(n6255) );
  XOR U5873 ( .A(n6258), .B(n6259), .Z(n6253) );
  AND U5874 ( .A(n1124), .B(n6260), .Z(n6259) );
  XOR U5875 ( .A(p_input[1588]), .B(n6258), .Z(n6260) );
  XOR U5876 ( .A(n6261), .B(n6262), .Z(n6258) );
  AND U5877 ( .A(n1128), .B(n6263), .Z(n6262) );
  XOR U5878 ( .A(n6264), .B(n6265), .Z(n6256) );
  AND U5879 ( .A(n1132), .B(n6263), .Z(n6265) );
  XNOR U5880 ( .A(n6264), .B(n6261), .Z(n6263) );
  XOR U5881 ( .A(n6266), .B(n6267), .Z(n6261) );
  AND U5882 ( .A(n1135), .B(n6268), .Z(n6267) );
  XOR U5883 ( .A(p_input[1604]), .B(n6266), .Z(n6268) );
  XOR U5884 ( .A(n6269), .B(n6270), .Z(n6266) );
  AND U5885 ( .A(n1139), .B(n6271), .Z(n6270) );
  XOR U5886 ( .A(n6272), .B(n6273), .Z(n6264) );
  AND U5887 ( .A(n1143), .B(n6271), .Z(n6273) );
  XNOR U5888 ( .A(n6272), .B(n6269), .Z(n6271) );
  XOR U5889 ( .A(n6274), .B(n6275), .Z(n6269) );
  AND U5890 ( .A(n1146), .B(n6276), .Z(n6275) );
  XOR U5891 ( .A(p_input[1620]), .B(n6274), .Z(n6276) );
  XOR U5892 ( .A(n6277), .B(n6278), .Z(n6274) );
  AND U5893 ( .A(n1150), .B(n6279), .Z(n6278) );
  XOR U5894 ( .A(n6280), .B(n6281), .Z(n6272) );
  AND U5895 ( .A(n1154), .B(n6279), .Z(n6281) );
  XNOR U5896 ( .A(n6280), .B(n6277), .Z(n6279) );
  XOR U5897 ( .A(n6282), .B(n6283), .Z(n6277) );
  AND U5898 ( .A(n1157), .B(n6284), .Z(n6283) );
  XOR U5899 ( .A(p_input[1636]), .B(n6282), .Z(n6284) );
  XOR U5900 ( .A(n6285), .B(n6286), .Z(n6282) );
  AND U5901 ( .A(n1161), .B(n6287), .Z(n6286) );
  XOR U5902 ( .A(n6288), .B(n6289), .Z(n6280) );
  AND U5903 ( .A(n1165), .B(n6287), .Z(n6289) );
  XNOR U5904 ( .A(n6288), .B(n6285), .Z(n6287) );
  XOR U5905 ( .A(n6290), .B(n6291), .Z(n6285) );
  AND U5906 ( .A(n1168), .B(n6292), .Z(n6291) );
  XOR U5907 ( .A(p_input[1652]), .B(n6290), .Z(n6292) );
  XOR U5908 ( .A(n6293), .B(n6294), .Z(n6290) );
  AND U5909 ( .A(n1172), .B(n6295), .Z(n6294) );
  XOR U5910 ( .A(n6296), .B(n6297), .Z(n6288) );
  AND U5911 ( .A(n1176), .B(n6295), .Z(n6297) );
  XNOR U5912 ( .A(n6296), .B(n6293), .Z(n6295) );
  XOR U5913 ( .A(n6298), .B(n6299), .Z(n6293) );
  AND U5914 ( .A(n1179), .B(n6300), .Z(n6299) );
  XOR U5915 ( .A(p_input[1668]), .B(n6298), .Z(n6300) );
  XOR U5916 ( .A(n6301), .B(n6302), .Z(n6298) );
  AND U5917 ( .A(n1183), .B(n6303), .Z(n6302) );
  XOR U5918 ( .A(n6304), .B(n6305), .Z(n6296) );
  AND U5919 ( .A(n1187), .B(n6303), .Z(n6305) );
  XNOR U5920 ( .A(n6304), .B(n6301), .Z(n6303) );
  XOR U5921 ( .A(n6306), .B(n6307), .Z(n6301) );
  AND U5922 ( .A(n1190), .B(n6308), .Z(n6307) );
  XOR U5923 ( .A(p_input[1684]), .B(n6306), .Z(n6308) );
  XOR U5924 ( .A(n6309), .B(n6310), .Z(n6306) );
  AND U5925 ( .A(n1194), .B(n6311), .Z(n6310) );
  XOR U5926 ( .A(n6312), .B(n6313), .Z(n6304) );
  AND U5927 ( .A(n1198), .B(n6311), .Z(n6313) );
  XNOR U5928 ( .A(n6312), .B(n6309), .Z(n6311) );
  XOR U5929 ( .A(n6314), .B(n6315), .Z(n6309) );
  AND U5930 ( .A(n1201), .B(n6316), .Z(n6315) );
  XOR U5931 ( .A(p_input[1700]), .B(n6314), .Z(n6316) );
  XOR U5932 ( .A(n6317), .B(n6318), .Z(n6314) );
  AND U5933 ( .A(n1205), .B(n6319), .Z(n6318) );
  XOR U5934 ( .A(n6320), .B(n6321), .Z(n6312) );
  AND U5935 ( .A(n1209), .B(n6319), .Z(n6321) );
  XNOR U5936 ( .A(n6320), .B(n6317), .Z(n6319) );
  XOR U5937 ( .A(n6322), .B(n6323), .Z(n6317) );
  AND U5938 ( .A(n1212), .B(n6324), .Z(n6323) );
  XOR U5939 ( .A(p_input[1716]), .B(n6322), .Z(n6324) );
  XOR U5940 ( .A(n6325), .B(n6326), .Z(n6322) );
  AND U5941 ( .A(n1216), .B(n6327), .Z(n6326) );
  XOR U5942 ( .A(n6328), .B(n6329), .Z(n6320) );
  AND U5943 ( .A(n1220), .B(n6327), .Z(n6329) );
  XNOR U5944 ( .A(n6328), .B(n6325), .Z(n6327) );
  XOR U5945 ( .A(n6330), .B(n6331), .Z(n6325) );
  AND U5946 ( .A(n1223), .B(n6332), .Z(n6331) );
  XOR U5947 ( .A(p_input[1732]), .B(n6330), .Z(n6332) );
  XOR U5948 ( .A(n6333), .B(n6334), .Z(n6330) );
  AND U5949 ( .A(n1227), .B(n6335), .Z(n6334) );
  XOR U5950 ( .A(n6336), .B(n6337), .Z(n6328) );
  AND U5951 ( .A(n1231), .B(n6335), .Z(n6337) );
  XNOR U5952 ( .A(n6336), .B(n6333), .Z(n6335) );
  XOR U5953 ( .A(n6338), .B(n6339), .Z(n6333) );
  AND U5954 ( .A(n1234), .B(n6340), .Z(n6339) );
  XOR U5955 ( .A(p_input[1748]), .B(n6338), .Z(n6340) );
  XOR U5956 ( .A(n6341), .B(n6342), .Z(n6338) );
  AND U5957 ( .A(n1238), .B(n6343), .Z(n6342) );
  XOR U5958 ( .A(n6344), .B(n6345), .Z(n6336) );
  AND U5959 ( .A(n1242), .B(n6343), .Z(n6345) );
  XNOR U5960 ( .A(n6344), .B(n6341), .Z(n6343) );
  XOR U5961 ( .A(n6346), .B(n6347), .Z(n6341) );
  AND U5962 ( .A(n1245), .B(n6348), .Z(n6347) );
  XOR U5963 ( .A(p_input[1764]), .B(n6346), .Z(n6348) );
  XOR U5964 ( .A(n6349), .B(n6350), .Z(n6346) );
  AND U5965 ( .A(n1249), .B(n6351), .Z(n6350) );
  XOR U5966 ( .A(n6352), .B(n6353), .Z(n6344) );
  AND U5967 ( .A(n1253), .B(n6351), .Z(n6353) );
  XNOR U5968 ( .A(n6352), .B(n6349), .Z(n6351) );
  XOR U5969 ( .A(n6354), .B(n6355), .Z(n6349) );
  AND U5970 ( .A(n1256), .B(n6356), .Z(n6355) );
  XOR U5971 ( .A(p_input[1780]), .B(n6354), .Z(n6356) );
  XOR U5972 ( .A(n6357), .B(n6358), .Z(n6354) );
  AND U5973 ( .A(n1260), .B(n6359), .Z(n6358) );
  XOR U5974 ( .A(n6360), .B(n6361), .Z(n6352) );
  AND U5975 ( .A(n1264), .B(n6359), .Z(n6361) );
  XNOR U5976 ( .A(n6360), .B(n6357), .Z(n6359) );
  XOR U5977 ( .A(n6362), .B(n6363), .Z(n6357) );
  AND U5978 ( .A(n1267), .B(n6364), .Z(n6363) );
  XOR U5979 ( .A(p_input[1796]), .B(n6362), .Z(n6364) );
  XOR U5980 ( .A(n6365), .B(n6366), .Z(n6362) );
  AND U5981 ( .A(n1271), .B(n6367), .Z(n6366) );
  XOR U5982 ( .A(n6368), .B(n6369), .Z(n6360) );
  AND U5983 ( .A(n1275), .B(n6367), .Z(n6369) );
  XNOR U5984 ( .A(n6368), .B(n6365), .Z(n6367) );
  XOR U5985 ( .A(n6370), .B(n6371), .Z(n6365) );
  AND U5986 ( .A(n1278), .B(n6372), .Z(n6371) );
  XOR U5987 ( .A(p_input[1812]), .B(n6370), .Z(n6372) );
  XOR U5988 ( .A(n6373), .B(n6374), .Z(n6370) );
  AND U5989 ( .A(n1282), .B(n6375), .Z(n6374) );
  XOR U5990 ( .A(n6376), .B(n6377), .Z(n6368) );
  AND U5991 ( .A(n1286), .B(n6375), .Z(n6377) );
  XNOR U5992 ( .A(n6376), .B(n6373), .Z(n6375) );
  XOR U5993 ( .A(n6378), .B(n6379), .Z(n6373) );
  AND U5994 ( .A(n1289), .B(n6380), .Z(n6379) );
  XOR U5995 ( .A(p_input[1828]), .B(n6378), .Z(n6380) );
  XOR U5996 ( .A(n6381), .B(n6382), .Z(n6378) );
  AND U5997 ( .A(n1293), .B(n6383), .Z(n6382) );
  XOR U5998 ( .A(n6384), .B(n6385), .Z(n6376) );
  AND U5999 ( .A(n1297), .B(n6383), .Z(n6385) );
  XNOR U6000 ( .A(n6384), .B(n6381), .Z(n6383) );
  XOR U6001 ( .A(n6386), .B(n6387), .Z(n6381) );
  AND U6002 ( .A(n1300), .B(n6388), .Z(n6387) );
  XOR U6003 ( .A(p_input[1844]), .B(n6386), .Z(n6388) );
  XOR U6004 ( .A(n6389), .B(n6390), .Z(n6386) );
  AND U6005 ( .A(n1304), .B(n6391), .Z(n6390) );
  XOR U6006 ( .A(n6392), .B(n6393), .Z(n6384) );
  AND U6007 ( .A(n1308), .B(n6391), .Z(n6393) );
  XNOR U6008 ( .A(n6392), .B(n6389), .Z(n6391) );
  XOR U6009 ( .A(n6394), .B(n6395), .Z(n6389) );
  AND U6010 ( .A(n1311), .B(n6396), .Z(n6395) );
  XOR U6011 ( .A(p_input[1860]), .B(n6394), .Z(n6396) );
  XOR U6012 ( .A(n6397), .B(n6398), .Z(n6394) );
  AND U6013 ( .A(n1315), .B(n6399), .Z(n6398) );
  XOR U6014 ( .A(n6400), .B(n6401), .Z(n6392) );
  AND U6015 ( .A(n1319), .B(n6399), .Z(n6401) );
  XNOR U6016 ( .A(n6400), .B(n6397), .Z(n6399) );
  XOR U6017 ( .A(n6402), .B(n6403), .Z(n6397) );
  AND U6018 ( .A(n1322), .B(n6404), .Z(n6403) );
  XOR U6019 ( .A(p_input[1876]), .B(n6402), .Z(n6404) );
  XOR U6020 ( .A(n6405), .B(n6406), .Z(n6402) );
  AND U6021 ( .A(n1326), .B(n6407), .Z(n6406) );
  XOR U6022 ( .A(n6408), .B(n6409), .Z(n6400) );
  AND U6023 ( .A(n1330), .B(n6407), .Z(n6409) );
  XNOR U6024 ( .A(n6408), .B(n6405), .Z(n6407) );
  XOR U6025 ( .A(n6410), .B(n6411), .Z(n6405) );
  AND U6026 ( .A(n1333), .B(n6412), .Z(n6411) );
  XOR U6027 ( .A(p_input[1892]), .B(n6410), .Z(n6412) );
  XOR U6028 ( .A(n6413), .B(n6414), .Z(n6410) );
  AND U6029 ( .A(n1337), .B(n6415), .Z(n6414) );
  XOR U6030 ( .A(n6416), .B(n6417), .Z(n6408) );
  AND U6031 ( .A(n1341), .B(n6415), .Z(n6417) );
  XNOR U6032 ( .A(n6416), .B(n6413), .Z(n6415) );
  XOR U6033 ( .A(n6418), .B(n6419), .Z(n6413) );
  AND U6034 ( .A(n1344), .B(n6420), .Z(n6419) );
  XOR U6035 ( .A(p_input[1908]), .B(n6418), .Z(n6420) );
  XOR U6036 ( .A(n6421), .B(n6422), .Z(n6418) );
  AND U6037 ( .A(n1348), .B(n6423), .Z(n6422) );
  XOR U6038 ( .A(n6424), .B(n6425), .Z(n6416) );
  AND U6039 ( .A(n1352), .B(n6423), .Z(n6425) );
  XNOR U6040 ( .A(n6424), .B(n6421), .Z(n6423) );
  XOR U6041 ( .A(n6426), .B(n6427), .Z(n6421) );
  AND U6042 ( .A(n1355), .B(n6428), .Z(n6427) );
  XOR U6043 ( .A(p_input[1924]), .B(n6426), .Z(n6428) );
  XOR U6044 ( .A(n6429), .B(n6430), .Z(n6426) );
  AND U6045 ( .A(n1359), .B(n6431), .Z(n6430) );
  XOR U6046 ( .A(n6432), .B(n6433), .Z(n6424) );
  AND U6047 ( .A(n1363), .B(n6431), .Z(n6433) );
  XNOR U6048 ( .A(n6432), .B(n6429), .Z(n6431) );
  XOR U6049 ( .A(n6434), .B(n6435), .Z(n6429) );
  AND U6050 ( .A(n1366), .B(n6436), .Z(n6435) );
  XOR U6051 ( .A(p_input[1940]), .B(n6434), .Z(n6436) );
  XOR U6052 ( .A(n6437), .B(n6438), .Z(n6434) );
  AND U6053 ( .A(n1370), .B(n6439), .Z(n6438) );
  XOR U6054 ( .A(n6440), .B(n6441), .Z(n6432) );
  AND U6055 ( .A(n1374), .B(n6439), .Z(n6441) );
  XNOR U6056 ( .A(n6440), .B(n6437), .Z(n6439) );
  XOR U6057 ( .A(n6442), .B(n6443), .Z(n6437) );
  AND U6058 ( .A(n1377), .B(n6444), .Z(n6443) );
  XOR U6059 ( .A(p_input[1956]), .B(n6442), .Z(n6444) );
  XOR U6060 ( .A(n6445), .B(n6446), .Z(n6442) );
  AND U6061 ( .A(n1381), .B(n6447), .Z(n6446) );
  XOR U6062 ( .A(n6448), .B(n6449), .Z(n6440) );
  AND U6063 ( .A(n1385), .B(n6447), .Z(n6449) );
  XNOR U6064 ( .A(n6448), .B(n6445), .Z(n6447) );
  XOR U6065 ( .A(n6450), .B(n6451), .Z(n6445) );
  AND U6066 ( .A(n1388), .B(n6452), .Z(n6451) );
  XOR U6067 ( .A(p_input[1972]), .B(n6450), .Z(n6452) );
  XOR U6068 ( .A(n6453), .B(n6454), .Z(n6450) );
  AND U6069 ( .A(n1392), .B(n6455), .Z(n6454) );
  XOR U6070 ( .A(n6456), .B(n6457), .Z(n6448) );
  AND U6071 ( .A(n1396), .B(n6455), .Z(n6457) );
  XNOR U6072 ( .A(n6456), .B(n6453), .Z(n6455) );
  XOR U6073 ( .A(n6458), .B(n6459), .Z(n6453) );
  AND U6074 ( .A(n1399), .B(n6460), .Z(n6459) );
  XOR U6075 ( .A(p_input[1988]), .B(n6458), .Z(n6460) );
  XOR U6076 ( .A(n6461), .B(n6462), .Z(n6458) );
  AND U6077 ( .A(n1403), .B(n6463), .Z(n6462) );
  XOR U6078 ( .A(n6464), .B(n6465), .Z(n6456) );
  AND U6079 ( .A(n1407), .B(n6463), .Z(n6465) );
  XNOR U6080 ( .A(n6464), .B(n6461), .Z(n6463) );
  XOR U6081 ( .A(n6466), .B(n6467), .Z(n6461) );
  AND U6082 ( .A(n1410), .B(n6468), .Z(n6467) );
  XOR U6083 ( .A(p_input[2004]), .B(n6466), .Z(n6468) );
  XNOR U6084 ( .A(n6469), .B(n6470), .Z(n6466) );
  AND U6085 ( .A(n1414), .B(n6471), .Z(n6470) );
  XNOR U6086 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n6472), .Z(n6464) );
  AND U6087 ( .A(n1417), .B(n6471), .Z(n6472) );
  XOR U6088 ( .A(n6473), .B(n6469), .Z(n6471) );
  IV U6089 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .Z(n6469) );
  IV U6090 ( .A(\knn_comb_/min_val_out[0][4] ), .Z(n6473) );
  XOR U6091 ( .A(n6474), .B(n6475), .Z(o[1]) );
  XOR U6092 ( .A(n13), .B(n6476), .Z(o[19]) );
  AND U6093 ( .A(n30), .B(n6477), .Z(n13) );
  XOR U6094 ( .A(n14), .B(n6476), .Z(n6477) );
  XOR U6095 ( .A(n6478), .B(n6479), .Z(n6476) );
  AND U6096 ( .A(n34), .B(n6480), .Z(n6479) );
  XOR U6097 ( .A(p_input[3]), .B(n6478), .Z(n6480) );
  XOR U6098 ( .A(n6481), .B(n6482), .Z(n6478) );
  AND U6099 ( .A(n38), .B(n6483), .Z(n6482) );
  XOR U6100 ( .A(n6484), .B(n6485), .Z(n14) );
  AND U6101 ( .A(n42), .B(n6483), .Z(n6485) );
  XNOR U6102 ( .A(n6486), .B(n6481), .Z(n6483) );
  XOR U6103 ( .A(n6487), .B(n6488), .Z(n6481) );
  AND U6104 ( .A(n46), .B(n6489), .Z(n6488) );
  XOR U6105 ( .A(p_input[19]), .B(n6487), .Z(n6489) );
  XOR U6106 ( .A(n6490), .B(n6491), .Z(n6487) );
  AND U6107 ( .A(n50), .B(n6492), .Z(n6491) );
  IV U6108 ( .A(n6484), .Z(n6486) );
  XNOR U6109 ( .A(n6493), .B(n6494), .Z(n6484) );
  AND U6110 ( .A(n54), .B(n6492), .Z(n6494) );
  XNOR U6111 ( .A(n6493), .B(n6490), .Z(n6492) );
  XOR U6112 ( .A(n6495), .B(n6496), .Z(n6490) );
  AND U6113 ( .A(n57), .B(n6497), .Z(n6496) );
  XOR U6114 ( .A(p_input[35]), .B(n6495), .Z(n6497) );
  XOR U6115 ( .A(n6498), .B(n6499), .Z(n6495) );
  AND U6116 ( .A(n61), .B(n6500), .Z(n6499) );
  XOR U6117 ( .A(n6501), .B(n6502), .Z(n6493) );
  AND U6118 ( .A(n65), .B(n6500), .Z(n6502) );
  XNOR U6119 ( .A(n6501), .B(n6498), .Z(n6500) );
  XOR U6120 ( .A(n6503), .B(n6504), .Z(n6498) );
  AND U6121 ( .A(n68), .B(n6505), .Z(n6504) );
  XOR U6122 ( .A(p_input[51]), .B(n6503), .Z(n6505) );
  XOR U6123 ( .A(n6506), .B(n6507), .Z(n6503) );
  AND U6124 ( .A(n72), .B(n6508), .Z(n6507) );
  XOR U6125 ( .A(n6509), .B(n6510), .Z(n6501) );
  AND U6126 ( .A(n76), .B(n6508), .Z(n6510) );
  XNOR U6127 ( .A(n6509), .B(n6506), .Z(n6508) );
  XOR U6128 ( .A(n6511), .B(n6512), .Z(n6506) );
  AND U6129 ( .A(n79), .B(n6513), .Z(n6512) );
  XOR U6130 ( .A(p_input[67]), .B(n6511), .Z(n6513) );
  XOR U6131 ( .A(n6514), .B(n6515), .Z(n6511) );
  AND U6132 ( .A(n83), .B(n6516), .Z(n6515) );
  XOR U6133 ( .A(n6517), .B(n6518), .Z(n6509) );
  AND U6134 ( .A(n87), .B(n6516), .Z(n6518) );
  XNOR U6135 ( .A(n6517), .B(n6514), .Z(n6516) );
  XOR U6136 ( .A(n6519), .B(n6520), .Z(n6514) );
  AND U6137 ( .A(n90), .B(n6521), .Z(n6520) );
  XOR U6138 ( .A(p_input[83]), .B(n6519), .Z(n6521) );
  XOR U6139 ( .A(n6522), .B(n6523), .Z(n6519) );
  AND U6140 ( .A(n94), .B(n6524), .Z(n6523) );
  XOR U6141 ( .A(n6525), .B(n6526), .Z(n6517) );
  AND U6142 ( .A(n98), .B(n6524), .Z(n6526) );
  XNOR U6143 ( .A(n6525), .B(n6522), .Z(n6524) );
  XOR U6144 ( .A(n6527), .B(n6528), .Z(n6522) );
  AND U6145 ( .A(n101), .B(n6529), .Z(n6528) );
  XOR U6146 ( .A(p_input[99]), .B(n6527), .Z(n6529) );
  XOR U6147 ( .A(n6530), .B(n6531), .Z(n6527) );
  AND U6148 ( .A(n105), .B(n6532), .Z(n6531) );
  XOR U6149 ( .A(n6533), .B(n6534), .Z(n6525) );
  AND U6150 ( .A(n109), .B(n6532), .Z(n6534) );
  XNOR U6151 ( .A(n6533), .B(n6530), .Z(n6532) );
  XOR U6152 ( .A(n6535), .B(n6536), .Z(n6530) );
  AND U6153 ( .A(n112), .B(n6537), .Z(n6536) );
  XOR U6154 ( .A(p_input[115]), .B(n6535), .Z(n6537) );
  XOR U6155 ( .A(n6538), .B(n6539), .Z(n6535) );
  AND U6156 ( .A(n116), .B(n6540), .Z(n6539) );
  XOR U6157 ( .A(n6541), .B(n6542), .Z(n6533) );
  AND U6158 ( .A(n120), .B(n6540), .Z(n6542) );
  XNOR U6159 ( .A(n6541), .B(n6538), .Z(n6540) );
  XOR U6160 ( .A(n6543), .B(n6544), .Z(n6538) );
  AND U6161 ( .A(n123), .B(n6545), .Z(n6544) );
  XOR U6162 ( .A(p_input[131]), .B(n6543), .Z(n6545) );
  XOR U6163 ( .A(n6546), .B(n6547), .Z(n6543) );
  AND U6164 ( .A(n127), .B(n6548), .Z(n6547) );
  XOR U6165 ( .A(n6549), .B(n6550), .Z(n6541) );
  AND U6166 ( .A(n131), .B(n6548), .Z(n6550) );
  XNOR U6167 ( .A(n6549), .B(n6546), .Z(n6548) );
  XOR U6168 ( .A(n6551), .B(n6552), .Z(n6546) );
  AND U6169 ( .A(n134), .B(n6553), .Z(n6552) );
  XOR U6170 ( .A(p_input[147]), .B(n6551), .Z(n6553) );
  XOR U6171 ( .A(n6554), .B(n6555), .Z(n6551) );
  AND U6172 ( .A(n138), .B(n6556), .Z(n6555) );
  XOR U6173 ( .A(n6557), .B(n6558), .Z(n6549) );
  AND U6174 ( .A(n142), .B(n6556), .Z(n6558) );
  XNOR U6175 ( .A(n6557), .B(n6554), .Z(n6556) );
  XOR U6176 ( .A(n6559), .B(n6560), .Z(n6554) );
  AND U6177 ( .A(n145), .B(n6561), .Z(n6560) );
  XOR U6178 ( .A(p_input[163]), .B(n6559), .Z(n6561) );
  XOR U6179 ( .A(n6562), .B(n6563), .Z(n6559) );
  AND U6180 ( .A(n149), .B(n6564), .Z(n6563) );
  XOR U6181 ( .A(n6565), .B(n6566), .Z(n6557) );
  AND U6182 ( .A(n153), .B(n6564), .Z(n6566) );
  XNOR U6183 ( .A(n6565), .B(n6562), .Z(n6564) );
  XOR U6184 ( .A(n6567), .B(n6568), .Z(n6562) );
  AND U6185 ( .A(n156), .B(n6569), .Z(n6568) );
  XOR U6186 ( .A(p_input[179]), .B(n6567), .Z(n6569) );
  XOR U6187 ( .A(n6570), .B(n6571), .Z(n6567) );
  AND U6188 ( .A(n160), .B(n6572), .Z(n6571) );
  XOR U6189 ( .A(n6573), .B(n6574), .Z(n6565) );
  AND U6190 ( .A(n164), .B(n6572), .Z(n6574) );
  XNOR U6191 ( .A(n6573), .B(n6570), .Z(n6572) );
  XOR U6192 ( .A(n6575), .B(n6576), .Z(n6570) );
  AND U6193 ( .A(n167), .B(n6577), .Z(n6576) );
  XOR U6194 ( .A(p_input[195]), .B(n6575), .Z(n6577) );
  XOR U6195 ( .A(n6578), .B(n6579), .Z(n6575) );
  AND U6196 ( .A(n171), .B(n6580), .Z(n6579) );
  XOR U6197 ( .A(n6581), .B(n6582), .Z(n6573) );
  AND U6198 ( .A(n175), .B(n6580), .Z(n6582) );
  XNOR U6199 ( .A(n6581), .B(n6578), .Z(n6580) );
  XOR U6200 ( .A(n6583), .B(n6584), .Z(n6578) );
  AND U6201 ( .A(n178), .B(n6585), .Z(n6584) );
  XOR U6202 ( .A(p_input[211]), .B(n6583), .Z(n6585) );
  XOR U6203 ( .A(n6586), .B(n6587), .Z(n6583) );
  AND U6204 ( .A(n182), .B(n6588), .Z(n6587) );
  XOR U6205 ( .A(n6589), .B(n6590), .Z(n6581) );
  AND U6206 ( .A(n186), .B(n6588), .Z(n6590) );
  XNOR U6207 ( .A(n6589), .B(n6586), .Z(n6588) );
  XOR U6208 ( .A(n6591), .B(n6592), .Z(n6586) );
  AND U6209 ( .A(n189), .B(n6593), .Z(n6592) );
  XOR U6210 ( .A(p_input[227]), .B(n6591), .Z(n6593) );
  XOR U6211 ( .A(n6594), .B(n6595), .Z(n6591) );
  AND U6212 ( .A(n193), .B(n6596), .Z(n6595) );
  XOR U6213 ( .A(n6597), .B(n6598), .Z(n6589) );
  AND U6214 ( .A(n197), .B(n6596), .Z(n6598) );
  XNOR U6215 ( .A(n6597), .B(n6594), .Z(n6596) );
  XOR U6216 ( .A(n6599), .B(n6600), .Z(n6594) );
  AND U6217 ( .A(n200), .B(n6601), .Z(n6600) );
  XOR U6218 ( .A(p_input[243]), .B(n6599), .Z(n6601) );
  XOR U6219 ( .A(n6602), .B(n6603), .Z(n6599) );
  AND U6220 ( .A(n204), .B(n6604), .Z(n6603) );
  XOR U6221 ( .A(n6605), .B(n6606), .Z(n6597) );
  AND U6222 ( .A(n208), .B(n6604), .Z(n6606) );
  XNOR U6223 ( .A(n6605), .B(n6602), .Z(n6604) );
  XOR U6224 ( .A(n6607), .B(n6608), .Z(n6602) );
  AND U6225 ( .A(n211), .B(n6609), .Z(n6608) );
  XOR U6226 ( .A(p_input[259]), .B(n6607), .Z(n6609) );
  XOR U6227 ( .A(n6610), .B(n6611), .Z(n6607) );
  AND U6228 ( .A(n215), .B(n6612), .Z(n6611) );
  XOR U6229 ( .A(n6613), .B(n6614), .Z(n6605) );
  AND U6230 ( .A(n219), .B(n6612), .Z(n6614) );
  XNOR U6231 ( .A(n6613), .B(n6610), .Z(n6612) );
  XOR U6232 ( .A(n6615), .B(n6616), .Z(n6610) );
  AND U6233 ( .A(n222), .B(n6617), .Z(n6616) );
  XOR U6234 ( .A(p_input[275]), .B(n6615), .Z(n6617) );
  XOR U6235 ( .A(n6618), .B(n6619), .Z(n6615) );
  AND U6236 ( .A(n226), .B(n6620), .Z(n6619) );
  XOR U6237 ( .A(n6621), .B(n6622), .Z(n6613) );
  AND U6238 ( .A(n230), .B(n6620), .Z(n6622) );
  XNOR U6239 ( .A(n6621), .B(n6618), .Z(n6620) );
  XOR U6240 ( .A(n6623), .B(n6624), .Z(n6618) );
  AND U6241 ( .A(n233), .B(n6625), .Z(n6624) );
  XOR U6242 ( .A(p_input[291]), .B(n6623), .Z(n6625) );
  XOR U6243 ( .A(n6626), .B(n6627), .Z(n6623) );
  AND U6244 ( .A(n237), .B(n6628), .Z(n6627) );
  XOR U6245 ( .A(n6629), .B(n6630), .Z(n6621) );
  AND U6246 ( .A(n241), .B(n6628), .Z(n6630) );
  XNOR U6247 ( .A(n6629), .B(n6626), .Z(n6628) );
  XOR U6248 ( .A(n6631), .B(n6632), .Z(n6626) );
  AND U6249 ( .A(n244), .B(n6633), .Z(n6632) );
  XOR U6250 ( .A(p_input[307]), .B(n6631), .Z(n6633) );
  XOR U6251 ( .A(n6634), .B(n6635), .Z(n6631) );
  AND U6252 ( .A(n248), .B(n6636), .Z(n6635) );
  XOR U6253 ( .A(n6637), .B(n6638), .Z(n6629) );
  AND U6254 ( .A(n252), .B(n6636), .Z(n6638) );
  XNOR U6255 ( .A(n6637), .B(n6634), .Z(n6636) );
  XOR U6256 ( .A(n6639), .B(n6640), .Z(n6634) );
  AND U6257 ( .A(n255), .B(n6641), .Z(n6640) );
  XOR U6258 ( .A(p_input[323]), .B(n6639), .Z(n6641) );
  XOR U6259 ( .A(n6642), .B(n6643), .Z(n6639) );
  AND U6260 ( .A(n259), .B(n6644), .Z(n6643) );
  XOR U6261 ( .A(n6645), .B(n6646), .Z(n6637) );
  AND U6262 ( .A(n263), .B(n6644), .Z(n6646) );
  XNOR U6263 ( .A(n6645), .B(n6642), .Z(n6644) );
  XOR U6264 ( .A(n6647), .B(n6648), .Z(n6642) );
  AND U6265 ( .A(n266), .B(n6649), .Z(n6648) );
  XOR U6266 ( .A(p_input[339]), .B(n6647), .Z(n6649) );
  XOR U6267 ( .A(n6650), .B(n6651), .Z(n6647) );
  AND U6268 ( .A(n270), .B(n6652), .Z(n6651) );
  XOR U6269 ( .A(n6653), .B(n6654), .Z(n6645) );
  AND U6270 ( .A(n274), .B(n6652), .Z(n6654) );
  XNOR U6271 ( .A(n6653), .B(n6650), .Z(n6652) );
  XOR U6272 ( .A(n6655), .B(n6656), .Z(n6650) );
  AND U6273 ( .A(n277), .B(n6657), .Z(n6656) );
  XOR U6274 ( .A(p_input[355]), .B(n6655), .Z(n6657) );
  XOR U6275 ( .A(n6658), .B(n6659), .Z(n6655) );
  AND U6276 ( .A(n281), .B(n6660), .Z(n6659) );
  XOR U6277 ( .A(n6661), .B(n6662), .Z(n6653) );
  AND U6278 ( .A(n285), .B(n6660), .Z(n6662) );
  XNOR U6279 ( .A(n6661), .B(n6658), .Z(n6660) );
  XOR U6280 ( .A(n6663), .B(n6664), .Z(n6658) );
  AND U6281 ( .A(n288), .B(n6665), .Z(n6664) );
  XOR U6282 ( .A(p_input[371]), .B(n6663), .Z(n6665) );
  XOR U6283 ( .A(n6666), .B(n6667), .Z(n6663) );
  AND U6284 ( .A(n292), .B(n6668), .Z(n6667) );
  XOR U6285 ( .A(n6669), .B(n6670), .Z(n6661) );
  AND U6286 ( .A(n296), .B(n6668), .Z(n6670) );
  XNOR U6287 ( .A(n6669), .B(n6666), .Z(n6668) );
  XOR U6288 ( .A(n6671), .B(n6672), .Z(n6666) );
  AND U6289 ( .A(n299), .B(n6673), .Z(n6672) );
  XOR U6290 ( .A(p_input[387]), .B(n6671), .Z(n6673) );
  XOR U6291 ( .A(n6674), .B(n6675), .Z(n6671) );
  AND U6292 ( .A(n303), .B(n6676), .Z(n6675) );
  XOR U6293 ( .A(n6677), .B(n6678), .Z(n6669) );
  AND U6294 ( .A(n307), .B(n6676), .Z(n6678) );
  XNOR U6295 ( .A(n6677), .B(n6674), .Z(n6676) );
  XOR U6296 ( .A(n6679), .B(n6680), .Z(n6674) );
  AND U6297 ( .A(n310), .B(n6681), .Z(n6680) );
  XOR U6298 ( .A(p_input[403]), .B(n6679), .Z(n6681) );
  XOR U6299 ( .A(n6682), .B(n6683), .Z(n6679) );
  AND U6300 ( .A(n314), .B(n6684), .Z(n6683) );
  XOR U6301 ( .A(n6685), .B(n6686), .Z(n6677) );
  AND U6302 ( .A(n318), .B(n6684), .Z(n6686) );
  XNOR U6303 ( .A(n6685), .B(n6682), .Z(n6684) );
  XOR U6304 ( .A(n6687), .B(n6688), .Z(n6682) );
  AND U6305 ( .A(n321), .B(n6689), .Z(n6688) );
  XOR U6306 ( .A(p_input[419]), .B(n6687), .Z(n6689) );
  XOR U6307 ( .A(n6690), .B(n6691), .Z(n6687) );
  AND U6308 ( .A(n325), .B(n6692), .Z(n6691) );
  XOR U6309 ( .A(n6693), .B(n6694), .Z(n6685) );
  AND U6310 ( .A(n329), .B(n6692), .Z(n6694) );
  XNOR U6311 ( .A(n6693), .B(n6690), .Z(n6692) );
  XOR U6312 ( .A(n6695), .B(n6696), .Z(n6690) );
  AND U6313 ( .A(n332), .B(n6697), .Z(n6696) );
  XOR U6314 ( .A(p_input[435]), .B(n6695), .Z(n6697) );
  XOR U6315 ( .A(n6698), .B(n6699), .Z(n6695) );
  AND U6316 ( .A(n336), .B(n6700), .Z(n6699) );
  XOR U6317 ( .A(n6701), .B(n6702), .Z(n6693) );
  AND U6318 ( .A(n340), .B(n6700), .Z(n6702) );
  XNOR U6319 ( .A(n6701), .B(n6698), .Z(n6700) );
  XOR U6320 ( .A(n6703), .B(n6704), .Z(n6698) );
  AND U6321 ( .A(n343), .B(n6705), .Z(n6704) );
  XOR U6322 ( .A(p_input[451]), .B(n6703), .Z(n6705) );
  XOR U6323 ( .A(n6706), .B(n6707), .Z(n6703) );
  AND U6324 ( .A(n347), .B(n6708), .Z(n6707) );
  XOR U6325 ( .A(n6709), .B(n6710), .Z(n6701) );
  AND U6326 ( .A(n351), .B(n6708), .Z(n6710) );
  XNOR U6327 ( .A(n6709), .B(n6706), .Z(n6708) );
  XOR U6328 ( .A(n6711), .B(n6712), .Z(n6706) );
  AND U6329 ( .A(n354), .B(n6713), .Z(n6712) );
  XOR U6330 ( .A(p_input[467]), .B(n6711), .Z(n6713) );
  XOR U6331 ( .A(n6714), .B(n6715), .Z(n6711) );
  AND U6332 ( .A(n358), .B(n6716), .Z(n6715) );
  XOR U6333 ( .A(n6717), .B(n6718), .Z(n6709) );
  AND U6334 ( .A(n362), .B(n6716), .Z(n6718) );
  XNOR U6335 ( .A(n6717), .B(n6714), .Z(n6716) );
  XOR U6336 ( .A(n6719), .B(n6720), .Z(n6714) );
  AND U6337 ( .A(n365), .B(n6721), .Z(n6720) );
  XOR U6338 ( .A(p_input[483]), .B(n6719), .Z(n6721) );
  XOR U6339 ( .A(n6722), .B(n6723), .Z(n6719) );
  AND U6340 ( .A(n369), .B(n6724), .Z(n6723) );
  XOR U6341 ( .A(n6725), .B(n6726), .Z(n6717) );
  AND U6342 ( .A(n373), .B(n6724), .Z(n6726) );
  XNOR U6343 ( .A(n6725), .B(n6722), .Z(n6724) );
  XOR U6344 ( .A(n6727), .B(n6728), .Z(n6722) );
  AND U6345 ( .A(n376), .B(n6729), .Z(n6728) );
  XOR U6346 ( .A(p_input[499]), .B(n6727), .Z(n6729) );
  XOR U6347 ( .A(n6730), .B(n6731), .Z(n6727) );
  AND U6348 ( .A(n380), .B(n6732), .Z(n6731) );
  XOR U6349 ( .A(n6733), .B(n6734), .Z(n6725) );
  AND U6350 ( .A(n384), .B(n6732), .Z(n6734) );
  XNOR U6351 ( .A(n6733), .B(n6730), .Z(n6732) );
  XOR U6352 ( .A(n6735), .B(n6736), .Z(n6730) );
  AND U6353 ( .A(n387), .B(n6737), .Z(n6736) );
  XOR U6354 ( .A(p_input[515]), .B(n6735), .Z(n6737) );
  XOR U6355 ( .A(n6738), .B(n6739), .Z(n6735) );
  AND U6356 ( .A(n391), .B(n6740), .Z(n6739) );
  XOR U6357 ( .A(n6741), .B(n6742), .Z(n6733) );
  AND U6358 ( .A(n395), .B(n6740), .Z(n6742) );
  XNOR U6359 ( .A(n6741), .B(n6738), .Z(n6740) );
  XOR U6360 ( .A(n6743), .B(n6744), .Z(n6738) );
  AND U6361 ( .A(n398), .B(n6745), .Z(n6744) );
  XOR U6362 ( .A(p_input[531]), .B(n6743), .Z(n6745) );
  XOR U6363 ( .A(n6746), .B(n6747), .Z(n6743) );
  AND U6364 ( .A(n402), .B(n6748), .Z(n6747) );
  XOR U6365 ( .A(n6749), .B(n6750), .Z(n6741) );
  AND U6366 ( .A(n406), .B(n6748), .Z(n6750) );
  XNOR U6367 ( .A(n6749), .B(n6746), .Z(n6748) );
  XOR U6368 ( .A(n6751), .B(n6752), .Z(n6746) );
  AND U6369 ( .A(n409), .B(n6753), .Z(n6752) );
  XOR U6370 ( .A(p_input[547]), .B(n6751), .Z(n6753) );
  XOR U6371 ( .A(n6754), .B(n6755), .Z(n6751) );
  AND U6372 ( .A(n413), .B(n6756), .Z(n6755) );
  XOR U6373 ( .A(n6757), .B(n6758), .Z(n6749) );
  AND U6374 ( .A(n417), .B(n6756), .Z(n6758) );
  XNOR U6375 ( .A(n6757), .B(n6754), .Z(n6756) );
  XOR U6376 ( .A(n6759), .B(n6760), .Z(n6754) );
  AND U6377 ( .A(n420), .B(n6761), .Z(n6760) );
  XOR U6378 ( .A(p_input[563]), .B(n6759), .Z(n6761) );
  XOR U6379 ( .A(n6762), .B(n6763), .Z(n6759) );
  AND U6380 ( .A(n424), .B(n6764), .Z(n6763) );
  XOR U6381 ( .A(n6765), .B(n6766), .Z(n6757) );
  AND U6382 ( .A(n428), .B(n6764), .Z(n6766) );
  XNOR U6383 ( .A(n6765), .B(n6762), .Z(n6764) );
  XOR U6384 ( .A(n6767), .B(n6768), .Z(n6762) );
  AND U6385 ( .A(n431), .B(n6769), .Z(n6768) );
  XOR U6386 ( .A(p_input[579]), .B(n6767), .Z(n6769) );
  XOR U6387 ( .A(n6770), .B(n6771), .Z(n6767) );
  AND U6388 ( .A(n435), .B(n6772), .Z(n6771) );
  XOR U6389 ( .A(n6773), .B(n6774), .Z(n6765) );
  AND U6390 ( .A(n439), .B(n6772), .Z(n6774) );
  XNOR U6391 ( .A(n6773), .B(n6770), .Z(n6772) );
  XOR U6392 ( .A(n6775), .B(n6776), .Z(n6770) );
  AND U6393 ( .A(n442), .B(n6777), .Z(n6776) );
  XOR U6394 ( .A(p_input[595]), .B(n6775), .Z(n6777) );
  XOR U6395 ( .A(n6778), .B(n6779), .Z(n6775) );
  AND U6396 ( .A(n446), .B(n6780), .Z(n6779) );
  XOR U6397 ( .A(n6781), .B(n6782), .Z(n6773) );
  AND U6398 ( .A(n450), .B(n6780), .Z(n6782) );
  XNOR U6399 ( .A(n6781), .B(n6778), .Z(n6780) );
  XOR U6400 ( .A(n6783), .B(n6784), .Z(n6778) );
  AND U6401 ( .A(n453), .B(n6785), .Z(n6784) );
  XOR U6402 ( .A(p_input[611]), .B(n6783), .Z(n6785) );
  XOR U6403 ( .A(n6786), .B(n6787), .Z(n6783) );
  AND U6404 ( .A(n457), .B(n6788), .Z(n6787) );
  XOR U6405 ( .A(n6789), .B(n6790), .Z(n6781) );
  AND U6406 ( .A(n461), .B(n6788), .Z(n6790) );
  XNOR U6407 ( .A(n6789), .B(n6786), .Z(n6788) );
  XOR U6408 ( .A(n6791), .B(n6792), .Z(n6786) );
  AND U6409 ( .A(n464), .B(n6793), .Z(n6792) );
  XOR U6410 ( .A(p_input[627]), .B(n6791), .Z(n6793) );
  XOR U6411 ( .A(n6794), .B(n6795), .Z(n6791) );
  AND U6412 ( .A(n468), .B(n6796), .Z(n6795) );
  XOR U6413 ( .A(n6797), .B(n6798), .Z(n6789) );
  AND U6414 ( .A(n472), .B(n6796), .Z(n6798) );
  XNOR U6415 ( .A(n6797), .B(n6794), .Z(n6796) );
  XOR U6416 ( .A(n6799), .B(n6800), .Z(n6794) );
  AND U6417 ( .A(n475), .B(n6801), .Z(n6800) );
  XOR U6418 ( .A(p_input[643]), .B(n6799), .Z(n6801) );
  XOR U6419 ( .A(n6802), .B(n6803), .Z(n6799) );
  AND U6420 ( .A(n479), .B(n6804), .Z(n6803) );
  XOR U6421 ( .A(n6805), .B(n6806), .Z(n6797) );
  AND U6422 ( .A(n483), .B(n6804), .Z(n6806) );
  XNOR U6423 ( .A(n6805), .B(n6802), .Z(n6804) );
  XOR U6424 ( .A(n6807), .B(n6808), .Z(n6802) );
  AND U6425 ( .A(n486), .B(n6809), .Z(n6808) );
  XOR U6426 ( .A(p_input[659]), .B(n6807), .Z(n6809) );
  XOR U6427 ( .A(n6810), .B(n6811), .Z(n6807) );
  AND U6428 ( .A(n490), .B(n6812), .Z(n6811) );
  XOR U6429 ( .A(n6813), .B(n6814), .Z(n6805) );
  AND U6430 ( .A(n494), .B(n6812), .Z(n6814) );
  XNOR U6431 ( .A(n6813), .B(n6810), .Z(n6812) );
  XOR U6432 ( .A(n6815), .B(n6816), .Z(n6810) );
  AND U6433 ( .A(n497), .B(n6817), .Z(n6816) );
  XOR U6434 ( .A(p_input[675]), .B(n6815), .Z(n6817) );
  XOR U6435 ( .A(n6818), .B(n6819), .Z(n6815) );
  AND U6436 ( .A(n501), .B(n6820), .Z(n6819) );
  XOR U6437 ( .A(n6821), .B(n6822), .Z(n6813) );
  AND U6438 ( .A(n505), .B(n6820), .Z(n6822) );
  XNOR U6439 ( .A(n6821), .B(n6818), .Z(n6820) );
  XOR U6440 ( .A(n6823), .B(n6824), .Z(n6818) );
  AND U6441 ( .A(n508), .B(n6825), .Z(n6824) );
  XOR U6442 ( .A(p_input[691]), .B(n6823), .Z(n6825) );
  XOR U6443 ( .A(n6826), .B(n6827), .Z(n6823) );
  AND U6444 ( .A(n512), .B(n6828), .Z(n6827) );
  XOR U6445 ( .A(n6829), .B(n6830), .Z(n6821) );
  AND U6446 ( .A(n516), .B(n6828), .Z(n6830) );
  XNOR U6447 ( .A(n6829), .B(n6826), .Z(n6828) );
  XOR U6448 ( .A(n6831), .B(n6832), .Z(n6826) );
  AND U6449 ( .A(n519), .B(n6833), .Z(n6832) );
  XOR U6450 ( .A(p_input[707]), .B(n6831), .Z(n6833) );
  XOR U6451 ( .A(n6834), .B(n6835), .Z(n6831) );
  AND U6452 ( .A(n523), .B(n6836), .Z(n6835) );
  XOR U6453 ( .A(n6837), .B(n6838), .Z(n6829) );
  AND U6454 ( .A(n527), .B(n6836), .Z(n6838) );
  XNOR U6455 ( .A(n6837), .B(n6834), .Z(n6836) );
  XOR U6456 ( .A(n6839), .B(n6840), .Z(n6834) );
  AND U6457 ( .A(n530), .B(n6841), .Z(n6840) );
  XOR U6458 ( .A(p_input[723]), .B(n6839), .Z(n6841) );
  XOR U6459 ( .A(n6842), .B(n6843), .Z(n6839) );
  AND U6460 ( .A(n534), .B(n6844), .Z(n6843) );
  XOR U6461 ( .A(n6845), .B(n6846), .Z(n6837) );
  AND U6462 ( .A(n538), .B(n6844), .Z(n6846) );
  XNOR U6463 ( .A(n6845), .B(n6842), .Z(n6844) );
  XOR U6464 ( .A(n6847), .B(n6848), .Z(n6842) );
  AND U6465 ( .A(n541), .B(n6849), .Z(n6848) );
  XOR U6466 ( .A(p_input[739]), .B(n6847), .Z(n6849) );
  XOR U6467 ( .A(n6850), .B(n6851), .Z(n6847) );
  AND U6468 ( .A(n545), .B(n6852), .Z(n6851) );
  XOR U6469 ( .A(n6853), .B(n6854), .Z(n6845) );
  AND U6470 ( .A(n549), .B(n6852), .Z(n6854) );
  XNOR U6471 ( .A(n6853), .B(n6850), .Z(n6852) );
  XOR U6472 ( .A(n6855), .B(n6856), .Z(n6850) );
  AND U6473 ( .A(n552), .B(n6857), .Z(n6856) );
  XOR U6474 ( .A(p_input[755]), .B(n6855), .Z(n6857) );
  XOR U6475 ( .A(n6858), .B(n6859), .Z(n6855) );
  AND U6476 ( .A(n556), .B(n6860), .Z(n6859) );
  XOR U6477 ( .A(n6861), .B(n6862), .Z(n6853) );
  AND U6478 ( .A(n560), .B(n6860), .Z(n6862) );
  XNOR U6479 ( .A(n6861), .B(n6858), .Z(n6860) );
  XOR U6480 ( .A(n6863), .B(n6864), .Z(n6858) );
  AND U6481 ( .A(n563), .B(n6865), .Z(n6864) );
  XOR U6482 ( .A(p_input[771]), .B(n6863), .Z(n6865) );
  XOR U6483 ( .A(n6866), .B(n6867), .Z(n6863) );
  AND U6484 ( .A(n567), .B(n6868), .Z(n6867) );
  XOR U6485 ( .A(n6869), .B(n6870), .Z(n6861) );
  AND U6486 ( .A(n571), .B(n6868), .Z(n6870) );
  XNOR U6487 ( .A(n6869), .B(n6866), .Z(n6868) );
  XOR U6488 ( .A(n6871), .B(n6872), .Z(n6866) );
  AND U6489 ( .A(n574), .B(n6873), .Z(n6872) );
  XOR U6490 ( .A(p_input[787]), .B(n6871), .Z(n6873) );
  XOR U6491 ( .A(n6874), .B(n6875), .Z(n6871) );
  AND U6492 ( .A(n578), .B(n6876), .Z(n6875) );
  XOR U6493 ( .A(n6877), .B(n6878), .Z(n6869) );
  AND U6494 ( .A(n582), .B(n6876), .Z(n6878) );
  XNOR U6495 ( .A(n6877), .B(n6874), .Z(n6876) );
  XOR U6496 ( .A(n6879), .B(n6880), .Z(n6874) );
  AND U6497 ( .A(n585), .B(n6881), .Z(n6880) );
  XOR U6498 ( .A(p_input[803]), .B(n6879), .Z(n6881) );
  XOR U6499 ( .A(n6882), .B(n6883), .Z(n6879) );
  AND U6500 ( .A(n589), .B(n6884), .Z(n6883) );
  XOR U6501 ( .A(n6885), .B(n6886), .Z(n6877) );
  AND U6502 ( .A(n593), .B(n6884), .Z(n6886) );
  XNOR U6503 ( .A(n6885), .B(n6882), .Z(n6884) );
  XOR U6504 ( .A(n6887), .B(n6888), .Z(n6882) );
  AND U6505 ( .A(n596), .B(n6889), .Z(n6888) );
  XOR U6506 ( .A(p_input[819]), .B(n6887), .Z(n6889) );
  XOR U6507 ( .A(n6890), .B(n6891), .Z(n6887) );
  AND U6508 ( .A(n600), .B(n6892), .Z(n6891) );
  XOR U6509 ( .A(n6893), .B(n6894), .Z(n6885) );
  AND U6510 ( .A(n604), .B(n6892), .Z(n6894) );
  XNOR U6511 ( .A(n6893), .B(n6890), .Z(n6892) );
  XOR U6512 ( .A(n6895), .B(n6896), .Z(n6890) );
  AND U6513 ( .A(n607), .B(n6897), .Z(n6896) );
  XOR U6514 ( .A(p_input[835]), .B(n6895), .Z(n6897) );
  XOR U6515 ( .A(n6898), .B(n6899), .Z(n6895) );
  AND U6516 ( .A(n611), .B(n6900), .Z(n6899) );
  XOR U6517 ( .A(n6901), .B(n6902), .Z(n6893) );
  AND U6518 ( .A(n615), .B(n6900), .Z(n6902) );
  XNOR U6519 ( .A(n6901), .B(n6898), .Z(n6900) );
  XOR U6520 ( .A(n6903), .B(n6904), .Z(n6898) );
  AND U6521 ( .A(n618), .B(n6905), .Z(n6904) );
  XOR U6522 ( .A(p_input[851]), .B(n6903), .Z(n6905) );
  XOR U6523 ( .A(n6906), .B(n6907), .Z(n6903) );
  AND U6524 ( .A(n622), .B(n6908), .Z(n6907) );
  XOR U6525 ( .A(n6909), .B(n6910), .Z(n6901) );
  AND U6526 ( .A(n626), .B(n6908), .Z(n6910) );
  XNOR U6527 ( .A(n6909), .B(n6906), .Z(n6908) );
  XOR U6528 ( .A(n6911), .B(n6912), .Z(n6906) );
  AND U6529 ( .A(n629), .B(n6913), .Z(n6912) );
  XOR U6530 ( .A(p_input[867]), .B(n6911), .Z(n6913) );
  XOR U6531 ( .A(n6914), .B(n6915), .Z(n6911) );
  AND U6532 ( .A(n633), .B(n6916), .Z(n6915) );
  XOR U6533 ( .A(n6917), .B(n6918), .Z(n6909) );
  AND U6534 ( .A(n637), .B(n6916), .Z(n6918) );
  XNOR U6535 ( .A(n6917), .B(n6914), .Z(n6916) );
  XOR U6536 ( .A(n6919), .B(n6920), .Z(n6914) );
  AND U6537 ( .A(n640), .B(n6921), .Z(n6920) );
  XOR U6538 ( .A(p_input[883]), .B(n6919), .Z(n6921) );
  XOR U6539 ( .A(n6922), .B(n6923), .Z(n6919) );
  AND U6540 ( .A(n644), .B(n6924), .Z(n6923) );
  XOR U6541 ( .A(n6925), .B(n6926), .Z(n6917) );
  AND U6542 ( .A(n648), .B(n6924), .Z(n6926) );
  XNOR U6543 ( .A(n6925), .B(n6922), .Z(n6924) );
  XOR U6544 ( .A(n6927), .B(n6928), .Z(n6922) );
  AND U6545 ( .A(n651), .B(n6929), .Z(n6928) );
  XOR U6546 ( .A(p_input[899]), .B(n6927), .Z(n6929) );
  XOR U6547 ( .A(n6930), .B(n6931), .Z(n6927) );
  AND U6548 ( .A(n655), .B(n6932), .Z(n6931) );
  XOR U6549 ( .A(n6933), .B(n6934), .Z(n6925) );
  AND U6550 ( .A(n659), .B(n6932), .Z(n6934) );
  XNOR U6551 ( .A(n6933), .B(n6930), .Z(n6932) );
  XOR U6552 ( .A(n6935), .B(n6936), .Z(n6930) );
  AND U6553 ( .A(n662), .B(n6937), .Z(n6936) );
  XOR U6554 ( .A(p_input[915]), .B(n6935), .Z(n6937) );
  XOR U6555 ( .A(n6938), .B(n6939), .Z(n6935) );
  AND U6556 ( .A(n666), .B(n6940), .Z(n6939) );
  XOR U6557 ( .A(n6941), .B(n6942), .Z(n6933) );
  AND U6558 ( .A(n670), .B(n6940), .Z(n6942) );
  XNOR U6559 ( .A(n6941), .B(n6938), .Z(n6940) );
  XOR U6560 ( .A(n6943), .B(n6944), .Z(n6938) );
  AND U6561 ( .A(n673), .B(n6945), .Z(n6944) );
  XOR U6562 ( .A(p_input[931]), .B(n6943), .Z(n6945) );
  XOR U6563 ( .A(n6946), .B(n6947), .Z(n6943) );
  AND U6564 ( .A(n677), .B(n6948), .Z(n6947) );
  XOR U6565 ( .A(n6949), .B(n6950), .Z(n6941) );
  AND U6566 ( .A(n681), .B(n6948), .Z(n6950) );
  XNOR U6567 ( .A(n6949), .B(n6946), .Z(n6948) );
  XOR U6568 ( .A(n6951), .B(n6952), .Z(n6946) );
  AND U6569 ( .A(n684), .B(n6953), .Z(n6952) );
  XOR U6570 ( .A(p_input[947]), .B(n6951), .Z(n6953) );
  XOR U6571 ( .A(n6954), .B(n6955), .Z(n6951) );
  AND U6572 ( .A(n688), .B(n6956), .Z(n6955) );
  XOR U6573 ( .A(n6957), .B(n6958), .Z(n6949) );
  AND U6574 ( .A(n692), .B(n6956), .Z(n6958) );
  XNOR U6575 ( .A(n6957), .B(n6954), .Z(n6956) );
  XOR U6576 ( .A(n6959), .B(n6960), .Z(n6954) );
  AND U6577 ( .A(n695), .B(n6961), .Z(n6960) );
  XOR U6578 ( .A(p_input[963]), .B(n6959), .Z(n6961) );
  XOR U6579 ( .A(n6962), .B(n6963), .Z(n6959) );
  AND U6580 ( .A(n699), .B(n6964), .Z(n6963) );
  XOR U6581 ( .A(n6965), .B(n6966), .Z(n6957) );
  AND U6582 ( .A(n703), .B(n6964), .Z(n6966) );
  XNOR U6583 ( .A(n6965), .B(n6962), .Z(n6964) );
  XOR U6584 ( .A(n6967), .B(n6968), .Z(n6962) );
  AND U6585 ( .A(n706), .B(n6969), .Z(n6968) );
  XOR U6586 ( .A(p_input[979]), .B(n6967), .Z(n6969) );
  XOR U6587 ( .A(n6970), .B(n6971), .Z(n6967) );
  AND U6588 ( .A(n710), .B(n6972), .Z(n6971) );
  XOR U6589 ( .A(n6973), .B(n6974), .Z(n6965) );
  AND U6590 ( .A(n714), .B(n6972), .Z(n6974) );
  XNOR U6591 ( .A(n6973), .B(n6970), .Z(n6972) );
  XOR U6592 ( .A(n6975), .B(n6976), .Z(n6970) );
  AND U6593 ( .A(n717), .B(n6977), .Z(n6976) );
  XOR U6594 ( .A(p_input[995]), .B(n6975), .Z(n6977) );
  XOR U6595 ( .A(n6978), .B(n6979), .Z(n6975) );
  AND U6596 ( .A(n721), .B(n6980), .Z(n6979) );
  XOR U6597 ( .A(n6981), .B(n6982), .Z(n6973) );
  AND U6598 ( .A(n725), .B(n6980), .Z(n6982) );
  XNOR U6599 ( .A(n6981), .B(n6978), .Z(n6980) );
  XOR U6600 ( .A(n6983), .B(n6984), .Z(n6978) );
  AND U6601 ( .A(n728), .B(n6985), .Z(n6984) );
  XOR U6602 ( .A(p_input[1011]), .B(n6983), .Z(n6985) );
  XOR U6603 ( .A(n6986), .B(n6987), .Z(n6983) );
  AND U6604 ( .A(n732), .B(n6988), .Z(n6987) );
  XOR U6605 ( .A(n6989), .B(n6990), .Z(n6981) );
  AND U6606 ( .A(n736), .B(n6988), .Z(n6990) );
  XNOR U6607 ( .A(n6989), .B(n6986), .Z(n6988) );
  XOR U6608 ( .A(n6991), .B(n6992), .Z(n6986) );
  AND U6609 ( .A(n739), .B(n6993), .Z(n6992) );
  XOR U6610 ( .A(p_input[1027]), .B(n6991), .Z(n6993) );
  XOR U6611 ( .A(n6994), .B(n6995), .Z(n6991) );
  AND U6612 ( .A(n743), .B(n6996), .Z(n6995) );
  XOR U6613 ( .A(n6997), .B(n6998), .Z(n6989) );
  AND U6614 ( .A(n747), .B(n6996), .Z(n6998) );
  XNOR U6615 ( .A(n6997), .B(n6994), .Z(n6996) );
  XOR U6616 ( .A(n6999), .B(n7000), .Z(n6994) );
  AND U6617 ( .A(n750), .B(n7001), .Z(n7000) );
  XOR U6618 ( .A(p_input[1043]), .B(n6999), .Z(n7001) );
  XOR U6619 ( .A(n7002), .B(n7003), .Z(n6999) );
  AND U6620 ( .A(n754), .B(n7004), .Z(n7003) );
  XOR U6621 ( .A(n7005), .B(n7006), .Z(n6997) );
  AND U6622 ( .A(n758), .B(n7004), .Z(n7006) );
  XNOR U6623 ( .A(n7005), .B(n7002), .Z(n7004) );
  XOR U6624 ( .A(n7007), .B(n7008), .Z(n7002) );
  AND U6625 ( .A(n761), .B(n7009), .Z(n7008) );
  XOR U6626 ( .A(p_input[1059]), .B(n7007), .Z(n7009) );
  XOR U6627 ( .A(n7010), .B(n7011), .Z(n7007) );
  AND U6628 ( .A(n765), .B(n7012), .Z(n7011) );
  XOR U6629 ( .A(n7013), .B(n7014), .Z(n7005) );
  AND U6630 ( .A(n769), .B(n7012), .Z(n7014) );
  XNOR U6631 ( .A(n7013), .B(n7010), .Z(n7012) );
  XOR U6632 ( .A(n7015), .B(n7016), .Z(n7010) );
  AND U6633 ( .A(n772), .B(n7017), .Z(n7016) );
  XOR U6634 ( .A(p_input[1075]), .B(n7015), .Z(n7017) );
  XOR U6635 ( .A(n7018), .B(n7019), .Z(n7015) );
  AND U6636 ( .A(n776), .B(n7020), .Z(n7019) );
  XOR U6637 ( .A(n7021), .B(n7022), .Z(n7013) );
  AND U6638 ( .A(n780), .B(n7020), .Z(n7022) );
  XNOR U6639 ( .A(n7021), .B(n7018), .Z(n7020) );
  XOR U6640 ( .A(n7023), .B(n7024), .Z(n7018) );
  AND U6641 ( .A(n783), .B(n7025), .Z(n7024) );
  XOR U6642 ( .A(p_input[1091]), .B(n7023), .Z(n7025) );
  XOR U6643 ( .A(n7026), .B(n7027), .Z(n7023) );
  AND U6644 ( .A(n787), .B(n7028), .Z(n7027) );
  XOR U6645 ( .A(n7029), .B(n7030), .Z(n7021) );
  AND U6646 ( .A(n791), .B(n7028), .Z(n7030) );
  XNOR U6647 ( .A(n7029), .B(n7026), .Z(n7028) );
  XOR U6648 ( .A(n7031), .B(n7032), .Z(n7026) );
  AND U6649 ( .A(n794), .B(n7033), .Z(n7032) );
  XOR U6650 ( .A(p_input[1107]), .B(n7031), .Z(n7033) );
  XOR U6651 ( .A(n7034), .B(n7035), .Z(n7031) );
  AND U6652 ( .A(n798), .B(n7036), .Z(n7035) );
  XOR U6653 ( .A(n7037), .B(n7038), .Z(n7029) );
  AND U6654 ( .A(n802), .B(n7036), .Z(n7038) );
  XNOR U6655 ( .A(n7037), .B(n7034), .Z(n7036) );
  XOR U6656 ( .A(n7039), .B(n7040), .Z(n7034) );
  AND U6657 ( .A(n805), .B(n7041), .Z(n7040) );
  XOR U6658 ( .A(p_input[1123]), .B(n7039), .Z(n7041) );
  XOR U6659 ( .A(n7042), .B(n7043), .Z(n7039) );
  AND U6660 ( .A(n809), .B(n7044), .Z(n7043) );
  XOR U6661 ( .A(n7045), .B(n7046), .Z(n7037) );
  AND U6662 ( .A(n813), .B(n7044), .Z(n7046) );
  XNOR U6663 ( .A(n7045), .B(n7042), .Z(n7044) );
  XOR U6664 ( .A(n7047), .B(n7048), .Z(n7042) );
  AND U6665 ( .A(n816), .B(n7049), .Z(n7048) );
  XOR U6666 ( .A(p_input[1139]), .B(n7047), .Z(n7049) );
  XOR U6667 ( .A(n7050), .B(n7051), .Z(n7047) );
  AND U6668 ( .A(n820), .B(n7052), .Z(n7051) );
  XOR U6669 ( .A(n7053), .B(n7054), .Z(n7045) );
  AND U6670 ( .A(n824), .B(n7052), .Z(n7054) );
  XNOR U6671 ( .A(n7053), .B(n7050), .Z(n7052) );
  XOR U6672 ( .A(n7055), .B(n7056), .Z(n7050) );
  AND U6673 ( .A(n827), .B(n7057), .Z(n7056) );
  XOR U6674 ( .A(p_input[1155]), .B(n7055), .Z(n7057) );
  XOR U6675 ( .A(n7058), .B(n7059), .Z(n7055) );
  AND U6676 ( .A(n831), .B(n7060), .Z(n7059) );
  XOR U6677 ( .A(n7061), .B(n7062), .Z(n7053) );
  AND U6678 ( .A(n835), .B(n7060), .Z(n7062) );
  XNOR U6679 ( .A(n7061), .B(n7058), .Z(n7060) );
  XOR U6680 ( .A(n7063), .B(n7064), .Z(n7058) );
  AND U6681 ( .A(n838), .B(n7065), .Z(n7064) );
  XOR U6682 ( .A(p_input[1171]), .B(n7063), .Z(n7065) );
  XOR U6683 ( .A(n7066), .B(n7067), .Z(n7063) );
  AND U6684 ( .A(n842), .B(n7068), .Z(n7067) );
  XOR U6685 ( .A(n7069), .B(n7070), .Z(n7061) );
  AND U6686 ( .A(n846), .B(n7068), .Z(n7070) );
  XNOR U6687 ( .A(n7069), .B(n7066), .Z(n7068) );
  XOR U6688 ( .A(n7071), .B(n7072), .Z(n7066) );
  AND U6689 ( .A(n849), .B(n7073), .Z(n7072) );
  XOR U6690 ( .A(p_input[1187]), .B(n7071), .Z(n7073) );
  XOR U6691 ( .A(n7074), .B(n7075), .Z(n7071) );
  AND U6692 ( .A(n853), .B(n7076), .Z(n7075) );
  XOR U6693 ( .A(n7077), .B(n7078), .Z(n7069) );
  AND U6694 ( .A(n857), .B(n7076), .Z(n7078) );
  XNOR U6695 ( .A(n7077), .B(n7074), .Z(n7076) );
  XOR U6696 ( .A(n7079), .B(n7080), .Z(n7074) );
  AND U6697 ( .A(n860), .B(n7081), .Z(n7080) );
  XOR U6698 ( .A(p_input[1203]), .B(n7079), .Z(n7081) );
  XOR U6699 ( .A(n7082), .B(n7083), .Z(n7079) );
  AND U6700 ( .A(n864), .B(n7084), .Z(n7083) );
  XOR U6701 ( .A(n7085), .B(n7086), .Z(n7077) );
  AND U6702 ( .A(n868), .B(n7084), .Z(n7086) );
  XNOR U6703 ( .A(n7085), .B(n7082), .Z(n7084) );
  XOR U6704 ( .A(n7087), .B(n7088), .Z(n7082) );
  AND U6705 ( .A(n871), .B(n7089), .Z(n7088) );
  XOR U6706 ( .A(p_input[1219]), .B(n7087), .Z(n7089) );
  XOR U6707 ( .A(n7090), .B(n7091), .Z(n7087) );
  AND U6708 ( .A(n875), .B(n7092), .Z(n7091) );
  XOR U6709 ( .A(n7093), .B(n7094), .Z(n7085) );
  AND U6710 ( .A(n879), .B(n7092), .Z(n7094) );
  XNOR U6711 ( .A(n7093), .B(n7090), .Z(n7092) );
  XOR U6712 ( .A(n7095), .B(n7096), .Z(n7090) );
  AND U6713 ( .A(n882), .B(n7097), .Z(n7096) );
  XOR U6714 ( .A(p_input[1235]), .B(n7095), .Z(n7097) );
  XOR U6715 ( .A(n7098), .B(n7099), .Z(n7095) );
  AND U6716 ( .A(n886), .B(n7100), .Z(n7099) );
  XOR U6717 ( .A(n7101), .B(n7102), .Z(n7093) );
  AND U6718 ( .A(n890), .B(n7100), .Z(n7102) );
  XNOR U6719 ( .A(n7101), .B(n7098), .Z(n7100) );
  XOR U6720 ( .A(n7103), .B(n7104), .Z(n7098) );
  AND U6721 ( .A(n893), .B(n7105), .Z(n7104) );
  XOR U6722 ( .A(p_input[1251]), .B(n7103), .Z(n7105) );
  XOR U6723 ( .A(n7106), .B(n7107), .Z(n7103) );
  AND U6724 ( .A(n897), .B(n7108), .Z(n7107) );
  XOR U6725 ( .A(n7109), .B(n7110), .Z(n7101) );
  AND U6726 ( .A(n901), .B(n7108), .Z(n7110) );
  XNOR U6727 ( .A(n7109), .B(n7106), .Z(n7108) );
  XOR U6728 ( .A(n7111), .B(n7112), .Z(n7106) );
  AND U6729 ( .A(n904), .B(n7113), .Z(n7112) );
  XOR U6730 ( .A(p_input[1267]), .B(n7111), .Z(n7113) );
  XOR U6731 ( .A(n7114), .B(n7115), .Z(n7111) );
  AND U6732 ( .A(n908), .B(n7116), .Z(n7115) );
  XOR U6733 ( .A(n7117), .B(n7118), .Z(n7109) );
  AND U6734 ( .A(n912), .B(n7116), .Z(n7118) );
  XNOR U6735 ( .A(n7117), .B(n7114), .Z(n7116) );
  XOR U6736 ( .A(n7119), .B(n7120), .Z(n7114) );
  AND U6737 ( .A(n915), .B(n7121), .Z(n7120) );
  XOR U6738 ( .A(p_input[1283]), .B(n7119), .Z(n7121) );
  XOR U6739 ( .A(n7122), .B(n7123), .Z(n7119) );
  AND U6740 ( .A(n919), .B(n7124), .Z(n7123) );
  XOR U6741 ( .A(n7125), .B(n7126), .Z(n7117) );
  AND U6742 ( .A(n923), .B(n7124), .Z(n7126) );
  XNOR U6743 ( .A(n7125), .B(n7122), .Z(n7124) );
  XOR U6744 ( .A(n7127), .B(n7128), .Z(n7122) );
  AND U6745 ( .A(n926), .B(n7129), .Z(n7128) );
  XOR U6746 ( .A(p_input[1299]), .B(n7127), .Z(n7129) );
  XOR U6747 ( .A(n7130), .B(n7131), .Z(n7127) );
  AND U6748 ( .A(n930), .B(n7132), .Z(n7131) );
  XOR U6749 ( .A(n7133), .B(n7134), .Z(n7125) );
  AND U6750 ( .A(n934), .B(n7132), .Z(n7134) );
  XNOR U6751 ( .A(n7133), .B(n7130), .Z(n7132) );
  XOR U6752 ( .A(n7135), .B(n7136), .Z(n7130) );
  AND U6753 ( .A(n937), .B(n7137), .Z(n7136) );
  XOR U6754 ( .A(p_input[1315]), .B(n7135), .Z(n7137) );
  XOR U6755 ( .A(n7138), .B(n7139), .Z(n7135) );
  AND U6756 ( .A(n941), .B(n7140), .Z(n7139) );
  XOR U6757 ( .A(n7141), .B(n7142), .Z(n7133) );
  AND U6758 ( .A(n945), .B(n7140), .Z(n7142) );
  XNOR U6759 ( .A(n7141), .B(n7138), .Z(n7140) );
  XOR U6760 ( .A(n7143), .B(n7144), .Z(n7138) );
  AND U6761 ( .A(n948), .B(n7145), .Z(n7144) );
  XOR U6762 ( .A(p_input[1331]), .B(n7143), .Z(n7145) );
  XOR U6763 ( .A(n7146), .B(n7147), .Z(n7143) );
  AND U6764 ( .A(n952), .B(n7148), .Z(n7147) );
  XOR U6765 ( .A(n7149), .B(n7150), .Z(n7141) );
  AND U6766 ( .A(n956), .B(n7148), .Z(n7150) );
  XNOR U6767 ( .A(n7149), .B(n7146), .Z(n7148) );
  XOR U6768 ( .A(n7151), .B(n7152), .Z(n7146) );
  AND U6769 ( .A(n959), .B(n7153), .Z(n7152) );
  XOR U6770 ( .A(p_input[1347]), .B(n7151), .Z(n7153) );
  XOR U6771 ( .A(n7154), .B(n7155), .Z(n7151) );
  AND U6772 ( .A(n963), .B(n7156), .Z(n7155) );
  XOR U6773 ( .A(n7157), .B(n7158), .Z(n7149) );
  AND U6774 ( .A(n967), .B(n7156), .Z(n7158) );
  XNOR U6775 ( .A(n7157), .B(n7154), .Z(n7156) );
  XOR U6776 ( .A(n7159), .B(n7160), .Z(n7154) );
  AND U6777 ( .A(n970), .B(n7161), .Z(n7160) );
  XOR U6778 ( .A(p_input[1363]), .B(n7159), .Z(n7161) );
  XOR U6779 ( .A(n7162), .B(n7163), .Z(n7159) );
  AND U6780 ( .A(n974), .B(n7164), .Z(n7163) );
  XOR U6781 ( .A(n7165), .B(n7166), .Z(n7157) );
  AND U6782 ( .A(n978), .B(n7164), .Z(n7166) );
  XNOR U6783 ( .A(n7165), .B(n7162), .Z(n7164) );
  XOR U6784 ( .A(n7167), .B(n7168), .Z(n7162) );
  AND U6785 ( .A(n981), .B(n7169), .Z(n7168) );
  XOR U6786 ( .A(p_input[1379]), .B(n7167), .Z(n7169) );
  XOR U6787 ( .A(n7170), .B(n7171), .Z(n7167) );
  AND U6788 ( .A(n985), .B(n7172), .Z(n7171) );
  XOR U6789 ( .A(n7173), .B(n7174), .Z(n7165) );
  AND U6790 ( .A(n989), .B(n7172), .Z(n7174) );
  XNOR U6791 ( .A(n7173), .B(n7170), .Z(n7172) );
  XOR U6792 ( .A(n7175), .B(n7176), .Z(n7170) );
  AND U6793 ( .A(n992), .B(n7177), .Z(n7176) );
  XOR U6794 ( .A(p_input[1395]), .B(n7175), .Z(n7177) );
  XOR U6795 ( .A(n7178), .B(n7179), .Z(n7175) );
  AND U6796 ( .A(n996), .B(n7180), .Z(n7179) );
  XOR U6797 ( .A(n7181), .B(n7182), .Z(n7173) );
  AND U6798 ( .A(n1000), .B(n7180), .Z(n7182) );
  XNOR U6799 ( .A(n7181), .B(n7178), .Z(n7180) );
  XOR U6800 ( .A(n7183), .B(n7184), .Z(n7178) );
  AND U6801 ( .A(n1003), .B(n7185), .Z(n7184) );
  XOR U6802 ( .A(p_input[1411]), .B(n7183), .Z(n7185) );
  XOR U6803 ( .A(n7186), .B(n7187), .Z(n7183) );
  AND U6804 ( .A(n1007), .B(n7188), .Z(n7187) );
  XOR U6805 ( .A(n7189), .B(n7190), .Z(n7181) );
  AND U6806 ( .A(n1011), .B(n7188), .Z(n7190) );
  XNOR U6807 ( .A(n7189), .B(n7186), .Z(n7188) );
  XOR U6808 ( .A(n7191), .B(n7192), .Z(n7186) );
  AND U6809 ( .A(n1014), .B(n7193), .Z(n7192) );
  XOR U6810 ( .A(p_input[1427]), .B(n7191), .Z(n7193) );
  XOR U6811 ( .A(n7194), .B(n7195), .Z(n7191) );
  AND U6812 ( .A(n1018), .B(n7196), .Z(n7195) );
  XOR U6813 ( .A(n7197), .B(n7198), .Z(n7189) );
  AND U6814 ( .A(n1022), .B(n7196), .Z(n7198) );
  XNOR U6815 ( .A(n7197), .B(n7194), .Z(n7196) );
  XOR U6816 ( .A(n7199), .B(n7200), .Z(n7194) );
  AND U6817 ( .A(n1025), .B(n7201), .Z(n7200) );
  XOR U6818 ( .A(p_input[1443]), .B(n7199), .Z(n7201) );
  XOR U6819 ( .A(n7202), .B(n7203), .Z(n7199) );
  AND U6820 ( .A(n1029), .B(n7204), .Z(n7203) );
  XOR U6821 ( .A(n7205), .B(n7206), .Z(n7197) );
  AND U6822 ( .A(n1033), .B(n7204), .Z(n7206) );
  XNOR U6823 ( .A(n7205), .B(n7202), .Z(n7204) );
  XOR U6824 ( .A(n7207), .B(n7208), .Z(n7202) );
  AND U6825 ( .A(n1036), .B(n7209), .Z(n7208) );
  XOR U6826 ( .A(p_input[1459]), .B(n7207), .Z(n7209) );
  XOR U6827 ( .A(n7210), .B(n7211), .Z(n7207) );
  AND U6828 ( .A(n1040), .B(n7212), .Z(n7211) );
  XOR U6829 ( .A(n7213), .B(n7214), .Z(n7205) );
  AND U6830 ( .A(n1044), .B(n7212), .Z(n7214) );
  XNOR U6831 ( .A(n7213), .B(n7210), .Z(n7212) );
  XOR U6832 ( .A(n7215), .B(n7216), .Z(n7210) );
  AND U6833 ( .A(n1047), .B(n7217), .Z(n7216) );
  XOR U6834 ( .A(p_input[1475]), .B(n7215), .Z(n7217) );
  XOR U6835 ( .A(n7218), .B(n7219), .Z(n7215) );
  AND U6836 ( .A(n1051), .B(n7220), .Z(n7219) );
  XOR U6837 ( .A(n7221), .B(n7222), .Z(n7213) );
  AND U6838 ( .A(n1055), .B(n7220), .Z(n7222) );
  XNOR U6839 ( .A(n7221), .B(n7218), .Z(n7220) );
  XOR U6840 ( .A(n7223), .B(n7224), .Z(n7218) );
  AND U6841 ( .A(n1058), .B(n7225), .Z(n7224) );
  XOR U6842 ( .A(p_input[1491]), .B(n7223), .Z(n7225) );
  XOR U6843 ( .A(n7226), .B(n7227), .Z(n7223) );
  AND U6844 ( .A(n1062), .B(n7228), .Z(n7227) );
  XOR U6845 ( .A(n7229), .B(n7230), .Z(n7221) );
  AND U6846 ( .A(n1066), .B(n7228), .Z(n7230) );
  XNOR U6847 ( .A(n7229), .B(n7226), .Z(n7228) );
  XOR U6848 ( .A(n7231), .B(n7232), .Z(n7226) );
  AND U6849 ( .A(n1069), .B(n7233), .Z(n7232) );
  XOR U6850 ( .A(p_input[1507]), .B(n7231), .Z(n7233) );
  XOR U6851 ( .A(n7234), .B(n7235), .Z(n7231) );
  AND U6852 ( .A(n1073), .B(n7236), .Z(n7235) );
  XOR U6853 ( .A(n7237), .B(n7238), .Z(n7229) );
  AND U6854 ( .A(n1077), .B(n7236), .Z(n7238) );
  XNOR U6855 ( .A(n7237), .B(n7234), .Z(n7236) );
  XOR U6856 ( .A(n7239), .B(n7240), .Z(n7234) );
  AND U6857 ( .A(n1080), .B(n7241), .Z(n7240) );
  XOR U6858 ( .A(p_input[1523]), .B(n7239), .Z(n7241) );
  XOR U6859 ( .A(n7242), .B(n7243), .Z(n7239) );
  AND U6860 ( .A(n1084), .B(n7244), .Z(n7243) );
  XOR U6861 ( .A(n7245), .B(n7246), .Z(n7237) );
  AND U6862 ( .A(n1088), .B(n7244), .Z(n7246) );
  XNOR U6863 ( .A(n7245), .B(n7242), .Z(n7244) );
  XOR U6864 ( .A(n7247), .B(n7248), .Z(n7242) );
  AND U6865 ( .A(n1091), .B(n7249), .Z(n7248) );
  XOR U6866 ( .A(p_input[1539]), .B(n7247), .Z(n7249) );
  XOR U6867 ( .A(n7250), .B(n7251), .Z(n7247) );
  AND U6868 ( .A(n1095), .B(n7252), .Z(n7251) );
  XOR U6869 ( .A(n7253), .B(n7254), .Z(n7245) );
  AND U6870 ( .A(n1099), .B(n7252), .Z(n7254) );
  XNOR U6871 ( .A(n7253), .B(n7250), .Z(n7252) );
  XOR U6872 ( .A(n7255), .B(n7256), .Z(n7250) );
  AND U6873 ( .A(n1102), .B(n7257), .Z(n7256) );
  XOR U6874 ( .A(p_input[1555]), .B(n7255), .Z(n7257) );
  XOR U6875 ( .A(n7258), .B(n7259), .Z(n7255) );
  AND U6876 ( .A(n1106), .B(n7260), .Z(n7259) );
  XOR U6877 ( .A(n7261), .B(n7262), .Z(n7253) );
  AND U6878 ( .A(n1110), .B(n7260), .Z(n7262) );
  XNOR U6879 ( .A(n7261), .B(n7258), .Z(n7260) );
  XOR U6880 ( .A(n7263), .B(n7264), .Z(n7258) );
  AND U6881 ( .A(n1113), .B(n7265), .Z(n7264) );
  XOR U6882 ( .A(p_input[1571]), .B(n7263), .Z(n7265) );
  XOR U6883 ( .A(n7266), .B(n7267), .Z(n7263) );
  AND U6884 ( .A(n1117), .B(n7268), .Z(n7267) );
  XOR U6885 ( .A(n7269), .B(n7270), .Z(n7261) );
  AND U6886 ( .A(n1121), .B(n7268), .Z(n7270) );
  XNOR U6887 ( .A(n7269), .B(n7266), .Z(n7268) );
  XOR U6888 ( .A(n7271), .B(n7272), .Z(n7266) );
  AND U6889 ( .A(n1124), .B(n7273), .Z(n7272) );
  XOR U6890 ( .A(p_input[1587]), .B(n7271), .Z(n7273) );
  XOR U6891 ( .A(n7274), .B(n7275), .Z(n7271) );
  AND U6892 ( .A(n1128), .B(n7276), .Z(n7275) );
  XOR U6893 ( .A(n7277), .B(n7278), .Z(n7269) );
  AND U6894 ( .A(n1132), .B(n7276), .Z(n7278) );
  XNOR U6895 ( .A(n7277), .B(n7274), .Z(n7276) );
  XOR U6896 ( .A(n7279), .B(n7280), .Z(n7274) );
  AND U6897 ( .A(n1135), .B(n7281), .Z(n7280) );
  XOR U6898 ( .A(p_input[1603]), .B(n7279), .Z(n7281) );
  XOR U6899 ( .A(n7282), .B(n7283), .Z(n7279) );
  AND U6900 ( .A(n1139), .B(n7284), .Z(n7283) );
  XOR U6901 ( .A(n7285), .B(n7286), .Z(n7277) );
  AND U6902 ( .A(n1143), .B(n7284), .Z(n7286) );
  XNOR U6903 ( .A(n7285), .B(n7282), .Z(n7284) );
  XOR U6904 ( .A(n7287), .B(n7288), .Z(n7282) );
  AND U6905 ( .A(n1146), .B(n7289), .Z(n7288) );
  XOR U6906 ( .A(p_input[1619]), .B(n7287), .Z(n7289) );
  XOR U6907 ( .A(n7290), .B(n7291), .Z(n7287) );
  AND U6908 ( .A(n1150), .B(n7292), .Z(n7291) );
  XOR U6909 ( .A(n7293), .B(n7294), .Z(n7285) );
  AND U6910 ( .A(n1154), .B(n7292), .Z(n7294) );
  XNOR U6911 ( .A(n7293), .B(n7290), .Z(n7292) );
  XOR U6912 ( .A(n7295), .B(n7296), .Z(n7290) );
  AND U6913 ( .A(n1157), .B(n7297), .Z(n7296) );
  XOR U6914 ( .A(p_input[1635]), .B(n7295), .Z(n7297) );
  XOR U6915 ( .A(n7298), .B(n7299), .Z(n7295) );
  AND U6916 ( .A(n1161), .B(n7300), .Z(n7299) );
  XOR U6917 ( .A(n7301), .B(n7302), .Z(n7293) );
  AND U6918 ( .A(n1165), .B(n7300), .Z(n7302) );
  XNOR U6919 ( .A(n7301), .B(n7298), .Z(n7300) );
  XOR U6920 ( .A(n7303), .B(n7304), .Z(n7298) );
  AND U6921 ( .A(n1168), .B(n7305), .Z(n7304) );
  XOR U6922 ( .A(p_input[1651]), .B(n7303), .Z(n7305) );
  XOR U6923 ( .A(n7306), .B(n7307), .Z(n7303) );
  AND U6924 ( .A(n1172), .B(n7308), .Z(n7307) );
  XOR U6925 ( .A(n7309), .B(n7310), .Z(n7301) );
  AND U6926 ( .A(n1176), .B(n7308), .Z(n7310) );
  XNOR U6927 ( .A(n7309), .B(n7306), .Z(n7308) );
  XOR U6928 ( .A(n7311), .B(n7312), .Z(n7306) );
  AND U6929 ( .A(n1179), .B(n7313), .Z(n7312) );
  XOR U6930 ( .A(p_input[1667]), .B(n7311), .Z(n7313) );
  XOR U6931 ( .A(n7314), .B(n7315), .Z(n7311) );
  AND U6932 ( .A(n1183), .B(n7316), .Z(n7315) );
  XOR U6933 ( .A(n7317), .B(n7318), .Z(n7309) );
  AND U6934 ( .A(n1187), .B(n7316), .Z(n7318) );
  XNOR U6935 ( .A(n7317), .B(n7314), .Z(n7316) );
  XOR U6936 ( .A(n7319), .B(n7320), .Z(n7314) );
  AND U6937 ( .A(n1190), .B(n7321), .Z(n7320) );
  XOR U6938 ( .A(p_input[1683]), .B(n7319), .Z(n7321) );
  XOR U6939 ( .A(n7322), .B(n7323), .Z(n7319) );
  AND U6940 ( .A(n1194), .B(n7324), .Z(n7323) );
  XOR U6941 ( .A(n7325), .B(n7326), .Z(n7317) );
  AND U6942 ( .A(n1198), .B(n7324), .Z(n7326) );
  XNOR U6943 ( .A(n7325), .B(n7322), .Z(n7324) );
  XOR U6944 ( .A(n7327), .B(n7328), .Z(n7322) );
  AND U6945 ( .A(n1201), .B(n7329), .Z(n7328) );
  XOR U6946 ( .A(p_input[1699]), .B(n7327), .Z(n7329) );
  XOR U6947 ( .A(n7330), .B(n7331), .Z(n7327) );
  AND U6948 ( .A(n1205), .B(n7332), .Z(n7331) );
  XOR U6949 ( .A(n7333), .B(n7334), .Z(n7325) );
  AND U6950 ( .A(n1209), .B(n7332), .Z(n7334) );
  XNOR U6951 ( .A(n7333), .B(n7330), .Z(n7332) );
  XOR U6952 ( .A(n7335), .B(n7336), .Z(n7330) );
  AND U6953 ( .A(n1212), .B(n7337), .Z(n7336) );
  XOR U6954 ( .A(p_input[1715]), .B(n7335), .Z(n7337) );
  XOR U6955 ( .A(n7338), .B(n7339), .Z(n7335) );
  AND U6956 ( .A(n1216), .B(n7340), .Z(n7339) );
  XOR U6957 ( .A(n7341), .B(n7342), .Z(n7333) );
  AND U6958 ( .A(n1220), .B(n7340), .Z(n7342) );
  XNOR U6959 ( .A(n7341), .B(n7338), .Z(n7340) );
  XOR U6960 ( .A(n7343), .B(n7344), .Z(n7338) );
  AND U6961 ( .A(n1223), .B(n7345), .Z(n7344) );
  XOR U6962 ( .A(p_input[1731]), .B(n7343), .Z(n7345) );
  XOR U6963 ( .A(n7346), .B(n7347), .Z(n7343) );
  AND U6964 ( .A(n1227), .B(n7348), .Z(n7347) );
  XOR U6965 ( .A(n7349), .B(n7350), .Z(n7341) );
  AND U6966 ( .A(n1231), .B(n7348), .Z(n7350) );
  XNOR U6967 ( .A(n7349), .B(n7346), .Z(n7348) );
  XOR U6968 ( .A(n7351), .B(n7352), .Z(n7346) );
  AND U6969 ( .A(n1234), .B(n7353), .Z(n7352) );
  XOR U6970 ( .A(p_input[1747]), .B(n7351), .Z(n7353) );
  XOR U6971 ( .A(n7354), .B(n7355), .Z(n7351) );
  AND U6972 ( .A(n1238), .B(n7356), .Z(n7355) );
  XOR U6973 ( .A(n7357), .B(n7358), .Z(n7349) );
  AND U6974 ( .A(n1242), .B(n7356), .Z(n7358) );
  XNOR U6975 ( .A(n7357), .B(n7354), .Z(n7356) );
  XOR U6976 ( .A(n7359), .B(n7360), .Z(n7354) );
  AND U6977 ( .A(n1245), .B(n7361), .Z(n7360) );
  XOR U6978 ( .A(p_input[1763]), .B(n7359), .Z(n7361) );
  XOR U6979 ( .A(n7362), .B(n7363), .Z(n7359) );
  AND U6980 ( .A(n1249), .B(n7364), .Z(n7363) );
  XOR U6981 ( .A(n7365), .B(n7366), .Z(n7357) );
  AND U6982 ( .A(n1253), .B(n7364), .Z(n7366) );
  XNOR U6983 ( .A(n7365), .B(n7362), .Z(n7364) );
  XOR U6984 ( .A(n7367), .B(n7368), .Z(n7362) );
  AND U6985 ( .A(n1256), .B(n7369), .Z(n7368) );
  XOR U6986 ( .A(p_input[1779]), .B(n7367), .Z(n7369) );
  XOR U6987 ( .A(n7370), .B(n7371), .Z(n7367) );
  AND U6988 ( .A(n1260), .B(n7372), .Z(n7371) );
  XOR U6989 ( .A(n7373), .B(n7374), .Z(n7365) );
  AND U6990 ( .A(n1264), .B(n7372), .Z(n7374) );
  XNOR U6991 ( .A(n7373), .B(n7370), .Z(n7372) );
  XOR U6992 ( .A(n7375), .B(n7376), .Z(n7370) );
  AND U6993 ( .A(n1267), .B(n7377), .Z(n7376) );
  XOR U6994 ( .A(p_input[1795]), .B(n7375), .Z(n7377) );
  XOR U6995 ( .A(n7378), .B(n7379), .Z(n7375) );
  AND U6996 ( .A(n1271), .B(n7380), .Z(n7379) );
  XOR U6997 ( .A(n7381), .B(n7382), .Z(n7373) );
  AND U6998 ( .A(n1275), .B(n7380), .Z(n7382) );
  XNOR U6999 ( .A(n7381), .B(n7378), .Z(n7380) );
  XOR U7000 ( .A(n7383), .B(n7384), .Z(n7378) );
  AND U7001 ( .A(n1278), .B(n7385), .Z(n7384) );
  XOR U7002 ( .A(p_input[1811]), .B(n7383), .Z(n7385) );
  XOR U7003 ( .A(n7386), .B(n7387), .Z(n7383) );
  AND U7004 ( .A(n1282), .B(n7388), .Z(n7387) );
  XOR U7005 ( .A(n7389), .B(n7390), .Z(n7381) );
  AND U7006 ( .A(n1286), .B(n7388), .Z(n7390) );
  XNOR U7007 ( .A(n7389), .B(n7386), .Z(n7388) );
  XOR U7008 ( .A(n7391), .B(n7392), .Z(n7386) );
  AND U7009 ( .A(n1289), .B(n7393), .Z(n7392) );
  XOR U7010 ( .A(p_input[1827]), .B(n7391), .Z(n7393) );
  XOR U7011 ( .A(n7394), .B(n7395), .Z(n7391) );
  AND U7012 ( .A(n1293), .B(n7396), .Z(n7395) );
  XOR U7013 ( .A(n7397), .B(n7398), .Z(n7389) );
  AND U7014 ( .A(n1297), .B(n7396), .Z(n7398) );
  XNOR U7015 ( .A(n7397), .B(n7394), .Z(n7396) );
  XOR U7016 ( .A(n7399), .B(n7400), .Z(n7394) );
  AND U7017 ( .A(n1300), .B(n7401), .Z(n7400) );
  XOR U7018 ( .A(p_input[1843]), .B(n7399), .Z(n7401) );
  XOR U7019 ( .A(n7402), .B(n7403), .Z(n7399) );
  AND U7020 ( .A(n1304), .B(n7404), .Z(n7403) );
  XOR U7021 ( .A(n7405), .B(n7406), .Z(n7397) );
  AND U7022 ( .A(n1308), .B(n7404), .Z(n7406) );
  XNOR U7023 ( .A(n7405), .B(n7402), .Z(n7404) );
  XOR U7024 ( .A(n7407), .B(n7408), .Z(n7402) );
  AND U7025 ( .A(n1311), .B(n7409), .Z(n7408) );
  XOR U7026 ( .A(p_input[1859]), .B(n7407), .Z(n7409) );
  XOR U7027 ( .A(n7410), .B(n7411), .Z(n7407) );
  AND U7028 ( .A(n1315), .B(n7412), .Z(n7411) );
  XOR U7029 ( .A(n7413), .B(n7414), .Z(n7405) );
  AND U7030 ( .A(n1319), .B(n7412), .Z(n7414) );
  XNOR U7031 ( .A(n7413), .B(n7410), .Z(n7412) );
  XOR U7032 ( .A(n7415), .B(n7416), .Z(n7410) );
  AND U7033 ( .A(n1322), .B(n7417), .Z(n7416) );
  XOR U7034 ( .A(p_input[1875]), .B(n7415), .Z(n7417) );
  XOR U7035 ( .A(n7418), .B(n7419), .Z(n7415) );
  AND U7036 ( .A(n1326), .B(n7420), .Z(n7419) );
  XOR U7037 ( .A(n7421), .B(n7422), .Z(n7413) );
  AND U7038 ( .A(n1330), .B(n7420), .Z(n7422) );
  XNOR U7039 ( .A(n7421), .B(n7418), .Z(n7420) );
  XOR U7040 ( .A(n7423), .B(n7424), .Z(n7418) );
  AND U7041 ( .A(n1333), .B(n7425), .Z(n7424) );
  XOR U7042 ( .A(p_input[1891]), .B(n7423), .Z(n7425) );
  XOR U7043 ( .A(n7426), .B(n7427), .Z(n7423) );
  AND U7044 ( .A(n1337), .B(n7428), .Z(n7427) );
  XOR U7045 ( .A(n7429), .B(n7430), .Z(n7421) );
  AND U7046 ( .A(n1341), .B(n7428), .Z(n7430) );
  XNOR U7047 ( .A(n7429), .B(n7426), .Z(n7428) );
  XOR U7048 ( .A(n7431), .B(n7432), .Z(n7426) );
  AND U7049 ( .A(n1344), .B(n7433), .Z(n7432) );
  XOR U7050 ( .A(p_input[1907]), .B(n7431), .Z(n7433) );
  XOR U7051 ( .A(n7434), .B(n7435), .Z(n7431) );
  AND U7052 ( .A(n1348), .B(n7436), .Z(n7435) );
  XOR U7053 ( .A(n7437), .B(n7438), .Z(n7429) );
  AND U7054 ( .A(n1352), .B(n7436), .Z(n7438) );
  XNOR U7055 ( .A(n7437), .B(n7434), .Z(n7436) );
  XOR U7056 ( .A(n7439), .B(n7440), .Z(n7434) );
  AND U7057 ( .A(n1355), .B(n7441), .Z(n7440) );
  XOR U7058 ( .A(p_input[1923]), .B(n7439), .Z(n7441) );
  XOR U7059 ( .A(n7442), .B(n7443), .Z(n7439) );
  AND U7060 ( .A(n1359), .B(n7444), .Z(n7443) );
  XOR U7061 ( .A(n7445), .B(n7446), .Z(n7437) );
  AND U7062 ( .A(n1363), .B(n7444), .Z(n7446) );
  XNOR U7063 ( .A(n7445), .B(n7442), .Z(n7444) );
  XOR U7064 ( .A(n7447), .B(n7448), .Z(n7442) );
  AND U7065 ( .A(n1366), .B(n7449), .Z(n7448) );
  XOR U7066 ( .A(p_input[1939]), .B(n7447), .Z(n7449) );
  XOR U7067 ( .A(n7450), .B(n7451), .Z(n7447) );
  AND U7068 ( .A(n1370), .B(n7452), .Z(n7451) );
  XOR U7069 ( .A(n7453), .B(n7454), .Z(n7445) );
  AND U7070 ( .A(n1374), .B(n7452), .Z(n7454) );
  XNOR U7071 ( .A(n7453), .B(n7450), .Z(n7452) );
  XOR U7072 ( .A(n7455), .B(n7456), .Z(n7450) );
  AND U7073 ( .A(n1377), .B(n7457), .Z(n7456) );
  XOR U7074 ( .A(p_input[1955]), .B(n7455), .Z(n7457) );
  XOR U7075 ( .A(n7458), .B(n7459), .Z(n7455) );
  AND U7076 ( .A(n1381), .B(n7460), .Z(n7459) );
  XOR U7077 ( .A(n7461), .B(n7462), .Z(n7453) );
  AND U7078 ( .A(n1385), .B(n7460), .Z(n7462) );
  XNOR U7079 ( .A(n7461), .B(n7458), .Z(n7460) );
  XOR U7080 ( .A(n7463), .B(n7464), .Z(n7458) );
  AND U7081 ( .A(n1388), .B(n7465), .Z(n7464) );
  XOR U7082 ( .A(p_input[1971]), .B(n7463), .Z(n7465) );
  XOR U7083 ( .A(n7466), .B(n7467), .Z(n7463) );
  AND U7084 ( .A(n1392), .B(n7468), .Z(n7467) );
  XOR U7085 ( .A(n7469), .B(n7470), .Z(n7461) );
  AND U7086 ( .A(n1396), .B(n7468), .Z(n7470) );
  XNOR U7087 ( .A(n7469), .B(n7466), .Z(n7468) );
  XOR U7088 ( .A(n7471), .B(n7472), .Z(n7466) );
  AND U7089 ( .A(n1399), .B(n7473), .Z(n7472) );
  XOR U7090 ( .A(p_input[1987]), .B(n7471), .Z(n7473) );
  XOR U7091 ( .A(n7474), .B(n7475), .Z(n7471) );
  AND U7092 ( .A(n1403), .B(n7476), .Z(n7475) );
  XOR U7093 ( .A(n7477), .B(n7478), .Z(n7469) );
  AND U7094 ( .A(n1407), .B(n7476), .Z(n7478) );
  XNOR U7095 ( .A(n7477), .B(n7474), .Z(n7476) );
  XOR U7096 ( .A(n7479), .B(n7480), .Z(n7474) );
  AND U7097 ( .A(n1410), .B(n7481), .Z(n7480) );
  XOR U7098 ( .A(p_input[2003]), .B(n7479), .Z(n7481) );
  XNOR U7099 ( .A(n7482), .B(n7483), .Z(n7479) );
  AND U7100 ( .A(n1414), .B(n7484), .Z(n7483) );
  XNOR U7101 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n7485), .Z(n7477) );
  AND U7102 ( .A(n1417), .B(n7484), .Z(n7485) );
  XOR U7103 ( .A(n7486), .B(n7482), .Z(n7484) );
  XOR U7104 ( .A(n19), .B(n7487), .Z(o[18]) );
  AND U7105 ( .A(n30), .B(n7488), .Z(n19) );
  XOR U7106 ( .A(n20), .B(n7487), .Z(n7488) );
  XOR U7107 ( .A(n7489), .B(n7490), .Z(n7487) );
  AND U7108 ( .A(n34), .B(n7491), .Z(n7490) );
  XOR U7109 ( .A(p_input[2]), .B(n7489), .Z(n7491) );
  XOR U7110 ( .A(n7492), .B(n7493), .Z(n7489) );
  AND U7111 ( .A(n38), .B(n7494), .Z(n7493) );
  XOR U7112 ( .A(n7495), .B(n7496), .Z(n20) );
  AND U7113 ( .A(n42), .B(n7494), .Z(n7496) );
  XNOR U7114 ( .A(n7497), .B(n7492), .Z(n7494) );
  XOR U7115 ( .A(n7498), .B(n7499), .Z(n7492) );
  AND U7116 ( .A(n46), .B(n7500), .Z(n7499) );
  XOR U7117 ( .A(p_input[18]), .B(n7498), .Z(n7500) );
  XOR U7118 ( .A(n7501), .B(n7502), .Z(n7498) );
  AND U7119 ( .A(n50), .B(n7503), .Z(n7502) );
  IV U7120 ( .A(n7495), .Z(n7497) );
  XNOR U7121 ( .A(n7504), .B(n7505), .Z(n7495) );
  AND U7122 ( .A(n54), .B(n7503), .Z(n7505) );
  XNOR U7123 ( .A(n7504), .B(n7501), .Z(n7503) );
  XOR U7124 ( .A(n7506), .B(n7507), .Z(n7501) );
  AND U7125 ( .A(n57), .B(n7508), .Z(n7507) );
  XOR U7126 ( .A(p_input[34]), .B(n7506), .Z(n7508) );
  XOR U7127 ( .A(n7509), .B(n7510), .Z(n7506) );
  AND U7128 ( .A(n61), .B(n7511), .Z(n7510) );
  XOR U7129 ( .A(n7512), .B(n7513), .Z(n7504) );
  AND U7130 ( .A(n65), .B(n7511), .Z(n7513) );
  XNOR U7131 ( .A(n7512), .B(n7509), .Z(n7511) );
  XOR U7132 ( .A(n7514), .B(n7515), .Z(n7509) );
  AND U7133 ( .A(n68), .B(n7516), .Z(n7515) );
  XOR U7134 ( .A(p_input[50]), .B(n7514), .Z(n7516) );
  XOR U7135 ( .A(n7517), .B(n7518), .Z(n7514) );
  AND U7136 ( .A(n72), .B(n7519), .Z(n7518) );
  XOR U7137 ( .A(n7520), .B(n7521), .Z(n7512) );
  AND U7138 ( .A(n76), .B(n7519), .Z(n7521) );
  XNOR U7139 ( .A(n7520), .B(n7517), .Z(n7519) );
  XOR U7140 ( .A(n7522), .B(n7523), .Z(n7517) );
  AND U7141 ( .A(n79), .B(n7524), .Z(n7523) );
  XOR U7142 ( .A(p_input[66]), .B(n7522), .Z(n7524) );
  XOR U7143 ( .A(n7525), .B(n7526), .Z(n7522) );
  AND U7144 ( .A(n83), .B(n7527), .Z(n7526) );
  XOR U7145 ( .A(n7528), .B(n7529), .Z(n7520) );
  AND U7146 ( .A(n87), .B(n7527), .Z(n7529) );
  XNOR U7147 ( .A(n7528), .B(n7525), .Z(n7527) );
  XOR U7148 ( .A(n7530), .B(n7531), .Z(n7525) );
  AND U7149 ( .A(n90), .B(n7532), .Z(n7531) );
  XOR U7150 ( .A(p_input[82]), .B(n7530), .Z(n7532) );
  XOR U7151 ( .A(n7533), .B(n7534), .Z(n7530) );
  AND U7152 ( .A(n94), .B(n7535), .Z(n7534) );
  XOR U7153 ( .A(n7536), .B(n7537), .Z(n7528) );
  AND U7154 ( .A(n98), .B(n7535), .Z(n7537) );
  XNOR U7155 ( .A(n7536), .B(n7533), .Z(n7535) );
  XOR U7156 ( .A(n7538), .B(n7539), .Z(n7533) );
  AND U7157 ( .A(n101), .B(n7540), .Z(n7539) );
  XOR U7158 ( .A(p_input[98]), .B(n7538), .Z(n7540) );
  XOR U7159 ( .A(n7541), .B(n7542), .Z(n7538) );
  AND U7160 ( .A(n105), .B(n7543), .Z(n7542) );
  XOR U7161 ( .A(n7544), .B(n7545), .Z(n7536) );
  AND U7162 ( .A(n109), .B(n7543), .Z(n7545) );
  XNOR U7163 ( .A(n7544), .B(n7541), .Z(n7543) );
  XOR U7164 ( .A(n7546), .B(n7547), .Z(n7541) );
  AND U7165 ( .A(n112), .B(n7548), .Z(n7547) );
  XOR U7166 ( .A(p_input[114]), .B(n7546), .Z(n7548) );
  XOR U7167 ( .A(n7549), .B(n7550), .Z(n7546) );
  AND U7168 ( .A(n116), .B(n7551), .Z(n7550) );
  XOR U7169 ( .A(n7552), .B(n7553), .Z(n7544) );
  AND U7170 ( .A(n120), .B(n7551), .Z(n7553) );
  XNOR U7171 ( .A(n7552), .B(n7549), .Z(n7551) );
  XOR U7172 ( .A(n7554), .B(n7555), .Z(n7549) );
  AND U7173 ( .A(n123), .B(n7556), .Z(n7555) );
  XOR U7174 ( .A(p_input[130]), .B(n7554), .Z(n7556) );
  XOR U7175 ( .A(n7557), .B(n7558), .Z(n7554) );
  AND U7176 ( .A(n127), .B(n7559), .Z(n7558) );
  XOR U7177 ( .A(n7560), .B(n7561), .Z(n7552) );
  AND U7178 ( .A(n131), .B(n7559), .Z(n7561) );
  XNOR U7179 ( .A(n7560), .B(n7557), .Z(n7559) );
  XOR U7180 ( .A(n7562), .B(n7563), .Z(n7557) );
  AND U7181 ( .A(n134), .B(n7564), .Z(n7563) );
  XOR U7182 ( .A(p_input[146]), .B(n7562), .Z(n7564) );
  XOR U7183 ( .A(n7565), .B(n7566), .Z(n7562) );
  AND U7184 ( .A(n138), .B(n7567), .Z(n7566) );
  XOR U7185 ( .A(n7568), .B(n7569), .Z(n7560) );
  AND U7186 ( .A(n142), .B(n7567), .Z(n7569) );
  XNOR U7187 ( .A(n7568), .B(n7565), .Z(n7567) );
  XOR U7188 ( .A(n7570), .B(n7571), .Z(n7565) );
  AND U7189 ( .A(n145), .B(n7572), .Z(n7571) );
  XOR U7190 ( .A(p_input[162]), .B(n7570), .Z(n7572) );
  XOR U7191 ( .A(n7573), .B(n7574), .Z(n7570) );
  AND U7192 ( .A(n149), .B(n7575), .Z(n7574) );
  XOR U7193 ( .A(n7576), .B(n7577), .Z(n7568) );
  AND U7194 ( .A(n153), .B(n7575), .Z(n7577) );
  XNOR U7195 ( .A(n7576), .B(n7573), .Z(n7575) );
  XOR U7196 ( .A(n7578), .B(n7579), .Z(n7573) );
  AND U7197 ( .A(n156), .B(n7580), .Z(n7579) );
  XOR U7198 ( .A(p_input[178]), .B(n7578), .Z(n7580) );
  XOR U7199 ( .A(n7581), .B(n7582), .Z(n7578) );
  AND U7200 ( .A(n160), .B(n7583), .Z(n7582) );
  XOR U7201 ( .A(n7584), .B(n7585), .Z(n7576) );
  AND U7202 ( .A(n164), .B(n7583), .Z(n7585) );
  XNOR U7203 ( .A(n7584), .B(n7581), .Z(n7583) );
  XOR U7204 ( .A(n7586), .B(n7587), .Z(n7581) );
  AND U7205 ( .A(n167), .B(n7588), .Z(n7587) );
  XOR U7206 ( .A(p_input[194]), .B(n7586), .Z(n7588) );
  XOR U7207 ( .A(n7589), .B(n7590), .Z(n7586) );
  AND U7208 ( .A(n171), .B(n7591), .Z(n7590) );
  XOR U7209 ( .A(n7592), .B(n7593), .Z(n7584) );
  AND U7210 ( .A(n175), .B(n7591), .Z(n7593) );
  XNOR U7211 ( .A(n7592), .B(n7589), .Z(n7591) );
  XOR U7212 ( .A(n7594), .B(n7595), .Z(n7589) );
  AND U7213 ( .A(n178), .B(n7596), .Z(n7595) );
  XOR U7214 ( .A(p_input[210]), .B(n7594), .Z(n7596) );
  XOR U7215 ( .A(n7597), .B(n7598), .Z(n7594) );
  AND U7216 ( .A(n182), .B(n7599), .Z(n7598) );
  XOR U7217 ( .A(n7600), .B(n7601), .Z(n7592) );
  AND U7218 ( .A(n186), .B(n7599), .Z(n7601) );
  XNOR U7219 ( .A(n7600), .B(n7597), .Z(n7599) );
  XOR U7220 ( .A(n7602), .B(n7603), .Z(n7597) );
  AND U7221 ( .A(n189), .B(n7604), .Z(n7603) );
  XOR U7222 ( .A(p_input[226]), .B(n7602), .Z(n7604) );
  XOR U7223 ( .A(n7605), .B(n7606), .Z(n7602) );
  AND U7224 ( .A(n193), .B(n7607), .Z(n7606) );
  XOR U7225 ( .A(n7608), .B(n7609), .Z(n7600) );
  AND U7226 ( .A(n197), .B(n7607), .Z(n7609) );
  XNOR U7227 ( .A(n7608), .B(n7605), .Z(n7607) );
  XOR U7228 ( .A(n7610), .B(n7611), .Z(n7605) );
  AND U7229 ( .A(n200), .B(n7612), .Z(n7611) );
  XOR U7230 ( .A(p_input[242]), .B(n7610), .Z(n7612) );
  XOR U7231 ( .A(n7613), .B(n7614), .Z(n7610) );
  AND U7232 ( .A(n204), .B(n7615), .Z(n7614) );
  XOR U7233 ( .A(n7616), .B(n7617), .Z(n7608) );
  AND U7234 ( .A(n208), .B(n7615), .Z(n7617) );
  XNOR U7235 ( .A(n7616), .B(n7613), .Z(n7615) );
  XOR U7236 ( .A(n7618), .B(n7619), .Z(n7613) );
  AND U7237 ( .A(n211), .B(n7620), .Z(n7619) );
  XOR U7238 ( .A(p_input[258]), .B(n7618), .Z(n7620) );
  XOR U7239 ( .A(n7621), .B(n7622), .Z(n7618) );
  AND U7240 ( .A(n215), .B(n7623), .Z(n7622) );
  XOR U7241 ( .A(n7624), .B(n7625), .Z(n7616) );
  AND U7242 ( .A(n219), .B(n7623), .Z(n7625) );
  XNOR U7243 ( .A(n7624), .B(n7621), .Z(n7623) );
  XOR U7244 ( .A(n7626), .B(n7627), .Z(n7621) );
  AND U7245 ( .A(n222), .B(n7628), .Z(n7627) );
  XOR U7246 ( .A(p_input[274]), .B(n7626), .Z(n7628) );
  XOR U7247 ( .A(n7629), .B(n7630), .Z(n7626) );
  AND U7248 ( .A(n226), .B(n7631), .Z(n7630) );
  XOR U7249 ( .A(n7632), .B(n7633), .Z(n7624) );
  AND U7250 ( .A(n230), .B(n7631), .Z(n7633) );
  XNOR U7251 ( .A(n7632), .B(n7629), .Z(n7631) );
  XOR U7252 ( .A(n7634), .B(n7635), .Z(n7629) );
  AND U7253 ( .A(n233), .B(n7636), .Z(n7635) );
  XOR U7254 ( .A(p_input[290]), .B(n7634), .Z(n7636) );
  XOR U7255 ( .A(n7637), .B(n7638), .Z(n7634) );
  AND U7256 ( .A(n237), .B(n7639), .Z(n7638) );
  XOR U7257 ( .A(n7640), .B(n7641), .Z(n7632) );
  AND U7258 ( .A(n241), .B(n7639), .Z(n7641) );
  XNOR U7259 ( .A(n7640), .B(n7637), .Z(n7639) );
  XOR U7260 ( .A(n7642), .B(n7643), .Z(n7637) );
  AND U7261 ( .A(n244), .B(n7644), .Z(n7643) );
  XOR U7262 ( .A(p_input[306]), .B(n7642), .Z(n7644) );
  XOR U7263 ( .A(n7645), .B(n7646), .Z(n7642) );
  AND U7264 ( .A(n248), .B(n7647), .Z(n7646) );
  XOR U7265 ( .A(n7648), .B(n7649), .Z(n7640) );
  AND U7266 ( .A(n252), .B(n7647), .Z(n7649) );
  XNOR U7267 ( .A(n7648), .B(n7645), .Z(n7647) );
  XOR U7268 ( .A(n7650), .B(n7651), .Z(n7645) );
  AND U7269 ( .A(n255), .B(n7652), .Z(n7651) );
  XOR U7270 ( .A(p_input[322]), .B(n7650), .Z(n7652) );
  XOR U7271 ( .A(n7653), .B(n7654), .Z(n7650) );
  AND U7272 ( .A(n259), .B(n7655), .Z(n7654) );
  XOR U7273 ( .A(n7656), .B(n7657), .Z(n7648) );
  AND U7274 ( .A(n263), .B(n7655), .Z(n7657) );
  XNOR U7275 ( .A(n7656), .B(n7653), .Z(n7655) );
  XOR U7276 ( .A(n7658), .B(n7659), .Z(n7653) );
  AND U7277 ( .A(n266), .B(n7660), .Z(n7659) );
  XOR U7278 ( .A(p_input[338]), .B(n7658), .Z(n7660) );
  XOR U7279 ( .A(n7661), .B(n7662), .Z(n7658) );
  AND U7280 ( .A(n270), .B(n7663), .Z(n7662) );
  XOR U7281 ( .A(n7664), .B(n7665), .Z(n7656) );
  AND U7282 ( .A(n274), .B(n7663), .Z(n7665) );
  XNOR U7283 ( .A(n7664), .B(n7661), .Z(n7663) );
  XOR U7284 ( .A(n7666), .B(n7667), .Z(n7661) );
  AND U7285 ( .A(n277), .B(n7668), .Z(n7667) );
  XOR U7286 ( .A(p_input[354]), .B(n7666), .Z(n7668) );
  XOR U7287 ( .A(n7669), .B(n7670), .Z(n7666) );
  AND U7288 ( .A(n281), .B(n7671), .Z(n7670) );
  XOR U7289 ( .A(n7672), .B(n7673), .Z(n7664) );
  AND U7290 ( .A(n285), .B(n7671), .Z(n7673) );
  XNOR U7291 ( .A(n7672), .B(n7669), .Z(n7671) );
  XOR U7292 ( .A(n7674), .B(n7675), .Z(n7669) );
  AND U7293 ( .A(n288), .B(n7676), .Z(n7675) );
  XOR U7294 ( .A(p_input[370]), .B(n7674), .Z(n7676) );
  XOR U7295 ( .A(n7677), .B(n7678), .Z(n7674) );
  AND U7296 ( .A(n292), .B(n7679), .Z(n7678) );
  XOR U7297 ( .A(n7680), .B(n7681), .Z(n7672) );
  AND U7298 ( .A(n296), .B(n7679), .Z(n7681) );
  XNOR U7299 ( .A(n7680), .B(n7677), .Z(n7679) );
  XOR U7300 ( .A(n7682), .B(n7683), .Z(n7677) );
  AND U7301 ( .A(n299), .B(n7684), .Z(n7683) );
  XOR U7302 ( .A(p_input[386]), .B(n7682), .Z(n7684) );
  XOR U7303 ( .A(n7685), .B(n7686), .Z(n7682) );
  AND U7304 ( .A(n303), .B(n7687), .Z(n7686) );
  XOR U7305 ( .A(n7688), .B(n7689), .Z(n7680) );
  AND U7306 ( .A(n307), .B(n7687), .Z(n7689) );
  XNOR U7307 ( .A(n7688), .B(n7685), .Z(n7687) );
  XOR U7308 ( .A(n7690), .B(n7691), .Z(n7685) );
  AND U7309 ( .A(n310), .B(n7692), .Z(n7691) );
  XOR U7310 ( .A(p_input[402]), .B(n7690), .Z(n7692) );
  XOR U7311 ( .A(n7693), .B(n7694), .Z(n7690) );
  AND U7312 ( .A(n314), .B(n7695), .Z(n7694) );
  XOR U7313 ( .A(n7696), .B(n7697), .Z(n7688) );
  AND U7314 ( .A(n318), .B(n7695), .Z(n7697) );
  XNOR U7315 ( .A(n7696), .B(n7693), .Z(n7695) );
  XOR U7316 ( .A(n7698), .B(n7699), .Z(n7693) );
  AND U7317 ( .A(n321), .B(n7700), .Z(n7699) );
  XOR U7318 ( .A(p_input[418]), .B(n7698), .Z(n7700) );
  XOR U7319 ( .A(n7701), .B(n7702), .Z(n7698) );
  AND U7320 ( .A(n325), .B(n7703), .Z(n7702) );
  XOR U7321 ( .A(n7704), .B(n7705), .Z(n7696) );
  AND U7322 ( .A(n329), .B(n7703), .Z(n7705) );
  XNOR U7323 ( .A(n7704), .B(n7701), .Z(n7703) );
  XOR U7324 ( .A(n7706), .B(n7707), .Z(n7701) );
  AND U7325 ( .A(n332), .B(n7708), .Z(n7707) );
  XOR U7326 ( .A(p_input[434]), .B(n7706), .Z(n7708) );
  XOR U7327 ( .A(n7709), .B(n7710), .Z(n7706) );
  AND U7328 ( .A(n336), .B(n7711), .Z(n7710) );
  XOR U7329 ( .A(n7712), .B(n7713), .Z(n7704) );
  AND U7330 ( .A(n340), .B(n7711), .Z(n7713) );
  XNOR U7331 ( .A(n7712), .B(n7709), .Z(n7711) );
  XOR U7332 ( .A(n7714), .B(n7715), .Z(n7709) );
  AND U7333 ( .A(n343), .B(n7716), .Z(n7715) );
  XOR U7334 ( .A(p_input[450]), .B(n7714), .Z(n7716) );
  XOR U7335 ( .A(n7717), .B(n7718), .Z(n7714) );
  AND U7336 ( .A(n347), .B(n7719), .Z(n7718) );
  XOR U7337 ( .A(n7720), .B(n7721), .Z(n7712) );
  AND U7338 ( .A(n351), .B(n7719), .Z(n7721) );
  XNOR U7339 ( .A(n7720), .B(n7717), .Z(n7719) );
  XOR U7340 ( .A(n7722), .B(n7723), .Z(n7717) );
  AND U7341 ( .A(n354), .B(n7724), .Z(n7723) );
  XOR U7342 ( .A(p_input[466]), .B(n7722), .Z(n7724) );
  XOR U7343 ( .A(n7725), .B(n7726), .Z(n7722) );
  AND U7344 ( .A(n358), .B(n7727), .Z(n7726) );
  XOR U7345 ( .A(n7728), .B(n7729), .Z(n7720) );
  AND U7346 ( .A(n362), .B(n7727), .Z(n7729) );
  XNOR U7347 ( .A(n7728), .B(n7725), .Z(n7727) );
  XOR U7348 ( .A(n7730), .B(n7731), .Z(n7725) );
  AND U7349 ( .A(n365), .B(n7732), .Z(n7731) );
  XOR U7350 ( .A(p_input[482]), .B(n7730), .Z(n7732) );
  XOR U7351 ( .A(n7733), .B(n7734), .Z(n7730) );
  AND U7352 ( .A(n369), .B(n7735), .Z(n7734) );
  XOR U7353 ( .A(n7736), .B(n7737), .Z(n7728) );
  AND U7354 ( .A(n373), .B(n7735), .Z(n7737) );
  XNOR U7355 ( .A(n7736), .B(n7733), .Z(n7735) );
  XOR U7356 ( .A(n7738), .B(n7739), .Z(n7733) );
  AND U7357 ( .A(n376), .B(n7740), .Z(n7739) );
  XOR U7358 ( .A(p_input[498]), .B(n7738), .Z(n7740) );
  XOR U7359 ( .A(n7741), .B(n7742), .Z(n7738) );
  AND U7360 ( .A(n380), .B(n7743), .Z(n7742) );
  XOR U7361 ( .A(n7744), .B(n7745), .Z(n7736) );
  AND U7362 ( .A(n384), .B(n7743), .Z(n7745) );
  XNOR U7363 ( .A(n7744), .B(n7741), .Z(n7743) );
  XOR U7364 ( .A(n7746), .B(n7747), .Z(n7741) );
  AND U7365 ( .A(n387), .B(n7748), .Z(n7747) );
  XOR U7366 ( .A(p_input[514]), .B(n7746), .Z(n7748) );
  XOR U7367 ( .A(n7749), .B(n7750), .Z(n7746) );
  AND U7368 ( .A(n391), .B(n7751), .Z(n7750) );
  XOR U7369 ( .A(n7752), .B(n7753), .Z(n7744) );
  AND U7370 ( .A(n395), .B(n7751), .Z(n7753) );
  XNOR U7371 ( .A(n7752), .B(n7749), .Z(n7751) );
  XOR U7372 ( .A(n7754), .B(n7755), .Z(n7749) );
  AND U7373 ( .A(n398), .B(n7756), .Z(n7755) );
  XOR U7374 ( .A(p_input[530]), .B(n7754), .Z(n7756) );
  XOR U7375 ( .A(n7757), .B(n7758), .Z(n7754) );
  AND U7376 ( .A(n402), .B(n7759), .Z(n7758) );
  XOR U7377 ( .A(n7760), .B(n7761), .Z(n7752) );
  AND U7378 ( .A(n406), .B(n7759), .Z(n7761) );
  XNOR U7379 ( .A(n7760), .B(n7757), .Z(n7759) );
  XOR U7380 ( .A(n7762), .B(n7763), .Z(n7757) );
  AND U7381 ( .A(n409), .B(n7764), .Z(n7763) );
  XOR U7382 ( .A(p_input[546]), .B(n7762), .Z(n7764) );
  XOR U7383 ( .A(n7765), .B(n7766), .Z(n7762) );
  AND U7384 ( .A(n413), .B(n7767), .Z(n7766) );
  XOR U7385 ( .A(n7768), .B(n7769), .Z(n7760) );
  AND U7386 ( .A(n417), .B(n7767), .Z(n7769) );
  XNOR U7387 ( .A(n7768), .B(n7765), .Z(n7767) );
  XOR U7388 ( .A(n7770), .B(n7771), .Z(n7765) );
  AND U7389 ( .A(n420), .B(n7772), .Z(n7771) );
  XOR U7390 ( .A(p_input[562]), .B(n7770), .Z(n7772) );
  XOR U7391 ( .A(n7773), .B(n7774), .Z(n7770) );
  AND U7392 ( .A(n424), .B(n7775), .Z(n7774) );
  XOR U7393 ( .A(n7776), .B(n7777), .Z(n7768) );
  AND U7394 ( .A(n428), .B(n7775), .Z(n7777) );
  XNOR U7395 ( .A(n7776), .B(n7773), .Z(n7775) );
  XOR U7396 ( .A(n7778), .B(n7779), .Z(n7773) );
  AND U7397 ( .A(n431), .B(n7780), .Z(n7779) );
  XOR U7398 ( .A(p_input[578]), .B(n7778), .Z(n7780) );
  XOR U7399 ( .A(n7781), .B(n7782), .Z(n7778) );
  AND U7400 ( .A(n435), .B(n7783), .Z(n7782) );
  XOR U7401 ( .A(n7784), .B(n7785), .Z(n7776) );
  AND U7402 ( .A(n439), .B(n7783), .Z(n7785) );
  XNOR U7403 ( .A(n7784), .B(n7781), .Z(n7783) );
  XOR U7404 ( .A(n7786), .B(n7787), .Z(n7781) );
  AND U7405 ( .A(n442), .B(n7788), .Z(n7787) );
  XOR U7406 ( .A(p_input[594]), .B(n7786), .Z(n7788) );
  XOR U7407 ( .A(n7789), .B(n7790), .Z(n7786) );
  AND U7408 ( .A(n446), .B(n7791), .Z(n7790) );
  XOR U7409 ( .A(n7792), .B(n7793), .Z(n7784) );
  AND U7410 ( .A(n450), .B(n7791), .Z(n7793) );
  XNOR U7411 ( .A(n7792), .B(n7789), .Z(n7791) );
  XOR U7412 ( .A(n7794), .B(n7795), .Z(n7789) );
  AND U7413 ( .A(n453), .B(n7796), .Z(n7795) );
  XOR U7414 ( .A(p_input[610]), .B(n7794), .Z(n7796) );
  XOR U7415 ( .A(n7797), .B(n7798), .Z(n7794) );
  AND U7416 ( .A(n457), .B(n7799), .Z(n7798) );
  XOR U7417 ( .A(n7800), .B(n7801), .Z(n7792) );
  AND U7418 ( .A(n461), .B(n7799), .Z(n7801) );
  XNOR U7419 ( .A(n7800), .B(n7797), .Z(n7799) );
  XOR U7420 ( .A(n7802), .B(n7803), .Z(n7797) );
  AND U7421 ( .A(n464), .B(n7804), .Z(n7803) );
  XOR U7422 ( .A(p_input[626]), .B(n7802), .Z(n7804) );
  XOR U7423 ( .A(n7805), .B(n7806), .Z(n7802) );
  AND U7424 ( .A(n468), .B(n7807), .Z(n7806) );
  XOR U7425 ( .A(n7808), .B(n7809), .Z(n7800) );
  AND U7426 ( .A(n472), .B(n7807), .Z(n7809) );
  XNOR U7427 ( .A(n7808), .B(n7805), .Z(n7807) );
  XOR U7428 ( .A(n7810), .B(n7811), .Z(n7805) );
  AND U7429 ( .A(n475), .B(n7812), .Z(n7811) );
  XOR U7430 ( .A(p_input[642]), .B(n7810), .Z(n7812) );
  XOR U7431 ( .A(n7813), .B(n7814), .Z(n7810) );
  AND U7432 ( .A(n479), .B(n7815), .Z(n7814) );
  XOR U7433 ( .A(n7816), .B(n7817), .Z(n7808) );
  AND U7434 ( .A(n483), .B(n7815), .Z(n7817) );
  XNOR U7435 ( .A(n7816), .B(n7813), .Z(n7815) );
  XOR U7436 ( .A(n7818), .B(n7819), .Z(n7813) );
  AND U7437 ( .A(n486), .B(n7820), .Z(n7819) );
  XOR U7438 ( .A(p_input[658]), .B(n7818), .Z(n7820) );
  XOR U7439 ( .A(n7821), .B(n7822), .Z(n7818) );
  AND U7440 ( .A(n490), .B(n7823), .Z(n7822) );
  XOR U7441 ( .A(n7824), .B(n7825), .Z(n7816) );
  AND U7442 ( .A(n494), .B(n7823), .Z(n7825) );
  XNOR U7443 ( .A(n7824), .B(n7821), .Z(n7823) );
  XOR U7444 ( .A(n7826), .B(n7827), .Z(n7821) );
  AND U7445 ( .A(n497), .B(n7828), .Z(n7827) );
  XOR U7446 ( .A(p_input[674]), .B(n7826), .Z(n7828) );
  XOR U7447 ( .A(n7829), .B(n7830), .Z(n7826) );
  AND U7448 ( .A(n501), .B(n7831), .Z(n7830) );
  XOR U7449 ( .A(n7832), .B(n7833), .Z(n7824) );
  AND U7450 ( .A(n505), .B(n7831), .Z(n7833) );
  XNOR U7451 ( .A(n7832), .B(n7829), .Z(n7831) );
  XOR U7452 ( .A(n7834), .B(n7835), .Z(n7829) );
  AND U7453 ( .A(n508), .B(n7836), .Z(n7835) );
  XOR U7454 ( .A(p_input[690]), .B(n7834), .Z(n7836) );
  XOR U7455 ( .A(n7837), .B(n7838), .Z(n7834) );
  AND U7456 ( .A(n512), .B(n7839), .Z(n7838) );
  XOR U7457 ( .A(n7840), .B(n7841), .Z(n7832) );
  AND U7458 ( .A(n516), .B(n7839), .Z(n7841) );
  XNOR U7459 ( .A(n7840), .B(n7837), .Z(n7839) );
  XOR U7460 ( .A(n7842), .B(n7843), .Z(n7837) );
  AND U7461 ( .A(n519), .B(n7844), .Z(n7843) );
  XOR U7462 ( .A(p_input[706]), .B(n7842), .Z(n7844) );
  XOR U7463 ( .A(n7845), .B(n7846), .Z(n7842) );
  AND U7464 ( .A(n523), .B(n7847), .Z(n7846) );
  XOR U7465 ( .A(n7848), .B(n7849), .Z(n7840) );
  AND U7466 ( .A(n527), .B(n7847), .Z(n7849) );
  XNOR U7467 ( .A(n7848), .B(n7845), .Z(n7847) );
  XOR U7468 ( .A(n7850), .B(n7851), .Z(n7845) );
  AND U7469 ( .A(n530), .B(n7852), .Z(n7851) );
  XOR U7470 ( .A(p_input[722]), .B(n7850), .Z(n7852) );
  XOR U7471 ( .A(n7853), .B(n7854), .Z(n7850) );
  AND U7472 ( .A(n534), .B(n7855), .Z(n7854) );
  XOR U7473 ( .A(n7856), .B(n7857), .Z(n7848) );
  AND U7474 ( .A(n538), .B(n7855), .Z(n7857) );
  XNOR U7475 ( .A(n7856), .B(n7853), .Z(n7855) );
  XOR U7476 ( .A(n7858), .B(n7859), .Z(n7853) );
  AND U7477 ( .A(n541), .B(n7860), .Z(n7859) );
  XOR U7478 ( .A(p_input[738]), .B(n7858), .Z(n7860) );
  XOR U7479 ( .A(n7861), .B(n7862), .Z(n7858) );
  AND U7480 ( .A(n545), .B(n7863), .Z(n7862) );
  XOR U7481 ( .A(n7864), .B(n7865), .Z(n7856) );
  AND U7482 ( .A(n549), .B(n7863), .Z(n7865) );
  XNOR U7483 ( .A(n7864), .B(n7861), .Z(n7863) );
  XOR U7484 ( .A(n7866), .B(n7867), .Z(n7861) );
  AND U7485 ( .A(n552), .B(n7868), .Z(n7867) );
  XOR U7486 ( .A(p_input[754]), .B(n7866), .Z(n7868) );
  XOR U7487 ( .A(n7869), .B(n7870), .Z(n7866) );
  AND U7488 ( .A(n556), .B(n7871), .Z(n7870) );
  XOR U7489 ( .A(n7872), .B(n7873), .Z(n7864) );
  AND U7490 ( .A(n560), .B(n7871), .Z(n7873) );
  XNOR U7491 ( .A(n7872), .B(n7869), .Z(n7871) );
  XOR U7492 ( .A(n7874), .B(n7875), .Z(n7869) );
  AND U7493 ( .A(n563), .B(n7876), .Z(n7875) );
  XOR U7494 ( .A(p_input[770]), .B(n7874), .Z(n7876) );
  XOR U7495 ( .A(n7877), .B(n7878), .Z(n7874) );
  AND U7496 ( .A(n567), .B(n7879), .Z(n7878) );
  XOR U7497 ( .A(n7880), .B(n7881), .Z(n7872) );
  AND U7498 ( .A(n571), .B(n7879), .Z(n7881) );
  XNOR U7499 ( .A(n7880), .B(n7877), .Z(n7879) );
  XOR U7500 ( .A(n7882), .B(n7883), .Z(n7877) );
  AND U7501 ( .A(n574), .B(n7884), .Z(n7883) );
  XOR U7502 ( .A(p_input[786]), .B(n7882), .Z(n7884) );
  XOR U7503 ( .A(n7885), .B(n7886), .Z(n7882) );
  AND U7504 ( .A(n578), .B(n7887), .Z(n7886) );
  XOR U7505 ( .A(n7888), .B(n7889), .Z(n7880) );
  AND U7506 ( .A(n582), .B(n7887), .Z(n7889) );
  XNOR U7507 ( .A(n7888), .B(n7885), .Z(n7887) );
  XOR U7508 ( .A(n7890), .B(n7891), .Z(n7885) );
  AND U7509 ( .A(n585), .B(n7892), .Z(n7891) );
  XOR U7510 ( .A(p_input[802]), .B(n7890), .Z(n7892) );
  XOR U7511 ( .A(n7893), .B(n7894), .Z(n7890) );
  AND U7512 ( .A(n589), .B(n7895), .Z(n7894) );
  XOR U7513 ( .A(n7896), .B(n7897), .Z(n7888) );
  AND U7514 ( .A(n593), .B(n7895), .Z(n7897) );
  XNOR U7515 ( .A(n7896), .B(n7893), .Z(n7895) );
  XOR U7516 ( .A(n7898), .B(n7899), .Z(n7893) );
  AND U7517 ( .A(n596), .B(n7900), .Z(n7899) );
  XOR U7518 ( .A(p_input[818]), .B(n7898), .Z(n7900) );
  XOR U7519 ( .A(n7901), .B(n7902), .Z(n7898) );
  AND U7520 ( .A(n600), .B(n7903), .Z(n7902) );
  XOR U7521 ( .A(n7904), .B(n7905), .Z(n7896) );
  AND U7522 ( .A(n604), .B(n7903), .Z(n7905) );
  XNOR U7523 ( .A(n7904), .B(n7901), .Z(n7903) );
  XOR U7524 ( .A(n7906), .B(n7907), .Z(n7901) );
  AND U7525 ( .A(n607), .B(n7908), .Z(n7907) );
  XOR U7526 ( .A(p_input[834]), .B(n7906), .Z(n7908) );
  XOR U7527 ( .A(n7909), .B(n7910), .Z(n7906) );
  AND U7528 ( .A(n611), .B(n7911), .Z(n7910) );
  XOR U7529 ( .A(n7912), .B(n7913), .Z(n7904) );
  AND U7530 ( .A(n615), .B(n7911), .Z(n7913) );
  XNOR U7531 ( .A(n7912), .B(n7909), .Z(n7911) );
  XOR U7532 ( .A(n7914), .B(n7915), .Z(n7909) );
  AND U7533 ( .A(n618), .B(n7916), .Z(n7915) );
  XOR U7534 ( .A(p_input[850]), .B(n7914), .Z(n7916) );
  XOR U7535 ( .A(n7917), .B(n7918), .Z(n7914) );
  AND U7536 ( .A(n622), .B(n7919), .Z(n7918) );
  XOR U7537 ( .A(n7920), .B(n7921), .Z(n7912) );
  AND U7538 ( .A(n626), .B(n7919), .Z(n7921) );
  XNOR U7539 ( .A(n7920), .B(n7917), .Z(n7919) );
  XOR U7540 ( .A(n7922), .B(n7923), .Z(n7917) );
  AND U7541 ( .A(n629), .B(n7924), .Z(n7923) );
  XOR U7542 ( .A(p_input[866]), .B(n7922), .Z(n7924) );
  XOR U7543 ( .A(n7925), .B(n7926), .Z(n7922) );
  AND U7544 ( .A(n633), .B(n7927), .Z(n7926) );
  XOR U7545 ( .A(n7928), .B(n7929), .Z(n7920) );
  AND U7546 ( .A(n637), .B(n7927), .Z(n7929) );
  XNOR U7547 ( .A(n7928), .B(n7925), .Z(n7927) );
  XOR U7548 ( .A(n7930), .B(n7931), .Z(n7925) );
  AND U7549 ( .A(n640), .B(n7932), .Z(n7931) );
  XOR U7550 ( .A(p_input[882]), .B(n7930), .Z(n7932) );
  XOR U7551 ( .A(n7933), .B(n7934), .Z(n7930) );
  AND U7552 ( .A(n644), .B(n7935), .Z(n7934) );
  XOR U7553 ( .A(n7936), .B(n7937), .Z(n7928) );
  AND U7554 ( .A(n648), .B(n7935), .Z(n7937) );
  XNOR U7555 ( .A(n7936), .B(n7933), .Z(n7935) );
  XOR U7556 ( .A(n7938), .B(n7939), .Z(n7933) );
  AND U7557 ( .A(n651), .B(n7940), .Z(n7939) );
  XOR U7558 ( .A(p_input[898]), .B(n7938), .Z(n7940) );
  XOR U7559 ( .A(n7941), .B(n7942), .Z(n7938) );
  AND U7560 ( .A(n655), .B(n7943), .Z(n7942) );
  XOR U7561 ( .A(n7944), .B(n7945), .Z(n7936) );
  AND U7562 ( .A(n659), .B(n7943), .Z(n7945) );
  XNOR U7563 ( .A(n7944), .B(n7941), .Z(n7943) );
  XOR U7564 ( .A(n7946), .B(n7947), .Z(n7941) );
  AND U7565 ( .A(n662), .B(n7948), .Z(n7947) );
  XOR U7566 ( .A(p_input[914]), .B(n7946), .Z(n7948) );
  XOR U7567 ( .A(n7949), .B(n7950), .Z(n7946) );
  AND U7568 ( .A(n666), .B(n7951), .Z(n7950) );
  XOR U7569 ( .A(n7952), .B(n7953), .Z(n7944) );
  AND U7570 ( .A(n670), .B(n7951), .Z(n7953) );
  XNOR U7571 ( .A(n7952), .B(n7949), .Z(n7951) );
  XOR U7572 ( .A(n7954), .B(n7955), .Z(n7949) );
  AND U7573 ( .A(n673), .B(n7956), .Z(n7955) );
  XOR U7574 ( .A(p_input[930]), .B(n7954), .Z(n7956) );
  XOR U7575 ( .A(n7957), .B(n7958), .Z(n7954) );
  AND U7576 ( .A(n677), .B(n7959), .Z(n7958) );
  XOR U7577 ( .A(n7960), .B(n7961), .Z(n7952) );
  AND U7578 ( .A(n681), .B(n7959), .Z(n7961) );
  XNOR U7579 ( .A(n7960), .B(n7957), .Z(n7959) );
  XOR U7580 ( .A(n7962), .B(n7963), .Z(n7957) );
  AND U7581 ( .A(n684), .B(n7964), .Z(n7963) );
  XOR U7582 ( .A(p_input[946]), .B(n7962), .Z(n7964) );
  XOR U7583 ( .A(n7965), .B(n7966), .Z(n7962) );
  AND U7584 ( .A(n688), .B(n7967), .Z(n7966) );
  XOR U7585 ( .A(n7968), .B(n7969), .Z(n7960) );
  AND U7586 ( .A(n692), .B(n7967), .Z(n7969) );
  XNOR U7587 ( .A(n7968), .B(n7965), .Z(n7967) );
  XOR U7588 ( .A(n7970), .B(n7971), .Z(n7965) );
  AND U7589 ( .A(n695), .B(n7972), .Z(n7971) );
  XOR U7590 ( .A(p_input[962]), .B(n7970), .Z(n7972) );
  XOR U7591 ( .A(n7973), .B(n7974), .Z(n7970) );
  AND U7592 ( .A(n699), .B(n7975), .Z(n7974) );
  XOR U7593 ( .A(n7976), .B(n7977), .Z(n7968) );
  AND U7594 ( .A(n703), .B(n7975), .Z(n7977) );
  XNOR U7595 ( .A(n7976), .B(n7973), .Z(n7975) );
  XOR U7596 ( .A(n7978), .B(n7979), .Z(n7973) );
  AND U7597 ( .A(n706), .B(n7980), .Z(n7979) );
  XOR U7598 ( .A(p_input[978]), .B(n7978), .Z(n7980) );
  XOR U7599 ( .A(n7981), .B(n7982), .Z(n7978) );
  AND U7600 ( .A(n710), .B(n7983), .Z(n7982) );
  XOR U7601 ( .A(n7984), .B(n7985), .Z(n7976) );
  AND U7602 ( .A(n714), .B(n7983), .Z(n7985) );
  XNOR U7603 ( .A(n7984), .B(n7981), .Z(n7983) );
  XOR U7604 ( .A(n7986), .B(n7987), .Z(n7981) );
  AND U7605 ( .A(n717), .B(n7988), .Z(n7987) );
  XOR U7606 ( .A(p_input[994]), .B(n7986), .Z(n7988) );
  XOR U7607 ( .A(n7989), .B(n7990), .Z(n7986) );
  AND U7608 ( .A(n721), .B(n7991), .Z(n7990) );
  XOR U7609 ( .A(n7992), .B(n7993), .Z(n7984) );
  AND U7610 ( .A(n725), .B(n7991), .Z(n7993) );
  XNOR U7611 ( .A(n7992), .B(n7989), .Z(n7991) );
  XOR U7612 ( .A(n7994), .B(n7995), .Z(n7989) );
  AND U7613 ( .A(n728), .B(n7996), .Z(n7995) );
  XOR U7614 ( .A(p_input[1010]), .B(n7994), .Z(n7996) );
  XOR U7615 ( .A(n7997), .B(n7998), .Z(n7994) );
  AND U7616 ( .A(n732), .B(n7999), .Z(n7998) );
  XOR U7617 ( .A(n8000), .B(n8001), .Z(n7992) );
  AND U7618 ( .A(n736), .B(n7999), .Z(n8001) );
  XNOR U7619 ( .A(n8000), .B(n7997), .Z(n7999) );
  XOR U7620 ( .A(n8002), .B(n8003), .Z(n7997) );
  AND U7621 ( .A(n739), .B(n8004), .Z(n8003) );
  XOR U7622 ( .A(p_input[1026]), .B(n8002), .Z(n8004) );
  XOR U7623 ( .A(n8005), .B(n8006), .Z(n8002) );
  AND U7624 ( .A(n743), .B(n8007), .Z(n8006) );
  XOR U7625 ( .A(n8008), .B(n8009), .Z(n8000) );
  AND U7626 ( .A(n747), .B(n8007), .Z(n8009) );
  XNOR U7627 ( .A(n8008), .B(n8005), .Z(n8007) );
  XOR U7628 ( .A(n8010), .B(n8011), .Z(n8005) );
  AND U7629 ( .A(n750), .B(n8012), .Z(n8011) );
  XOR U7630 ( .A(p_input[1042]), .B(n8010), .Z(n8012) );
  XOR U7631 ( .A(n8013), .B(n8014), .Z(n8010) );
  AND U7632 ( .A(n754), .B(n8015), .Z(n8014) );
  XOR U7633 ( .A(n8016), .B(n8017), .Z(n8008) );
  AND U7634 ( .A(n758), .B(n8015), .Z(n8017) );
  XNOR U7635 ( .A(n8016), .B(n8013), .Z(n8015) );
  XOR U7636 ( .A(n8018), .B(n8019), .Z(n8013) );
  AND U7637 ( .A(n761), .B(n8020), .Z(n8019) );
  XOR U7638 ( .A(p_input[1058]), .B(n8018), .Z(n8020) );
  XOR U7639 ( .A(n8021), .B(n8022), .Z(n8018) );
  AND U7640 ( .A(n765), .B(n8023), .Z(n8022) );
  XOR U7641 ( .A(n8024), .B(n8025), .Z(n8016) );
  AND U7642 ( .A(n769), .B(n8023), .Z(n8025) );
  XNOR U7643 ( .A(n8024), .B(n8021), .Z(n8023) );
  XOR U7644 ( .A(n8026), .B(n8027), .Z(n8021) );
  AND U7645 ( .A(n772), .B(n8028), .Z(n8027) );
  XOR U7646 ( .A(p_input[1074]), .B(n8026), .Z(n8028) );
  XOR U7647 ( .A(n8029), .B(n8030), .Z(n8026) );
  AND U7648 ( .A(n776), .B(n8031), .Z(n8030) );
  XOR U7649 ( .A(n8032), .B(n8033), .Z(n8024) );
  AND U7650 ( .A(n780), .B(n8031), .Z(n8033) );
  XNOR U7651 ( .A(n8032), .B(n8029), .Z(n8031) );
  XOR U7652 ( .A(n8034), .B(n8035), .Z(n8029) );
  AND U7653 ( .A(n783), .B(n8036), .Z(n8035) );
  XOR U7654 ( .A(p_input[1090]), .B(n8034), .Z(n8036) );
  XOR U7655 ( .A(n8037), .B(n8038), .Z(n8034) );
  AND U7656 ( .A(n787), .B(n8039), .Z(n8038) );
  XOR U7657 ( .A(n8040), .B(n8041), .Z(n8032) );
  AND U7658 ( .A(n791), .B(n8039), .Z(n8041) );
  XNOR U7659 ( .A(n8040), .B(n8037), .Z(n8039) );
  XOR U7660 ( .A(n8042), .B(n8043), .Z(n8037) );
  AND U7661 ( .A(n794), .B(n8044), .Z(n8043) );
  XOR U7662 ( .A(p_input[1106]), .B(n8042), .Z(n8044) );
  XOR U7663 ( .A(n8045), .B(n8046), .Z(n8042) );
  AND U7664 ( .A(n798), .B(n8047), .Z(n8046) );
  XOR U7665 ( .A(n8048), .B(n8049), .Z(n8040) );
  AND U7666 ( .A(n802), .B(n8047), .Z(n8049) );
  XNOR U7667 ( .A(n8048), .B(n8045), .Z(n8047) );
  XOR U7668 ( .A(n8050), .B(n8051), .Z(n8045) );
  AND U7669 ( .A(n805), .B(n8052), .Z(n8051) );
  XOR U7670 ( .A(p_input[1122]), .B(n8050), .Z(n8052) );
  XOR U7671 ( .A(n8053), .B(n8054), .Z(n8050) );
  AND U7672 ( .A(n809), .B(n8055), .Z(n8054) );
  XOR U7673 ( .A(n8056), .B(n8057), .Z(n8048) );
  AND U7674 ( .A(n813), .B(n8055), .Z(n8057) );
  XNOR U7675 ( .A(n8056), .B(n8053), .Z(n8055) );
  XOR U7676 ( .A(n8058), .B(n8059), .Z(n8053) );
  AND U7677 ( .A(n816), .B(n8060), .Z(n8059) );
  XOR U7678 ( .A(p_input[1138]), .B(n8058), .Z(n8060) );
  XOR U7679 ( .A(n8061), .B(n8062), .Z(n8058) );
  AND U7680 ( .A(n820), .B(n8063), .Z(n8062) );
  XOR U7681 ( .A(n8064), .B(n8065), .Z(n8056) );
  AND U7682 ( .A(n824), .B(n8063), .Z(n8065) );
  XNOR U7683 ( .A(n8064), .B(n8061), .Z(n8063) );
  XOR U7684 ( .A(n8066), .B(n8067), .Z(n8061) );
  AND U7685 ( .A(n827), .B(n8068), .Z(n8067) );
  XOR U7686 ( .A(p_input[1154]), .B(n8066), .Z(n8068) );
  XOR U7687 ( .A(n8069), .B(n8070), .Z(n8066) );
  AND U7688 ( .A(n831), .B(n8071), .Z(n8070) );
  XOR U7689 ( .A(n8072), .B(n8073), .Z(n8064) );
  AND U7690 ( .A(n835), .B(n8071), .Z(n8073) );
  XNOR U7691 ( .A(n8072), .B(n8069), .Z(n8071) );
  XOR U7692 ( .A(n8074), .B(n8075), .Z(n8069) );
  AND U7693 ( .A(n838), .B(n8076), .Z(n8075) );
  XOR U7694 ( .A(p_input[1170]), .B(n8074), .Z(n8076) );
  XOR U7695 ( .A(n8077), .B(n8078), .Z(n8074) );
  AND U7696 ( .A(n842), .B(n8079), .Z(n8078) );
  XOR U7697 ( .A(n8080), .B(n8081), .Z(n8072) );
  AND U7698 ( .A(n846), .B(n8079), .Z(n8081) );
  XNOR U7699 ( .A(n8080), .B(n8077), .Z(n8079) );
  XOR U7700 ( .A(n8082), .B(n8083), .Z(n8077) );
  AND U7701 ( .A(n849), .B(n8084), .Z(n8083) );
  XOR U7702 ( .A(p_input[1186]), .B(n8082), .Z(n8084) );
  XOR U7703 ( .A(n8085), .B(n8086), .Z(n8082) );
  AND U7704 ( .A(n853), .B(n8087), .Z(n8086) );
  XOR U7705 ( .A(n8088), .B(n8089), .Z(n8080) );
  AND U7706 ( .A(n857), .B(n8087), .Z(n8089) );
  XNOR U7707 ( .A(n8088), .B(n8085), .Z(n8087) );
  XOR U7708 ( .A(n8090), .B(n8091), .Z(n8085) );
  AND U7709 ( .A(n860), .B(n8092), .Z(n8091) );
  XOR U7710 ( .A(p_input[1202]), .B(n8090), .Z(n8092) );
  XOR U7711 ( .A(n8093), .B(n8094), .Z(n8090) );
  AND U7712 ( .A(n864), .B(n8095), .Z(n8094) );
  XOR U7713 ( .A(n8096), .B(n8097), .Z(n8088) );
  AND U7714 ( .A(n868), .B(n8095), .Z(n8097) );
  XNOR U7715 ( .A(n8096), .B(n8093), .Z(n8095) );
  XOR U7716 ( .A(n8098), .B(n8099), .Z(n8093) );
  AND U7717 ( .A(n871), .B(n8100), .Z(n8099) );
  XOR U7718 ( .A(p_input[1218]), .B(n8098), .Z(n8100) );
  XOR U7719 ( .A(n8101), .B(n8102), .Z(n8098) );
  AND U7720 ( .A(n875), .B(n8103), .Z(n8102) );
  XOR U7721 ( .A(n8104), .B(n8105), .Z(n8096) );
  AND U7722 ( .A(n879), .B(n8103), .Z(n8105) );
  XNOR U7723 ( .A(n8104), .B(n8101), .Z(n8103) );
  XOR U7724 ( .A(n8106), .B(n8107), .Z(n8101) );
  AND U7725 ( .A(n882), .B(n8108), .Z(n8107) );
  XOR U7726 ( .A(p_input[1234]), .B(n8106), .Z(n8108) );
  XOR U7727 ( .A(n8109), .B(n8110), .Z(n8106) );
  AND U7728 ( .A(n886), .B(n8111), .Z(n8110) );
  XOR U7729 ( .A(n8112), .B(n8113), .Z(n8104) );
  AND U7730 ( .A(n890), .B(n8111), .Z(n8113) );
  XNOR U7731 ( .A(n8112), .B(n8109), .Z(n8111) );
  XOR U7732 ( .A(n8114), .B(n8115), .Z(n8109) );
  AND U7733 ( .A(n893), .B(n8116), .Z(n8115) );
  XOR U7734 ( .A(p_input[1250]), .B(n8114), .Z(n8116) );
  XOR U7735 ( .A(n8117), .B(n8118), .Z(n8114) );
  AND U7736 ( .A(n897), .B(n8119), .Z(n8118) );
  XOR U7737 ( .A(n8120), .B(n8121), .Z(n8112) );
  AND U7738 ( .A(n901), .B(n8119), .Z(n8121) );
  XNOR U7739 ( .A(n8120), .B(n8117), .Z(n8119) );
  XOR U7740 ( .A(n8122), .B(n8123), .Z(n8117) );
  AND U7741 ( .A(n904), .B(n8124), .Z(n8123) );
  XOR U7742 ( .A(p_input[1266]), .B(n8122), .Z(n8124) );
  XOR U7743 ( .A(n8125), .B(n8126), .Z(n8122) );
  AND U7744 ( .A(n908), .B(n8127), .Z(n8126) );
  XOR U7745 ( .A(n8128), .B(n8129), .Z(n8120) );
  AND U7746 ( .A(n912), .B(n8127), .Z(n8129) );
  XNOR U7747 ( .A(n8128), .B(n8125), .Z(n8127) );
  XOR U7748 ( .A(n8130), .B(n8131), .Z(n8125) );
  AND U7749 ( .A(n915), .B(n8132), .Z(n8131) );
  XOR U7750 ( .A(p_input[1282]), .B(n8130), .Z(n8132) );
  XOR U7751 ( .A(n8133), .B(n8134), .Z(n8130) );
  AND U7752 ( .A(n919), .B(n8135), .Z(n8134) );
  XOR U7753 ( .A(n8136), .B(n8137), .Z(n8128) );
  AND U7754 ( .A(n923), .B(n8135), .Z(n8137) );
  XNOR U7755 ( .A(n8136), .B(n8133), .Z(n8135) );
  XOR U7756 ( .A(n8138), .B(n8139), .Z(n8133) );
  AND U7757 ( .A(n926), .B(n8140), .Z(n8139) );
  XOR U7758 ( .A(p_input[1298]), .B(n8138), .Z(n8140) );
  XOR U7759 ( .A(n8141), .B(n8142), .Z(n8138) );
  AND U7760 ( .A(n930), .B(n8143), .Z(n8142) );
  XOR U7761 ( .A(n8144), .B(n8145), .Z(n8136) );
  AND U7762 ( .A(n934), .B(n8143), .Z(n8145) );
  XNOR U7763 ( .A(n8144), .B(n8141), .Z(n8143) );
  XOR U7764 ( .A(n8146), .B(n8147), .Z(n8141) );
  AND U7765 ( .A(n937), .B(n8148), .Z(n8147) );
  XOR U7766 ( .A(p_input[1314]), .B(n8146), .Z(n8148) );
  XOR U7767 ( .A(n8149), .B(n8150), .Z(n8146) );
  AND U7768 ( .A(n941), .B(n8151), .Z(n8150) );
  XOR U7769 ( .A(n8152), .B(n8153), .Z(n8144) );
  AND U7770 ( .A(n945), .B(n8151), .Z(n8153) );
  XNOR U7771 ( .A(n8152), .B(n8149), .Z(n8151) );
  XOR U7772 ( .A(n8154), .B(n8155), .Z(n8149) );
  AND U7773 ( .A(n948), .B(n8156), .Z(n8155) );
  XOR U7774 ( .A(p_input[1330]), .B(n8154), .Z(n8156) );
  XOR U7775 ( .A(n8157), .B(n8158), .Z(n8154) );
  AND U7776 ( .A(n952), .B(n8159), .Z(n8158) );
  XOR U7777 ( .A(n8160), .B(n8161), .Z(n8152) );
  AND U7778 ( .A(n956), .B(n8159), .Z(n8161) );
  XNOR U7779 ( .A(n8160), .B(n8157), .Z(n8159) );
  XOR U7780 ( .A(n8162), .B(n8163), .Z(n8157) );
  AND U7781 ( .A(n959), .B(n8164), .Z(n8163) );
  XOR U7782 ( .A(p_input[1346]), .B(n8162), .Z(n8164) );
  XOR U7783 ( .A(n8165), .B(n8166), .Z(n8162) );
  AND U7784 ( .A(n963), .B(n8167), .Z(n8166) );
  XOR U7785 ( .A(n8168), .B(n8169), .Z(n8160) );
  AND U7786 ( .A(n967), .B(n8167), .Z(n8169) );
  XNOR U7787 ( .A(n8168), .B(n8165), .Z(n8167) );
  XOR U7788 ( .A(n8170), .B(n8171), .Z(n8165) );
  AND U7789 ( .A(n970), .B(n8172), .Z(n8171) );
  XOR U7790 ( .A(p_input[1362]), .B(n8170), .Z(n8172) );
  XOR U7791 ( .A(n8173), .B(n8174), .Z(n8170) );
  AND U7792 ( .A(n974), .B(n8175), .Z(n8174) );
  XOR U7793 ( .A(n8176), .B(n8177), .Z(n8168) );
  AND U7794 ( .A(n978), .B(n8175), .Z(n8177) );
  XNOR U7795 ( .A(n8176), .B(n8173), .Z(n8175) );
  XOR U7796 ( .A(n8178), .B(n8179), .Z(n8173) );
  AND U7797 ( .A(n981), .B(n8180), .Z(n8179) );
  XOR U7798 ( .A(p_input[1378]), .B(n8178), .Z(n8180) );
  XOR U7799 ( .A(n8181), .B(n8182), .Z(n8178) );
  AND U7800 ( .A(n985), .B(n8183), .Z(n8182) );
  XOR U7801 ( .A(n8184), .B(n8185), .Z(n8176) );
  AND U7802 ( .A(n989), .B(n8183), .Z(n8185) );
  XNOR U7803 ( .A(n8184), .B(n8181), .Z(n8183) );
  XOR U7804 ( .A(n8186), .B(n8187), .Z(n8181) );
  AND U7805 ( .A(n992), .B(n8188), .Z(n8187) );
  XOR U7806 ( .A(p_input[1394]), .B(n8186), .Z(n8188) );
  XOR U7807 ( .A(n8189), .B(n8190), .Z(n8186) );
  AND U7808 ( .A(n996), .B(n8191), .Z(n8190) );
  XOR U7809 ( .A(n8192), .B(n8193), .Z(n8184) );
  AND U7810 ( .A(n1000), .B(n8191), .Z(n8193) );
  XNOR U7811 ( .A(n8192), .B(n8189), .Z(n8191) );
  XOR U7812 ( .A(n8194), .B(n8195), .Z(n8189) );
  AND U7813 ( .A(n1003), .B(n8196), .Z(n8195) );
  XOR U7814 ( .A(p_input[1410]), .B(n8194), .Z(n8196) );
  XOR U7815 ( .A(n8197), .B(n8198), .Z(n8194) );
  AND U7816 ( .A(n1007), .B(n8199), .Z(n8198) );
  XOR U7817 ( .A(n8200), .B(n8201), .Z(n8192) );
  AND U7818 ( .A(n1011), .B(n8199), .Z(n8201) );
  XNOR U7819 ( .A(n8200), .B(n8197), .Z(n8199) );
  XOR U7820 ( .A(n8202), .B(n8203), .Z(n8197) );
  AND U7821 ( .A(n1014), .B(n8204), .Z(n8203) );
  XOR U7822 ( .A(p_input[1426]), .B(n8202), .Z(n8204) );
  XOR U7823 ( .A(n8205), .B(n8206), .Z(n8202) );
  AND U7824 ( .A(n1018), .B(n8207), .Z(n8206) );
  XOR U7825 ( .A(n8208), .B(n8209), .Z(n8200) );
  AND U7826 ( .A(n1022), .B(n8207), .Z(n8209) );
  XNOR U7827 ( .A(n8208), .B(n8205), .Z(n8207) );
  XOR U7828 ( .A(n8210), .B(n8211), .Z(n8205) );
  AND U7829 ( .A(n1025), .B(n8212), .Z(n8211) );
  XOR U7830 ( .A(p_input[1442]), .B(n8210), .Z(n8212) );
  XOR U7831 ( .A(n8213), .B(n8214), .Z(n8210) );
  AND U7832 ( .A(n1029), .B(n8215), .Z(n8214) );
  XOR U7833 ( .A(n8216), .B(n8217), .Z(n8208) );
  AND U7834 ( .A(n1033), .B(n8215), .Z(n8217) );
  XNOR U7835 ( .A(n8216), .B(n8213), .Z(n8215) );
  XOR U7836 ( .A(n8218), .B(n8219), .Z(n8213) );
  AND U7837 ( .A(n1036), .B(n8220), .Z(n8219) );
  XOR U7838 ( .A(p_input[1458]), .B(n8218), .Z(n8220) );
  XOR U7839 ( .A(n8221), .B(n8222), .Z(n8218) );
  AND U7840 ( .A(n1040), .B(n8223), .Z(n8222) );
  XOR U7841 ( .A(n8224), .B(n8225), .Z(n8216) );
  AND U7842 ( .A(n1044), .B(n8223), .Z(n8225) );
  XNOR U7843 ( .A(n8224), .B(n8221), .Z(n8223) );
  XOR U7844 ( .A(n8226), .B(n8227), .Z(n8221) );
  AND U7845 ( .A(n1047), .B(n8228), .Z(n8227) );
  XOR U7846 ( .A(p_input[1474]), .B(n8226), .Z(n8228) );
  XOR U7847 ( .A(n8229), .B(n8230), .Z(n8226) );
  AND U7848 ( .A(n1051), .B(n8231), .Z(n8230) );
  XOR U7849 ( .A(n8232), .B(n8233), .Z(n8224) );
  AND U7850 ( .A(n1055), .B(n8231), .Z(n8233) );
  XNOR U7851 ( .A(n8232), .B(n8229), .Z(n8231) );
  XOR U7852 ( .A(n8234), .B(n8235), .Z(n8229) );
  AND U7853 ( .A(n1058), .B(n8236), .Z(n8235) );
  XOR U7854 ( .A(p_input[1490]), .B(n8234), .Z(n8236) );
  XOR U7855 ( .A(n8237), .B(n8238), .Z(n8234) );
  AND U7856 ( .A(n1062), .B(n8239), .Z(n8238) );
  XOR U7857 ( .A(n8240), .B(n8241), .Z(n8232) );
  AND U7858 ( .A(n1066), .B(n8239), .Z(n8241) );
  XNOR U7859 ( .A(n8240), .B(n8237), .Z(n8239) );
  XOR U7860 ( .A(n8242), .B(n8243), .Z(n8237) );
  AND U7861 ( .A(n1069), .B(n8244), .Z(n8243) );
  XOR U7862 ( .A(p_input[1506]), .B(n8242), .Z(n8244) );
  XOR U7863 ( .A(n8245), .B(n8246), .Z(n8242) );
  AND U7864 ( .A(n1073), .B(n8247), .Z(n8246) );
  XOR U7865 ( .A(n8248), .B(n8249), .Z(n8240) );
  AND U7866 ( .A(n1077), .B(n8247), .Z(n8249) );
  XNOR U7867 ( .A(n8248), .B(n8245), .Z(n8247) );
  XOR U7868 ( .A(n8250), .B(n8251), .Z(n8245) );
  AND U7869 ( .A(n1080), .B(n8252), .Z(n8251) );
  XOR U7870 ( .A(p_input[1522]), .B(n8250), .Z(n8252) );
  XOR U7871 ( .A(n8253), .B(n8254), .Z(n8250) );
  AND U7872 ( .A(n1084), .B(n8255), .Z(n8254) );
  XOR U7873 ( .A(n8256), .B(n8257), .Z(n8248) );
  AND U7874 ( .A(n1088), .B(n8255), .Z(n8257) );
  XNOR U7875 ( .A(n8256), .B(n8253), .Z(n8255) );
  XOR U7876 ( .A(n8258), .B(n8259), .Z(n8253) );
  AND U7877 ( .A(n1091), .B(n8260), .Z(n8259) );
  XOR U7878 ( .A(p_input[1538]), .B(n8258), .Z(n8260) );
  XOR U7879 ( .A(n8261), .B(n8262), .Z(n8258) );
  AND U7880 ( .A(n1095), .B(n8263), .Z(n8262) );
  XOR U7881 ( .A(n8264), .B(n8265), .Z(n8256) );
  AND U7882 ( .A(n1099), .B(n8263), .Z(n8265) );
  XNOR U7883 ( .A(n8264), .B(n8261), .Z(n8263) );
  XOR U7884 ( .A(n8266), .B(n8267), .Z(n8261) );
  AND U7885 ( .A(n1102), .B(n8268), .Z(n8267) );
  XOR U7886 ( .A(p_input[1554]), .B(n8266), .Z(n8268) );
  XOR U7887 ( .A(n8269), .B(n8270), .Z(n8266) );
  AND U7888 ( .A(n1106), .B(n8271), .Z(n8270) );
  XOR U7889 ( .A(n8272), .B(n8273), .Z(n8264) );
  AND U7890 ( .A(n1110), .B(n8271), .Z(n8273) );
  XNOR U7891 ( .A(n8272), .B(n8269), .Z(n8271) );
  XOR U7892 ( .A(n8274), .B(n8275), .Z(n8269) );
  AND U7893 ( .A(n1113), .B(n8276), .Z(n8275) );
  XOR U7894 ( .A(p_input[1570]), .B(n8274), .Z(n8276) );
  XOR U7895 ( .A(n8277), .B(n8278), .Z(n8274) );
  AND U7896 ( .A(n1117), .B(n8279), .Z(n8278) );
  XOR U7897 ( .A(n8280), .B(n8281), .Z(n8272) );
  AND U7898 ( .A(n1121), .B(n8279), .Z(n8281) );
  XNOR U7899 ( .A(n8280), .B(n8277), .Z(n8279) );
  XOR U7900 ( .A(n8282), .B(n8283), .Z(n8277) );
  AND U7901 ( .A(n1124), .B(n8284), .Z(n8283) );
  XOR U7902 ( .A(p_input[1586]), .B(n8282), .Z(n8284) );
  XOR U7903 ( .A(n8285), .B(n8286), .Z(n8282) );
  AND U7904 ( .A(n1128), .B(n8287), .Z(n8286) );
  XOR U7905 ( .A(n8288), .B(n8289), .Z(n8280) );
  AND U7906 ( .A(n1132), .B(n8287), .Z(n8289) );
  XNOR U7907 ( .A(n8288), .B(n8285), .Z(n8287) );
  XOR U7908 ( .A(n8290), .B(n8291), .Z(n8285) );
  AND U7909 ( .A(n1135), .B(n8292), .Z(n8291) );
  XOR U7910 ( .A(p_input[1602]), .B(n8290), .Z(n8292) );
  XOR U7911 ( .A(n8293), .B(n8294), .Z(n8290) );
  AND U7912 ( .A(n1139), .B(n8295), .Z(n8294) );
  XOR U7913 ( .A(n8296), .B(n8297), .Z(n8288) );
  AND U7914 ( .A(n1143), .B(n8295), .Z(n8297) );
  XNOR U7915 ( .A(n8296), .B(n8293), .Z(n8295) );
  XOR U7916 ( .A(n8298), .B(n8299), .Z(n8293) );
  AND U7917 ( .A(n1146), .B(n8300), .Z(n8299) );
  XOR U7918 ( .A(p_input[1618]), .B(n8298), .Z(n8300) );
  XOR U7919 ( .A(n8301), .B(n8302), .Z(n8298) );
  AND U7920 ( .A(n1150), .B(n8303), .Z(n8302) );
  XOR U7921 ( .A(n8304), .B(n8305), .Z(n8296) );
  AND U7922 ( .A(n1154), .B(n8303), .Z(n8305) );
  XNOR U7923 ( .A(n8304), .B(n8301), .Z(n8303) );
  XOR U7924 ( .A(n8306), .B(n8307), .Z(n8301) );
  AND U7925 ( .A(n1157), .B(n8308), .Z(n8307) );
  XOR U7926 ( .A(p_input[1634]), .B(n8306), .Z(n8308) );
  XOR U7927 ( .A(n8309), .B(n8310), .Z(n8306) );
  AND U7928 ( .A(n1161), .B(n8311), .Z(n8310) );
  XOR U7929 ( .A(n8312), .B(n8313), .Z(n8304) );
  AND U7930 ( .A(n1165), .B(n8311), .Z(n8313) );
  XNOR U7931 ( .A(n8312), .B(n8309), .Z(n8311) );
  XOR U7932 ( .A(n8314), .B(n8315), .Z(n8309) );
  AND U7933 ( .A(n1168), .B(n8316), .Z(n8315) );
  XOR U7934 ( .A(p_input[1650]), .B(n8314), .Z(n8316) );
  XOR U7935 ( .A(n8317), .B(n8318), .Z(n8314) );
  AND U7936 ( .A(n1172), .B(n8319), .Z(n8318) );
  XOR U7937 ( .A(n8320), .B(n8321), .Z(n8312) );
  AND U7938 ( .A(n1176), .B(n8319), .Z(n8321) );
  XNOR U7939 ( .A(n8320), .B(n8317), .Z(n8319) );
  XOR U7940 ( .A(n8322), .B(n8323), .Z(n8317) );
  AND U7941 ( .A(n1179), .B(n8324), .Z(n8323) );
  XOR U7942 ( .A(p_input[1666]), .B(n8322), .Z(n8324) );
  XOR U7943 ( .A(n8325), .B(n8326), .Z(n8322) );
  AND U7944 ( .A(n1183), .B(n8327), .Z(n8326) );
  XOR U7945 ( .A(n8328), .B(n8329), .Z(n8320) );
  AND U7946 ( .A(n1187), .B(n8327), .Z(n8329) );
  XNOR U7947 ( .A(n8328), .B(n8325), .Z(n8327) );
  XOR U7948 ( .A(n8330), .B(n8331), .Z(n8325) );
  AND U7949 ( .A(n1190), .B(n8332), .Z(n8331) );
  XOR U7950 ( .A(p_input[1682]), .B(n8330), .Z(n8332) );
  XOR U7951 ( .A(n8333), .B(n8334), .Z(n8330) );
  AND U7952 ( .A(n1194), .B(n8335), .Z(n8334) );
  XOR U7953 ( .A(n8336), .B(n8337), .Z(n8328) );
  AND U7954 ( .A(n1198), .B(n8335), .Z(n8337) );
  XNOR U7955 ( .A(n8336), .B(n8333), .Z(n8335) );
  XOR U7956 ( .A(n8338), .B(n8339), .Z(n8333) );
  AND U7957 ( .A(n1201), .B(n8340), .Z(n8339) );
  XOR U7958 ( .A(p_input[1698]), .B(n8338), .Z(n8340) );
  XOR U7959 ( .A(n8341), .B(n8342), .Z(n8338) );
  AND U7960 ( .A(n1205), .B(n8343), .Z(n8342) );
  XOR U7961 ( .A(n8344), .B(n8345), .Z(n8336) );
  AND U7962 ( .A(n1209), .B(n8343), .Z(n8345) );
  XNOR U7963 ( .A(n8344), .B(n8341), .Z(n8343) );
  XOR U7964 ( .A(n8346), .B(n8347), .Z(n8341) );
  AND U7965 ( .A(n1212), .B(n8348), .Z(n8347) );
  XOR U7966 ( .A(p_input[1714]), .B(n8346), .Z(n8348) );
  XOR U7967 ( .A(n8349), .B(n8350), .Z(n8346) );
  AND U7968 ( .A(n1216), .B(n8351), .Z(n8350) );
  XOR U7969 ( .A(n8352), .B(n8353), .Z(n8344) );
  AND U7970 ( .A(n1220), .B(n8351), .Z(n8353) );
  XNOR U7971 ( .A(n8352), .B(n8349), .Z(n8351) );
  XOR U7972 ( .A(n8354), .B(n8355), .Z(n8349) );
  AND U7973 ( .A(n1223), .B(n8356), .Z(n8355) );
  XOR U7974 ( .A(p_input[1730]), .B(n8354), .Z(n8356) );
  XOR U7975 ( .A(n8357), .B(n8358), .Z(n8354) );
  AND U7976 ( .A(n1227), .B(n8359), .Z(n8358) );
  XOR U7977 ( .A(n8360), .B(n8361), .Z(n8352) );
  AND U7978 ( .A(n1231), .B(n8359), .Z(n8361) );
  XNOR U7979 ( .A(n8360), .B(n8357), .Z(n8359) );
  XOR U7980 ( .A(n8362), .B(n8363), .Z(n8357) );
  AND U7981 ( .A(n1234), .B(n8364), .Z(n8363) );
  XOR U7982 ( .A(p_input[1746]), .B(n8362), .Z(n8364) );
  XOR U7983 ( .A(n8365), .B(n8366), .Z(n8362) );
  AND U7984 ( .A(n1238), .B(n8367), .Z(n8366) );
  XOR U7985 ( .A(n8368), .B(n8369), .Z(n8360) );
  AND U7986 ( .A(n1242), .B(n8367), .Z(n8369) );
  XNOR U7987 ( .A(n8368), .B(n8365), .Z(n8367) );
  XOR U7988 ( .A(n8370), .B(n8371), .Z(n8365) );
  AND U7989 ( .A(n1245), .B(n8372), .Z(n8371) );
  XOR U7990 ( .A(p_input[1762]), .B(n8370), .Z(n8372) );
  XOR U7991 ( .A(n8373), .B(n8374), .Z(n8370) );
  AND U7992 ( .A(n1249), .B(n8375), .Z(n8374) );
  XOR U7993 ( .A(n8376), .B(n8377), .Z(n8368) );
  AND U7994 ( .A(n1253), .B(n8375), .Z(n8377) );
  XNOR U7995 ( .A(n8376), .B(n8373), .Z(n8375) );
  XOR U7996 ( .A(n8378), .B(n8379), .Z(n8373) );
  AND U7997 ( .A(n1256), .B(n8380), .Z(n8379) );
  XOR U7998 ( .A(p_input[1778]), .B(n8378), .Z(n8380) );
  XOR U7999 ( .A(n8381), .B(n8382), .Z(n8378) );
  AND U8000 ( .A(n1260), .B(n8383), .Z(n8382) );
  XOR U8001 ( .A(n8384), .B(n8385), .Z(n8376) );
  AND U8002 ( .A(n1264), .B(n8383), .Z(n8385) );
  XNOR U8003 ( .A(n8384), .B(n8381), .Z(n8383) );
  XOR U8004 ( .A(n8386), .B(n8387), .Z(n8381) );
  AND U8005 ( .A(n1267), .B(n8388), .Z(n8387) );
  XOR U8006 ( .A(p_input[1794]), .B(n8386), .Z(n8388) );
  XOR U8007 ( .A(n8389), .B(n8390), .Z(n8386) );
  AND U8008 ( .A(n1271), .B(n8391), .Z(n8390) );
  XOR U8009 ( .A(n8392), .B(n8393), .Z(n8384) );
  AND U8010 ( .A(n1275), .B(n8391), .Z(n8393) );
  XNOR U8011 ( .A(n8392), .B(n8389), .Z(n8391) );
  XOR U8012 ( .A(n8394), .B(n8395), .Z(n8389) );
  AND U8013 ( .A(n1278), .B(n8396), .Z(n8395) );
  XOR U8014 ( .A(p_input[1810]), .B(n8394), .Z(n8396) );
  XOR U8015 ( .A(n8397), .B(n8398), .Z(n8394) );
  AND U8016 ( .A(n1282), .B(n8399), .Z(n8398) );
  XOR U8017 ( .A(n8400), .B(n8401), .Z(n8392) );
  AND U8018 ( .A(n1286), .B(n8399), .Z(n8401) );
  XNOR U8019 ( .A(n8400), .B(n8397), .Z(n8399) );
  XOR U8020 ( .A(n8402), .B(n8403), .Z(n8397) );
  AND U8021 ( .A(n1289), .B(n8404), .Z(n8403) );
  XOR U8022 ( .A(p_input[1826]), .B(n8402), .Z(n8404) );
  XOR U8023 ( .A(n8405), .B(n8406), .Z(n8402) );
  AND U8024 ( .A(n1293), .B(n8407), .Z(n8406) );
  XOR U8025 ( .A(n8408), .B(n8409), .Z(n8400) );
  AND U8026 ( .A(n1297), .B(n8407), .Z(n8409) );
  XNOR U8027 ( .A(n8408), .B(n8405), .Z(n8407) );
  XOR U8028 ( .A(n8410), .B(n8411), .Z(n8405) );
  AND U8029 ( .A(n1300), .B(n8412), .Z(n8411) );
  XOR U8030 ( .A(p_input[1842]), .B(n8410), .Z(n8412) );
  XOR U8031 ( .A(n8413), .B(n8414), .Z(n8410) );
  AND U8032 ( .A(n1304), .B(n8415), .Z(n8414) );
  XOR U8033 ( .A(n8416), .B(n8417), .Z(n8408) );
  AND U8034 ( .A(n1308), .B(n8415), .Z(n8417) );
  XNOR U8035 ( .A(n8416), .B(n8413), .Z(n8415) );
  XOR U8036 ( .A(n8418), .B(n8419), .Z(n8413) );
  AND U8037 ( .A(n1311), .B(n8420), .Z(n8419) );
  XOR U8038 ( .A(p_input[1858]), .B(n8418), .Z(n8420) );
  XOR U8039 ( .A(n8421), .B(n8422), .Z(n8418) );
  AND U8040 ( .A(n1315), .B(n8423), .Z(n8422) );
  XOR U8041 ( .A(n8424), .B(n8425), .Z(n8416) );
  AND U8042 ( .A(n1319), .B(n8423), .Z(n8425) );
  XNOR U8043 ( .A(n8424), .B(n8421), .Z(n8423) );
  XOR U8044 ( .A(n8426), .B(n8427), .Z(n8421) );
  AND U8045 ( .A(n1322), .B(n8428), .Z(n8427) );
  XOR U8046 ( .A(p_input[1874]), .B(n8426), .Z(n8428) );
  XOR U8047 ( .A(n8429), .B(n8430), .Z(n8426) );
  AND U8048 ( .A(n1326), .B(n8431), .Z(n8430) );
  XOR U8049 ( .A(n8432), .B(n8433), .Z(n8424) );
  AND U8050 ( .A(n1330), .B(n8431), .Z(n8433) );
  XNOR U8051 ( .A(n8432), .B(n8429), .Z(n8431) );
  XOR U8052 ( .A(n8434), .B(n8435), .Z(n8429) );
  AND U8053 ( .A(n1333), .B(n8436), .Z(n8435) );
  XOR U8054 ( .A(p_input[1890]), .B(n8434), .Z(n8436) );
  XOR U8055 ( .A(n8437), .B(n8438), .Z(n8434) );
  AND U8056 ( .A(n1337), .B(n8439), .Z(n8438) );
  XOR U8057 ( .A(n8440), .B(n8441), .Z(n8432) );
  AND U8058 ( .A(n1341), .B(n8439), .Z(n8441) );
  XNOR U8059 ( .A(n8440), .B(n8437), .Z(n8439) );
  XOR U8060 ( .A(n8442), .B(n8443), .Z(n8437) );
  AND U8061 ( .A(n1344), .B(n8444), .Z(n8443) );
  XOR U8062 ( .A(p_input[1906]), .B(n8442), .Z(n8444) );
  XOR U8063 ( .A(n8445), .B(n8446), .Z(n8442) );
  AND U8064 ( .A(n1348), .B(n8447), .Z(n8446) );
  XOR U8065 ( .A(n8448), .B(n8449), .Z(n8440) );
  AND U8066 ( .A(n1352), .B(n8447), .Z(n8449) );
  XNOR U8067 ( .A(n8448), .B(n8445), .Z(n8447) );
  XOR U8068 ( .A(n8450), .B(n8451), .Z(n8445) );
  AND U8069 ( .A(n1355), .B(n8452), .Z(n8451) );
  XOR U8070 ( .A(p_input[1922]), .B(n8450), .Z(n8452) );
  XOR U8071 ( .A(n8453), .B(n8454), .Z(n8450) );
  AND U8072 ( .A(n1359), .B(n8455), .Z(n8454) );
  XOR U8073 ( .A(n8456), .B(n8457), .Z(n8448) );
  AND U8074 ( .A(n1363), .B(n8455), .Z(n8457) );
  XNOR U8075 ( .A(n8456), .B(n8453), .Z(n8455) );
  XOR U8076 ( .A(n8458), .B(n8459), .Z(n8453) );
  AND U8077 ( .A(n1366), .B(n8460), .Z(n8459) );
  XOR U8078 ( .A(p_input[1938]), .B(n8458), .Z(n8460) );
  XOR U8079 ( .A(n8461), .B(n8462), .Z(n8458) );
  AND U8080 ( .A(n1370), .B(n8463), .Z(n8462) );
  XOR U8081 ( .A(n8464), .B(n8465), .Z(n8456) );
  AND U8082 ( .A(n1374), .B(n8463), .Z(n8465) );
  XNOR U8083 ( .A(n8464), .B(n8461), .Z(n8463) );
  XOR U8084 ( .A(n8466), .B(n8467), .Z(n8461) );
  AND U8085 ( .A(n1377), .B(n8468), .Z(n8467) );
  XOR U8086 ( .A(p_input[1954]), .B(n8466), .Z(n8468) );
  XOR U8087 ( .A(n8469), .B(n8470), .Z(n8466) );
  AND U8088 ( .A(n1381), .B(n8471), .Z(n8470) );
  XOR U8089 ( .A(n8472), .B(n8473), .Z(n8464) );
  AND U8090 ( .A(n1385), .B(n8471), .Z(n8473) );
  XNOR U8091 ( .A(n8472), .B(n8469), .Z(n8471) );
  XOR U8092 ( .A(n8474), .B(n8475), .Z(n8469) );
  AND U8093 ( .A(n1388), .B(n8476), .Z(n8475) );
  XOR U8094 ( .A(p_input[1970]), .B(n8474), .Z(n8476) );
  XOR U8095 ( .A(n8477), .B(n8478), .Z(n8474) );
  AND U8096 ( .A(n1392), .B(n8479), .Z(n8478) );
  XOR U8097 ( .A(n8480), .B(n8481), .Z(n8472) );
  AND U8098 ( .A(n1396), .B(n8479), .Z(n8481) );
  XNOR U8099 ( .A(n8480), .B(n8477), .Z(n8479) );
  XOR U8100 ( .A(n8482), .B(n8483), .Z(n8477) );
  AND U8101 ( .A(n1399), .B(n8484), .Z(n8483) );
  XOR U8102 ( .A(p_input[1986]), .B(n8482), .Z(n8484) );
  XOR U8103 ( .A(n8485), .B(n8486), .Z(n8482) );
  AND U8104 ( .A(n1403), .B(n8487), .Z(n8486) );
  XOR U8105 ( .A(n8488), .B(n8489), .Z(n8480) );
  AND U8106 ( .A(n1407), .B(n8487), .Z(n8489) );
  XNOR U8107 ( .A(n8488), .B(n8485), .Z(n8487) );
  XOR U8108 ( .A(n8490), .B(n8491), .Z(n8485) );
  AND U8109 ( .A(n1410), .B(n8492), .Z(n8491) );
  XOR U8110 ( .A(p_input[2002]), .B(n8490), .Z(n8492) );
  XNOR U8111 ( .A(n8493), .B(n8494), .Z(n8490) );
  AND U8112 ( .A(n1414), .B(n8495), .Z(n8494) );
  XNOR U8113 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n8496), .Z(n8488) );
  AND U8114 ( .A(n1417), .B(n8495), .Z(n8496) );
  XOR U8115 ( .A(n8497), .B(n8493), .Z(n8495) );
  XOR U8116 ( .A(n6474), .B(n8498), .Z(o[17]) );
  AND U8117 ( .A(n30), .B(n8499), .Z(n6474) );
  XOR U8118 ( .A(n6475), .B(n8498), .Z(n8499) );
  XOR U8119 ( .A(n8500), .B(n8501), .Z(n8498) );
  AND U8120 ( .A(n34), .B(n8502), .Z(n8501) );
  XOR U8121 ( .A(p_input[1]), .B(n8500), .Z(n8502) );
  XOR U8122 ( .A(n8503), .B(n8504), .Z(n8500) );
  AND U8123 ( .A(n38), .B(n8505), .Z(n8504) );
  XOR U8124 ( .A(n8506), .B(n8507), .Z(n6475) );
  AND U8125 ( .A(n42), .B(n8505), .Z(n8507) );
  XNOR U8126 ( .A(n8508), .B(n8503), .Z(n8505) );
  XOR U8127 ( .A(n8509), .B(n8510), .Z(n8503) );
  AND U8128 ( .A(n46), .B(n8511), .Z(n8510) );
  XOR U8129 ( .A(p_input[17]), .B(n8509), .Z(n8511) );
  XOR U8130 ( .A(n8512), .B(n8513), .Z(n8509) );
  AND U8131 ( .A(n50), .B(n8514), .Z(n8513) );
  IV U8132 ( .A(n8506), .Z(n8508) );
  XNOR U8133 ( .A(n8515), .B(n8516), .Z(n8506) );
  AND U8134 ( .A(n54), .B(n8514), .Z(n8516) );
  XNOR U8135 ( .A(n8515), .B(n8512), .Z(n8514) );
  XOR U8136 ( .A(n8517), .B(n8518), .Z(n8512) );
  AND U8137 ( .A(n57), .B(n8519), .Z(n8518) );
  XOR U8138 ( .A(p_input[33]), .B(n8517), .Z(n8519) );
  XOR U8139 ( .A(n8520), .B(n8521), .Z(n8517) );
  AND U8140 ( .A(n61), .B(n8522), .Z(n8521) );
  XOR U8141 ( .A(n8523), .B(n8524), .Z(n8515) );
  AND U8142 ( .A(n65), .B(n8522), .Z(n8524) );
  XNOR U8143 ( .A(n8523), .B(n8520), .Z(n8522) );
  XOR U8144 ( .A(n8525), .B(n8526), .Z(n8520) );
  AND U8145 ( .A(n68), .B(n8527), .Z(n8526) );
  XOR U8146 ( .A(p_input[49]), .B(n8525), .Z(n8527) );
  XOR U8147 ( .A(n8528), .B(n8529), .Z(n8525) );
  AND U8148 ( .A(n72), .B(n8530), .Z(n8529) );
  XOR U8149 ( .A(n8531), .B(n8532), .Z(n8523) );
  AND U8150 ( .A(n76), .B(n8530), .Z(n8532) );
  XNOR U8151 ( .A(n8531), .B(n8528), .Z(n8530) );
  XOR U8152 ( .A(n8533), .B(n8534), .Z(n8528) );
  AND U8153 ( .A(n79), .B(n8535), .Z(n8534) );
  XOR U8154 ( .A(p_input[65]), .B(n8533), .Z(n8535) );
  XOR U8155 ( .A(n8536), .B(n8537), .Z(n8533) );
  AND U8156 ( .A(n83), .B(n8538), .Z(n8537) );
  XOR U8157 ( .A(n8539), .B(n8540), .Z(n8531) );
  AND U8158 ( .A(n87), .B(n8538), .Z(n8540) );
  XNOR U8159 ( .A(n8539), .B(n8536), .Z(n8538) );
  XOR U8160 ( .A(n8541), .B(n8542), .Z(n8536) );
  AND U8161 ( .A(n90), .B(n8543), .Z(n8542) );
  XOR U8162 ( .A(p_input[81]), .B(n8541), .Z(n8543) );
  XOR U8163 ( .A(n8544), .B(n8545), .Z(n8541) );
  AND U8164 ( .A(n94), .B(n8546), .Z(n8545) );
  XOR U8165 ( .A(n8547), .B(n8548), .Z(n8539) );
  AND U8166 ( .A(n98), .B(n8546), .Z(n8548) );
  XNOR U8167 ( .A(n8547), .B(n8544), .Z(n8546) );
  XOR U8168 ( .A(n8549), .B(n8550), .Z(n8544) );
  AND U8169 ( .A(n101), .B(n8551), .Z(n8550) );
  XOR U8170 ( .A(p_input[97]), .B(n8549), .Z(n8551) );
  XOR U8171 ( .A(n8552), .B(n8553), .Z(n8549) );
  AND U8172 ( .A(n105), .B(n8554), .Z(n8553) );
  XOR U8173 ( .A(n8555), .B(n8556), .Z(n8547) );
  AND U8174 ( .A(n109), .B(n8554), .Z(n8556) );
  XNOR U8175 ( .A(n8555), .B(n8552), .Z(n8554) );
  XOR U8176 ( .A(n8557), .B(n8558), .Z(n8552) );
  AND U8177 ( .A(n112), .B(n8559), .Z(n8558) );
  XOR U8178 ( .A(p_input[113]), .B(n8557), .Z(n8559) );
  XOR U8179 ( .A(n8560), .B(n8561), .Z(n8557) );
  AND U8180 ( .A(n116), .B(n8562), .Z(n8561) );
  XOR U8181 ( .A(n8563), .B(n8564), .Z(n8555) );
  AND U8182 ( .A(n120), .B(n8562), .Z(n8564) );
  XNOR U8183 ( .A(n8563), .B(n8560), .Z(n8562) );
  XOR U8184 ( .A(n8565), .B(n8566), .Z(n8560) );
  AND U8185 ( .A(n123), .B(n8567), .Z(n8566) );
  XOR U8186 ( .A(p_input[129]), .B(n8565), .Z(n8567) );
  XOR U8187 ( .A(n8568), .B(n8569), .Z(n8565) );
  AND U8188 ( .A(n127), .B(n8570), .Z(n8569) );
  XOR U8189 ( .A(n8571), .B(n8572), .Z(n8563) );
  AND U8190 ( .A(n131), .B(n8570), .Z(n8572) );
  XNOR U8191 ( .A(n8571), .B(n8568), .Z(n8570) );
  XOR U8192 ( .A(n8573), .B(n8574), .Z(n8568) );
  AND U8193 ( .A(n134), .B(n8575), .Z(n8574) );
  XOR U8194 ( .A(p_input[145]), .B(n8573), .Z(n8575) );
  XOR U8195 ( .A(n8576), .B(n8577), .Z(n8573) );
  AND U8196 ( .A(n138), .B(n8578), .Z(n8577) );
  XOR U8197 ( .A(n8579), .B(n8580), .Z(n8571) );
  AND U8198 ( .A(n142), .B(n8578), .Z(n8580) );
  XNOR U8199 ( .A(n8579), .B(n8576), .Z(n8578) );
  XOR U8200 ( .A(n8581), .B(n8582), .Z(n8576) );
  AND U8201 ( .A(n145), .B(n8583), .Z(n8582) );
  XOR U8202 ( .A(p_input[161]), .B(n8581), .Z(n8583) );
  XOR U8203 ( .A(n8584), .B(n8585), .Z(n8581) );
  AND U8204 ( .A(n149), .B(n8586), .Z(n8585) );
  XOR U8205 ( .A(n8587), .B(n8588), .Z(n8579) );
  AND U8206 ( .A(n153), .B(n8586), .Z(n8588) );
  XNOR U8207 ( .A(n8587), .B(n8584), .Z(n8586) );
  XOR U8208 ( .A(n8589), .B(n8590), .Z(n8584) );
  AND U8209 ( .A(n156), .B(n8591), .Z(n8590) );
  XOR U8210 ( .A(p_input[177]), .B(n8589), .Z(n8591) );
  XOR U8211 ( .A(n8592), .B(n8593), .Z(n8589) );
  AND U8212 ( .A(n160), .B(n8594), .Z(n8593) );
  XOR U8213 ( .A(n8595), .B(n8596), .Z(n8587) );
  AND U8214 ( .A(n164), .B(n8594), .Z(n8596) );
  XNOR U8215 ( .A(n8595), .B(n8592), .Z(n8594) );
  XOR U8216 ( .A(n8597), .B(n8598), .Z(n8592) );
  AND U8217 ( .A(n167), .B(n8599), .Z(n8598) );
  XOR U8218 ( .A(p_input[193]), .B(n8597), .Z(n8599) );
  XOR U8219 ( .A(n8600), .B(n8601), .Z(n8597) );
  AND U8220 ( .A(n171), .B(n8602), .Z(n8601) );
  XOR U8221 ( .A(n8603), .B(n8604), .Z(n8595) );
  AND U8222 ( .A(n175), .B(n8602), .Z(n8604) );
  XNOR U8223 ( .A(n8603), .B(n8600), .Z(n8602) );
  XOR U8224 ( .A(n8605), .B(n8606), .Z(n8600) );
  AND U8225 ( .A(n178), .B(n8607), .Z(n8606) );
  XOR U8226 ( .A(p_input[209]), .B(n8605), .Z(n8607) );
  XOR U8227 ( .A(n8608), .B(n8609), .Z(n8605) );
  AND U8228 ( .A(n182), .B(n8610), .Z(n8609) );
  XOR U8229 ( .A(n8611), .B(n8612), .Z(n8603) );
  AND U8230 ( .A(n186), .B(n8610), .Z(n8612) );
  XNOR U8231 ( .A(n8611), .B(n8608), .Z(n8610) );
  XOR U8232 ( .A(n8613), .B(n8614), .Z(n8608) );
  AND U8233 ( .A(n189), .B(n8615), .Z(n8614) );
  XOR U8234 ( .A(p_input[225]), .B(n8613), .Z(n8615) );
  XOR U8235 ( .A(n8616), .B(n8617), .Z(n8613) );
  AND U8236 ( .A(n193), .B(n8618), .Z(n8617) );
  XOR U8237 ( .A(n8619), .B(n8620), .Z(n8611) );
  AND U8238 ( .A(n197), .B(n8618), .Z(n8620) );
  XNOR U8239 ( .A(n8619), .B(n8616), .Z(n8618) );
  XOR U8240 ( .A(n8621), .B(n8622), .Z(n8616) );
  AND U8241 ( .A(n200), .B(n8623), .Z(n8622) );
  XOR U8242 ( .A(p_input[241]), .B(n8621), .Z(n8623) );
  XOR U8243 ( .A(n8624), .B(n8625), .Z(n8621) );
  AND U8244 ( .A(n204), .B(n8626), .Z(n8625) );
  XOR U8245 ( .A(n8627), .B(n8628), .Z(n8619) );
  AND U8246 ( .A(n208), .B(n8626), .Z(n8628) );
  XNOR U8247 ( .A(n8627), .B(n8624), .Z(n8626) );
  XOR U8248 ( .A(n8629), .B(n8630), .Z(n8624) );
  AND U8249 ( .A(n211), .B(n8631), .Z(n8630) );
  XOR U8250 ( .A(p_input[257]), .B(n8629), .Z(n8631) );
  XOR U8251 ( .A(n8632), .B(n8633), .Z(n8629) );
  AND U8252 ( .A(n215), .B(n8634), .Z(n8633) );
  XOR U8253 ( .A(n8635), .B(n8636), .Z(n8627) );
  AND U8254 ( .A(n219), .B(n8634), .Z(n8636) );
  XNOR U8255 ( .A(n8635), .B(n8632), .Z(n8634) );
  XOR U8256 ( .A(n8637), .B(n8638), .Z(n8632) );
  AND U8257 ( .A(n222), .B(n8639), .Z(n8638) );
  XOR U8258 ( .A(p_input[273]), .B(n8637), .Z(n8639) );
  XOR U8259 ( .A(n8640), .B(n8641), .Z(n8637) );
  AND U8260 ( .A(n226), .B(n8642), .Z(n8641) );
  XOR U8261 ( .A(n8643), .B(n8644), .Z(n8635) );
  AND U8262 ( .A(n230), .B(n8642), .Z(n8644) );
  XNOR U8263 ( .A(n8643), .B(n8640), .Z(n8642) );
  XOR U8264 ( .A(n8645), .B(n8646), .Z(n8640) );
  AND U8265 ( .A(n233), .B(n8647), .Z(n8646) );
  XOR U8266 ( .A(p_input[289]), .B(n8645), .Z(n8647) );
  XOR U8267 ( .A(n8648), .B(n8649), .Z(n8645) );
  AND U8268 ( .A(n237), .B(n8650), .Z(n8649) );
  XOR U8269 ( .A(n8651), .B(n8652), .Z(n8643) );
  AND U8270 ( .A(n241), .B(n8650), .Z(n8652) );
  XNOR U8271 ( .A(n8651), .B(n8648), .Z(n8650) );
  XOR U8272 ( .A(n8653), .B(n8654), .Z(n8648) );
  AND U8273 ( .A(n244), .B(n8655), .Z(n8654) );
  XOR U8274 ( .A(p_input[305]), .B(n8653), .Z(n8655) );
  XOR U8275 ( .A(n8656), .B(n8657), .Z(n8653) );
  AND U8276 ( .A(n248), .B(n8658), .Z(n8657) );
  XOR U8277 ( .A(n8659), .B(n8660), .Z(n8651) );
  AND U8278 ( .A(n252), .B(n8658), .Z(n8660) );
  XNOR U8279 ( .A(n8659), .B(n8656), .Z(n8658) );
  XOR U8280 ( .A(n8661), .B(n8662), .Z(n8656) );
  AND U8281 ( .A(n255), .B(n8663), .Z(n8662) );
  XOR U8282 ( .A(p_input[321]), .B(n8661), .Z(n8663) );
  XOR U8283 ( .A(n8664), .B(n8665), .Z(n8661) );
  AND U8284 ( .A(n259), .B(n8666), .Z(n8665) );
  XOR U8285 ( .A(n8667), .B(n8668), .Z(n8659) );
  AND U8286 ( .A(n263), .B(n8666), .Z(n8668) );
  XNOR U8287 ( .A(n8667), .B(n8664), .Z(n8666) );
  XOR U8288 ( .A(n8669), .B(n8670), .Z(n8664) );
  AND U8289 ( .A(n266), .B(n8671), .Z(n8670) );
  XOR U8290 ( .A(p_input[337]), .B(n8669), .Z(n8671) );
  XOR U8291 ( .A(n8672), .B(n8673), .Z(n8669) );
  AND U8292 ( .A(n270), .B(n8674), .Z(n8673) );
  XOR U8293 ( .A(n8675), .B(n8676), .Z(n8667) );
  AND U8294 ( .A(n274), .B(n8674), .Z(n8676) );
  XNOR U8295 ( .A(n8675), .B(n8672), .Z(n8674) );
  XOR U8296 ( .A(n8677), .B(n8678), .Z(n8672) );
  AND U8297 ( .A(n277), .B(n8679), .Z(n8678) );
  XOR U8298 ( .A(p_input[353]), .B(n8677), .Z(n8679) );
  XOR U8299 ( .A(n8680), .B(n8681), .Z(n8677) );
  AND U8300 ( .A(n281), .B(n8682), .Z(n8681) );
  XOR U8301 ( .A(n8683), .B(n8684), .Z(n8675) );
  AND U8302 ( .A(n285), .B(n8682), .Z(n8684) );
  XNOR U8303 ( .A(n8683), .B(n8680), .Z(n8682) );
  XOR U8304 ( .A(n8685), .B(n8686), .Z(n8680) );
  AND U8305 ( .A(n288), .B(n8687), .Z(n8686) );
  XOR U8306 ( .A(p_input[369]), .B(n8685), .Z(n8687) );
  XOR U8307 ( .A(n8688), .B(n8689), .Z(n8685) );
  AND U8308 ( .A(n292), .B(n8690), .Z(n8689) );
  XOR U8309 ( .A(n8691), .B(n8692), .Z(n8683) );
  AND U8310 ( .A(n296), .B(n8690), .Z(n8692) );
  XNOR U8311 ( .A(n8691), .B(n8688), .Z(n8690) );
  XOR U8312 ( .A(n8693), .B(n8694), .Z(n8688) );
  AND U8313 ( .A(n299), .B(n8695), .Z(n8694) );
  XOR U8314 ( .A(p_input[385]), .B(n8693), .Z(n8695) );
  XOR U8315 ( .A(n8696), .B(n8697), .Z(n8693) );
  AND U8316 ( .A(n303), .B(n8698), .Z(n8697) );
  XOR U8317 ( .A(n8699), .B(n8700), .Z(n8691) );
  AND U8318 ( .A(n307), .B(n8698), .Z(n8700) );
  XNOR U8319 ( .A(n8699), .B(n8696), .Z(n8698) );
  XOR U8320 ( .A(n8701), .B(n8702), .Z(n8696) );
  AND U8321 ( .A(n310), .B(n8703), .Z(n8702) );
  XOR U8322 ( .A(p_input[401]), .B(n8701), .Z(n8703) );
  XOR U8323 ( .A(n8704), .B(n8705), .Z(n8701) );
  AND U8324 ( .A(n314), .B(n8706), .Z(n8705) );
  XOR U8325 ( .A(n8707), .B(n8708), .Z(n8699) );
  AND U8326 ( .A(n318), .B(n8706), .Z(n8708) );
  XNOR U8327 ( .A(n8707), .B(n8704), .Z(n8706) );
  XOR U8328 ( .A(n8709), .B(n8710), .Z(n8704) );
  AND U8329 ( .A(n321), .B(n8711), .Z(n8710) );
  XOR U8330 ( .A(p_input[417]), .B(n8709), .Z(n8711) );
  XOR U8331 ( .A(n8712), .B(n8713), .Z(n8709) );
  AND U8332 ( .A(n325), .B(n8714), .Z(n8713) );
  XOR U8333 ( .A(n8715), .B(n8716), .Z(n8707) );
  AND U8334 ( .A(n329), .B(n8714), .Z(n8716) );
  XNOR U8335 ( .A(n8715), .B(n8712), .Z(n8714) );
  XOR U8336 ( .A(n8717), .B(n8718), .Z(n8712) );
  AND U8337 ( .A(n332), .B(n8719), .Z(n8718) );
  XOR U8338 ( .A(p_input[433]), .B(n8717), .Z(n8719) );
  XOR U8339 ( .A(n8720), .B(n8721), .Z(n8717) );
  AND U8340 ( .A(n336), .B(n8722), .Z(n8721) );
  XOR U8341 ( .A(n8723), .B(n8724), .Z(n8715) );
  AND U8342 ( .A(n340), .B(n8722), .Z(n8724) );
  XNOR U8343 ( .A(n8723), .B(n8720), .Z(n8722) );
  XOR U8344 ( .A(n8725), .B(n8726), .Z(n8720) );
  AND U8345 ( .A(n343), .B(n8727), .Z(n8726) );
  XOR U8346 ( .A(p_input[449]), .B(n8725), .Z(n8727) );
  XOR U8347 ( .A(n8728), .B(n8729), .Z(n8725) );
  AND U8348 ( .A(n347), .B(n8730), .Z(n8729) );
  XOR U8349 ( .A(n8731), .B(n8732), .Z(n8723) );
  AND U8350 ( .A(n351), .B(n8730), .Z(n8732) );
  XNOR U8351 ( .A(n8731), .B(n8728), .Z(n8730) );
  XOR U8352 ( .A(n8733), .B(n8734), .Z(n8728) );
  AND U8353 ( .A(n354), .B(n8735), .Z(n8734) );
  XOR U8354 ( .A(p_input[465]), .B(n8733), .Z(n8735) );
  XOR U8355 ( .A(n8736), .B(n8737), .Z(n8733) );
  AND U8356 ( .A(n358), .B(n8738), .Z(n8737) );
  XOR U8357 ( .A(n8739), .B(n8740), .Z(n8731) );
  AND U8358 ( .A(n362), .B(n8738), .Z(n8740) );
  XNOR U8359 ( .A(n8739), .B(n8736), .Z(n8738) );
  XOR U8360 ( .A(n8741), .B(n8742), .Z(n8736) );
  AND U8361 ( .A(n365), .B(n8743), .Z(n8742) );
  XOR U8362 ( .A(p_input[481]), .B(n8741), .Z(n8743) );
  XOR U8363 ( .A(n8744), .B(n8745), .Z(n8741) );
  AND U8364 ( .A(n369), .B(n8746), .Z(n8745) );
  XOR U8365 ( .A(n8747), .B(n8748), .Z(n8739) );
  AND U8366 ( .A(n373), .B(n8746), .Z(n8748) );
  XNOR U8367 ( .A(n8747), .B(n8744), .Z(n8746) );
  XOR U8368 ( .A(n8749), .B(n8750), .Z(n8744) );
  AND U8369 ( .A(n376), .B(n8751), .Z(n8750) );
  XOR U8370 ( .A(p_input[497]), .B(n8749), .Z(n8751) );
  XOR U8371 ( .A(n8752), .B(n8753), .Z(n8749) );
  AND U8372 ( .A(n380), .B(n8754), .Z(n8753) );
  XOR U8373 ( .A(n8755), .B(n8756), .Z(n8747) );
  AND U8374 ( .A(n384), .B(n8754), .Z(n8756) );
  XNOR U8375 ( .A(n8755), .B(n8752), .Z(n8754) );
  XOR U8376 ( .A(n8757), .B(n8758), .Z(n8752) );
  AND U8377 ( .A(n387), .B(n8759), .Z(n8758) );
  XOR U8378 ( .A(p_input[513]), .B(n8757), .Z(n8759) );
  XOR U8379 ( .A(n8760), .B(n8761), .Z(n8757) );
  AND U8380 ( .A(n391), .B(n8762), .Z(n8761) );
  XOR U8381 ( .A(n8763), .B(n8764), .Z(n8755) );
  AND U8382 ( .A(n395), .B(n8762), .Z(n8764) );
  XNOR U8383 ( .A(n8763), .B(n8760), .Z(n8762) );
  XOR U8384 ( .A(n8765), .B(n8766), .Z(n8760) );
  AND U8385 ( .A(n398), .B(n8767), .Z(n8766) );
  XOR U8386 ( .A(p_input[529]), .B(n8765), .Z(n8767) );
  XOR U8387 ( .A(n8768), .B(n8769), .Z(n8765) );
  AND U8388 ( .A(n402), .B(n8770), .Z(n8769) );
  XOR U8389 ( .A(n8771), .B(n8772), .Z(n8763) );
  AND U8390 ( .A(n406), .B(n8770), .Z(n8772) );
  XNOR U8391 ( .A(n8771), .B(n8768), .Z(n8770) );
  XOR U8392 ( .A(n8773), .B(n8774), .Z(n8768) );
  AND U8393 ( .A(n409), .B(n8775), .Z(n8774) );
  XOR U8394 ( .A(p_input[545]), .B(n8773), .Z(n8775) );
  XOR U8395 ( .A(n8776), .B(n8777), .Z(n8773) );
  AND U8396 ( .A(n413), .B(n8778), .Z(n8777) );
  XOR U8397 ( .A(n8779), .B(n8780), .Z(n8771) );
  AND U8398 ( .A(n417), .B(n8778), .Z(n8780) );
  XNOR U8399 ( .A(n8779), .B(n8776), .Z(n8778) );
  XOR U8400 ( .A(n8781), .B(n8782), .Z(n8776) );
  AND U8401 ( .A(n420), .B(n8783), .Z(n8782) );
  XOR U8402 ( .A(p_input[561]), .B(n8781), .Z(n8783) );
  XOR U8403 ( .A(n8784), .B(n8785), .Z(n8781) );
  AND U8404 ( .A(n424), .B(n8786), .Z(n8785) );
  XOR U8405 ( .A(n8787), .B(n8788), .Z(n8779) );
  AND U8406 ( .A(n428), .B(n8786), .Z(n8788) );
  XNOR U8407 ( .A(n8787), .B(n8784), .Z(n8786) );
  XOR U8408 ( .A(n8789), .B(n8790), .Z(n8784) );
  AND U8409 ( .A(n431), .B(n8791), .Z(n8790) );
  XOR U8410 ( .A(p_input[577]), .B(n8789), .Z(n8791) );
  XOR U8411 ( .A(n8792), .B(n8793), .Z(n8789) );
  AND U8412 ( .A(n435), .B(n8794), .Z(n8793) );
  XOR U8413 ( .A(n8795), .B(n8796), .Z(n8787) );
  AND U8414 ( .A(n439), .B(n8794), .Z(n8796) );
  XNOR U8415 ( .A(n8795), .B(n8792), .Z(n8794) );
  XOR U8416 ( .A(n8797), .B(n8798), .Z(n8792) );
  AND U8417 ( .A(n442), .B(n8799), .Z(n8798) );
  XOR U8418 ( .A(p_input[593]), .B(n8797), .Z(n8799) );
  XOR U8419 ( .A(n8800), .B(n8801), .Z(n8797) );
  AND U8420 ( .A(n446), .B(n8802), .Z(n8801) );
  XOR U8421 ( .A(n8803), .B(n8804), .Z(n8795) );
  AND U8422 ( .A(n450), .B(n8802), .Z(n8804) );
  XNOR U8423 ( .A(n8803), .B(n8800), .Z(n8802) );
  XOR U8424 ( .A(n8805), .B(n8806), .Z(n8800) );
  AND U8425 ( .A(n453), .B(n8807), .Z(n8806) );
  XOR U8426 ( .A(p_input[609]), .B(n8805), .Z(n8807) );
  XOR U8427 ( .A(n8808), .B(n8809), .Z(n8805) );
  AND U8428 ( .A(n457), .B(n8810), .Z(n8809) );
  XOR U8429 ( .A(n8811), .B(n8812), .Z(n8803) );
  AND U8430 ( .A(n461), .B(n8810), .Z(n8812) );
  XNOR U8431 ( .A(n8811), .B(n8808), .Z(n8810) );
  XOR U8432 ( .A(n8813), .B(n8814), .Z(n8808) );
  AND U8433 ( .A(n464), .B(n8815), .Z(n8814) );
  XOR U8434 ( .A(p_input[625]), .B(n8813), .Z(n8815) );
  XOR U8435 ( .A(n8816), .B(n8817), .Z(n8813) );
  AND U8436 ( .A(n468), .B(n8818), .Z(n8817) );
  XOR U8437 ( .A(n8819), .B(n8820), .Z(n8811) );
  AND U8438 ( .A(n472), .B(n8818), .Z(n8820) );
  XNOR U8439 ( .A(n8819), .B(n8816), .Z(n8818) );
  XOR U8440 ( .A(n8821), .B(n8822), .Z(n8816) );
  AND U8441 ( .A(n475), .B(n8823), .Z(n8822) );
  XOR U8442 ( .A(p_input[641]), .B(n8821), .Z(n8823) );
  XOR U8443 ( .A(n8824), .B(n8825), .Z(n8821) );
  AND U8444 ( .A(n479), .B(n8826), .Z(n8825) );
  XOR U8445 ( .A(n8827), .B(n8828), .Z(n8819) );
  AND U8446 ( .A(n483), .B(n8826), .Z(n8828) );
  XNOR U8447 ( .A(n8827), .B(n8824), .Z(n8826) );
  XOR U8448 ( .A(n8829), .B(n8830), .Z(n8824) );
  AND U8449 ( .A(n486), .B(n8831), .Z(n8830) );
  XOR U8450 ( .A(p_input[657]), .B(n8829), .Z(n8831) );
  XOR U8451 ( .A(n8832), .B(n8833), .Z(n8829) );
  AND U8452 ( .A(n490), .B(n8834), .Z(n8833) );
  XOR U8453 ( .A(n8835), .B(n8836), .Z(n8827) );
  AND U8454 ( .A(n494), .B(n8834), .Z(n8836) );
  XNOR U8455 ( .A(n8835), .B(n8832), .Z(n8834) );
  XOR U8456 ( .A(n8837), .B(n8838), .Z(n8832) );
  AND U8457 ( .A(n497), .B(n8839), .Z(n8838) );
  XOR U8458 ( .A(p_input[673]), .B(n8837), .Z(n8839) );
  XOR U8459 ( .A(n8840), .B(n8841), .Z(n8837) );
  AND U8460 ( .A(n501), .B(n8842), .Z(n8841) );
  XOR U8461 ( .A(n8843), .B(n8844), .Z(n8835) );
  AND U8462 ( .A(n505), .B(n8842), .Z(n8844) );
  XNOR U8463 ( .A(n8843), .B(n8840), .Z(n8842) );
  XOR U8464 ( .A(n8845), .B(n8846), .Z(n8840) );
  AND U8465 ( .A(n508), .B(n8847), .Z(n8846) );
  XOR U8466 ( .A(p_input[689]), .B(n8845), .Z(n8847) );
  XOR U8467 ( .A(n8848), .B(n8849), .Z(n8845) );
  AND U8468 ( .A(n512), .B(n8850), .Z(n8849) );
  XOR U8469 ( .A(n8851), .B(n8852), .Z(n8843) );
  AND U8470 ( .A(n516), .B(n8850), .Z(n8852) );
  XNOR U8471 ( .A(n8851), .B(n8848), .Z(n8850) );
  XOR U8472 ( .A(n8853), .B(n8854), .Z(n8848) );
  AND U8473 ( .A(n519), .B(n8855), .Z(n8854) );
  XOR U8474 ( .A(p_input[705]), .B(n8853), .Z(n8855) );
  XOR U8475 ( .A(n8856), .B(n8857), .Z(n8853) );
  AND U8476 ( .A(n523), .B(n8858), .Z(n8857) );
  XOR U8477 ( .A(n8859), .B(n8860), .Z(n8851) );
  AND U8478 ( .A(n527), .B(n8858), .Z(n8860) );
  XNOR U8479 ( .A(n8859), .B(n8856), .Z(n8858) );
  XOR U8480 ( .A(n8861), .B(n8862), .Z(n8856) );
  AND U8481 ( .A(n530), .B(n8863), .Z(n8862) );
  XOR U8482 ( .A(p_input[721]), .B(n8861), .Z(n8863) );
  XOR U8483 ( .A(n8864), .B(n8865), .Z(n8861) );
  AND U8484 ( .A(n534), .B(n8866), .Z(n8865) );
  XOR U8485 ( .A(n8867), .B(n8868), .Z(n8859) );
  AND U8486 ( .A(n538), .B(n8866), .Z(n8868) );
  XNOR U8487 ( .A(n8867), .B(n8864), .Z(n8866) );
  XOR U8488 ( .A(n8869), .B(n8870), .Z(n8864) );
  AND U8489 ( .A(n541), .B(n8871), .Z(n8870) );
  XOR U8490 ( .A(p_input[737]), .B(n8869), .Z(n8871) );
  XOR U8491 ( .A(n8872), .B(n8873), .Z(n8869) );
  AND U8492 ( .A(n545), .B(n8874), .Z(n8873) );
  XOR U8493 ( .A(n8875), .B(n8876), .Z(n8867) );
  AND U8494 ( .A(n549), .B(n8874), .Z(n8876) );
  XNOR U8495 ( .A(n8875), .B(n8872), .Z(n8874) );
  XOR U8496 ( .A(n8877), .B(n8878), .Z(n8872) );
  AND U8497 ( .A(n552), .B(n8879), .Z(n8878) );
  XOR U8498 ( .A(p_input[753]), .B(n8877), .Z(n8879) );
  XOR U8499 ( .A(n8880), .B(n8881), .Z(n8877) );
  AND U8500 ( .A(n556), .B(n8882), .Z(n8881) );
  XOR U8501 ( .A(n8883), .B(n8884), .Z(n8875) );
  AND U8502 ( .A(n560), .B(n8882), .Z(n8884) );
  XNOR U8503 ( .A(n8883), .B(n8880), .Z(n8882) );
  XOR U8504 ( .A(n8885), .B(n8886), .Z(n8880) );
  AND U8505 ( .A(n563), .B(n8887), .Z(n8886) );
  XOR U8506 ( .A(p_input[769]), .B(n8885), .Z(n8887) );
  XOR U8507 ( .A(n8888), .B(n8889), .Z(n8885) );
  AND U8508 ( .A(n567), .B(n8890), .Z(n8889) );
  XOR U8509 ( .A(n8891), .B(n8892), .Z(n8883) );
  AND U8510 ( .A(n571), .B(n8890), .Z(n8892) );
  XNOR U8511 ( .A(n8891), .B(n8888), .Z(n8890) );
  XOR U8512 ( .A(n8893), .B(n8894), .Z(n8888) );
  AND U8513 ( .A(n574), .B(n8895), .Z(n8894) );
  XOR U8514 ( .A(p_input[785]), .B(n8893), .Z(n8895) );
  XOR U8515 ( .A(n8896), .B(n8897), .Z(n8893) );
  AND U8516 ( .A(n578), .B(n8898), .Z(n8897) );
  XOR U8517 ( .A(n8899), .B(n8900), .Z(n8891) );
  AND U8518 ( .A(n582), .B(n8898), .Z(n8900) );
  XNOR U8519 ( .A(n8899), .B(n8896), .Z(n8898) );
  XOR U8520 ( .A(n8901), .B(n8902), .Z(n8896) );
  AND U8521 ( .A(n585), .B(n8903), .Z(n8902) );
  XOR U8522 ( .A(p_input[801]), .B(n8901), .Z(n8903) );
  XOR U8523 ( .A(n8904), .B(n8905), .Z(n8901) );
  AND U8524 ( .A(n589), .B(n8906), .Z(n8905) );
  XOR U8525 ( .A(n8907), .B(n8908), .Z(n8899) );
  AND U8526 ( .A(n593), .B(n8906), .Z(n8908) );
  XNOR U8527 ( .A(n8907), .B(n8904), .Z(n8906) );
  XOR U8528 ( .A(n8909), .B(n8910), .Z(n8904) );
  AND U8529 ( .A(n596), .B(n8911), .Z(n8910) );
  XOR U8530 ( .A(p_input[817]), .B(n8909), .Z(n8911) );
  XOR U8531 ( .A(n8912), .B(n8913), .Z(n8909) );
  AND U8532 ( .A(n600), .B(n8914), .Z(n8913) );
  XOR U8533 ( .A(n8915), .B(n8916), .Z(n8907) );
  AND U8534 ( .A(n604), .B(n8914), .Z(n8916) );
  XNOR U8535 ( .A(n8915), .B(n8912), .Z(n8914) );
  XOR U8536 ( .A(n8917), .B(n8918), .Z(n8912) );
  AND U8537 ( .A(n607), .B(n8919), .Z(n8918) );
  XOR U8538 ( .A(p_input[833]), .B(n8917), .Z(n8919) );
  XOR U8539 ( .A(n8920), .B(n8921), .Z(n8917) );
  AND U8540 ( .A(n611), .B(n8922), .Z(n8921) );
  XOR U8541 ( .A(n8923), .B(n8924), .Z(n8915) );
  AND U8542 ( .A(n615), .B(n8922), .Z(n8924) );
  XNOR U8543 ( .A(n8923), .B(n8920), .Z(n8922) );
  XOR U8544 ( .A(n8925), .B(n8926), .Z(n8920) );
  AND U8545 ( .A(n618), .B(n8927), .Z(n8926) );
  XOR U8546 ( .A(p_input[849]), .B(n8925), .Z(n8927) );
  XOR U8547 ( .A(n8928), .B(n8929), .Z(n8925) );
  AND U8548 ( .A(n622), .B(n8930), .Z(n8929) );
  XOR U8549 ( .A(n8931), .B(n8932), .Z(n8923) );
  AND U8550 ( .A(n626), .B(n8930), .Z(n8932) );
  XNOR U8551 ( .A(n8931), .B(n8928), .Z(n8930) );
  XOR U8552 ( .A(n8933), .B(n8934), .Z(n8928) );
  AND U8553 ( .A(n629), .B(n8935), .Z(n8934) );
  XOR U8554 ( .A(p_input[865]), .B(n8933), .Z(n8935) );
  XOR U8555 ( .A(n8936), .B(n8937), .Z(n8933) );
  AND U8556 ( .A(n633), .B(n8938), .Z(n8937) );
  XOR U8557 ( .A(n8939), .B(n8940), .Z(n8931) );
  AND U8558 ( .A(n637), .B(n8938), .Z(n8940) );
  XNOR U8559 ( .A(n8939), .B(n8936), .Z(n8938) );
  XOR U8560 ( .A(n8941), .B(n8942), .Z(n8936) );
  AND U8561 ( .A(n640), .B(n8943), .Z(n8942) );
  XOR U8562 ( .A(p_input[881]), .B(n8941), .Z(n8943) );
  XOR U8563 ( .A(n8944), .B(n8945), .Z(n8941) );
  AND U8564 ( .A(n644), .B(n8946), .Z(n8945) );
  XOR U8565 ( .A(n8947), .B(n8948), .Z(n8939) );
  AND U8566 ( .A(n648), .B(n8946), .Z(n8948) );
  XNOR U8567 ( .A(n8947), .B(n8944), .Z(n8946) );
  XOR U8568 ( .A(n8949), .B(n8950), .Z(n8944) );
  AND U8569 ( .A(n651), .B(n8951), .Z(n8950) );
  XOR U8570 ( .A(p_input[897]), .B(n8949), .Z(n8951) );
  XOR U8571 ( .A(n8952), .B(n8953), .Z(n8949) );
  AND U8572 ( .A(n655), .B(n8954), .Z(n8953) );
  XOR U8573 ( .A(n8955), .B(n8956), .Z(n8947) );
  AND U8574 ( .A(n659), .B(n8954), .Z(n8956) );
  XNOR U8575 ( .A(n8955), .B(n8952), .Z(n8954) );
  XOR U8576 ( .A(n8957), .B(n8958), .Z(n8952) );
  AND U8577 ( .A(n662), .B(n8959), .Z(n8958) );
  XOR U8578 ( .A(p_input[913]), .B(n8957), .Z(n8959) );
  XOR U8579 ( .A(n8960), .B(n8961), .Z(n8957) );
  AND U8580 ( .A(n666), .B(n8962), .Z(n8961) );
  XOR U8581 ( .A(n8963), .B(n8964), .Z(n8955) );
  AND U8582 ( .A(n670), .B(n8962), .Z(n8964) );
  XNOR U8583 ( .A(n8963), .B(n8960), .Z(n8962) );
  XOR U8584 ( .A(n8965), .B(n8966), .Z(n8960) );
  AND U8585 ( .A(n673), .B(n8967), .Z(n8966) );
  XOR U8586 ( .A(p_input[929]), .B(n8965), .Z(n8967) );
  XOR U8587 ( .A(n8968), .B(n8969), .Z(n8965) );
  AND U8588 ( .A(n677), .B(n8970), .Z(n8969) );
  XOR U8589 ( .A(n8971), .B(n8972), .Z(n8963) );
  AND U8590 ( .A(n681), .B(n8970), .Z(n8972) );
  XNOR U8591 ( .A(n8971), .B(n8968), .Z(n8970) );
  XOR U8592 ( .A(n8973), .B(n8974), .Z(n8968) );
  AND U8593 ( .A(n684), .B(n8975), .Z(n8974) );
  XOR U8594 ( .A(p_input[945]), .B(n8973), .Z(n8975) );
  XOR U8595 ( .A(n8976), .B(n8977), .Z(n8973) );
  AND U8596 ( .A(n688), .B(n8978), .Z(n8977) );
  XOR U8597 ( .A(n8979), .B(n8980), .Z(n8971) );
  AND U8598 ( .A(n692), .B(n8978), .Z(n8980) );
  XNOR U8599 ( .A(n8979), .B(n8976), .Z(n8978) );
  XOR U8600 ( .A(n8981), .B(n8982), .Z(n8976) );
  AND U8601 ( .A(n695), .B(n8983), .Z(n8982) );
  XOR U8602 ( .A(p_input[961]), .B(n8981), .Z(n8983) );
  XOR U8603 ( .A(n8984), .B(n8985), .Z(n8981) );
  AND U8604 ( .A(n699), .B(n8986), .Z(n8985) );
  XOR U8605 ( .A(n8987), .B(n8988), .Z(n8979) );
  AND U8606 ( .A(n703), .B(n8986), .Z(n8988) );
  XNOR U8607 ( .A(n8987), .B(n8984), .Z(n8986) );
  XOR U8608 ( .A(n8989), .B(n8990), .Z(n8984) );
  AND U8609 ( .A(n706), .B(n8991), .Z(n8990) );
  XOR U8610 ( .A(p_input[977]), .B(n8989), .Z(n8991) );
  XOR U8611 ( .A(n8992), .B(n8993), .Z(n8989) );
  AND U8612 ( .A(n710), .B(n8994), .Z(n8993) );
  XOR U8613 ( .A(n8995), .B(n8996), .Z(n8987) );
  AND U8614 ( .A(n714), .B(n8994), .Z(n8996) );
  XNOR U8615 ( .A(n8995), .B(n8992), .Z(n8994) );
  XOR U8616 ( .A(n8997), .B(n8998), .Z(n8992) );
  AND U8617 ( .A(n717), .B(n8999), .Z(n8998) );
  XOR U8618 ( .A(p_input[993]), .B(n8997), .Z(n8999) );
  XOR U8619 ( .A(n9000), .B(n9001), .Z(n8997) );
  AND U8620 ( .A(n721), .B(n9002), .Z(n9001) );
  XOR U8621 ( .A(n9003), .B(n9004), .Z(n8995) );
  AND U8622 ( .A(n725), .B(n9002), .Z(n9004) );
  XNOR U8623 ( .A(n9003), .B(n9000), .Z(n9002) );
  XOR U8624 ( .A(n9005), .B(n9006), .Z(n9000) );
  AND U8625 ( .A(n728), .B(n9007), .Z(n9006) );
  XOR U8626 ( .A(p_input[1009]), .B(n9005), .Z(n9007) );
  XOR U8627 ( .A(n9008), .B(n9009), .Z(n9005) );
  AND U8628 ( .A(n732), .B(n9010), .Z(n9009) );
  XOR U8629 ( .A(n9011), .B(n9012), .Z(n9003) );
  AND U8630 ( .A(n736), .B(n9010), .Z(n9012) );
  XNOR U8631 ( .A(n9011), .B(n9008), .Z(n9010) );
  XOR U8632 ( .A(n9013), .B(n9014), .Z(n9008) );
  AND U8633 ( .A(n739), .B(n9015), .Z(n9014) );
  XOR U8634 ( .A(p_input[1025]), .B(n9013), .Z(n9015) );
  XOR U8635 ( .A(n9016), .B(n9017), .Z(n9013) );
  AND U8636 ( .A(n743), .B(n9018), .Z(n9017) );
  XOR U8637 ( .A(n9019), .B(n9020), .Z(n9011) );
  AND U8638 ( .A(n747), .B(n9018), .Z(n9020) );
  XNOR U8639 ( .A(n9019), .B(n9016), .Z(n9018) );
  XOR U8640 ( .A(n9021), .B(n9022), .Z(n9016) );
  AND U8641 ( .A(n750), .B(n9023), .Z(n9022) );
  XOR U8642 ( .A(p_input[1041]), .B(n9021), .Z(n9023) );
  XOR U8643 ( .A(n9024), .B(n9025), .Z(n9021) );
  AND U8644 ( .A(n754), .B(n9026), .Z(n9025) );
  XOR U8645 ( .A(n9027), .B(n9028), .Z(n9019) );
  AND U8646 ( .A(n758), .B(n9026), .Z(n9028) );
  XNOR U8647 ( .A(n9027), .B(n9024), .Z(n9026) );
  XOR U8648 ( .A(n9029), .B(n9030), .Z(n9024) );
  AND U8649 ( .A(n761), .B(n9031), .Z(n9030) );
  XOR U8650 ( .A(p_input[1057]), .B(n9029), .Z(n9031) );
  XOR U8651 ( .A(n9032), .B(n9033), .Z(n9029) );
  AND U8652 ( .A(n765), .B(n9034), .Z(n9033) );
  XOR U8653 ( .A(n9035), .B(n9036), .Z(n9027) );
  AND U8654 ( .A(n769), .B(n9034), .Z(n9036) );
  XNOR U8655 ( .A(n9035), .B(n9032), .Z(n9034) );
  XOR U8656 ( .A(n9037), .B(n9038), .Z(n9032) );
  AND U8657 ( .A(n772), .B(n9039), .Z(n9038) );
  XOR U8658 ( .A(p_input[1073]), .B(n9037), .Z(n9039) );
  XOR U8659 ( .A(n9040), .B(n9041), .Z(n9037) );
  AND U8660 ( .A(n776), .B(n9042), .Z(n9041) );
  XOR U8661 ( .A(n9043), .B(n9044), .Z(n9035) );
  AND U8662 ( .A(n780), .B(n9042), .Z(n9044) );
  XNOR U8663 ( .A(n9043), .B(n9040), .Z(n9042) );
  XOR U8664 ( .A(n9045), .B(n9046), .Z(n9040) );
  AND U8665 ( .A(n783), .B(n9047), .Z(n9046) );
  XOR U8666 ( .A(p_input[1089]), .B(n9045), .Z(n9047) );
  XOR U8667 ( .A(n9048), .B(n9049), .Z(n9045) );
  AND U8668 ( .A(n787), .B(n9050), .Z(n9049) );
  XOR U8669 ( .A(n9051), .B(n9052), .Z(n9043) );
  AND U8670 ( .A(n791), .B(n9050), .Z(n9052) );
  XNOR U8671 ( .A(n9051), .B(n9048), .Z(n9050) );
  XOR U8672 ( .A(n9053), .B(n9054), .Z(n9048) );
  AND U8673 ( .A(n794), .B(n9055), .Z(n9054) );
  XOR U8674 ( .A(p_input[1105]), .B(n9053), .Z(n9055) );
  XOR U8675 ( .A(n9056), .B(n9057), .Z(n9053) );
  AND U8676 ( .A(n798), .B(n9058), .Z(n9057) );
  XOR U8677 ( .A(n9059), .B(n9060), .Z(n9051) );
  AND U8678 ( .A(n802), .B(n9058), .Z(n9060) );
  XNOR U8679 ( .A(n9059), .B(n9056), .Z(n9058) );
  XOR U8680 ( .A(n9061), .B(n9062), .Z(n9056) );
  AND U8681 ( .A(n805), .B(n9063), .Z(n9062) );
  XOR U8682 ( .A(p_input[1121]), .B(n9061), .Z(n9063) );
  XOR U8683 ( .A(n9064), .B(n9065), .Z(n9061) );
  AND U8684 ( .A(n809), .B(n9066), .Z(n9065) );
  XOR U8685 ( .A(n9067), .B(n9068), .Z(n9059) );
  AND U8686 ( .A(n813), .B(n9066), .Z(n9068) );
  XNOR U8687 ( .A(n9067), .B(n9064), .Z(n9066) );
  XOR U8688 ( .A(n9069), .B(n9070), .Z(n9064) );
  AND U8689 ( .A(n816), .B(n9071), .Z(n9070) );
  XOR U8690 ( .A(p_input[1137]), .B(n9069), .Z(n9071) );
  XOR U8691 ( .A(n9072), .B(n9073), .Z(n9069) );
  AND U8692 ( .A(n820), .B(n9074), .Z(n9073) );
  XOR U8693 ( .A(n9075), .B(n9076), .Z(n9067) );
  AND U8694 ( .A(n824), .B(n9074), .Z(n9076) );
  XNOR U8695 ( .A(n9075), .B(n9072), .Z(n9074) );
  XOR U8696 ( .A(n9077), .B(n9078), .Z(n9072) );
  AND U8697 ( .A(n827), .B(n9079), .Z(n9078) );
  XOR U8698 ( .A(p_input[1153]), .B(n9077), .Z(n9079) );
  XOR U8699 ( .A(n9080), .B(n9081), .Z(n9077) );
  AND U8700 ( .A(n831), .B(n9082), .Z(n9081) );
  XOR U8701 ( .A(n9083), .B(n9084), .Z(n9075) );
  AND U8702 ( .A(n835), .B(n9082), .Z(n9084) );
  XNOR U8703 ( .A(n9083), .B(n9080), .Z(n9082) );
  XOR U8704 ( .A(n9085), .B(n9086), .Z(n9080) );
  AND U8705 ( .A(n838), .B(n9087), .Z(n9086) );
  XOR U8706 ( .A(p_input[1169]), .B(n9085), .Z(n9087) );
  XOR U8707 ( .A(n9088), .B(n9089), .Z(n9085) );
  AND U8708 ( .A(n842), .B(n9090), .Z(n9089) );
  XOR U8709 ( .A(n9091), .B(n9092), .Z(n9083) );
  AND U8710 ( .A(n846), .B(n9090), .Z(n9092) );
  XNOR U8711 ( .A(n9091), .B(n9088), .Z(n9090) );
  XOR U8712 ( .A(n9093), .B(n9094), .Z(n9088) );
  AND U8713 ( .A(n849), .B(n9095), .Z(n9094) );
  XOR U8714 ( .A(p_input[1185]), .B(n9093), .Z(n9095) );
  XOR U8715 ( .A(n9096), .B(n9097), .Z(n9093) );
  AND U8716 ( .A(n853), .B(n9098), .Z(n9097) );
  XOR U8717 ( .A(n9099), .B(n9100), .Z(n9091) );
  AND U8718 ( .A(n857), .B(n9098), .Z(n9100) );
  XNOR U8719 ( .A(n9099), .B(n9096), .Z(n9098) );
  XOR U8720 ( .A(n9101), .B(n9102), .Z(n9096) );
  AND U8721 ( .A(n860), .B(n9103), .Z(n9102) );
  XOR U8722 ( .A(p_input[1201]), .B(n9101), .Z(n9103) );
  XOR U8723 ( .A(n9104), .B(n9105), .Z(n9101) );
  AND U8724 ( .A(n864), .B(n9106), .Z(n9105) );
  XOR U8725 ( .A(n9107), .B(n9108), .Z(n9099) );
  AND U8726 ( .A(n868), .B(n9106), .Z(n9108) );
  XNOR U8727 ( .A(n9107), .B(n9104), .Z(n9106) );
  XOR U8728 ( .A(n9109), .B(n9110), .Z(n9104) );
  AND U8729 ( .A(n871), .B(n9111), .Z(n9110) );
  XOR U8730 ( .A(p_input[1217]), .B(n9109), .Z(n9111) );
  XOR U8731 ( .A(n9112), .B(n9113), .Z(n9109) );
  AND U8732 ( .A(n875), .B(n9114), .Z(n9113) );
  XOR U8733 ( .A(n9115), .B(n9116), .Z(n9107) );
  AND U8734 ( .A(n879), .B(n9114), .Z(n9116) );
  XNOR U8735 ( .A(n9115), .B(n9112), .Z(n9114) );
  XOR U8736 ( .A(n9117), .B(n9118), .Z(n9112) );
  AND U8737 ( .A(n882), .B(n9119), .Z(n9118) );
  XOR U8738 ( .A(p_input[1233]), .B(n9117), .Z(n9119) );
  XOR U8739 ( .A(n9120), .B(n9121), .Z(n9117) );
  AND U8740 ( .A(n886), .B(n9122), .Z(n9121) );
  XOR U8741 ( .A(n9123), .B(n9124), .Z(n9115) );
  AND U8742 ( .A(n890), .B(n9122), .Z(n9124) );
  XNOR U8743 ( .A(n9123), .B(n9120), .Z(n9122) );
  XOR U8744 ( .A(n9125), .B(n9126), .Z(n9120) );
  AND U8745 ( .A(n893), .B(n9127), .Z(n9126) );
  XOR U8746 ( .A(p_input[1249]), .B(n9125), .Z(n9127) );
  XOR U8747 ( .A(n9128), .B(n9129), .Z(n9125) );
  AND U8748 ( .A(n897), .B(n9130), .Z(n9129) );
  XOR U8749 ( .A(n9131), .B(n9132), .Z(n9123) );
  AND U8750 ( .A(n901), .B(n9130), .Z(n9132) );
  XNOR U8751 ( .A(n9131), .B(n9128), .Z(n9130) );
  XOR U8752 ( .A(n9133), .B(n9134), .Z(n9128) );
  AND U8753 ( .A(n904), .B(n9135), .Z(n9134) );
  XOR U8754 ( .A(p_input[1265]), .B(n9133), .Z(n9135) );
  XOR U8755 ( .A(n9136), .B(n9137), .Z(n9133) );
  AND U8756 ( .A(n908), .B(n9138), .Z(n9137) );
  XOR U8757 ( .A(n9139), .B(n9140), .Z(n9131) );
  AND U8758 ( .A(n912), .B(n9138), .Z(n9140) );
  XNOR U8759 ( .A(n9139), .B(n9136), .Z(n9138) );
  XOR U8760 ( .A(n9141), .B(n9142), .Z(n9136) );
  AND U8761 ( .A(n915), .B(n9143), .Z(n9142) );
  XOR U8762 ( .A(p_input[1281]), .B(n9141), .Z(n9143) );
  XOR U8763 ( .A(n9144), .B(n9145), .Z(n9141) );
  AND U8764 ( .A(n919), .B(n9146), .Z(n9145) );
  XOR U8765 ( .A(n9147), .B(n9148), .Z(n9139) );
  AND U8766 ( .A(n923), .B(n9146), .Z(n9148) );
  XNOR U8767 ( .A(n9147), .B(n9144), .Z(n9146) );
  XOR U8768 ( .A(n9149), .B(n9150), .Z(n9144) );
  AND U8769 ( .A(n926), .B(n9151), .Z(n9150) );
  XOR U8770 ( .A(p_input[1297]), .B(n9149), .Z(n9151) );
  XOR U8771 ( .A(n9152), .B(n9153), .Z(n9149) );
  AND U8772 ( .A(n930), .B(n9154), .Z(n9153) );
  XOR U8773 ( .A(n9155), .B(n9156), .Z(n9147) );
  AND U8774 ( .A(n934), .B(n9154), .Z(n9156) );
  XNOR U8775 ( .A(n9155), .B(n9152), .Z(n9154) );
  XOR U8776 ( .A(n9157), .B(n9158), .Z(n9152) );
  AND U8777 ( .A(n937), .B(n9159), .Z(n9158) );
  XOR U8778 ( .A(p_input[1313]), .B(n9157), .Z(n9159) );
  XOR U8779 ( .A(n9160), .B(n9161), .Z(n9157) );
  AND U8780 ( .A(n941), .B(n9162), .Z(n9161) );
  XOR U8781 ( .A(n9163), .B(n9164), .Z(n9155) );
  AND U8782 ( .A(n945), .B(n9162), .Z(n9164) );
  XNOR U8783 ( .A(n9163), .B(n9160), .Z(n9162) );
  XOR U8784 ( .A(n9165), .B(n9166), .Z(n9160) );
  AND U8785 ( .A(n948), .B(n9167), .Z(n9166) );
  XOR U8786 ( .A(p_input[1329]), .B(n9165), .Z(n9167) );
  XOR U8787 ( .A(n9168), .B(n9169), .Z(n9165) );
  AND U8788 ( .A(n952), .B(n9170), .Z(n9169) );
  XOR U8789 ( .A(n9171), .B(n9172), .Z(n9163) );
  AND U8790 ( .A(n956), .B(n9170), .Z(n9172) );
  XNOR U8791 ( .A(n9171), .B(n9168), .Z(n9170) );
  XOR U8792 ( .A(n9173), .B(n9174), .Z(n9168) );
  AND U8793 ( .A(n959), .B(n9175), .Z(n9174) );
  XOR U8794 ( .A(p_input[1345]), .B(n9173), .Z(n9175) );
  XOR U8795 ( .A(n9176), .B(n9177), .Z(n9173) );
  AND U8796 ( .A(n963), .B(n9178), .Z(n9177) );
  XOR U8797 ( .A(n9179), .B(n9180), .Z(n9171) );
  AND U8798 ( .A(n967), .B(n9178), .Z(n9180) );
  XNOR U8799 ( .A(n9179), .B(n9176), .Z(n9178) );
  XOR U8800 ( .A(n9181), .B(n9182), .Z(n9176) );
  AND U8801 ( .A(n970), .B(n9183), .Z(n9182) );
  XOR U8802 ( .A(p_input[1361]), .B(n9181), .Z(n9183) );
  XOR U8803 ( .A(n9184), .B(n9185), .Z(n9181) );
  AND U8804 ( .A(n974), .B(n9186), .Z(n9185) );
  XOR U8805 ( .A(n9187), .B(n9188), .Z(n9179) );
  AND U8806 ( .A(n978), .B(n9186), .Z(n9188) );
  XNOR U8807 ( .A(n9187), .B(n9184), .Z(n9186) );
  XOR U8808 ( .A(n9189), .B(n9190), .Z(n9184) );
  AND U8809 ( .A(n981), .B(n9191), .Z(n9190) );
  XOR U8810 ( .A(p_input[1377]), .B(n9189), .Z(n9191) );
  XOR U8811 ( .A(n9192), .B(n9193), .Z(n9189) );
  AND U8812 ( .A(n985), .B(n9194), .Z(n9193) );
  XOR U8813 ( .A(n9195), .B(n9196), .Z(n9187) );
  AND U8814 ( .A(n989), .B(n9194), .Z(n9196) );
  XNOR U8815 ( .A(n9195), .B(n9192), .Z(n9194) );
  XOR U8816 ( .A(n9197), .B(n9198), .Z(n9192) );
  AND U8817 ( .A(n992), .B(n9199), .Z(n9198) );
  XOR U8818 ( .A(p_input[1393]), .B(n9197), .Z(n9199) );
  XOR U8819 ( .A(n9200), .B(n9201), .Z(n9197) );
  AND U8820 ( .A(n996), .B(n9202), .Z(n9201) );
  XOR U8821 ( .A(n9203), .B(n9204), .Z(n9195) );
  AND U8822 ( .A(n1000), .B(n9202), .Z(n9204) );
  XNOR U8823 ( .A(n9203), .B(n9200), .Z(n9202) );
  XOR U8824 ( .A(n9205), .B(n9206), .Z(n9200) );
  AND U8825 ( .A(n1003), .B(n9207), .Z(n9206) );
  XOR U8826 ( .A(p_input[1409]), .B(n9205), .Z(n9207) );
  XOR U8827 ( .A(n9208), .B(n9209), .Z(n9205) );
  AND U8828 ( .A(n1007), .B(n9210), .Z(n9209) );
  XOR U8829 ( .A(n9211), .B(n9212), .Z(n9203) );
  AND U8830 ( .A(n1011), .B(n9210), .Z(n9212) );
  XNOR U8831 ( .A(n9211), .B(n9208), .Z(n9210) );
  XOR U8832 ( .A(n9213), .B(n9214), .Z(n9208) );
  AND U8833 ( .A(n1014), .B(n9215), .Z(n9214) );
  XOR U8834 ( .A(p_input[1425]), .B(n9213), .Z(n9215) );
  XOR U8835 ( .A(n9216), .B(n9217), .Z(n9213) );
  AND U8836 ( .A(n1018), .B(n9218), .Z(n9217) );
  XOR U8837 ( .A(n9219), .B(n9220), .Z(n9211) );
  AND U8838 ( .A(n1022), .B(n9218), .Z(n9220) );
  XNOR U8839 ( .A(n9219), .B(n9216), .Z(n9218) );
  XOR U8840 ( .A(n9221), .B(n9222), .Z(n9216) );
  AND U8841 ( .A(n1025), .B(n9223), .Z(n9222) );
  XOR U8842 ( .A(p_input[1441]), .B(n9221), .Z(n9223) );
  XOR U8843 ( .A(n9224), .B(n9225), .Z(n9221) );
  AND U8844 ( .A(n1029), .B(n9226), .Z(n9225) );
  XOR U8845 ( .A(n9227), .B(n9228), .Z(n9219) );
  AND U8846 ( .A(n1033), .B(n9226), .Z(n9228) );
  XNOR U8847 ( .A(n9227), .B(n9224), .Z(n9226) );
  XOR U8848 ( .A(n9229), .B(n9230), .Z(n9224) );
  AND U8849 ( .A(n1036), .B(n9231), .Z(n9230) );
  XOR U8850 ( .A(p_input[1457]), .B(n9229), .Z(n9231) );
  XOR U8851 ( .A(n9232), .B(n9233), .Z(n9229) );
  AND U8852 ( .A(n1040), .B(n9234), .Z(n9233) );
  XOR U8853 ( .A(n9235), .B(n9236), .Z(n9227) );
  AND U8854 ( .A(n1044), .B(n9234), .Z(n9236) );
  XNOR U8855 ( .A(n9235), .B(n9232), .Z(n9234) );
  XOR U8856 ( .A(n9237), .B(n9238), .Z(n9232) );
  AND U8857 ( .A(n1047), .B(n9239), .Z(n9238) );
  XOR U8858 ( .A(p_input[1473]), .B(n9237), .Z(n9239) );
  XOR U8859 ( .A(n9240), .B(n9241), .Z(n9237) );
  AND U8860 ( .A(n1051), .B(n9242), .Z(n9241) );
  XOR U8861 ( .A(n9243), .B(n9244), .Z(n9235) );
  AND U8862 ( .A(n1055), .B(n9242), .Z(n9244) );
  XNOR U8863 ( .A(n9243), .B(n9240), .Z(n9242) );
  XOR U8864 ( .A(n9245), .B(n9246), .Z(n9240) );
  AND U8865 ( .A(n1058), .B(n9247), .Z(n9246) );
  XOR U8866 ( .A(p_input[1489]), .B(n9245), .Z(n9247) );
  XOR U8867 ( .A(n9248), .B(n9249), .Z(n9245) );
  AND U8868 ( .A(n1062), .B(n9250), .Z(n9249) );
  XOR U8869 ( .A(n9251), .B(n9252), .Z(n9243) );
  AND U8870 ( .A(n1066), .B(n9250), .Z(n9252) );
  XNOR U8871 ( .A(n9251), .B(n9248), .Z(n9250) );
  XOR U8872 ( .A(n9253), .B(n9254), .Z(n9248) );
  AND U8873 ( .A(n1069), .B(n9255), .Z(n9254) );
  XOR U8874 ( .A(p_input[1505]), .B(n9253), .Z(n9255) );
  XOR U8875 ( .A(n9256), .B(n9257), .Z(n9253) );
  AND U8876 ( .A(n1073), .B(n9258), .Z(n9257) );
  XOR U8877 ( .A(n9259), .B(n9260), .Z(n9251) );
  AND U8878 ( .A(n1077), .B(n9258), .Z(n9260) );
  XNOR U8879 ( .A(n9259), .B(n9256), .Z(n9258) );
  XOR U8880 ( .A(n9261), .B(n9262), .Z(n9256) );
  AND U8881 ( .A(n1080), .B(n9263), .Z(n9262) );
  XOR U8882 ( .A(p_input[1521]), .B(n9261), .Z(n9263) );
  XOR U8883 ( .A(n9264), .B(n9265), .Z(n9261) );
  AND U8884 ( .A(n1084), .B(n9266), .Z(n9265) );
  XOR U8885 ( .A(n9267), .B(n9268), .Z(n9259) );
  AND U8886 ( .A(n1088), .B(n9266), .Z(n9268) );
  XNOR U8887 ( .A(n9267), .B(n9264), .Z(n9266) );
  XOR U8888 ( .A(n9269), .B(n9270), .Z(n9264) );
  AND U8889 ( .A(n1091), .B(n9271), .Z(n9270) );
  XOR U8890 ( .A(p_input[1537]), .B(n9269), .Z(n9271) );
  XOR U8891 ( .A(n9272), .B(n9273), .Z(n9269) );
  AND U8892 ( .A(n1095), .B(n9274), .Z(n9273) );
  XOR U8893 ( .A(n9275), .B(n9276), .Z(n9267) );
  AND U8894 ( .A(n1099), .B(n9274), .Z(n9276) );
  XNOR U8895 ( .A(n9275), .B(n9272), .Z(n9274) );
  XOR U8896 ( .A(n9277), .B(n9278), .Z(n9272) );
  AND U8897 ( .A(n1102), .B(n9279), .Z(n9278) );
  XOR U8898 ( .A(p_input[1553]), .B(n9277), .Z(n9279) );
  XOR U8899 ( .A(n9280), .B(n9281), .Z(n9277) );
  AND U8900 ( .A(n1106), .B(n9282), .Z(n9281) );
  XOR U8901 ( .A(n9283), .B(n9284), .Z(n9275) );
  AND U8902 ( .A(n1110), .B(n9282), .Z(n9284) );
  XNOR U8903 ( .A(n9283), .B(n9280), .Z(n9282) );
  XOR U8904 ( .A(n9285), .B(n9286), .Z(n9280) );
  AND U8905 ( .A(n1113), .B(n9287), .Z(n9286) );
  XOR U8906 ( .A(p_input[1569]), .B(n9285), .Z(n9287) );
  XOR U8907 ( .A(n9288), .B(n9289), .Z(n9285) );
  AND U8908 ( .A(n1117), .B(n9290), .Z(n9289) );
  XOR U8909 ( .A(n9291), .B(n9292), .Z(n9283) );
  AND U8910 ( .A(n1121), .B(n9290), .Z(n9292) );
  XNOR U8911 ( .A(n9291), .B(n9288), .Z(n9290) );
  XOR U8912 ( .A(n9293), .B(n9294), .Z(n9288) );
  AND U8913 ( .A(n1124), .B(n9295), .Z(n9294) );
  XOR U8914 ( .A(p_input[1585]), .B(n9293), .Z(n9295) );
  XOR U8915 ( .A(n9296), .B(n9297), .Z(n9293) );
  AND U8916 ( .A(n1128), .B(n9298), .Z(n9297) );
  XOR U8917 ( .A(n9299), .B(n9300), .Z(n9291) );
  AND U8918 ( .A(n1132), .B(n9298), .Z(n9300) );
  XNOR U8919 ( .A(n9299), .B(n9296), .Z(n9298) );
  XOR U8920 ( .A(n9301), .B(n9302), .Z(n9296) );
  AND U8921 ( .A(n1135), .B(n9303), .Z(n9302) );
  XOR U8922 ( .A(p_input[1601]), .B(n9301), .Z(n9303) );
  XOR U8923 ( .A(n9304), .B(n9305), .Z(n9301) );
  AND U8924 ( .A(n1139), .B(n9306), .Z(n9305) );
  XOR U8925 ( .A(n9307), .B(n9308), .Z(n9299) );
  AND U8926 ( .A(n1143), .B(n9306), .Z(n9308) );
  XNOR U8927 ( .A(n9307), .B(n9304), .Z(n9306) );
  XOR U8928 ( .A(n9309), .B(n9310), .Z(n9304) );
  AND U8929 ( .A(n1146), .B(n9311), .Z(n9310) );
  XOR U8930 ( .A(p_input[1617]), .B(n9309), .Z(n9311) );
  XOR U8931 ( .A(n9312), .B(n9313), .Z(n9309) );
  AND U8932 ( .A(n1150), .B(n9314), .Z(n9313) );
  XOR U8933 ( .A(n9315), .B(n9316), .Z(n9307) );
  AND U8934 ( .A(n1154), .B(n9314), .Z(n9316) );
  XNOR U8935 ( .A(n9315), .B(n9312), .Z(n9314) );
  XOR U8936 ( .A(n9317), .B(n9318), .Z(n9312) );
  AND U8937 ( .A(n1157), .B(n9319), .Z(n9318) );
  XOR U8938 ( .A(p_input[1633]), .B(n9317), .Z(n9319) );
  XOR U8939 ( .A(n9320), .B(n9321), .Z(n9317) );
  AND U8940 ( .A(n1161), .B(n9322), .Z(n9321) );
  XOR U8941 ( .A(n9323), .B(n9324), .Z(n9315) );
  AND U8942 ( .A(n1165), .B(n9322), .Z(n9324) );
  XNOR U8943 ( .A(n9323), .B(n9320), .Z(n9322) );
  XOR U8944 ( .A(n9325), .B(n9326), .Z(n9320) );
  AND U8945 ( .A(n1168), .B(n9327), .Z(n9326) );
  XOR U8946 ( .A(p_input[1649]), .B(n9325), .Z(n9327) );
  XOR U8947 ( .A(n9328), .B(n9329), .Z(n9325) );
  AND U8948 ( .A(n1172), .B(n9330), .Z(n9329) );
  XOR U8949 ( .A(n9331), .B(n9332), .Z(n9323) );
  AND U8950 ( .A(n1176), .B(n9330), .Z(n9332) );
  XNOR U8951 ( .A(n9331), .B(n9328), .Z(n9330) );
  XOR U8952 ( .A(n9333), .B(n9334), .Z(n9328) );
  AND U8953 ( .A(n1179), .B(n9335), .Z(n9334) );
  XOR U8954 ( .A(p_input[1665]), .B(n9333), .Z(n9335) );
  XOR U8955 ( .A(n9336), .B(n9337), .Z(n9333) );
  AND U8956 ( .A(n1183), .B(n9338), .Z(n9337) );
  XOR U8957 ( .A(n9339), .B(n9340), .Z(n9331) );
  AND U8958 ( .A(n1187), .B(n9338), .Z(n9340) );
  XNOR U8959 ( .A(n9339), .B(n9336), .Z(n9338) );
  XOR U8960 ( .A(n9341), .B(n9342), .Z(n9336) );
  AND U8961 ( .A(n1190), .B(n9343), .Z(n9342) );
  XOR U8962 ( .A(p_input[1681]), .B(n9341), .Z(n9343) );
  XOR U8963 ( .A(n9344), .B(n9345), .Z(n9341) );
  AND U8964 ( .A(n1194), .B(n9346), .Z(n9345) );
  XOR U8965 ( .A(n9347), .B(n9348), .Z(n9339) );
  AND U8966 ( .A(n1198), .B(n9346), .Z(n9348) );
  XNOR U8967 ( .A(n9347), .B(n9344), .Z(n9346) );
  XOR U8968 ( .A(n9349), .B(n9350), .Z(n9344) );
  AND U8969 ( .A(n1201), .B(n9351), .Z(n9350) );
  XOR U8970 ( .A(p_input[1697]), .B(n9349), .Z(n9351) );
  XOR U8971 ( .A(n9352), .B(n9353), .Z(n9349) );
  AND U8972 ( .A(n1205), .B(n9354), .Z(n9353) );
  XOR U8973 ( .A(n9355), .B(n9356), .Z(n9347) );
  AND U8974 ( .A(n1209), .B(n9354), .Z(n9356) );
  XNOR U8975 ( .A(n9355), .B(n9352), .Z(n9354) );
  XOR U8976 ( .A(n9357), .B(n9358), .Z(n9352) );
  AND U8977 ( .A(n1212), .B(n9359), .Z(n9358) );
  XOR U8978 ( .A(p_input[1713]), .B(n9357), .Z(n9359) );
  XOR U8979 ( .A(n9360), .B(n9361), .Z(n9357) );
  AND U8980 ( .A(n1216), .B(n9362), .Z(n9361) );
  XOR U8981 ( .A(n9363), .B(n9364), .Z(n9355) );
  AND U8982 ( .A(n1220), .B(n9362), .Z(n9364) );
  XNOR U8983 ( .A(n9363), .B(n9360), .Z(n9362) );
  XOR U8984 ( .A(n9365), .B(n9366), .Z(n9360) );
  AND U8985 ( .A(n1223), .B(n9367), .Z(n9366) );
  XOR U8986 ( .A(p_input[1729]), .B(n9365), .Z(n9367) );
  XOR U8987 ( .A(n9368), .B(n9369), .Z(n9365) );
  AND U8988 ( .A(n1227), .B(n9370), .Z(n9369) );
  XOR U8989 ( .A(n9371), .B(n9372), .Z(n9363) );
  AND U8990 ( .A(n1231), .B(n9370), .Z(n9372) );
  XNOR U8991 ( .A(n9371), .B(n9368), .Z(n9370) );
  XOR U8992 ( .A(n9373), .B(n9374), .Z(n9368) );
  AND U8993 ( .A(n1234), .B(n9375), .Z(n9374) );
  XOR U8994 ( .A(p_input[1745]), .B(n9373), .Z(n9375) );
  XOR U8995 ( .A(n9376), .B(n9377), .Z(n9373) );
  AND U8996 ( .A(n1238), .B(n9378), .Z(n9377) );
  XOR U8997 ( .A(n9379), .B(n9380), .Z(n9371) );
  AND U8998 ( .A(n1242), .B(n9378), .Z(n9380) );
  XNOR U8999 ( .A(n9379), .B(n9376), .Z(n9378) );
  XOR U9000 ( .A(n9381), .B(n9382), .Z(n9376) );
  AND U9001 ( .A(n1245), .B(n9383), .Z(n9382) );
  XOR U9002 ( .A(p_input[1761]), .B(n9381), .Z(n9383) );
  XOR U9003 ( .A(n9384), .B(n9385), .Z(n9381) );
  AND U9004 ( .A(n1249), .B(n9386), .Z(n9385) );
  XOR U9005 ( .A(n9387), .B(n9388), .Z(n9379) );
  AND U9006 ( .A(n1253), .B(n9386), .Z(n9388) );
  XNOR U9007 ( .A(n9387), .B(n9384), .Z(n9386) );
  XOR U9008 ( .A(n9389), .B(n9390), .Z(n9384) );
  AND U9009 ( .A(n1256), .B(n9391), .Z(n9390) );
  XOR U9010 ( .A(p_input[1777]), .B(n9389), .Z(n9391) );
  XOR U9011 ( .A(n9392), .B(n9393), .Z(n9389) );
  AND U9012 ( .A(n1260), .B(n9394), .Z(n9393) );
  XOR U9013 ( .A(n9395), .B(n9396), .Z(n9387) );
  AND U9014 ( .A(n1264), .B(n9394), .Z(n9396) );
  XNOR U9015 ( .A(n9395), .B(n9392), .Z(n9394) );
  XOR U9016 ( .A(n9397), .B(n9398), .Z(n9392) );
  AND U9017 ( .A(n1267), .B(n9399), .Z(n9398) );
  XOR U9018 ( .A(p_input[1793]), .B(n9397), .Z(n9399) );
  XOR U9019 ( .A(n9400), .B(n9401), .Z(n9397) );
  AND U9020 ( .A(n1271), .B(n9402), .Z(n9401) );
  XOR U9021 ( .A(n9403), .B(n9404), .Z(n9395) );
  AND U9022 ( .A(n1275), .B(n9402), .Z(n9404) );
  XNOR U9023 ( .A(n9403), .B(n9400), .Z(n9402) );
  XOR U9024 ( .A(n9405), .B(n9406), .Z(n9400) );
  AND U9025 ( .A(n1278), .B(n9407), .Z(n9406) );
  XOR U9026 ( .A(p_input[1809]), .B(n9405), .Z(n9407) );
  XOR U9027 ( .A(n9408), .B(n9409), .Z(n9405) );
  AND U9028 ( .A(n1282), .B(n9410), .Z(n9409) );
  XOR U9029 ( .A(n9411), .B(n9412), .Z(n9403) );
  AND U9030 ( .A(n1286), .B(n9410), .Z(n9412) );
  XNOR U9031 ( .A(n9411), .B(n9408), .Z(n9410) );
  XOR U9032 ( .A(n9413), .B(n9414), .Z(n9408) );
  AND U9033 ( .A(n1289), .B(n9415), .Z(n9414) );
  XOR U9034 ( .A(p_input[1825]), .B(n9413), .Z(n9415) );
  XOR U9035 ( .A(n9416), .B(n9417), .Z(n9413) );
  AND U9036 ( .A(n1293), .B(n9418), .Z(n9417) );
  XOR U9037 ( .A(n9419), .B(n9420), .Z(n9411) );
  AND U9038 ( .A(n1297), .B(n9418), .Z(n9420) );
  XNOR U9039 ( .A(n9419), .B(n9416), .Z(n9418) );
  XOR U9040 ( .A(n9421), .B(n9422), .Z(n9416) );
  AND U9041 ( .A(n1300), .B(n9423), .Z(n9422) );
  XOR U9042 ( .A(p_input[1841]), .B(n9421), .Z(n9423) );
  XOR U9043 ( .A(n9424), .B(n9425), .Z(n9421) );
  AND U9044 ( .A(n1304), .B(n9426), .Z(n9425) );
  XOR U9045 ( .A(n9427), .B(n9428), .Z(n9419) );
  AND U9046 ( .A(n1308), .B(n9426), .Z(n9428) );
  XNOR U9047 ( .A(n9427), .B(n9424), .Z(n9426) );
  XOR U9048 ( .A(n9429), .B(n9430), .Z(n9424) );
  AND U9049 ( .A(n1311), .B(n9431), .Z(n9430) );
  XOR U9050 ( .A(p_input[1857]), .B(n9429), .Z(n9431) );
  XOR U9051 ( .A(n9432), .B(n9433), .Z(n9429) );
  AND U9052 ( .A(n1315), .B(n9434), .Z(n9433) );
  XOR U9053 ( .A(n9435), .B(n9436), .Z(n9427) );
  AND U9054 ( .A(n1319), .B(n9434), .Z(n9436) );
  XNOR U9055 ( .A(n9435), .B(n9432), .Z(n9434) );
  XOR U9056 ( .A(n9437), .B(n9438), .Z(n9432) );
  AND U9057 ( .A(n1322), .B(n9439), .Z(n9438) );
  XOR U9058 ( .A(p_input[1873]), .B(n9437), .Z(n9439) );
  XOR U9059 ( .A(n9440), .B(n9441), .Z(n9437) );
  AND U9060 ( .A(n1326), .B(n9442), .Z(n9441) );
  XOR U9061 ( .A(n9443), .B(n9444), .Z(n9435) );
  AND U9062 ( .A(n1330), .B(n9442), .Z(n9444) );
  XNOR U9063 ( .A(n9443), .B(n9440), .Z(n9442) );
  XOR U9064 ( .A(n9445), .B(n9446), .Z(n9440) );
  AND U9065 ( .A(n1333), .B(n9447), .Z(n9446) );
  XOR U9066 ( .A(p_input[1889]), .B(n9445), .Z(n9447) );
  XOR U9067 ( .A(n9448), .B(n9449), .Z(n9445) );
  AND U9068 ( .A(n1337), .B(n9450), .Z(n9449) );
  XOR U9069 ( .A(n9451), .B(n9452), .Z(n9443) );
  AND U9070 ( .A(n1341), .B(n9450), .Z(n9452) );
  XNOR U9071 ( .A(n9451), .B(n9448), .Z(n9450) );
  XOR U9072 ( .A(n9453), .B(n9454), .Z(n9448) );
  AND U9073 ( .A(n1344), .B(n9455), .Z(n9454) );
  XOR U9074 ( .A(p_input[1905]), .B(n9453), .Z(n9455) );
  XOR U9075 ( .A(n9456), .B(n9457), .Z(n9453) );
  AND U9076 ( .A(n1348), .B(n9458), .Z(n9457) );
  XOR U9077 ( .A(n9459), .B(n9460), .Z(n9451) );
  AND U9078 ( .A(n1352), .B(n9458), .Z(n9460) );
  XNOR U9079 ( .A(n9459), .B(n9456), .Z(n9458) );
  XOR U9080 ( .A(n9461), .B(n9462), .Z(n9456) );
  AND U9081 ( .A(n1355), .B(n9463), .Z(n9462) );
  XOR U9082 ( .A(p_input[1921]), .B(n9461), .Z(n9463) );
  XOR U9083 ( .A(n9464), .B(n9465), .Z(n9461) );
  AND U9084 ( .A(n1359), .B(n9466), .Z(n9465) );
  XOR U9085 ( .A(n9467), .B(n9468), .Z(n9459) );
  AND U9086 ( .A(n1363), .B(n9466), .Z(n9468) );
  XNOR U9087 ( .A(n9467), .B(n9464), .Z(n9466) );
  XOR U9088 ( .A(n9469), .B(n9470), .Z(n9464) );
  AND U9089 ( .A(n1366), .B(n9471), .Z(n9470) );
  XOR U9090 ( .A(p_input[1937]), .B(n9469), .Z(n9471) );
  XOR U9091 ( .A(n9472), .B(n9473), .Z(n9469) );
  AND U9092 ( .A(n1370), .B(n9474), .Z(n9473) );
  XOR U9093 ( .A(n9475), .B(n9476), .Z(n9467) );
  AND U9094 ( .A(n1374), .B(n9474), .Z(n9476) );
  XNOR U9095 ( .A(n9475), .B(n9472), .Z(n9474) );
  XOR U9096 ( .A(n9477), .B(n9478), .Z(n9472) );
  AND U9097 ( .A(n1377), .B(n9479), .Z(n9478) );
  XOR U9098 ( .A(p_input[1953]), .B(n9477), .Z(n9479) );
  XOR U9099 ( .A(n9480), .B(n9481), .Z(n9477) );
  AND U9100 ( .A(n1381), .B(n9482), .Z(n9481) );
  XOR U9101 ( .A(n9483), .B(n9484), .Z(n9475) );
  AND U9102 ( .A(n1385), .B(n9482), .Z(n9484) );
  XNOR U9103 ( .A(n9483), .B(n9480), .Z(n9482) );
  XOR U9104 ( .A(n9485), .B(n9486), .Z(n9480) );
  AND U9105 ( .A(n1388), .B(n9487), .Z(n9486) );
  XOR U9106 ( .A(p_input[1969]), .B(n9485), .Z(n9487) );
  XOR U9107 ( .A(n9488), .B(n9489), .Z(n9485) );
  AND U9108 ( .A(n1392), .B(n9490), .Z(n9489) );
  XOR U9109 ( .A(n9491), .B(n9492), .Z(n9483) );
  AND U9110 ( .A(n1396), .B(n9490), .Z(n9492) );
  XNOR U9111 ( .A(n9491), .B(n9488), .Z(n9490) );
  XOR U9112 ( .A(n9493), .B(n9494), .Z(n9488) );
  AND U9113 ( .A(n1399), .B(n9495), .Z(n9494) );
  XOR U9114 ( .A(p_input[1985]), .B(n9493), .Z(n9495) );
  XOR U9115 ( .A(n9496), .B(n9497), .Z(n9493) );
  AND U9116 ( .A(n1403), .B(n9498), .Z(n9497) );
  XOR U9117 ( .A(n9499), .B(n9500), .Z(n9491) );
  AND U9118 ( .A(n1407), .B(n9498), .Z(n9500) );
  XNOR U9119 ( .A(n9499), .B(n9496), .Z(n9498) );
  XOR U9120 ( .A(n9501), .B(n9502), .Z(n9496) );
  AND U9121 ( .A(n1410), .B(n9503), .Z(n9502) );
  XOR U9122 ( .A(p_input[2001]), .B(n9501), .Z(n9503) );
  XNOR U9123 ( .A(n9504), .B(n9505), .Z(n9501) );
  AND U9124 ( .A(n1414), .B(n9506), .Z(n9505) );
  XNOR U9125 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n9507), .Z(n9499) );
  AND U9126 ( .A(n1417), .B(n9506), .Z(n9507) );
  XOR U9127 ( .A(n9508), .B(n9504), .Z(n9506) );
  XOR U9128 ( .A(n9509), .B(n9510), .Z(o[16]) );
  XOR U9129 ( .A(n15), .B(n9511), .Z(o[15]) );
  AND U9130 ( .A(n30), .B(n9512), .Z(n15) );
  XOR U9131 ( .A(n16), .B(n9511), .Z(n9512) );
  XOR U9132 ( .A(n9513), .B(n9514), .Z(n9511) );
  AND U9133 ( .A(n42), .B(n9515), .Z(n9514) );
  XOR U9134 ( .A(n9516), .B(n9517), .Z(n16) );
  AND U9135 ( .A(n34), .B(n9518), .Z(n9517) );
  XOR U9136 ( .A(p_input[15]), .B(n9516), .Z(n9518) );
  XNOR U9137 ( .A(n9519), .B(n9520), .Z(n9516) );
  AND U9138 ( .A(n38), .B(n9515), .Z(n9520) );
  XNOR U9139 ( .A(n9519), .B(n9513), .Z(n9515) );
  XOR U9140 ( .A(n9521), .B(n9522), .Z(n9513) );
  AND U9141 ( .A(n54), .B(n9523), .Z(n9522) );
  XNOR U9142 ( .A(n9524), .B(n9525), .Z(n9519) );
  AND U9143 ( .A(n46), .B(n9526), .Z(n9525) );
  XOR U9144 ( .A(p_input[31]), .B(n9524), .Z(n9526) );
  XNOR U9145 ( .A(n9527), .B(n9528), .Z(n9524) );
  AND U9146 ( .A(n50), .B(n9523), .Z(n9528) );
  XNOR U9147 ( .A(n9527), .B(n9521), .Z(n9523) );
  XOR U9148 ( .A(n9529), .B(n9530), .Z(n9521) );
  AND U9149 ( .A(n65), .B(n9531), .Z(n9530) );
  XNOR U9150 ( .A(n9532), .B(n9533), .Z(n9527) );
  AND U9151 ( .A(n57), .B(n9534), .Z(n9533) );
  XOR U9152 ( .A(p_input[47]), .B(n9532), .Z(n9534) );
  XNOR U9153 ( .A(n9535), .B(n9536), .Z(n9532) );
  AND U9154 ( .A(n61), .B(n9531), .Z(n9536) );
  XNOR U9155 ( .A(n9535), .B(n9529), .Z(n9531) );
  XOR U9156 ( .A(n9537), .B(n9538), .Z(n9529) );
  AND U9157 ( .A(n76), .B(n9539), .Z(n9538) );
  XNOR U9158 ( .A(n9540), .B(n9541), .Z(n9535) );
  AND U9159 ( .A(n68), .B(n9542), .Z(n9541) );
  XOR U9160 ( .A(p_input[63]), .B(n9540), .Z(n9542) );
  XNOR U9161 ( .A(n9543), .B(n9544), .Z(n9540) );
  AND U9162 ( .A(n72), .B(n9539), .Z(n9544) );
  XNOR U9163 ( .A(n9543), .B(n9537), .Z(n9539) );
  XOR U9164 ( .A(n9545), .B(n9546), .Z(n9537) );
  AND U9165 ( .A(n87), .B(n9547), .Z(n9546) );
  XNOR U9166 ( .A(n9548), .B(n9549), .Z(n9543) );
  AND U9167 ( .A(n79), .B(n9550), .Z(n9549) );
  XOR U9168 ( .A(p_input[79]), .B(n9548), .Z(n9550) );
  XNOR U9169 ( .A(n9551), .B(n9552), .Z(n9548) );
  AND U9170 ( .A(n83), .B(n9547), .Z(n9552) );
  XNOR U9171 ( .A(n9551), .B(n9545), .Z(n9547) );
  XOR U9172 ( .A(n9553), .B(n9554), .Z(n9545) );
  AND U9173 ( .A(n98), .B(n9555), .Z(n9554) );
  XNOR U9174 ( .A(n9556), .B(n9557), .Z(n9551) );
  AND U9175 ( .A(n90), .B(n9558), .Z(n9557) );
  XOR U9176 ( .A(p_input[95]), .B(n9556), .Z(n9558) );
  XNOR U9177 ( .A(n9559), .B(n9560), .Z(n9556) );
  AND U9178 ( .A(n94), .B(n9555), .Z(n9560) );
  XNOR U9179 ( .A(n9559), .B(n9553), .Z(n9555) );
  XOR U9180 ( .A(n9561), .B(n9562), .Z(n9553) );
  AND U9181 ( .A(n109), .B(n9563), .Z(n9562) );
  XNOR U9182 ( .A(n9564), .B(n9565), .Z(n9559) );
  AND U9183 ( .A(n101), .B(n9566), .Z(n9565) );
  XOR U9184 ( .A(p_input[111]), .B(n9564), .Z(n9566) );
  XNOR U9185 ( .A(n9567), .B(n9568), .Z(n9564) );
  AND U9186 ( .A(n105), .B(n9563), .Z(n9568) );
  XNOR U9187 ( .A(n9567), .B(n9561), .Z(n9563) );
  XOR U9188 ( .A(n9569), .B(n9570), .Z(n9561) );
  AND U9189 ( .A(n120), .B(n9571), .Z(n9570) );
  XNOR U9190 ( .A(n9572), .B(n9573), .Z(n9567) );
  AND U9191 ( .A(n112), .B(n9574), .Z(n9573) );
  XOR U9192 ( .A(p_input[127]), .B(n9572), .Z(n9574) );
  XNOR U9193 ( .A(n9575), .B(n9576), .Z(n9572) );
  AND U9194 ( .A(n116), .B(n9571), .Z(n9576) );
  XNOR U9195 ( .A(n9575), .B(n9569), .Z(n9571) );
  XOR U9196 ( .A(n9577), .B(n9578), .Z(n9569) );
  AND U9197 ( .A(n131), .B(n9579), .Z(n9578) );
  XNOR U9198 ( .A(n9580), .B(n9581), .Z(n9575) );
  AND U9199 ( .A(n123), .B(n9582), .Z(n9581) );
  XOR U9200 ( .A(p_input[143]), .B(n9580), .Z(n9582) );
  XNOR U9201 ( .A(n9583), .B(n9584), .Z(n9580) );
  AND U9202 ( .A(n127), .B(n9579), .Z(n9584) );
  XNOR U9203 ( .A(n9583), .B(n9577), .Z(n9579) );
  XOR U9204 ( .A(n9585), .B(n9586), .Z(n9577) );
  AND U9205 ( .A(n142), .B(n9587), .Z(n9586) );
  XNOR U9206 ( .A(n9588), .B(n9589), .Z(n9583) );
  AND U9207 ( .A(n134), .B(n9590), .Z(n9589) );
  XOR U9208 ( .A(p_input[159]), .B(n9588), .Z(n9590) );
  XNOR U9209 ( .A(n9591), .B(n9592), .Z(n9588) );
  AND U9210 ( .A(n138), .B(n9587), .Z(n9592) );
  XNOR U9211 ( .A(n9591), .B(n9585), .Z(n9587) );
  XOR U9212 ( .A(n9593), .B(n9594), .Z(n9585) );
  AND U9213 ( .A(n153), .B(n9595), .Z(n9594) );
  XNOR U9214 ( .A(n9596), .B(n9597), .Z(n9591) );
  AND U9215 ( .A(n145), .B(n9598), .Z(n9597) );
  XOR U9216 ( .A(p_input[175]), .B(n9596), .Z(n9598) );
  XNOR U9217 ( .A(n9599), .B(n9600), .Z(n9596) );
  AND U9218 ( .A(n149), .B(n9595), .Z(n9600) );
  XNOR U9219 ( .A(n9599), .B(n9593), .Z(n9595) );
  XOR U9220 ( .A(n9601), .B(n9602), .Z(n9593) );
  AND U9221 ( .A(n164), .B(n9603), .Z(n9602) );
  XNOR U9222 ( .A(n9604), .B(n9605), .Z(n9599) );
  AND U9223 ( .A(n156), .B(n9606), .Z(n9605) );
  XOR U9224 ( .A(p_input[191]), .B(n9604), .Z(n9606) );
  XNOR U9225 ( .A(n9607), .B(n9608), .Z(n9604) );
  AND U9226 ( .A(n160), .B(n9603), .Z(n9608) );
  XNOR U9227 ( .A(n9607), .B(n9601), .Z(n9603) );
  XOR U9228 ( .A(n9609), .B(n9610), .Z(n9601) );
  AND U9229 ( .A(n175), .B(n9611), .Z(n9610) );
  XNOR U9230 ( .A(n9612), .B(n9613), .Z(n9607) );
  AND U9231 ( .A(n167), .B(n9614), .Z(n9613) );
  XOR U9232 ( .A(p_input[207]), .B(n9612), .Z(n9614) );
  XNOR U9233 ( .A(n9615), .B(n9616), .Z(n9612) );
  AND U9234 ( .A(n171), .B(n9611), .Z(n9616) );
  XNOR U9235 ( .A(n9615), .B(n9609), .Z(n9611) );
  XOR U9236 ( .A(n9617), .B(n9618), .Z(n9609) );
  AND U9237 ( .A(n186), .B(n9619), .Z(n9618) );
  XNOR U9238 ( .A(n9620), .B(n9621), .Z(n9615) );
  AND U9239 ( .A(n178), .B(n9622), .Z(n9621) );
  XOR U9240 ( .A(p_input[223]), .B(n9620), .Z(n9622) );
  XNOR U9241 ( .A(n9623), .B(n9624), .Z(n9620) );
  AND U9242 ( .A(n182), .B(n9619), .Z(n9624) );
  XNOR U9243 ( .A(n9623), .B(n9617), .Z(n9619) );
  XOR U9244 ( .A(n9625), .B(n9626), .Z(n9617) );
  AND U9245 ( .A(n197), .B(n9627), .Z(n9626) );
  XNOR U9246 ( .A(n9628), .B(n9629), .Z(n9623) );
  AND U9247 ( .A(n189), .B(n9630), .Z(n9629) );
  XOR U9248 ( .A(p_input[239]), .B(n9628), .Z(n9630) );
  XNOR U9249 ( .A(n9631), .B(n9632), .Z(n9628) );
  AND U9250 ( .A(n193), .B(n9627), .Z(n9632) );
  XNOR U9251 ( .A(n9631), .B(n9625), .Z(n9627) );
  XOR U9252 ( .A(n9633), .B(n9634), .Z(n9625) );
  AND U9253 ( .A(n208), .B(n9635), .Z(n9634) );
  XNOR U9254 ( .A(n9636), .B(n9637), .Z(n9631) );
  AND U9255 ( .A(n200), .B(n9638), .Z(n9637) );
  XOR U9256 ( .A(p_input[255]), .B(n9636), .Z(n9638) );
  XNOR U9257 ( .A(n9639), .B(n9640), .Z(n9636) );
  AND U9258 ( .A(n204), .B(n9635), .Z(n9640) );
  XNOR U9259 ( .A(n9639), .B(n9633), .Z(n9635) );
  XOR U9260 ( .A(n9641), .B(n9642), .Z(n9633) );
  AND U9261 ( .A(n219), .B(n9643), .Z(n9642) );
  XNOR U9262 ( .A(n9644), .B(n9645), .Z(n9639) );
  AND U9263 ( .A(n211), .B(n9646), .Z(n9645) );
  XOR U9264 ( .A(p_input[271]), .B(n9644), .Z(n9646) );
  XNOR U9265 ( .A(n9647), .B(n9648), .Z(n9644) );
  AND U9266 ( .A(n215), .B(n9643), .Z(n9648) );
  XNOR U9267 ( .A(n9647), .B(n9641), .Z(n9643) );
  XOR U9268 ( .A(n9649), .B(n9650), .Z(n9641) );
  AND U9269 ( .A(n230), .B(n9651), .Z(n9650) );
  XNOR U9270 ( .A(n9652), .B(n9653), .Z(n9647) );
  AND U9271 ( .A(n222), .B(n9654), .Z(n9653) );
  XOR U9272 ( .A(p_input[287]), .B(n9652), .Z(n9654) );
  XNOR U9273 ( .A(n9655), .B(n9656), .Z(n9652) );
  AND U9274 ( .A(n226), .B(n9651), .Z(n9656) );
  XNOR U9275 ( .A(n9655), .B(n9649), .Z(n9651) );
  XOR U9276 ( .A(n9657), .B(n9658), .Z(n9649) );
  AND U9277 ( .A(n241), .B(n9659), .Z(n9658) );
  XNOR U9278 ( .A(n9660), .B(n9661), .Z(n9655) );
  AND U9279 ( .A(n233), .B(n9662), .Z(n9661) );
  XOR U9280 ( .A(p_input[303]), .B(n9660), .Z(n9662) );
  XNOR U9281 ( .A(n9663), .B(n9664), .Z(n9660) );
  AND U9282 ( .A(n237), .B(n9659), .Z(n9664) );
  XNOR U9283 ( .A(n9663), .B(n9657), .Z(n9659) );
  XOR U9284 ( .A(n9665), .B(n9666), .Z(n9657) );
  AND U9285 ( .A(n252), .B(n9667), .Z(n9666) );
  XNOR U9286 ( .A(n9668), .B(n9669), .Z(n9663) );
  AND U9287 ( .A(n244), .B(n9670), .Z(n9669) );
  XOR U9288 ( .A(p_input[319]), .B(n9668), .Z(n9670) );
  XNOR U9289 ( .A(n9671), .B(n9672), .Z(n9668) );
  AND U9290 ( .A(n248), .B(n9667), .Z(n9672) );
  XNOR U9291 ( .A(n9671), .B(n9665), .Z(n9667) );
  XOR U9292 ( .A(n9673), .B(n9674), .Z(n9665) );
  AND U9293 ( .A(n263), .B(n9675), .Z(n9674) );
  XNOR U9294 ( .A(n9676), .B(n9677), .Z(n9671) );
  AND U9295 ( .A(n255), .B(n9678), .Z(n9677) );
  XOR U9296 ( .A(p_input[335]), .B(n9676), .Z(n9678) );
  XNOR U9297 ( .A(n9679), .B(n9680), .Z(n9676) );
  AND U9298 ( .A(n259), .B(n9675), .Z(n9680) );
  XNOR U9299 ( .A(n9679), .B(n9673), .Z(n9675) );
  XOR U9300 ( .A(n9681), .B(n9682), .Z(n9673) );
  AND U9301 ( .A(n274), .B(n9683), .Z(n9682) );
  XNOR U9302 ( .A(n9684), .B(n9685), .Z(n9679) );
  AND U9303 ( .A(n266), .B(n9686), .Z(n9685) );
  XOR U9304 ( .A(p_input[351]), .B(n9684), .Z(n9686) );
  XNOR U9305 ( .A(n9687), .B(n9688), .Z(n9684) );
  AND U9306 ( .A(n270), .B(n9683), .Z(n9688) );
  XNOR U9307 ( .A(n9687), .B(n9681), .Z(n9683) );
  XOR U9308 ( .A(n9689), .B(n9690), .Z(n9681) );
  AND U9309 ( .A(n285), .B(n9691), .Z(n9690) );
  XNOR U9310 ( .A(n9692), .B(n9693), .Z(n9687) );
  AND U9311 ( .A(n277), .B(n9694), .Z(n9693) );
  XOR U9312 ( .A(p_input[367]), .B(n9692), .Z(n9694) );
  XNOR U9313 ( .A(n9695), .B(n9696), .Z(n9692) );
  AND U9314 ( .A(n281), .B(n9691), .Z(n9696) );
  XNOR U9315 ( .A(n9695), .B(n9689), .Z(n9691) );
  XOR U9316 ( .A(n9697), .B(n9698), .Z(n9689) );
  AND U9317 ( .A(n296), .B(n9699), .Z(n9698) );
  XNOR U9318 ( .A(n9700), .B(n9701), .Z(n9695) );
  AND U9319 ( .A(n288), .B(n9702), .Z(n9701) );
  XOR U9320 ( .A(p_input[383]), .B(n9700), .Z(n9702) );
  XNOR U9321 ( .A(n9703), .B(n9704), .Z(n9700) );
  AND U9322 ( .A(n292), .B(n9699), .Z(n9704) );
  XNOR U9323 ( .A(n9703), .B(n9697), .Z(n9699) );
  XOR U9324 ( .A(n9705), .B(n9706), .Z(n9697) );
  AND U9325 ( .A(n307), .B(n9707), .Z(n9706) );
  XNOR U9326 ( .A(n9708), .B(n9709), .Z(n9703) );
  AND U9327 ( .A(n299), .B(n9710), .Z(n9709) );
  XOR U9328 ( .A(p_input[399]), .B(n9708), .Z(n9710) );
  XNOR U9329 ( .A(n9711), .B(n9712), .Z(n9708) );
  AND U9330 ( .A(n303), .B(n9707), .Z(n9712) );
  XNOR U9331 ( .A(n9711), .B(n9705), .Z(n9707) );
  XOR U9332 ( .A(n9713), .B(n9714), .Z(n9705) );
  AND U9333 ( .A(n318), .B(n9715), .Z(n9714) );
  XNOR U9334 ( .A(n9716), .B(n9717), .Z(n9711) );
  AND U9335 ( .A(n310), .B(n9718), .Z(n9717) );
  XOR U9336 ( .A(p_input[415]), .B(n9716), .Z(n9718) );
  XNOR U9337 ( .A(n9719), .B(n9720), .Z(n9716) );
  AND U9338 ( .A(n314), .B(n9715), .Z(n9720) );
  XNOR U9339 ( .A(n9719), .B(n9713), .Z(n9715) );
  XOR U9340 ( .A(n9721), .B(n9722), .Z(n9713) );
  AND U9341 ( .A(n329), .B(n9723), .Z(n9722) );
  XNOR U9342 ( .A(n9724), .B(n9725), .Z(n9719) );
  AND U9343 ( .A(n321), .B(n9726), .Z(n9725) );
  XOR U9344 ( .A(p_input[431]), .B(n9724), .Z(n9726) );
  XNOR U9345 ( .A(n9727), .B(n9728), .Z(n9724) );
  AND U9346 ( .A(n325), .B(n9723), .Z(n9728) );
  XNOR U9347 ( .A(n9727), .B(n9721), .Z(n9723) );
  XOR U9348 ( .A(n9729), .B(n9730), .Z(n9721) );
  AND U9349 ( .A(n340), .B(n9731), .Z(n9730) );
  XNOR U9350 ( .A(n9732), .B(n9733), .Z(n9727) );
  AND U9351 ( .A(n332), .B(n9734), .Z(n9733) );
  XOR U9352 ( .A(p_input[447]), .B(n9732), .Z(n9734) );
  XNOR U9353 ( .A(n9735), .B(n9736), .Z(n9732) );
  AND U9354 ( .A(n336), .B(n9731), .Z(n9736) );
  XNOR U9355 ( .A(n9735), .B(n9729), .Z(n9731) );
  XOR U9356 ( .A(n9737), .B(n9738), .Z(n9729) );
  AND U9357 ( .A(n351), .B(n9739), .Z(n9738) );
  XNOR U9358 ( .A(n9740), .B(n9741), .Z(n9735) );
  AND U9359 ( .A(n343), .B(n9742), .Z(n9741) );
  XOR U9360 ( .A(p_input[463]), .B(n9740), .Z(n9742) );
  XNOR U9361 ( .A(n9743), .B(n9744), .Z(n9740) );
  AND U9362 ( .A(n347), .B(n9739), .Z(n9744) );
  XNOR U9363 ( .A(n9743), .B(n9737), .Z(n9739) );
  XOR U9364 ( .A(n9745), .B(n9746), .Z(n9737) );
  AND U9365 ( .A(n362), .B(n9747), .Z(n9746) );
  XNOR U9366 ( .A(n9748), .B(n9749), .Z(n9743) );
  AND U9367 ( .A(n354), .B(n9750), .Z(n9749) );
  XOR U9368 ( .A(p_input[479]), .B(n9748), .Z(n9750) );
  XNOR U9369 ( .A(n9751), .B(n9752), .Z(n9748) );
  AND U9370 ( .A(n358), .B(n9747), .Z(n9752) );
  XNOR U9371 ( .A(n9751), .B(n9745), .Z(n9747) );
  XOR U9372 ( .A(n9753), .B(n9754), .Z(n9745) );
  AND U9373 ( .A(n373), .B(n9755), .Z(n9754) );
  XNOR U9374 ( .A(n9756), .B(n9757), .Z(n9751) );
  AND U9375 ( .A(n365), .B(n9758), .Z(n9757) );
  XOR U9376 ( .A(p_input[495]), .B(n9756), .Z(n9758) );
  XNOR U9377 ( .A(n9759), .B(n9760), .Z(n9756) );
  AND U9378 ( .A(n369), .B(n9755), .Z(n9760) );
  XNOR U9379 ( .A(n9759), .B(n9753), .Z(n9755) );
  XOR U9380 ( .A(n9761), .B(n9762), .Z(n9753) );
  AND U9381 ( .A(n384), .B(n9763), .Z(n9762) );
  XNOR U9382 ( .A(n9764), .B(n9765), .Z(n9759) );
  AND U9383 ( .A(n376), .B(n9766), .Z(n9765) );
  XOR U9384 ( .A(p_input[511]), .B(n9764), .Z(n9766) );
  XNOR U9385 ( .A(n9767), .B(n9768), .Z(n9764) );
  AND U9386 ( .A(n380), .B(n9763), .Z(n9768) );
  XNOR U9387 ( .A(n9767), .B(n9761), .Z(n9763) );
  XOR U9388 ( .A(n9769), .B(n9770), .Z(n9761) );
  AND U9389 ( .A(n395), .B(n9771), .Z(n9770) );
  XNOR U9390 ( .A(n9772), .B(n9773), .Z(n9767) );
  AND U9391 ( .A(n387), .B(n9774), .Z(n9773) );
  XOR U9392 ( .A(p_input[527]), .B(n9772), .Z(n9774) );
  XNOR U9393 ( .A(n9775), .B(n9776), .Z(n9772) );
  AND U9394 ( .A(n391), .B(n9771), .Z(n9776) );
  XNOR U9395 ( .A(n9775), .B(n9769), .Z(n9771) );
  XOR U9396 ( .A(n9777), .B(n9778), .Z(n9769) );
  AND U9397 ( .A(n406), .B(n9779), .Z(n9778) );
  XNOR U9398 ( .A(n9780), .B(n9781), .Z(n9775) );
  AND U9399 ( .A(n398), .B(n9782), .Z(n9781) );
  XOR U9400 ( .A(p_input[543]), .B(n9780), .Z(n9782) );
  XNOR U9401 ( .A(n9783), .B(n9784), .Z(n9780) );
  AND U9402 ( .A(n402), .B(n9779), .Z(n9784) );
  XNOR U9403 ( .A(n9783), .B(n9777), .Z(n9779) );
  XOR U9404 ( .A(n9785), .B(n9786), .Z(n9777) );
  AND U9405 ( .A(n417), .B(n9787), .Z(n9786) );
  XNOR U9406 ( .A(n9788), .B(n9789), .Z(n9783) );
  AND U9407 ( .A(n409), .B(n9790), .Z(n9789) );
  XOR U9408 ( .A(p_input[559]), .B(n9788), .Z(n9790) );
  XNOR U9409 ( .A(n9791), .B(n9792), .Z(n9788) );
  AND U9410 ( .A(n413), .B(n9787), .Z(n9792) );
  XNOR U9411 ( .A(n9791), .B(n9785), .Z(n9787) );
  XOR U9412 ( .A(n9793), .B(n9794), .Z(n9785) );
  AND U9413 ( .A(n428), .B(n9795), .Z(n9794) );
  XNOR U9414 ( .A(n9796), .B(n9797), .Z(n9791) );
  AND U9415 ( .A(n420), .B(n9798), .Z(n9797) );
  XOR U9416 ( .A(p_input[575]), .B(n9796), .Z(n9798) );
  XNOR U9417 ( .A(n9799), .B(n9800), .Z(n9796) );
  AND U9418 ( .A(n424), .B(n9795), .Z(n9800) );
  XNOR U9419 ( .A(n9799), .B(n9793), .Z(n9795) );
  XOR U9420 ( .A(n9801), .B(n9802), .Z(n9793) );
  AND U9421 ( .A(n439), .B(n9803), .Z(n9802) );
  XNOR U9422 ( .A(n9804), .B(n9805), .Z(n9799) );
  AND U9423 ( .A(n431), .B(n9806), .Z(n9805) );
  XOR U9424 ( .A(p_input[591]), .B(n9804), .Z(n9806) );
  XNOR U9425 ( .A(n9807), .B(n9808), .Z(n9804) );
  AND U9426 ( .A(n435), .B(n9803), .Z(n9808) );
  XNOR U9427 ( .A(n9807), .B(n9801), .Z(n9803) );
  XOR U9428 ( .A(n9809), .B(n9810), .Z(n9801) );
  AND U9429 ( .A(n450), .B(n9811), .Z(n9810) );
  XNOR U9430 ( .A(n9812), .B(n9813), .Z(n9807) );
  AND U9431 ( .A(n442), .B(n9814), .Z(n9813) );
  XOR U9432 ( .A(p_input[607]), .B(n9812), .Z(n9814) );
  XNOR U9433 ( .A(n9815), .B(n9816), .Z(n9812) );
  AND U9434 ( .A(n446), .B(n9811), .Z(n9816) );
  XNOR U9435 ( .A(n9815), .B(n9809), .Z(n9811) );
  XOR U9436 ( .A(n9817), .B(n9818), .Z(n9809) );
  AND U9437 ( .A(n461), .B(n9819), .Z(n9818) );
  XNOR U9438 ( .A(n9820), .B(n9821), .Z(n9815) );
  AND U9439 ( .A(n453), .B(n9822), .Z(n9821) );
  XOR U9440 ( .A(p_input[623]), .B(n9820), .Z(n9822) );
  XNOR U9441 ( .A(n9823), .B(n9824), .Z(n9820) );
  AND U9442 ( .A(n457), .B(n9819), .Z(n9824) );
  XNOR U9443 ( .A(n9823), .B(n9817), .Z(n9819) );
  XOR U9444 ( .A(n9825), .B(n9826), .Z(n9817) );
  AND U9445 ( .A(n472), .B(n9827), .Z(n9826) );
  XNOR U9446 ( .A(n9828), .B(n9829), .Z(n9823) );
  AND U9447 ( .A(n464), .B(n9830), .Z(n9829) );
  XOR U9448 ( .A(p_input[639]), .B(n9828), .Z(n9830) );
  XNOR U9449 ( .A(n9831), .B(n9832), .Z(n9828) );
  AND U9450 ( .A(n468), .B(n9827), .Z(n9832) );
  XNOR U9451 ( .A(n9831), .B(n9825), .Z(n9827) );
  XOR U9452 ( .A(n9833), .B(n9834), .Z(n9825) );
  AND U9453 ( .A(n483), .B(n9835), .Z(n9834) );
  XNOR U9454 ( .A(n9836), .B(n9837), .Z(n9831) );
  AND U9455 ( .A(n475), .B(n9838), .Z(n9837) );
  XOR U9456 ( .A(p_input[655]), .B(n9836), .Z(n9838) );
  XNOR U9457 ( .A(n9839), .B(n9840), .Z(n9836) );
  AND U9458 ( .A(n479), .B(n9835), .Z(n9840) );
  XNOR U9459 ( .A(n9839), .B(n9833), .Z(n9835) );
  XOR U9460 ( .A(n9841), .B(n9842), .Z(n9833) );
  AND U9461 ( .A(n494), .B(n9843), .Z(n9842) );
  XNOR U9462 ( .A(n9844), .B(n9845), .Z(n9839) );
  AND U9463 ( .A(n486), .B(n9846), .Z(n9845) );
  XOR U9464 ( .A(p_input[671]), .B(n9844), .Z(n9846) );
  XNOR U9465 ( .A(n9847), .B(n9848), .Z(n9844) );
  AND U9466 ( .A(n490), .B(n9843), .Z(n9848) );
  XNOR U9467 ( .A(n9847), .B(n9841), .Z(n9843) );
  XOR U9468 ( .A(n9849), .B(n9850), .Z(n9841) );
  AND U9469 ( .A(n505), .B(n9851), .Z(n9850) );
  XNOR U9470 ( .A(n9852), .B(n9853), .Z(n9847) );
  AND U9471 ( .A(n497), .B(n9854), .Z(n9853) );
  XOR U9472 ( .A(p_input[687]), .B(n9852), .Z(n9854) );
  XNOR U9473 ( .A(n9855), .B(n9856), .Z(n9852) );
  AND U9474 ( .A(n501), .B(n9851), .Z(n9856) );
  XNOR U9475 ( .A(n9855), .B(n9849), .Z(n9851) );
  XOR U9476 ( .A(n9857), .B(n9858), .Z(n9849) );
  AND U9477 ( .A(n516), .B(n9859), .Z(n9858) );
  XNOR U9478 ( .A(n9860), .B(n9861), .Z(n9855) );
  AND U9479 ( .A(n508), .B(n9862), .Z(n9861) );
  XOR U9480 ( .A(p_input[703]), .B(n9860), .Z(n9862) );
  XNOR U9481 ( .A(n9863), .B(n9864), .Z(n9860) );
  AND U9482 ( .A(n512), .B(n9859), .Z(n9864) );
  XNOR U9483 ( .A(n9863), .B(n9857), .Z(n9859) );
  XOR U9484 ( .A(n9865), .B(n9866), .Z(n9857) );
  AND U9485 ( .A(n527), .B(n9867), .Z(n9866) );
  XNOR U9486 ( .A(n9868), .B(n9869), .Z(n9863) );
  AND U9487 ( .A(n519), .B(n9870), .Z(n9869) );
  XOR U9488 ( .A(p_input[719]), .B(n9868), .Z(n9870) );
  XNOR U9489 ( .A(n9871), .B(n9872), .Z(n9868) );
  AND U9490 ( .A(n523), .B(n9867), .Z(n9872) );
  XNOR U9491 ( .A(n9871), .B(n9865), .Z(n9867) );
  XOR U9492 ( .A(n9873), .B(n9874), .Z(n9865) );
  AND U9493 ( .A(n538), .B(n9875), .Z(n9874) );
  XNOR U9494 ( .A(n9876), .B(n9877), .Z(n9871) );
  AND U9495 ( .A(n530), .B(n9878), .Z(n9877) );
  XOR U9496 ( .A(p_input[735]), .B(n9876), .Z(n9878) );
  XNOR U9497 ( .A(n9879), .B(n9880), .Z(n9876) );
  AND U9498 ( .A(n534), .B(n9875), .Z(n9880) );
  XNOR U9499 ( .A(n9879), .B(n9873), .Z(n9875) );
  XOR U9500 ( .A(n9881), .B(n9882), .Z(n9873) );
  AND U9501 ( .A(n549), .B(n9883), .Z(n9882) );
  XNOR U9502 ( .A(n9884), .B(n9885), .Z(n9879) );
  AND U9503 ( .A(n541), .B(n9886), .Z(n9885) );
  XOR U9504 ( .A(p_input[751]), .B(n9884), .Z(n9886) );
  XNOR U9505 ( .A(n9887), .B(n9888), .Z(n9884) );
  AND U9506 ( .A(n545), .B(n9883), .Z(n9888) );
  XNOR U9507 ( .A(n9887), .B(n9881), .Z(n9883) );
  XOR U9508 ( .A(n9889), .B(n9890), .Z(n9881) );
  AND U9509 ( .A(n560), .B(n9891), .Z(n9890) );
  XNOR U9510 ( .A(n9892), .B(n9893), .Z(n9887) );
  AND U9511 ( .A(n552), .B(n9894), .Z(n9893) );
  XOR U9512 ( .A(p_input[767]), .B(n9892), .Z(n9894) );
  XNOR U9513 ( .A(n9895), .B(n9896), .Z(n9892) );
  AND U9514 ( .A(n556), .B(n9891), .Z(n9896) );
  XNOR U9515 ( .A(n9895), .B(n9889), .Z(n9891) );
  XOR U9516 ( .A(n9897), .B(n9898), .Z(n9889) );
  AND U9517 ( .A(n571), .B(n9899), .Z(n9898) );
  XNOR U9518 ( .A(n9900), .B(n9901), .Z(n9895) );
  AND U9519 ( .A(n563), .B(n9902), .Z(n9901) );
  XOR U9520 ( .A(p_input[783]), .B(n9900), .Z(n9902) );
  XNOR U9521 ( .A(n9903), .B(n9904), .Z(n9900) );
  AND U9522 ( .A(n567), .B(n9899), .Z(n9904) );
  XNOR U9523 ( .A(n9903), .B(n9897), .Z(n9899) );
  XOR U9524 ( .A(n9905), .B(n9906), .Z(n9897) );
  AND U9525 ( .A(n582), .B(n9907), .Z(n9906) );
  XNOR U9526 ( .A(n9908), .B(n9909), .Z(n9903) );
  AND U9527 ( .A(n574), .B(n9910), .Z(n9909) );
  XOR U9528 ( .A(p_input[799]), .B(n9908), .Z(n9910) );
  XNOR U9529 ( .A(n9911), .B(n9912), .Z(n9908) );
  AND U9530 ( .A(n578), .B(n9907), .Z(n9912) );
  XNOR U9531 ( .A(n9911), .B(n9905), .Z(n9907) );
  XOR U9532 ( .A(n9913), .B(n9914), .Z(n9905) );
  AND U9533 ( .A(n593), .B(n9915), .Z(n9914) );
  XNOR U9534 ( .A(n9916), .B(n9917), .Z(n9911) );
  AND U9535 ( .A(n585), .B(n9918), .Z(n9917) );
  XOR U9536 ( .A(p_input[815]), .B(n9916), .Z(n9918) );
  XNOR U9537 ( .A(n9919), .B(n9920), .Z(n9916) );
  AND U9538 ( .A(n589), .B(n9915), .Z(n9920) );
  XNOR U9539 ( .A(n9919), .B(n9913), .Z(n9915) );
  XOR U9540 ( .A(n9921), .B(n9922), .Z(n9913) );
  AND U9541 ( .A(n604), .B(n9923), .Z(n9922) );
  XNOR U9542 ( .A(n9924), .B(n9925), .Z(n9919) );
  AND U9543 ( .A(n596), .B(n9926), .Z(n9925) );
  XOR U9544 ( .A(p_input[831]), .B(n9924), .Z(n9926) );
  XNOR U9545 ( .A(n9927), .B(n9928), .Z(n9924) );
  AND U9546 ( .A(n600), .B(n9923), .Z(n9928) );
  XNOR U9547 ( .A(n9927), .B(n9921), .Z(n9923) );
  XOR U9548 ( .A(n9929), .B(n9930), .Z(n9921) );
  AND U9549 ( .A(n615), .B(n9931), .Z(n9930) );
  XNOR U9550 ( .A(n9932), .B(n9933), .Z(n9927) );
  AND U9551 ( .A(n607), .B(n9934), .Z(n9933) );
  XOR U9552 ( .A(p_input[847]), .B(n9932), .Z(n9934) );
  XNOR U9553 ( .A(n9935), .B(n9936), .Z(n9932) );
  AND U9554 ( .A(n611), .B(n9931), .Z(n9936) );
  XNOR U9555 ( .A(n9935), .B(n9929), .Z(n9931) );
  XOR U9556 ( .A(n9937), .B(n9938), .Z(n9929) );
  AND U9557 ( .A(n626), .B(n9939), .Z(n9938) );
  XNOR U9558 ( .A(n9940), .B(n9941), .Z(n9935) );
  AND U9559 ( .A(n618), .B(n9942), .Z(n9941) );
  XOR U9560 ( .A(p_input[863]), .B(n9940), .Z(n9942) );
  XNOR U9561 ( .A(n9943), .B(n9944), .Z(n9940) );
  AND U9562 ( .A(n622), .B(n9939), .Z(n9944) );
  XNOR U9563 ( .A(n9943), .B(n9937), .Z(n9939) );
  XOR U9564 ( .A(n9945), .B(n9946), .Z(n9937) );
  AND U9565 ( .A(n637), .B(n9947), .Z(n9946) );
  XNOR U9566 ( .A(n9948), .B(n9949), .Z(n9943) );
  AND U9567 ( .A(n629), .B(n9950), .Z(n9949) );
  XOR U9568 ( .A(p_input[879]), .B(n9948), .Z(n9950) );
  XNOR U9569 ( .A(n9951), .B(n9952), .Z(n9948) );
  AND U9570 ( .A(n633), .B(n9947), .Z(n9952) );
  XNOR U9571 ( .A(n9951), .B(n9945), .Z(n9947) );
  XOR U9572 ( .A(n9953), .B(n9954), .Z(n9945) );
  AND U9573 ( .A(n648), .B(n9955), .Z(n9954) );
  XNOR U9574 ( .A(n9956), .B(n9957), .Z(n9951) );
  AND U9575 ( .A(n640), .B(n9958), .Z(n9957) );
  XOR U9576 ( .A(p_input[895]), .B(n9956), .Z(n9958) );
  XNOR U9577 ( .A(n9959), .B(n9960), .Z(n9956) );
  AND U9578 ( .A(n644), .B(n9955), .Z(n9960) );
  XNOR U9579 ( .A(n9959), .B(n9953), .Z(n9955) );
  XOR U9580 ( .A(n9961), .B(n9962), .Z(n9953) );
  AND U9581 ( .A(n659), .B(n9963), .Z(n9962) );
  XNOR U9582 ( .A(n9964), .B(n9965), .Z(n9959) );
  AND U9583 ( .A(n651), .B(n9966), .Z(n9965) );
  XOR U9584 ( .A(p_input[911]), .B(n9964), .Z(n9966) );
  XNOR U9585 ( .A(n9967), .B(n9968), .Z(n9964) );
  AND U9586 ( .A(n655), .B(n9963), .Z(n9968) );
  XNOR U9587 ( .A(n9967), .B(n9961), .Z(n9963) );
  XOR U9588 ( .A(n9969), .B(n9970), .Z(n9961) );
  AND U9589 ( .A(n670), .B(n9971), .Z(n9970) );
  XNOR U9590 ( .A(n9972), .B(n9973), .Z(n9967) );
  AND U9591 ( .A(n662), .B(n9974), .Z(n9973) );
  XOR U9592 ( .A(p_input[927]), .B(n9972), .Z(n9974) );
  XNOR U9593 ( .A(n9975), .B(n9976), .Z(n9972) );
  AND U9594 ( .A(n666), .B(n9971), .Z(n9976) );
  XNOR U9595 ( .A(n9975), .B(n9969), .Z(n9971) );
  XOR U9596 ( .A(n9977), .B(n9978), .Z(n9969) );
  AND U9597 ( .A(n681), .B(n9979), .Z(n9978) );
  XNOR U9598 ( .A(n9980), .B(n9981), .Z(n9975) );
  AND U9599 ( .A(n673), .B(n9982), .Z(n9981) );
  XOR U9600 ( .A(p_input[943]), .B(n9980), .Z(n9982) );
  XNOR U9601 ( .A(n9983), .B(n9984), .Z(n9980) );
  AND U9602 ( .A(n677), .B(n9979), .Z(n9984) );
  XNOR U9603 ( .A(n9983), .B(n9977), .Z(n9979) );
  XOR U9604 ( .A(n9985), .B(n9986), .Z(n9977) );
  AND U9605 ( .A(n692), .B(n9987), .Z(n9986) );
  XNOR U9606 ( .A(n9988), .B(n9989), .Z(n9983) );
  AND U9607 ( .A(n684), .B(n9990), .Z(n9989) );
  XOR U9608 ( .A(p_input[959]), .B(n9988), .Z(n9990) );
  XNOR U9609 ( .A(n9991), .B(n9992), .Z(n9988) );
  AND U9610 ( .A(n688), .B(n9987), .Z(n9992) );
  XNOR U9611 ( .A(n9991), .B(n9985), .Z(n9987) );
  XOR U9612 ( .A(n9993), .B(n9994), .Z(n9985) );
  AND U9613 ( .A(n703), .B(n9995), .Z(n9994) );
  XNOR U9614 ( .A(n9996), .B(n9997), .Z(n9991) );
  AND U9615 ( .A(n695), .B(n9998), .Z(n9997) );
  XOR U9616 ( .A(p_input[975]), .B(n9996), .Z(n9998) );
  XNOR U9617 ( .A(n9999), .B(n10000), .Z(n9996) );
  AND U9618 ( .A(n699), .B(n9995), .Z(n10000) );
  XNOR U9619 ( .A(n9999), .B(n9993), .Z(n9995) );
  XOR U9620 ( .A(n10001), .B(n10002), .Z(n9993) );
  AND U9621 ( .A(n714), .B(n10003), .Z(n10002) );
  XNOR U9622 ( .A(n10004), .B(n10005), .Z(n9999) );
  AND U9623 ( .A(n706), .B(n10006), .Z(n10005) );
  XOR U9624 ( .A(p_input[991]), .B(n10004), .Z(n10006) );
  XNOR U9625 ( .A(n10007), .B(n10008), .Z(n10004) );
  AND U9626 ( .A(n710), .B(n10003), .Z(n10008) );
  XNOR U9627 ( .A(n10007), .B(n10001), .Z(n10003) );
  XOR U9628 ( .A(n10009), .B(n10010), .Z(n10001) );
  AND U9629 ( .A(n725), .B(n10011), .Z(n10010) );
  XNOR U9630 ( .A(n10012), .B(n10013), .Z(n10007) );
  AND U9631 ( .A(n717), .B(n10014), .Z(n10013) );
  XOR U9632 ( .A(p_input[1007]), .B(n10012), .Z(n10014) );
  XNOR U9633 ( .A(n10015), .B(n10016), .Z(n10012) );
  AND U9634 ( .A(n721), .B(n10011), .Z(n10016) );
  XNOR U9635 ( .A(n10015), .B(n10009), .Z(n10011) );
  XOR U9636 ( .A(n10017), .B(n10018), .Z(n10009) );
  AND U9637 ( .A(n736), .B(n10019), .Z(n10018) );
  XNOR U9638 ( .A(n10020), .B(n10021), .Z(n10015) );
  AND U9639 ( .A(n728), .B(n10022), .Z(n10021) );
  XOR U9640 ( .A(p_input[1023]), .B(n10020), .Z(n10022) );
  XNOR U9641 ( .A(n10023), .B(n10024), .Z(n10020) );
  AND U9642 ( .A(n732), .B(n10019), .Z(n10024) );
  XNOR U9643 ( .A(n10023), .B(n10017), .Z(n10019) );
  XOR U9644 ( .A(n10025), .B(n10026), .Z(n10017) );
  AND U9645 ( .A(n747), .B(n10027), .Z(n10026) );
  XNOR U9646 ( .A(n10028), .B(n10029), .Z(n10023) );
  AND U9647 ( .A(n739), .B(n10030), .Z(n10029) );
  XOR U9648 ( .A(p_input[1039]), .B(n10028), .Z(n10030) );
  XNOR U9649 ( .A(n10031), .B(n10032), .Z(n10028) );
  AND U9650 ( .A(n743), .B(n10027), .Z(n10032) );
  XNOR U9651 ( .A(n10031), .B(n10025), .Z(n10027) );
  XOR U9652 ( .A(n10033), .B(n10034), .Z(n10025) );
  AND U9653 ( .A(n758), .B(n10035), .Z(n10034) );
  XNOR U9654 ( .A(n10036), .B(n10037), .Z(n10031) );
  AND U9655 ( .A(n750), .B(n10038), .Z(n10037) );
  XOR U9656 ( .A(p_input[1055]), .B(n10036), .Z(n10038) );
  XNOR U9657 ( .A(n10039), .B(n10040), .Z(n10036) );
  AND U9658 ( .A(n754), .B(n10035), .Z(n10040) );
  XNOR U9659 ( .A(n10039), .B(n10033), .Z(n10035) );
  XOR U9660 ( .A(n10041), .B(n10042), .Z(n10033) );
  AND U9661 ( .A(n769), .B(n10043), .Z(n10042) );
  XNOR U9662 ( .A(n10044), .B(n10045), .Z(n10039) );
  AND U9663 ( .A(n761), .B(n10046), .Z(n10045) );
  XOR U9664 ( .A(p_input[1071]), .B(n10044), .Z(n10046) );
  XNOR U9665 ( .A(n10047), .B(n10048), .Z(n10044) );
  AND U9666 ( .A(n765), .B(n10043), .Z(n10048) );
  XNOR U9667 ( .A(n10047), .B(n10041), .Z(n10043) );
  XOR U9668 ( .A(n10049), .B(n10050), .Z(n10041) );
  AND U9669 ( .A(n780), .B(n10051), .Z(n10050) );
  XNOR U9670 ( .A(n10052), .B(n10053), .Z(n10047) );
  AND U9671 ( .A(n772), .B(n10054), .Z(n10053) );
  XOR U9672 ( .A(p_input[1087]), .B(n10052), .Z(n10054) );
  XNOR U9673 ( .A(n10055), .B(n10056), .Z(n10052) );
  AND U9674 ( .A(n776), .B(n10051), .Z(n10056) );
  XNOR U9675 ( .A(n10055), .B(n10049), .Z(n10051) );
  XOR U9676 ( .A(n10057), .B(n10058), .Z(n10049) );
  AND U9677 ( .A(n791), .B(n10059), .Z(n10058) );
  XNOR U9678 ( .A(n10060), .B(n10061), .Z(n10055) );
  AND U9679 ( .A(n783), .B(n10062), .Z(n10061) );
  XOR U9680 ( .A(p_input[1103]), .B(n10060), .Z(n10062) );
  XNOR U9681 ( .A(n10063), .B(n10064), .Z(n10060) );
  AND U9682 ( .A(n787), .B(n10059), .Z(n10064) );
  XNOR U9683 ( .A(n10063), .B(n10057), .Z(n10059) );
  XOR U9684 ( .A(n10065), .B(n10066), .Z(n10057) );
  AND U9685 ( .A(n802), .B(n10067), .Z(n10066) );
  XNOR U9686 ( .A(n10068), .B(n10069), .Z(n10063) );
  AND U9687 ( .A(n794), .B(n10070), .Z(n10069) );
  XOR U9688 ( .A(p_input[1119]), .B(n10068), .Z(n10070) );
  XNOR U9689 ( .A(n10071), .B(n10072), .Z(n10068) );
  AND U9690 ( .A(n798), .B(n10067), .Z(n10072) );
  XNOR U9691 ( .A(n10071), .B(n10065), .Z(n10067) );
  XOR U9692 ( .A(n10073), .B(n10074), .Z(n10065) );
  AND U9693 ( .A(n813), .B(n10075), .Z(n10074) );
  XNOR U9694 ( .A(n10076), .B(n10077), .Z(n10071) );
  AND U9695 ( .A(n805), .B(n10078), .Z(n10077) );
  XOR U9696 ( .A(p_input[1135]), .B(n10076), .Z(n10078) );
  XNOR U9697 ( .A(n10079), .B(n10080), .Z(n10076) );
  AND U9698 ( .A(n809), .B(n10075), .Z(n10080) );
  XNOR U9699 ( .A(n10079), .B(n10073), .Z(n10075) );
  XOR U9700 ( .A(n10081), .B(n10082), .Z(n10073) );
  AND U9701 ( .A(n824), .B(n10083), .Z(n10082) );
  XNOR U9702 ( .A(n10084), .B(n10085), .Z(n10079) );
  AND U9703 ( .A(n816), .B(n10086), .Z(n10085) );
  XOR U9704 ( .A(p_input[1151]), .B(n10084), .Z(n10086) );
  XNOR U9705 ( .A(n10087), .B(n10088), .Z(n10084) );
  AND U9706 ( .A(n820), .B(n10083), .Z(n10088) );
  XNOR U9707 ( .A(n10087), .B(n10081), .Z(n10083) );
  XOR U9708 ( .A(n10089), .B(n10090), .Z(n10081) );
  AND U9709 ( .A(n835), .B(n10091), .Z(n10090) );
  XNOR U9710 ( .A(n10092), .B(n10093), .Z(n10087) );
  AND U9711 ( .A(n827), .B(n10094), .Z(n10093) );
  XOR U9712 ( .A(p_input[1167]), .B(n10092), .Z(n10094) );
  XNOR U9713 ( .A(n10095), .B(n10096), .Z(n10092) );
  AND U9714 ( .A(n831), .B(n10091), .Z(n10096) );
  XNOR U9715 ( .A(n10095), .B(n10089), .Z(n10091) );
  XOR U9716 ( .A(n10097), .B(n10098), .Z(n10089) );
  AND U9717 ( .A(n846), .B(n10099), .Z(n10098) );
  XNOR U9718 ( .A(n10100), .B(n10101), .Z(n10095) );
  AND U9719 ( .A(n838), .B(n10102), .Z(n10101) );
  XOR U9720 ( .A(p_input[1183]), .B(n10100), .Z(n10102) );
  XNOR U9721 ( .A(n10103), .B(n10104), .Z(n10100) );
  AND U9722 ( .A(n842), .B(n10099), .Z(n10104) );
  XNOR U9723 ( .A(n10103), .B(n10097), .Z(n10099) );
  XOR U9724 ( .A(n10105), .B(n10106), .Z(n10097) );
  AND U9725 ( .A(n857), .B(n10107), .Z(n10106) );
  XNOR U9726 ( .A(n10108), .B(n10109), .Z(n10103) );
  AND U9727 ( .A(n849), .B(n10110), .Z(n10109) );
  XOR U9728 ( .A(p_input[1199]), .B(n10108), .Z(n10110) );
  XNOR U9729 ( .A(n10111), .B(n10112), .Z(n10108) );
  AND U9730 ( .A(n853), .B(n10107), .Z(n10112) );
  XNOR U9731 ( .A(n10111), .B(n10105), .Z(n10107) );
  XOR U9732 ( .A(n10113), .B(n10114), .Z(n10105) );
  AND U9733 ( .A(n868), .B(n10115), .Z(n10114) );
  XNOR U9734 ( .A(n10116), .B(n10117), .Z(n10111) );
  AND U9735 ( .A(n860), .B(n10118), .Z(n10117) );
  XOR U9736 ( .A(p_input[1215]), .B(n10116), .Z(n10118) );
  XNOR U9737 ( .A(n10119), .B(n10120), .Z(n10116) );
  AND U9738 ( .A(n864), .B(n10115), .Z(n10120) );
  XNOR U9739 ( .A(n10119), .B(n10113), .Z(n10115) );
  XOR U9740 ( .A(n10121), .B(n10122), .Z(n10113) );
  AND U9741 ( .A(n879), .B(n10123), .Z(n10122) );
  XNOR U9742 ( .A(n10124), .B(n10125), .Z(n10119) );
  AND U9743 ( .A(n871), .B(n10126), .Z(n10125) );
  XOR U9744 ( .A(p_input[1231]), .B(n10124), .Z(n10126) );
  XNOR U9745 ( .A(n10127), .B(n10128), .Z(n10124) );
  AND U9746 ( .A(n875), .B(n10123), .Z(n10128) );
  XNOR U9747 ( .A(n10127), .B(n10121), .Z(n10123) );
  XOR U9748 ( .A(n10129), .B(n10130), .Z(n10121) );
  AND U9749 ( .A(n890), .B(n10131), .Z(n10130) );
  XNOR U9750 ( .A(n10132), .B(n10133), .Z(n10127) );
  AND U9751 ( .A(n882), .B(n10134), .Z(n10133) );
  XOR U9752 ( .A(p_input[1247]), .B(n10132), .Z(n10134) );
  XNOR U9753 ( .A(n10135), .B(n10136), .Z(n10132) );
  AND U9754 ( .A(n886), .B(n10131), .Z(n10136) );
  XNOR U9755 ( .A(n10135), .B(n10129), .Z(n10131) );
  XOR U9756 ( .A(n10137), .B(n10138), .Z(n10129) );
  AND U9757 ( .A(n901), .B(n10139), .Z(n10138) );
  XNOR U9758 ( .A(n10140), .B(n10141), .Z(n10135) );
  AND U9759 ( .A(n893), .B(n10142), .Z(n10141) );
  XOR U9760 ( .A(p_input[1263]), .B(n10140), .Z(n10142) );
  XNOR U9761 ( .A(n10143), .B(n10144), .Z(n10140) );
  AND U9762 ( .A(n897), .B(n10139), .Z(n10144) );
  XNOR U9763 ( .A(n10143), .B(n10137), .Z(n10139) );
  XOR U9764 ( .A(n10145), .B(n10146), .Z(n10137) );
  AND U9765 ( .A(n912), .B(n10147), .Z(n10146) );
  XNOR U9766 ( .A(n10148), .B(n10149), .Z(n10143) );
  AND U9767 ( .A(n904), .B(n10150), .Z(n10149) );
  XOR U9768 ( .A(p_input[1279]), .B(n10148), .Z(n10150) );
  XNOR U9769 ( .A(n10151), .B(n10152), .Z(n10148) );
  AND U9770 ( .A(n908), .B(n10147), .Z(n10152) );
  XNOR U9771 ( .A(n10151), .B(n10145), .Z(n10147) );
  XOR U9772 ( .A(n10153), .B(n10154), .Z(n10145) );
  AND U9773 ( .A(n923), .B(n10155), .Z(n10154) );
  XNOR U9774 ( .A(n10156), .B(n10157), .Z(n10151) );
  AND U9775 ( .A(n915), .B(n10158), .Z(n10157) );
  XOR U9776 ( .A(p_input[1295]), .B(n10156), .Z(n10158) );
  XNOR U9777 ( .A(n10159), .B(n10160), .Z(n10156) );
  AND U9778 ( .A(n919), .B(n10155), .Z(n10160) );
  XNOR U9779 ( .A(n10159), .B(n10153), .Z(n10155) );
  XOR U9780 ( .A(n10161), .B(n10162), .Z(n10153) );
  AND U9781 ( .A(n934), .B(n10163), .Z(n10162) );
  XNOR U9782 ( .A(n10164), .B(n10165), .Z(n10159) );
  AND U9783 ( .A(n926), .B(n10166), .Z(n10165) );
  XOR U9784 ( .A(p_input[1311]), .B(n10164), .Z(n10166) );
  XNOR U9785 ( .A(n10167), .B(n10168), .Z(n10164) );
  AND U9786 ( .A(n930), .B(n10163), .Z(n10168) );
  XNOR U9787 ( .A(n10167), .B(n10161), .Z(n10163) );
  XOR U9788 ( .A(n10169), .B(n10170), .Z(n10161) );
  AND U9789 ( .A(n945), .B(n10171), .Z(n10170) );
  XNOR U9790 ( .A(n10172), .B(n10173), .Z(n10167) );
  AND U9791 ( .A(n937), .B(n10174), .Z(n10173) );
  XOR U9792 ( .A(p_input[1327]), .B(n10172), .Z(n10174) );
  XNOR U9793 ( .A(n10175), .B(n10176), .Z(n10172) );
  AND U9794 ( .A(n941), .B(n10171), .Z(n10176) );
  XNOR U9795 ( .A(n10175), .B(n10169), .Z(n10171) );
  XOR U9796 ( .A(n10177), .B(n10178), .Z(n10169) );
  AND U9797 ( .A(n956), .B(n10179), .Z(n10178) );
  XNOR U9798 ( .A(n10180), .B(n10181), .Z(n10175) );
  AND U9799 ( .A(n948), .B(n10182), .Z(n10181) );
  XOR U9800 ( .A(p_input[1343]), .B(n10180), .Z(n10182) );
  XNOR U9801 ( .A(n10183), .B(n10184), .Z(n10180) );
  AND U9802 ( .A(n952), .B(n10179), .Z(n10184) );
  XNOR U9803 ( .A(n10183), .B(n10177), .Z(n10179) );
  XOR U9804 ( .A(n10185), .B(n10186), .Z(n10177) );
  AND U9805 ( .A(n967), .B(n10187), .Z(n10186) );
  XNOR U9806 ( .A(n10188), .B(n10189), .Z(n10183) );
  AND U9807 ( .A(n959), .B(n10190), .Z(n10189) );
  XOR U9808 ( .A(p_input[1359]), .B(n10188), .Z(n10190) );
  XNOR U9809 ( .A(n10191), .B(n10192), .Z(n10188) );
  AND U9810 ( .A(n963), .B(n10187), .Z(n10192) );
  XNOR U9811 ( .A(n10191), .B(n10185), .Z(n10187) );
  XOR U9812 ( .A(n10193), .B(n10194), .Z(n10185) );
  AND U9813 ( .A(n978), .B(n10195), .Z(n10194) );
  XNOR U9814 ( .A(n10196), .B(n10197), .Z(n10191) );
  AND U9815 ( .A(n970), .B(n10198), .Z(n10197) );
  XOR U9816 ( .A(p_input[1375]), .B(n10196), .Z(n10198) );
  XNOR U9817 ( .A(n10199), .B(n10200), .Z(n10196) );
  AND U9818 ( .A(n974), .B(n10195), .Z(n10200) );
  XNOR U9819 ( .A(n10199), .B(n10193), .Z(n10195) );
  XOR U9820 ( .A(n10201), .B(n10202), .Z(n10193) );
  AND U9821 ( .A(n989), .B(n10203), .Z(n10202) );
  XNOR U9822 ( .A(n10204), .B(n10205), .Z(n10199) );
  AND U9823 ( .A(n981), .B(n10206), .Z(n10205) );
  XOR U9824 ( .A(p_input[1391]), .B(n10204), .Z(n10206) );
  XNOR U9825 ( .A(n10207), .B(n10208), .Z(n10204) );
  AND U9826 ( .A(n985), .B(n10203), .Z(n10208) );
  XNOR U9827 ( .A(n10207), .B(n10201), .Z(n10203) );
  XOR U9828 ( .A(n10209), .B(n10210), .Z(n10201) );
  AND U9829 ( .A(n1000), .B(n10211), .Z(n10210) );
  XNOR U9830 ( .A(n10212), .B(n10213), .Z(n10207) );
  AND U9831 ( .A(n992), .B(n10214), .Z(n10213) );
  XOR U9832 ( .A(p_input[1407]), .B(n10212), .Z(n10214) );
  XNOR U9833 ( .A(n10215), .B(n10216), .Z(n10212) );
  AND U9834 ( .A(n996), .B(n10211), .Z(n10216) );
  XNOR U9835 ( .A(n10215), .B(n10209), .Z(n10211) );
  XOR U9836 ( .A(n10217), .B(n10218), .Z(n10209) );
  AND U9837 ( .A(n1011), .B(n10219), .Z(n10218) );
  XNOR U9838 ( .A(n10220), .B(n10221), .Z(n10215) );
  AND U9839 ( .A(n1003), .B(n10222), .Z(n10221) );
  XOR U9840 ( .A(p_input[1423]), .B(n10220), .Z(n10222) );
  XNOR U9841 ( .A(n10223), .B(n10224), .Z(n10220) );
  AND U9842 ( .A(n1007), .B(n10219), .Z(n10224) );
  XNOR U9843 ( .A(n10223), .B(n10217), .Z(n10219) );
  XOR U9844 ( .A(n10225), .B(n10226), .Z(n10217) );
  AND U9845 ( .A(n1022), .B(n10227), .Z(n10226) );
  XNOR U9846 ( .A(n10228), .B(n10229), .Z(n10223) );
  AND U9847 ( .A(n1014), .B(n10230), .Z(n10229) );
  XOR U9848 ( .A(p_input[1439]), .B(n10228), .Z(n10230) );
  XNOR U9849 ( .A(n10231), .B(n10232), .Z(n10228) );
  AND U9850 ( .A(n1018), .B(n10227), .Z(n10232) );
  XNOR U9851 ( .A(n10231), .B(n10225), .Z(n10227) );
  XOR U9852 ( .A(n10233), .B(n10234), .Z(n10225) );
  AND U9853 ( .A(n1033), .B(n10235), .Z(n10234) );
  XNOR U9854 ( .A(n10236), .B(n10237), .Z(n10231) );
  AND U9855 ( .A(n1025), .B(n10238), .Z(n10237) );
  XOR U9856 ( .A(p_input[1455]), .B(n10236), .Z(n10238) );
  XNOR U9857 ( .A(n10239), .B(n10240), .Z(n10236) );
  AND U9858 ( .A(n1029), .B(n10235), .Z(n10240) );
  XNOR U9859 ( .A(n10239), .B(n10233), .Z(n10235) );
  XOR U9860 ( .A(n10241), .B(n10242), .Z(n10233) );
  AND U9861 ( .A(n1044), .B(n10243), .Z(n10242) );
  XNOR U9862 ( .A(n10244), .B(n10245), .Z(n10239) );
  AND U9863 ( .A(n1036), .B(n10246), .Z(n10245) );
  XOR U9864 ( .A(p_input[1471]), .B(n10244), .Z(n10246) );
  XNOR U9865 ( .A(n10247), .B(n10248), .Z(n10244) );
  AND U9866 ( .A(n1040), .B(n10243), .Z(n10248) );
  XNOR U9867 ( .A(n10247), .B(n10241), .Z(n10243) );
  XOR U9868 ( .A(n10249), .B(n10250), .Z(n10241) );
  AND U9869 ( .A(n1055), .B(n10251), .Z(n10250) );
  XNOR U9870 ( .A(n10252), .B(n10253), .Z(n10247) );
  AND U9871 ( .A(n1047), .B(n10254), .Z(n10253) );
  XOR U9872 ( .A(p_input[1487]), .B(n10252), .Z(n10254) );
  XNOR U9873 ( .A(n10255), .B(n10256), .Z(n10252) );
  AND U9874 ( .A(n1051), .B(n10251), .Z(n10256) );
  XNOR U9875 ( .A(n10255), .B(n10249), .Z(n10251) );
  XOR U9876 ( .A(n10257), .B(n10258), .Z(n10249) );
  AND U9877 ( .A(n1066), .B(n10259), .Z(n10258) );
  XNOR U9878 ( .A(n10260), .B(n10261), .Z(n10255) );
  AND U9879 ( .A(n1058), .B(n10262), .Z(n10261) );
  XOR U9880 ( .A(p_input[1503]), .B(n10260), .Z(n10262) );
  XNOR U9881 ( .A(n10263), .B(n10264), .Z(n10260) );
  AND U9882 ( .A(n1062), .B(n10259), .Z(n10264) );
  XNOR U9883 ( .A(n10263), .B(n10257), .Z(n10259) );
  XOR U9884 ( .A(n10265), .B(n10266), .Z(n10257) );
  AND U9885 ( .A(n1077), .B(n10267), .Z(n10266) );
  XNOR U9886 ( .A(n10268), .B(n10269), .Z(n10263) );
  AND U9887 ( .A(n1069), .B(n10270), .Z(n10269) );
  XOR U9888 ( .A(p_input[1519]), .B(n10268), .Z(n10270) );
  XNOR U9889 ( .A(n10271), .B(n10272), .Z(n10268) );
  AND U9890 ( .A(n1073), .B(n10267), .Z(n10272) );
  XNOR U9891 ( .A(n10271), .B(n10265), .Z(n10267) );
  XOR U9892 ( .A(n10273), .B(n10274), .Z(n10265) );
  AND U9893 ( .A(n1088), .B(n10275), .Z(n10274) );
  XNOR U9894 ( .A(n10276), .B(n10277), .Z(n10271) );
  AND U9895 ( .A(n1080), .B(n10278), .Z(n10277) );
  XOR U9896 ( .A(p_input[1535]), .B(n10276), .Z(n10278) );
  XNOR U9897 ( .A(n10279), .B(n10280), .Z(n10276) );
  AND U9898 ( .A(n1084), .B(n10275), .Z(n10280) );
  XNOR U9899 ( .A(n10279), .B(n10273), .Z(n10275) );
  XOR U9900 ( .A(n10281), .B(n10282), .Z(n10273) );
  AND U9901 ( .A(n1099), .B(n10283), .Z(n10282) );
  XNOR U9902 ( .A(n10284), .B(n10285), .Z(n10279) );
  AND U9903 ( .A(n1091), .B(n10286), .Z(n10285) );
  XOR U9904 ( .A(p_input[1551]), .B(n10284), .Z(n10286) );
  XNOR U9905 ( .A(n10287), .B(n10288), .Z(n10284) );
  AND U9906 ( .A(n1095), .B(n10283), .Z(n10288) );
  XNOR U9907 ( .A(n10287), .B(n10281), .Z(n10283) );
  XOR U9908 ( .A(n10289), .B(n10290), .Z(n10281) );
  AND U9909 ( .A(n1110), .B(n10291), .Z(n10290) );
  XNOR U9910 ( .A(n10292), .B(n10293), .Z(n10287) );
  AND U9911 ( .A(n1102), .B(n10294), .Z(n10293) );
  XOR U9912 ( .A(p_input[1567]), .B(n10292), .Z(n10294) );
  XNOR U9913 ( .A(n10295), .B(n10296), .Z(n10292) );
  AND U9914 ( .A(n1106), .B(n10291), .Z(n10296) );
  XNOR U9915 ( .A(n10295), .B(n10289), .Z(n10291) );
  XOR U9916 ( .A(n10297), .B(n10298), .Z(n10289) );
  AND U9917 ( .A(n1121), .B(n10299), .Z(n10298) );
  XNOR U9918 ( .A(n10300), .B(n10301), .Z(n10295) );
  AND U9919 ( .A(n1113), .B(n10302), .Z(n10301) );
  XOR U9920 ( .A(p_input[1583]), .B(n10300), .Z(n10302) );
  XNOR U9921 ( .A(n10303), .B(n10304), .Z(n10300) );
  AND U9922 ( .A(n1117), .B(n10299), .Z(n10304) );
  XNOR U9923 ( .A(n10303), .B(n10297), .Z(n10299) );
  XOR U9924 ( .A(n10305), .B(n10306), .Z(n10297) );
  AND U9925 ( .A(n1132), .B(n10307), .Z(n10306) );
  XNOR U9926 ( .A(n10308), .B(n10309), .Z(n10303) );
  AND U9927 ( .A(n1124), .B(n10310), .Z(n10309) );
  XOR U9928 ( .A(p_input[1599]), .B(n10308), .Z(n10310) );
  XNOR U9929 ( .A(n10311), .B(n10312), .Z(n10308) );
  AND U9930 ( .A(n1128), .B(n10307), .Z(n10312) );
  XNOR U9931 ( .A(n10311), .B(n10305), .Z(n10307) );
  XOR U9932 ( .A(n10313), .B(n10314), .Z(n10305) );
  AND U9933 ( .A(n1143), .B(n10315), .Z(n10314) );
  XNOR U9934 ( .A(n10316), .B(n10317), .Z(n10311) );
  AND U9935 ( .A(n1135), .B(n10318), .Z(n10317) );
  XOR U9936 ( .A(p_input[1615]), .B(n10316), .Z(n10318) );
  XNOR U9937 ( .A(n10319), .B(n10320), .Z(n10316) );
  AND U9938 ( .A(n1139), .B(n10315), .Z(n10320) );
  XNOR U9939 ( .A(n10319), .B(n10313), .Z(n10315) );
  XOR U9940 ( .A(n10321), .B(n10322), .Z(n10313) );
  AND U9941 ( .A(n1154), .B(n10323), .Z(n10322) );
  XNOR U9942 ( .A(n10324), .B(n10325), .Z(n10319) );
  AND U9943 ( .A(n1146), .B(n10326), .Z(n10325) );
  XOR U9944 ( .A(p_input[1631]), .B(n10324), .Z(n10326) );
  XNOR U9945 ( .A(n10327), .B(n10328), .Z(n10324) );
  AND U9946 ( .A(n1150), .B(n10323), .Z(n10328) );
  XNOR U9947 ( .A(n10327), .B(n10321), .Z(n10323) );
  XOR U9948 ( .A(n10329), .B(n10330), .Z(n10321) );
  AND U9949 ( .A(n1165), .B(n10331), .Z(n10330) );
  XNOR U9950 ( .A(n10332), .B(n10333), .Z(n10327) );
  AND U9951 ( .A(n1157), .B(n10334), .Z(n10333) );
  XOR U9952 ( .A(p_input[1647]), .B(n10332), .Z(n10334) );
  XNOR U9953 ( .A(n10335), .B(n10336), .Z(n10332) );
  AND U9954 ( .A(n1161), .B(n10331), .Z(n10336) );
  XNOR U9955 ( .A(n10335), .B(n10329), .Z(n10331) );
  XOR U9956 ( .A(n10337), .B(n10338), .Z(n10329) );
  AND U9957 ( .A(n1176), .B(n10339), .Z(n10338) );
  XNOR U9958 ( .A(n10340), .B(n10341), .Z(n10335) );
  AND U9959 ( .A(n1168), .B(n10342), .Z(n10341) );
  XOR U9960 ( .A(p_input[1663]), .B(n10340), .Z(n10342) );
  XNOR U9961 ( .A(n10343), .B(n10344), .Z(n10340) );
  AND U9962 ( .A(n1172), .B(n10339), .Z(n10344) );
  XNOR U9963 ( .A(n10343), .B(n10337), .Z(n10339) );
  XOR U9964 ( .A(n10345), .B(n10346), .Z(n10337) );
  AND U9965 ( .A(n1187), .B(n10347), .Z(n10346) );
  XNOR U9966 ( .A(n10348), .B(n10349), .Z(n10343) );
  AND U9967 ( .A(n1179), .B(n10350), .Z(n10349) );
  XOR U9968 ( .A(p_input[1679]), .B(n10348), .Z(n10350) );
  XNOR U9969 ( .A(n10351), .B(n10352), .Z(n10348) );
  AND U9970 ( .A(n1183), .B(n10347), .Z(n10352) );
  XNOR U9971 ( .A(n10351), .B(n10345), .Z(n10347) );
  XOR U9972 ( .A(n10353), .B(n10354), .Z(n10345) );
  AND U9973 ( .A(n1198), .B(n10355), .Z(n10354) );
  XNOR U9974 ( .A(n10356), .B(n10357), .Z(n10351) );
  AND U9975 ( .A(n1190), .B(n10358), .Z(n10357) );
  XOR U9976 ( .A(p_input[1695]), .B(n10356), .Z(n10358) );
  XNOR U9977 ( .A(n10359), .B(n10360), .Z(n10356) );
  AND U9978 ( .A(n1194), .B(n10355), .Z(n10360) );
  XNOR U9979 ( .A(n10359), .B(n10353), .Z(n10355) );
  XOR U9980 ( .A(n10361), .B(n10362), .Z(n10353) );
  AND U9981 ( .A(n1209), .B(n10363), .Z(n10362) );
  XNOR U9982 ( .A(n10364), .B(n10365), .Z(n10359) );
  AND U9983 ( .A(n1201), .B(n10366), .Z(n10365) );
  XOR U9984 ( .A(p_input[1711]), .B(n10364), .Z(n10366) );
  XNOR U9985 ( .A(n10367), .B(n10368), .Z(n10364) );
  AND U9986 ( .A(n1205), .B(n10363), .Z(n10368) );
  XNOR U9987 ( .A(n10367), .B(n10361), .Z(n10363) );
  XOR U9988 ( .A(n10369), .B(n10370), .Z(n10361) );
  AND U9989 ( .A(n1220), .B(n10371), .Z(n10370) );
  XNOR U9990 ( .A(n10372), .B(n10373), .Z(n10367) );
  AND U9991 ( .A(n1212), .B(n10374), .Z(n10373) );
  XOR U9992 ( .A(p_input[1727]), .B(n10372), .Z(n10374) );
  XNOR U9993 ( .A(n10375), .B(n10376), .Z(n10372) );
  AND U9994 ( .A(n1216), .B(n10371), .Z(n10376) );
  XNOR U9995 ( .A(n10375), .B(n10369), .Z(n10371) );
  XOR U9996 ( .A(n10377), .B(n10378), .Z(n10369) );
  AND U9997 ( .A(n1231), .B(n10379), .Z(n10378) );
  XNOR U9998 ( .A(n10380), .B(n10381), .Z(n10375) );
  AND U9999 ( .A(n1223), .B(n10382), .Z(n10381) );
  XOR U10000 ( .A(p_input[1743]), .B(n10380), .Z(n10382) );
  XNOR U10001 ( .A(n10383), .B(n10384), .Z(n10380) );
  AND U10002 ( .A(n1227), .B(n10379), .Z(n10384) );
  XNOR U10003 ( .A(n10383), .B(n10377), .Z(n10379) );
  XOR U10004 ( .A(n10385), .B(n10386), .Z(n10377) );
  AND U10005 ( .A(n1242), .B(n10387), .Z(n10386) );
  XNOR U10006 ( .A(n10388), .B(n10389), .Z(n10383) );
  AND U10007 ( .A(n1234), .B(n10390), .Z(n10389) );
  XOR U10008 ( .A(p_input[1759]), .B(n10388), .Z(n10390) );
  XNOR U10009 ( .A(n10391), .B(n10392), .Z(n10388) );
  AND U10010 ( .A(n1238), .B(n10387), .Z(n10392) );
  XNOR U10011 ( .A(n10391), .B(n10385), .Z(n10387) );
  XOR U10012 ( .A(n10393), .B(n10394), .Z(n10385) );
  AND U10013 ( .A(n1253), .B(n10395), .Z(n10394) );
  XNOR U10014 ( .A(n10396), .B(n10397), .Z(n10391) );
  AND U10015 ( .A(n1245), .B(n10398), .Z(n10397) );
  XOR U10016 ( .A(p_input[1775]), .B(n10396), .Z(n10398) );
  XNOR U10017 ( .A(n10399), .B(n10400), .Z(n10396) );
  AND U10018 ( .A(n1249), .B(n10395), .Z(n10400) );
  XNOR U10019 ( .A(n10399), .B(n10393), .Z(n10395) );
  XOR U10020 ( .A(n10401), .B(n10402), .Z(n10393) );
  AND U10021 ( .A(n1264), .B(n10403), .Z(n10402) );
  XNOR U10022 ( .A(n10404), .B(n10405), .Z(n10399) );
  AND U10023 ( .A(n1256), .B(n10406), .Z(n10405) );
  XOR U10024 ( .A(p_input[1791]), .B(n10404), .Z(n10406) );
  XNOR U10025 ( .A(n10407), .B(n10408), .Z(n10404) );
  AND U10026 ( .A(n1260), .B(n10403), .Z(n10408) );
  XNOR U10027 ( .A(n10407), .B(n10401), .Z(n10403) );
  XOR U10028 ( .A(n10409), .B(n10410), .Z(n10401) );
  AND U10029 ( .A(n1275), .B(n10411), .Z(n10410) );
  XNOR U10030 ( .A(n10412), .B(n10413), .Z(n10407) );
  AND U10031 ( .A(n1267), .B(n10414), .Z(n10413) );
  XOR U10032 ( .A(p_input[1807]), .B(n10412), .Z(n10414) );
  XNOR U10033 ( .A(n10415), .B(n10416), .Z(n10412) );
  AND U10034 ( .A(n1271), .B(n10411), .Z(n10416) );
  XNOR U10035 ( .A(n10415), .B(n10409), .Z(n10411) );
  XOR U10036 ( .A(n10417), .B(n10418), .Z(n10409) );
  AND U10037 ( .A(n1286), .B(n10419), .Z(n10418) );
  XNOR U10038 ( .A(n10420), .B(n10421), .Z(n10415) );
  AND U10039 ( .A(n1278), .B(n10422), .Z(n10421) );
  XOR U10040 ( .A(p_input[1823]), .B(n10420), .Z(n10422) );
  XNOR U10041 ( .A(n10423), .B(n10424), .Z(n10420) );
  AND U10042 ( .A(n1282), .B(n10419), .Z(n10424) );
  XNOR U10043 ( .A(n10423), .B(n10417), .Z(n10419) );
  XOR U10044 ( .A(n10425), .B(n10426), .Z(n10417) );
  AND U10045 ( .A(n1297), .B(n10427), .Z(n10426) );
  XNOR U10046 ( .A(n10428), .B(n10429), .Z(n10423) );
  AND U10047 ( .A(n1289), .B(n10430), .Z(n10429) );
  XOR U10048 ( .A(p_input[1839]), .B(n10428), .Z(n10430) );
  XNOR U10049 ( .A(n10431), .B(n10432), .Z(n10428) );
  AND U10050 ( .A(n1293), .B(n10427), .Z(n10432) );
  XNOR U10051 ( .A(n10431), .B(n10425), .Z(n10427) );
  XOR U10052 ( .A(n10433), .B(n10434), .Z(n10425) );
  AND U10053 ( .A(n1308), .B(n10435), .Z(n10434) );
  XNOR U10054 ( .A(n10436), .B(n10437), .Z(n10431) );
  AND U10055 ( .A(n1300), .B(n10438), .Z(n10437) );
  XOR U10056 ( .A(p_input[1855]), .B(n10436), .Z(n10438) );
  XNOR U10057 ( .A(n10439), .B(n10440), .Z(n10436) );
  AND U10058 ( .A(n1304), .B(n10435), .Z(n10440) );
  XNOR U10059 ( .A(n10439), .B(n10433), .Z(n10435) );
  XOR U10060 ( .A(n10441), .B(n10442), .Z(n10433) );
  AND U10061 ( .A(n1319), .B(n10443), .Z(n10442) );
  XNOR U10062 ( .A(n10444), .B(n10445), .Z(n10439) );
  AND U10063 ( .A(n1311), .B(n10446), .Z(n10445) );
  XOR U10064 ( .A(p_input[1871]), .B(n10444), .Z(n10446) );
  XNOR U10065 ( .A(n10447), .B(n10448), .Z(n10444) );
  AND U10066 ( .A(n1315), .B(n10443), .Z(n10448) );
  XNOR U10067 ( .A(n10447), .B(n10441), .Z(n10443) );
  XOR U10068 ( .A(n10449), .B(n10450), .Z(n10441) );
  AND U10069 ( .A(n1330), .B(n10451), .Z(n10450) );
  XNOR U10070 ( .A(n10452), .B(n10453), .Z(n10447) );
  AND U10071 ( .A(n1322), .B(n10454), .Z(n10453) );
  XOR U10072 ( .A(p_input[1887]), .B(n10452), .Z(n10454) );
  XNOR U10073 ( .A(n10455), .B(n10456), .Z(n10452) );
  AND U10074 ( .A(n1326), .B(n10451), .Z(n10456) );
  XNOR U10075 ( .A(n10455), .B(n10449), .Z(n10451) );
  XOR U10076 ( .A(n10457), .B(n10458), .Z(n10449) );
  AND U10077 ( .A(n1341), .B(n10459), .Z(n10458) );
  XNOR U10078 ( .A(n10460), .B(n10461), .Z(n10455) );
  AND U10079 ( .A(n1333), .B(n10462), .Z(n10461) );
  XOR U10080 ( .A(p_input[1903]), .B(n10460), .Z(n10462) );
  XNOR U10081 ( .A(n10463), .B(n10464), .Z(n10460) );
  AND U10082 ( .A(n1337), .B(n10459), .Z(n10464) );
  XNOR U10083 ( .A(n10463), .B(n10457), .Z(n10459) );
  XOR U10084 ( .A(n10465), .B(n10466), .Z(n10457) );
  AND U10085 ( .A(n1352), .B(n10467), .Z(n10466) );
  XNOR U10086 ( .A(n10468), .B(n10469), .Z(n10463) );
  AND U10087 ( .A(n1344), .B(n10470), .Z(n10469) );
  XOR U10088 ( .A(p_input[1919]), .B(n10468), .Z(n10470) );
  XNOR U10089 ( .A(n10471), .B(n10472), .Z(n10468) );
  AND U10090 ( .A(n1348), .B(n10467), .Z(n10472) );
  XNOR U10091 ( .A(n10471), .B(n10465), .Z(n10467) );
  XOR U10092 ( .A(n10473), .B(n10474), .Z(n10465) );
  AND U10093 ( .A(n1363), .B(n10475), .Z(n10474) );
  XNOR U10094 ( .A(n10476), .B(n10477), .Z(n10471) );
  AND U10095 ( .A(n1355), .B(n10478), .Z(n10477) );
  XOR U10096 ( .A(p_input[1935]), .B(n10476), .Z(n10478) );
  XNOR U10097 ( .A(n10479), .B(n10480), .Z(n10476) );
  AND U10098 ( .A(n1359), .B(n10475), .Z(n10480) );
  XNOR U10099 ( .A(n10479), .B(n10473), .Z(n10475) );
  XOR U10100 ( .A(n10481), .B(n10482), .Z(n10473) );
  AND U10101 ( .A(n1374), .B(n10483), .Z(n10482) );
  XNOR U10102 ( .A(n10484), .B(n10485), .Z(n10479) );
  AND U10103 ( .A(n1366), .B(n10486), .Z(n10485) );
  XOR U10104 ( .A(p_input[1951]), .B(n10484), .Z(n10486) );
  XNOR U10105 ( .A(n10487), .B(n10488), .Z(n10484) );
  AND U10106 ( .A(n1370), .B(n10483), .Z(n10488) );
  XNOR U10107 ( .A(n10487), .B(n10481), .Z(n10483) );
  XOR U10108 ( .A(n10489), .B(n10490), .Z(n10481) );
  AND U10109 ( .A(n1385), .B(n10491), .Z(n10490) );
  XNOR U10110 ( .A(n10492), .B(n10493), .Z(n10487) );
  AND U10111 ( .A(n1377), .B(n10494), .Z(n10493) );
  XOR U10112 ( .A(p_input[1967]), .B(n10492), .Z(n10494) );
  XNOR U10113 ( .A(n10495), .B(n10496), .Z(n10492) );
  AND U10114 ( .A(n1381), .B(n10491), .Z(n10496) );
  XNOR U10115 ( .A(n10495), .B(n10489), .Z(n10491) );
  XOR U10116 ( .A(n10497), .B(n10498), .Z(n10489) );
  AND U10117 ( .A(n1396), .B(n10499), .Z(n10498) );
  XNOR U10118 ( .A(n10500), .B(n10501), .Z(n10495) );
  AND U10119 ( .A(n1388), .B(n10502), .Z(n10501) );
  XOR U10120 ( .A(p_input[1983]), .B(n10500), .Z(n10502) );
  XNOR U10121 ( .A(n10503), .B(n10504), .Z(n10500) );
  AND U10122 ( .A(n1392), .B(n10499), .Z(n10504) );
  XNOR U10123 ( .A(n10503), .B(n10497), .Z(n10499) );
  XOR U10124 ( .A(n10505), .B(n10506), .Z(n10497) );
  AND U10125 ( .A(n1407), .B(n10507), .Z(n10506) );
  XNOR U10126 ( .A(n10508), .B(n10509), .Z(n10503) );
  AND U10127 ( .A(n1399), .B(n10510), .Z(n10509) );
  XOR U10128 ( .A(p_input[1999]), .B(n10508), .Z(n10510) );
  XNOR U10129 ( .A(n10511), .B(n10512), .Z(n10508) );
  AND U10130 ( .A(n1403), .B(n10507), .Z(n10512) );
  XNOR U10131 ( .A(n10511), .B(n10505), .Z(n10507) );
  XOR U10132 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n10513), .Z(n10505) );
  AND U10133 ( .A(n1417), .B(n10514), .Z(n10513) );
  XNOR U10134 ( .A(n10515), .B(n10516), .Z(n10511) );
  AND U10135 ( .A(n1410), .B(n10517), .Z(n10516) );
  XOR U10136 ( .A(p_input[2015]), .B(n10515), .Z(n10517) );
  XNOR U10137 ( .A(n10518), .B(n10519), .Z(n10515) );
  AND U10138 ( .A(n1414), .B(n10514), .Z(n10519) );
  XOR U10139 ( .A(n10520), .B(n10518), .Z(n10514) );
  IV U10140 ( .A(\knn_comb_/min_val_out[0][15] ), .Z(n10520) );
  IV U10141 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .Z(n10518)
         );
  XOR U10142 ( .A(n17), .B(n10521), .Z(o[14]) );
  AND U10143 ( .A(n30), .B(n10522), .Z(n17) );
  XOR U10144 ( .A(n18), .B(n10521), .Z(n10522) );
  XOR U10145 ( .A(n10523), .B(n10524), .Z(n10521) );
  AND U10146 ( .A(n42), .B(n10525), .Z(n10524) );
  XOR U10147 ( .A(n10526), .B(n10527), .Z(n18) );
  AND U10148 ( .A(n34), .B(n10528), .Z(n10527) );
  XOR U10149 ( .A(p_input[14]), .B(n10526), .Z(n10528) );
  XNOR U10150 ( .A(n10529), .B(n10530), .Z(n10526) );
  AND U10151 ( .A(n38), .B(n10525), .Z(n10530) );
  XNOR U10152 ( .A(n10529), .B(n10523), .Z(n10525) );
  XOR U10153 ( .A(n10531), .B(n10532), .Z(n10523) );
  AND U10154 ( .A(n54), .B(n10533), .Z(n10532) );
  XNOR U10155 ( .A(n10534), .B(n10535), .Z(n10529) );
  AND U10156 ( .A(n46), .B(n10536), .Z(n10535) );
  XOR U10157 ( .A(p_input[30]), .B(n10534), .Z(n10536) );
  XNOR U10158 ( .A(n10537), .B(n10538), .Z(n10534) );
  AND U10159 ( .A(n50), .B(n10533), .Z(n10538) );
  XNOR U10160 ( .A(n10537), .B(n10531), .Z(n10533) );
  XOR U10161 ( .A(n10539), .B(n10540), .Z(n10531) );
  AND U10162 ( .A(n65), .B(n10541), .Z(n10540) );
  XNOR U10163 ( .A(n10542), .B(n10543), .Z(n10537) );
  AND U10164 ( .A(n57), .B(n10544), .Z(n10543) );
  XOR U10165 ( .A(p_input[46]), .B(n10542), .Z(n10544) );
  XNOR U10166 ( .A(n10545), .B(n10546), .Z(n10542) );
  AND U10167 ( .A(n61), .B(n10541), .Z(n10546) );
  XNOR U10168 ( .A(n10545), .B(n10539), .Z(n10541) );
  XOR U10169 ( .A(n10547), .B(n10548), .Z(n10539) );
  AND U10170 ( .A(n76), .B(n10549), .Z(n10548) );
  XNOR U10171 ( .A(n10550), .B(n10551), .Z(n10545) );
  AND U10172 ( .A(n68), .B(n10552), .Z(n10551) );
  XOR U10173 ( .A(p_input[62]), .B(n10550), .Z(n10552) );
  XNOR U10174 ( .A(n10553), .B(n10554), .Z(n10550) );
  AND U10175 ( .A(n72), .B(n10549), .Z(n10554) );
  XNOR U10176 ( .A(n10553), .B(n10547), .Z(n10549) );
  XOR U10177 ( .A(n10555), .B(n10556), .Z(n10547) );
  AND U10178 ( .A(n87), .B(n10557), .Z(n10556) );
  XNOR U10179 ( .A(n10558), .B(n10559), .Z(n10553) );
  AND U10180 ( .A(n79), .B(n10560), .Z(n10559) );
  XOR U10181 ( .A(p_input[78]), .B(n10558), .Z(n10560) );
  XNOR U10182 ( .A(n10561), .B(n10562), .Z(n10558) );
  AND U10183 ( .A(n83), .B(n10557), .Z(n10562) );
  XNOR U10184 ( .A(n10561), .B(n10555), .Z(n10557) );
  XOR U10185 ( .A(n10563), .B(n10564), .Z(n10555) );
  AND U10186 ( .A(n98), .B(n10565), .Z(n10564) );
  XNOR U10187 ( .A(n10566), .B(n10567), .Z(n10561) );
  AND U10188 ( .A(n90), .B(n10568), .Z(n10567) );
  XOR U10189 ( .A(p_input[94]), .B(n10566), .Z(n10568) );
  XNOR U10190 ( .A(n10569), .B(n10570), .Z(n10566) );
  AND U10191 ( .A(n94), .B(n10565), .Z(n10570) );
  XNOR U10192 ( .A(n10569), .B(n10563), .Z(n10565) );
  XOR U10193 ( .A(n10571), .B(n10572), .Z(n10563) );
  AND U10194 ( .A(n109), .B(n10573), .Z(n10572) );
  XNOR U10195 ( .A(n10574), .B(n10575), .Z(n10569) );
  AND U10196 ( .A(n101), .B(n10576), .Z(n10575) );
  XOR U10197 ( .A(p_input[110]), .B(n10574), .Z(n10576) );
  XNOR U10198 ( .A(n10577), .B(n10578), .Z(n10574) );
  AND U10199 ( .A(n105), .B(n10573), .Z(n10578) );
  XNOR U10200 ( .A(n10577), .B(n10571), .Z(n10573) );
  XOR U10201 ( .A(n10579), .B(n10580), .Z(n10571) );
  AND U10202 ( .A(n120), .B(n10581), .Z(n10580) );
  XNOR U10203 ( .A(n10582), .B(n10583), .Z(n10577) );
  AND U10204 ( .A(n112), .B(n10584), .Z(n10583) );
  XOR U10205 ( .A(p_input[126]), .B(n10582), .Z(n10584) );
  XNOR U10206 ( .A(n10585), .B(n10586), .Z(n10582) );
  AND U10207 ( .A(n116), .B(n10581), .Z(n10586) );
  XNOR U10208 ( .A(n10585), .B(n10579), .Z(n10581) );
  XOR U10209 ( .A(n10587), .B(n10588), .Z(n10579) );
  AND U10210 ( .A(n131), .B(n10589), .Z(n10588) );
  XNOR U10211 ( .A(n10590), .B(n10591), .Z(n10585) );
  AND U10212 ( .A(n123), .B(n10592), .Z(n10591) );
  XOR U10213 ( .A(p_input[142]), .B(n10590), .Z(n10592) );
  XNOR U10214 ( .A(n10593), .B(n10594), .Z(n10590) );
  AND U10215 ( .A(n127), .B(n10589), .Z(n10594) );
  XNOR U10216 ( .A(n10593), .B(n10587), .Z(n10589) );
  XOR U10217 ( .A(n10595), .B(n10596), .Z(n10587) );
  AND U10218 ( .A(n142), .B(n10597), .Z(n10596) );
  XNOR U10219 ( .A(n10598), .B(n10599), .Z(n10593) );
  AND U10220 ( .A(n134), .B(n10600), .Z(n10599) );
  XOR U10221 ( .A(p_input[158]), .B(n10598), .Z(n10600) );
  XNOR U10222 ( .A(n10601), .B(n10602), .Z(n10598) );
  AND U10223 ( .A(n138), .B(n10597), .Z(n10602) );
  XNOR U10224 ( .A(n10601), .B(n10595), .Z(n10597) );
  XOR U10225 ( .A(n10603), .B(n10604), .Z(n10595) );
  AND U10226 ( .A(n153), .B(n10605), .Z(n10604) );
  XNOR U10227 ( .A(n10606), .B(n10607), .Z(n10601) );
  AND U10228 ( .A(n145), .B(n10608), .Z(n10607) );
  XOR U10229 ( .A(p_input[174]), .B(n10606), .Z(n10608) );
  XNOR U10230 ( .A(n10609), .B(n10610), .Z(n10606) );
  AND U10231 ( .A(n149), .B(n10605), .Z(n10610) );
  XNOR U10232 ( .A(n10609), .B(n10603), .Z(n10605) );
  XOR U10233 ( .A(n10611), .B(n10612), .Z(n10603) );
  AND U10234 ( .A(n164), .B(n10613), .Z(n10612) );
  XNOR U10235 ( .A(n10614), .B(n10615), .Z(n10609) );
  AND U10236 ( .A(n156), .B(n10616), .Z(n10615) );
  XOR U10237 ( .A(p_input[190]), .B(n10614), .Z(n10616) );
  XNOR U10238 ( .A(n10617), .B(n10618), .Z(n10614) );
  AND U10239 ( .A(n160), .B(n10613), .Z(n10618) );
  XNOR U10240 ( .A(n10617), .B(n10611), .Z(n10613) );
  XOR U10241 ( .A(n10619), .B(n10620), .Z(n10611) );
  AND U10242 ( .A(n175), .B(n10621), .Z(n10620) );
  XNOR U10243 ( .A(n10622), .B(n10623), .Z(n10617) );
  AND U10244 ( .A(n167), .B(n10624), .Z(n10623) );
  XOR U10245 ( .A(p_input[206]), .B(n10622), .Z(n10624) );
  XNOR U10246 ( .A(n10625), .B(n10626), .Z(n10622) );
  AND U10247 ( .A(n171), .B(n10621), .Z(n10626) );
  XNOR U10248 ( .A(n10625), .B(n10619), .Z(n10621) );
  XOR U10249 ( .A(n10627), .B(n10628), .Z(n10619) );
  AND U10250 ( .A(n186), .B(n10629), .Z(n10628) );
  XNOR U10251 ( .A(n10630), .B(n10631), .Z(n10625) );
  AND U10252 ( .A(n178), .B(n10632), .Z(n10631) );
  XOR U10253 ( .A(p_input[222]), .B(n10630), .Z(n10632) );
  XNOR U10254 ( .A(n10633), .B(n10634), .Z(n10630) );
  AND U10255 ( .A(n182), .B(n10629), .Z(n10634) );
  XNOR U10256 ( .A(n10633), .B(n10627), .Z(n10629) );
  XOR U10257 ( .A(n10635), .B(n10636), .Z(n10627) );
  AND U10258 ( .A(n197), .B(n10637), .Z(n10636) );
  XNOR U10259 ( .A(n10638), .B(n10639), .Z(n10633) );
  AND U10260 ( .A(n189), .B(n10640), .Z(n10639) );
  XOR U10261 ( .A(p_input[238]), .B(n10638), .Z(n10640) );
  XNOR U10262 ( .A(n10641), .B(n10642), .Z(n10638) );
  AND U10263 ( .A(n193), .B(n10637), .Z(n10642) );
  XNOR U10264 ( .A(n10641), .B(n10635), .Z(n10637) );
  XOR U10265 ( .A(n10643), .B(n10644), .Z(n10635) );
  AND U10266 ( .A(n208), .B(n10645), .Z(n10644) );
  XNOR U10267 ( .A(n10646), .B(n10647), .Z(n10641) );
  AND U10268 ( .A(n200), .B(n10648), .Z(n10647) );
  XOR U10269 ( .A(p_input[254]), .B(n10646), .Z(n10648) );
  XNOR U10270 ( .A(n10649), .B(n10650), .Z(n10646) );
  AND U10271 ( .A(n204), .B(n10645), .Z(n10650) );
  XNOR U10272 ( .A(n10649), .B(n10643), .Z(n10645) );
  XOR U10273 ( .A(n10651), .B(n10652), .Z(n10643) );
  AND U10274 ( .A(n219), .B(n10653), .Z(n10652) );
  XNOR U10275 ( .A(n10654), .B(n10655), .Z(n10649) );
  AND U10276 ( .A(n211), .B(n10656), .Z(n10655) );
  XOR U10277 ( .A(p_input[270]), .B(n10654), .Z(n10656) );
  XNOR U10278 ( .A(n10657), .B(n10658), .Z(n10654) );
  AND U10279 ( .A(n215), .B(n10653), .Z(n10658) );
  XNOR U10280 ( .A(n10657), .B(n10651), .Z(n10653) );
  XOR U10281 ( .A(n10659), .B(n10660), .Z(n10651) );
  AND U10282 ( .A(n230), .B(n10661), .Z(n10660) );
  XNOR U10283 ( .A(n10662), .B(n10663), .Z(n10657) );
  AND U10284 ( .A(n222), .B(n10664), .Z(n10663) );
  XOR U10285 ( .A(p_input[286]), .B(n10662), .Z(n10664) );
  XNOR U10286 ( .A(n10665), .B(n10666), .Z(n10662) );
  AND U10287 ( .A(n226), .B(n10661), .Z(n10666) );
  XNOR U10288 ( .A(n10665), .B(n10659), .Z(n10661) );
  XOR U10289 ( .A(n10667), .B(n10668), .Z(n10659) );
  AND U10290 ( .A(n241), .B(n10669), .Z(n10668) );
  XNOR U10291 ( .A(n10670), .B(n10671), .Z(n10665) );
  AND U10292 ( .A(n233), .B(n10672), .Z(n10671) );
  XOR U10293 ( .A(p_input[302]), .B(n10670), .Z(n10672) );
  XNOR U10294 ( .A(n10673), .B(n10674), .Z(n10670) );
  AND U10295 ( .A(n237), .B(n10669), .Z(n10674) );
  XNOR U10296 ( .A(n10673), .B(n10667), .Z(n10669) );
  XOR U10297 ( .A(n10675), .B(n10676), .Z(n10667) );
  AND U10298 ( .A(n252), .B(n10677), .Z(n10676) );
  XNOR U10299 ( .A(n10678), .B(n10679), .Z(n10673) );
  AND U10300 ( .A(n244), .B(n10680), .Z(n10679) );
  XOR U10301 ( .A(p_input[318]), .B(n10678), .Z(n10680) );
  XNOR U10302 ( .A(n10681), .B(n10682), .Z(n10678) );
  AND U10303 ( .A(n248), .B(n10677), .Z(n10682) );
  XNOR U10304 ( .A(n10681), .B(n10675), .Z(n10677) );
  XOR U10305 ( .A(n10683), .B(n10684), .Z(n10675) );
  AND U10306 ( .A(n263), .B(n10685), .Z(n10684) );
  XNOR U10307 ( .A(n10686), .B(n10687), .Z(n10681) );
  AND U10308 ( .A(n255), .B(n10688), .Z(n10687) );
  XOR U10309 ( .A(p_input[334]), .B(n10686), .Z(n10688) );
  XNOR U10310 ( .A(n10689), .B(n10690), .Z(n10686) );
  AND U10311 ( .A(n259), .B(n10685), .Z(n10690) );
  XNOR U10312 ( .A(n10689), .B(n10683), .Z(n10685) );
  XOR U10313 ( .A(n10691), .B(n10692), .Z(n10683) );
  AND U10314 ( .A(n274), .B(n10693), .Z(n10692) );
  XNOR U10315 ( .A(n10694), .B(n10695), .Z(n10689) );
  AND U10316 ( .A(n266), .B(n10696), .Z(n10695) );
  XOR U10317 ( .A(p_input[350]), .B(n10694), .Z(n10696) );
  XNOR U10318 ( .A(n10697), .B(n10698), .Z(n10694) );
  AND U10319 ( .A(n270), .B(n10693), .Z(n10698) );
  XNOR U10320 ( .A(n10697), .B(n10691), .Z(n10693) );
  XOR U10321 ( .A(n10699), .B(n10700), .Z(n10691) );
  AND U10322 ( .A(n285), .B(n10701), .Z(n10700) );
  XNOR U10323 ( .A(n10702), .B(n10703), .Z(n10697) );
  AND U10324 ( .A(n277), .B(n10704), .Z(n10703) );
  XOR U10325 ( .A(p_input[366]), .B(n10702), .Z(n10704) );
  XNOR U10326 ( .A(n10705), .B(n10706), .Z(n10702) );
  AND U10327 ( .A(n281), .B(n10701), .Z(n10706) );
  XNOR U10328 ( .A(n10705), .B(n10699), .Z(n10701) );
  XOR U10329 ( .A(n10707), .B(n10708), .Z(n10699) );
  AND U10330 ( .A(n296), .B(n10709), .Z(n10708) );
  XNOR U10331 ( .A(n10710), .B(n10711), .Z(n10705) );
  AND U10332 ( .A(n288), .B(n10712), .Z(n10711) );
  XOR U10333 ( .A(p_input[382]), .B(n10710), .Z(n10712) );
  XNOR U10334 ( .A(n10713), .B(n10714), .Z(n10710) );
  AND U10335 ( .A(n292), .B(n10709), .Z(n10714) );
  XNOR U10336 ( .A(n10713), .B(n10707), .Z(n10709) );
  XOR U10337 ( .A(n10715), .B(n10716), .Z(n10707) );
  AND U10338 ( .A(n307), .B(n10717), .Z(n10716) );
  XNOR U10339 ( .A(n10718), .B(n10719), .Z(n10713) );
  AND U10340 ( .A(n299), .B(n10720), .Z(n10719) );
  XOR U10341 ( .A(p_input[398]), .B(n10718), .Z(n10720) );
  XNOR U10342 ( .A(n10721), .B(n10722), .Z(n10718) );
  AND U10343 ( .A(n303), .B(n10717), .Z(n10722) );
  XNOR U10344 ( .A(n10721), .B(n10715), .Z(n10717) );
  XOR U10345 ( .A(n10723), .B(n10724), .Z(n10715) );
  AND U10346 ( .A(n318), .B(n10725), .Z(n10724) );
  XNOR U10347 ( .A(n10726), .B(n10727), .Z(n10721) );
  AND U10348 ( .A(n310), .B(n10728), .Z(n10727) );
  XOR U10349 ( .A(p_input[414]), .B(n10726), .Z(n10728) );
  XNOR U10350 ( .A(n10729), .B(n10730), .Z(n10726) );
  AND U10351 ( .A(n314), .B(n10725), .Z(n10730) );
  XNOR U10352 ( .A(n10729), .B(n10723), .Z(n10725) );
  XOR U10353 ( .A(n10731), .B(n10732), .Z(n10723) );
  AND U10354 ( .A(n329), .B(n10733), .Z(n10732) );
  XNOR U10355 ( .A(n10734), .B(n10735), .Z(n10729) );
  AND U10356 ( .A(n321), .B(n10736), .Z(n10735) );
  XOR U10357 ( .A(p_input[430]), .B(n10734), .Z(n10736) );
  XNOR U10358 ( .A(n10737), .B(n10738), .Z(n10734) );
  AND U10359 ( .A(n325), .B(n10733), .Z(n10738) );
  XNOR U10360 ( .A(n10737), .B(n10731), .Z(n10733) );
  XOR U10361 ( .A(n10739), .B(n10740), .Z(n10731) );
  AND U10362 ( .A(n340), .B(n10741), .Z(n10740) );
  XNOR U10363 ( .A(n10742), .B(n10743), .Z(n10737) );
  AND U10364 ( .A(n332), .B(n10744), .Z(n10743) );
  XOR U10365 ( .A(p_input[446]), .B(n10742), .Z(n10744) );
  XNOR U10366 ( .A(n10745), .B(n10746), .Z(n10742) );
  AND U10367 ( .A(n336), .B(n10741), .Z(n10746) );
  XNOR U10368 ( .A(n10745), .B(n10739), .Z(n10741) );
  XOR U10369 ( .A(n10747), .B(n10748), .Z(n10739) );
  AND U10370 ( .A(n351), .B(n10749), .Z(n10748) );
  XNOR U10371 ( .A(n10750), .B(n10751), .Z(n10745) );
  AND U10372 ( .A(n343), .B(n10752), .Z(n10751) );
  XOR U10373 ( .A(p_input[462]), .B(n10750), .Z(n10752) );
  XNOR U10374 ( .A(n10753), .B(n10754), .Z(n10750) );
  AND U10375 ( .A(n347), .B(n10749), .Z(n10754) );
  XNOR U10376 ( .A(n10753), .B(n10747), .Z(n10749) );
  XOR U10377 ( .A(n10755), .B(n10756), .Z(n10747) );
  AND U10378 ( .A(n362), .B(n10757), .Z(n10756) );
  XNOR U10379 ( .A(n10758), .B(n10759), .Z(n10753) );
  AND U10380 ( .A(n354), .B(n10760), .Z(n10759) );
  XOR U10381 ( .A(p_input[478]), .B(n10758), .Z(n10760) );
  XNOR U10382 ( .A(n10761), .B(n10762), .Z(n10758) );
  AND U10383 ( .A(n358), .B(n10757), .Z(n10762) );
  XNOR U10384 ( .A(n10761), .B(n10755), .Z(n10757) );
  XOR U10385 ( .A(n10763), .B(n10764), .Z(n10755) );
  AND U10386 ( .A(n373), .B(n10765), .Z(n10764) );
  XNOR U10387 ( .A(n10766), .B(n10767), .Z(n10761) );
  AND U10388 ( .A(n365), .B(n10768), .Z(n10767) );
  XOR U10389 ( .A(p_input[494]), .B(n10766), .Z(n10768) );
  XNOR U10390 ( .A(n10769), .B(n10770), .Z(n10766) );
  AND U10391 ( .A(n369), .B(n10765), .Z(n10770) );
  XNOR U10392 ( .A(n10769), .B(n10763), .Z(n10765) );
  XOR U10393 ( .A(n10771), .B(n10772), .Z(n10763) );
  AND U10394 ( .A(n384), .B(n10773), .Z(n10772) );
  XNOR U10395 ( .A(n10774), .B(n10775), .Z(n10769) );
  AND U10396 ( .A(n376), .B(n10776), .Z(n10775) );
  XOR U10397 ( .A(p_input[510]), .B(n10774), .Z(n10776) );
  XNOR U10398 ( .A(n10777), .B(n10778), .Z(n10774) );
  AND U10399 ( .A(n380), .B(n10773), .Z(n10778) );
  XNOR U10400 ( .A(n10777), .B(n10771), .Z(n10773) );
  XOR U10401 ( .A(n10779), .B(n10780), .Z(n10771) );
  AND U10402 ( .A(n395), .B(n10781), .Z(n10780) );
  XNOR U10403 ( .A(n10782), .B(n10783), .Z(n10777) );
  AND U10404 ( .A(n387), .B(n10784), .Z(n10783) );
  XOR U10405 ( .A(p_input[526]), .B(n10782), .Z(n10784) );
  XNOR U10406 ( .A(n10785), .B(n10786), .Z(n10782) );
  AND U10407 ( .A(n391), .B(n10781), .Z(n10786) );
  XNOR U10408 ( .A(n10785), .B(n10779), .Z(n10781) );
  XOR U10409 ( .A(n10787), .B(n10788), .Z(n10779) );
  AND U10410 ( .A(n406), .B(n10789), .Z(n10788) );
  XNOR U10411 ( .A(n10790), .B(n10791), .Z(n10785) );
  AND U10412 ( .A(n398), .B(n10792), .Z(n10791) );
  XOR U10413 ( .A(p_input[542]), .B(n10790), .Z(n10792) );
  XNOR U10414 ( .A(n10793), .B(n10794), .Z(n10790) );
  AND U10415 ( .A(n402), .B(n10789), .Z(n10794) );
  XNOR U10416 ( .A(n10793), .B(n10787), .Z(n10789) );
  XOR U10417 ( .A(n10795), .B(n10796), .Z(n10787) );
  AND U10418 ( .A(n417), .B(n10797), .Z(n10796) );
  XNOR U10419 ( .A(n10798), .B(n10799), .Z(n10793) );
  AND U10420 ( .A(n409), .B(n10800), .Z(n10799) );
  XOR U10421 ( .A(p_input[558]), .B(n10798), .Z(n10800) );
  XNOR U10422 ( .A(n10801), .B(n10802), .Z(n10798) );
  AND U10423 ( .A(n413), .B(n10797), .Z(n10802) );
  XNOR U10424 ( .A(n10801), .B(n10795), .Z(n10797) );
  XOR U10425 ( .A(n10803), .B(n10804), .Z(n10795) );
  AND U10426 ( .A(n428), .B(n10805), .Z(n10804) );
  XNOR U10427 ( .A(n10806), .B(n10807), .Z(n10801) );
  AND U10428 ( .A(n420), .B(n10808), .Z(n10807) );
  XOR U10429 ( .A(p_input[574]), .B(n10806), .Z(n10808) );
  XNOR U10430 ( .A(n10809), .B(n10810), .Z(n10806) );
  AND U10431 ( .A(n424), .B(n10805), .Z(n10810) );
  XNOR U10432 ( .A(n10809), .B(n10803), .Z(n10805) );
  XOR U10433 ( .A(n10811), .B(n10812), .Z(n10803) );
  AND U10434 ( .A(n439), .B(n10813), .Z(n10812) );
  XNOR U10435 ( .A(n10814), .B(n10815), .Z(n10809) );
  AND U10436 ( .A(n431), .B(n10816), .Z(n10815) );
  XOR U10437 ( .A(p_input[590]), .B(n10814), .Z(n10816) );
  XNOR U10438 ( .A(n10817), .B(n10818), .Z(n10814) );
  AND U10439 ( .A(n435), .B(n10813), .Z(n10818) );
  XNOR U10440 ( .A(n10817), .B(n10811), .Z(n10813) );
  XOR U10441 ( .A(n10819), .B(n10820), .Z(n10811) );
  AND U10442 ( .A(n450), .B(n10821), .Z(n10820) );
  XNOR U10443 ( .A(n10822), .B(n10823), .Z(n10817) );
  AND U10444 ( .A(n442), .B(n10824), .Z(n10823) );
  XOR U10445 ( .A(p_input[606]), .B(n10822), .Z(n10824) );
  XNOR U10446 ( .A(n10825), .B(n10826), .Z(n10822) );
  AND U10447 ( .A(n446), .B(n10821), .Z(n10826) );
  XNOR U10448 ( .A(n10825), .B(n10819), .Z(n10821) );
  XOR U10449 ( .A(n10827), .B(n10828), .Z(n10819) );
  AND U10450 ( .A(n461), .B(n10829), .Z(n10828) );
  XNOR U10451 ( .A(n10830), .B(n10831), .Z(n10825) );
  AND U10452 ( .A(n453), .B(n10832), .Z(n10831) );
  XOR U10453 ( .A(p_input[622]), .B(n10830), .Z(n10832) );
  XNOR U10454 ( .A(n10833), .B(n10834), .Z(n10830) );
  AND U10455 ( .A(n457), .B(n10829), .Z(n10834) );
  XNOR U10456 ( .A(n10833), .B(n10827), .Z(n10829) );
  XOR U10457 ( .A(n10835), .B(n10836), .Z(n10827) );
  AND U10458 ( .A(n472), .B(n10837), .Z(n10836) );
  XNOR U10459 ( .A(n10838), .B(n10839), .Z(n10833) );
  AND U10460 ( .A(n464), .B(n10840), .Z(n10839) );
  XOR U10461 ( .A(p_input[638]), .B(n10838), .Z(n10840) );
  XNOR U10462 ( .A(n10841), .B(n10842), .Z(n10838) );
  AND U10463 ( .A(n468), .B(n10837), .Z(n10842) );
  XNOR U10464 ( .A(n10841), .B(n10835), .Z(n10837) );
  XOR U10465 ( .A(n10843), .B(n10844), .Z(n10835) );
  AND U10466 ( .A(n483), .B(n10845), .Z(n10844) );
  XNOR U10467 ( .A(n10846), .B(n10847), .Z(n10841) );
  AND U10468 ( .A(n475), .B(n10848), .Z(n10847) );
  XOR U10469 ( .A(p_input[654]), .B(n10846), .Z(n10848) );
  XNOR U10470 ( .A(n10849), .B(n10850), .Z(n10846) );
  AND U10471 ( .A(n479), .B(n10845), .Z(n10850) );
  XNOR U10472 ( .A(n10849), .B(n10843), .Z(n10845) );
  XOR U10473 ( .A(n10851), .B(n10852), .Z(n10843) );
  AND U10474 ( .A(n494), .B(n10853), .Z(n10852) );
  XNOR U10475 ( .A(n10854), .B(n10855), .Z(n10849) );
  AND U10476 ( .A(n486), .B(n10856), .Z(n10855) );
  XOR U10477 ( .A(p_input[670]), .B(n10854), .Z(n10856) );
  XNOR U10478 ( .A(n10857), .B(n10858), .Z(n10854) );
  AND U10479 ( .A(n490), .B(n10853), .Z(n10858) );
  XNOR U10480 ( .A(n10857), .B(n10851), .Z(n10853) );
  XOR U10481 ( .A(n10859), .B(n10860), .Z(n10851) );
  AND U10482 ( .A(n505), .B(n10861), .Z(n10860) );
  XNOR U10483 ( .A(n10862), .B(n10863), .Z(n10857) );
  AND U10484 ( .A(n497), .B(n10864), .Z(n10863) );
  XOR U10485 ( .A(p_input[686]), .B(n10862), .Z(n10864) );
  XNOR U10486 ( .A(n10865), .B(n10866), .Z(n10862) );
  AND U10487 ( .A(n501), .B(n10861), .Z(n10866) );
  XNOR U10488 ( .A(n10865), .B(n10859), .Z(n10861) );
  XOR U10489 ( .A(n10867), .B(n10868), .Z(n10859) );
  AND U10490 ( .A(n516), .B(n10869), .Z(n10868) );
  XNOR U10491 ( .A(n10870), .B(n10871), .Z(n10865) );
  AND U10492 ( .A(n508), .B(n10872), .Z(n10871) );
  XOR U10493 ( .A(p_input[702]), .B(n10870), .Z(n10872) );
  XNOR U10494 ( .A(n10873), .B(n10874), .Z(n10870) );
  AND U10495 ( .A(n512), .B(n10869), .Z(n10874) );
  XNOR U10496 ( .A(n10873), .B(n10867), .Z(n10869) );
  XOR U10497 ( .A(n10875), .B(n10876), .Z(n10867) );
  AND U10498 ( .A(n527), .B(n10877), .Z(n10876) );
  XNOR U10499 ( .A(n10878), .B(n10879), .Z(n10873) );
  AND U10500 ( .A(n519), .B(n10880), .Z(n10879) );
  XOR U10501 ( .A(p_input[718]), .B(n10878), .Z(n10880) );
  XNOR U10502 ( .A(n10881), .B(n10882), .Z(n10878) );
  AND U10503 ( .A(n523), .B(n10877), .Z(n10882) );
  XNOR U10504 ( .A(n10881), .B(n10875), .Z(n10877) );
  XOR U10505 ( .A(n10883), .B(n10884), .Z(n10875) );
  AND U10506 ( .A(n538), .B(n10885), .Z(n10884) );
  XNOR U10507 ( .A(n10886), .B(n10887), .Z(n10881) );
  AND U10508 ( .A(n530), .B(n10888), .Z(n10887) );
  XOR U10509 ( .A(p_input[734]), .B(n10886), .Z(n10888) );
  XNOR U10510 ( .A(n10889), .B(n10890), .Z(n10886) );
  AND U10511 ( .A(n534), .B(n10885), .Z(n10890) );
  XNOR U10512 ( .A(n10889), .B(n10883), .Z(n10885) );
  XOR U10513 ( .A(n10891), .B(n10892), .Z(n10883) );
  AND U10514 ( .A(n549), .B(n10893), .Z(n10892) );
  XNOR U10515 ( .A(n10894), .B(n10895), .Z(n10889) );
  AND U10516 ( .A(n541), .B(n10896), .Z(n10895) );
  XOR U10517 ( .A(p_input[750]), .B(n10894), .Z(n10896) );
  XNOR U10518 ( .A(n10897), .B(n10898), .Z(n10894) );
  AND U10519 ( .A(n545), .B(n10893), .Z(n10898) );
  XNOR U10520 ( .A(n10897), .B(n10891), .Z(n10893) );
  XOR U10521 ( .A(n10899), .B(n10900), .Z(n10891) );
  AND U10522 ( .A(n560), .B(n10901), .Z(n10900) );
  XNOR U10523 ( .A(n10902), .B(n10903), .Z(n10897) );
  AND U10524 ( .A(n552), .B(n10904), .Z(n10903) );
  XOR U10525 ( .A(p_input[766]), .B(n10902), .Z(n10904) );
  XNOR U10526 ( .A(n10905), .B(n10906), .Z(n10902) );
  AND U10527 ( .A(n556), .B(n10901), .Z(n10906) );
  XNOR U10528 ( .A(n10905), .B(n10899), .Z(n10901) );
  XOR U10529 ( .A(n10907), .B(n10908), .Z(n10899) );
  AND U10530 ( .A(n571), .B(n10909), .Z(n10908) );
  XNOR U10531 ( .A(n10910), .B(n10911), .Z(n10905) );
  AND U10532 ( .A(n563), .B(n10912), .Z(n10911) );
  XOR U10533 ( .A(p_input[782]), .B(n10910), .Z(n10912) );
  XNOR U10534 ( .A(n10913), .B(n10914), .Z(n10910) );
  AND U10535 ( .A(n567), .B(n10909), .Z(n10914) );
  XNOR U10536 ( .A(n10913), .B(n10907), .Z(n10909) );
  XOR U10537 ( .A(n10915), .B(n10916), .Z(n10907) );
  AND U10538 ( .A(n582), .B(n10917), .Z(n10916) );
  XNOR U10539 ( .A(n10918), .B(n10919), .Z(n10913) );
  AND U10540 ( .A(n574), .B(n10920), .Z(n10919) );
  XOR U10541 ( .A(p_input[798]), .B(n10918), .Z(n10920) );
  XNOR U10542 ( .A(n10921), .B(n10922), .Z(n10918) );
  AND U10543 ( .A(n578), .B(n10917), .Z(n10922) );
  XNOR U10544 ( .A(n10921), .B(n10915), .Z(n10917) );
  XOR U10545 ( .A(n10923), .B(n10924), .Z(n10915) );
  AND U10546 ( .A(n593), .B(n10925), .Z(n10924) );
  XNOR U10547 ( .A(n10926), .B(n10927), .Z(n10921) );
  AND U10548 ( .A(n585), .B(n10928), .Z(n10927) );
  XOR U10549 ( .A(p_input[814]), .B(n10926), .Z(n10928) );
  XNOR U10550 ( .A(n10929), .B(n10930), .Z(n10926) );
  AND U10551 ( .A(n589), .B(n10925), .Z(n10930) );
  XNOR U10552 ( .A(n10929), .B(n10923), .Z(n10925) );
  XOR U10553 ( .A(n10931), .B(n10932), .Z(n10923) );
  AND U10554 ( .A(n604), .B(n10933), .Z(n10932) );
  XNOR U10555 ( .A(n10934), .B(n10935), .Z(n10929) );
  AND U10556 ( .A(n596), .B(n10936), .Z(n10935) );
  XOR U10557 ( .A(p_input[830]), .B(n10934), .Z(n10936) );
  XNOR U10558 ( .A(n10937), .B(n10938), .Z(n10934) );
  AND U10559 ( .A(n600), .B(n10933), .Z(n10938) );
  XNOR U10560 ( .A(n10937), .B(n10931), .Z(n10933) );
  XOR U10561 ( .A(n10939), .B(n10940), .Z(n10931) );
  AND U10562 ( .A(n615), .B(n10941), .Z(n10940) );
  XNOR U10563 ( .A(n10942), .B(n10943), .Z(n10937) );
  AND U10564 ( .A(n607), .B(n10944), .Z(n10943) );
  XOR U10565 ( .A(p_input[846]), .B(n10942), .Z(n10944) );
  XNOR U10566 ( .A(n10945), .B(n10946), .Z(n10942) );
  AND U10567 ( .A(n611), .B(n10941), .Z(n10946) );
  XNOR U10568 ( .A(n10945), .B(n10939), .Z(n10941) );
  XOR U10569 ( .A(n10947), .B(n10948), .Z(n10939) );
  AND U10570 ( .A(n626), .B(n10949), .Z(n10948) );
  XNOR U10571 ( .A(n10950), .B(n10951), .Z(n10945) );
  AND U10572 ( .A(n618), .B(n10952), .Z(n10951) );
  XOR U10573 ( .A(p_input[862]), .B(n10950), .Z(n10952) );
  XNOR U10574 ( .A(n10953), .B(n10954), .Z(n10950) );
  AND U10575 ( .A(n622), .B(n10949), .Z(n10954) );
  XNOR U10576 ( .A(n10953), .B(n10947), .Z(n10949) );
  XOR U10577 ( .A(n10955), .B(n10956), .Z(n10947) );
  AND U10578 ( .A(n637), .B(n10957), .Z(n10956) );
  XNOR U10579 ( .A(n10958), .B(n10959), .Z(n10953) );
  AND U10580 ( .A(n629), .B(n10960), .Z(n10959) );
  XOR U10581 ( .A(p_input[878]), .B(n10958), .Z(n10960) );
  XNOR U10582 ( .A(n10961), .B(n10962), .Z(n10958) );
  AND U10583 ( .A(n633), .B(n10957), .Z(n10962) );
  XNOR U10584 ( .A(n10961), .B(n10955), .Z(n10957) );
  XOR U10585 ( .A(n10963), .B(n10964), .Z(n10955) );
  AND U10586 ( .A(n648), .B(n10965), .Z(n10964) );
  XNOR U10587 ( .A(n10966), .B(n10967), .Z(n10961) );
  AND U10588 ( .A(n640), .B(n10968), .Z(n10967) );
  XOR U10589 ( .A(p_input[894]), .B(n10966), .Z(n10968) );
  XNOR U10590 ( .A(n10969), .B(n10970), .Z(n10966) );
  AND U10591 ( .A(n644), .B(n10965), .Z(n10970) );
  XNOR U10592 ( .A(n10969), .B(n10963), .Z(n10965) );
  XOR U10593 ( .A(n10971), .B(n10972), .Z(n10963) );
  AND U10594 ( .A(n659), .B(n10973), .Z(n10972) );
  XNOR U10595 ( .A(n10974), .B(n10975), .Z(n10969) );
  AND U10596 ( .A(n651), .B(n10976), .Z(n10975) );
  XOR U10597 ( .A(p_input[910]), .B(n10974), .Z(n10976) );
  XNOR U10598 ( .A(n10977), .B(n10978), .Z(n10974) );
  AND U10599 ( .A(n655), .B(n10973), .Z(n10978) );
  XNOR U10600 ( .A(n10977), .B(n10971), .Z(n10973) );
  XOR U10601 ( .A(n10979), .B(n10980), .Z(n10971) );
  AND U10602 ( .A(n670), .B(n10981), .Z(n10980) );
  XNOR U10603 ( .A(n10982), .B(n10983), .Z(n10977) );
  AND U10604 ( .A(n662), .B(n10984), .Z(n10983) );
  XOR U10605 ( .A(p_input[926]), .B(n10982), .Z(n10984) );
  XNOR U10606 ( .A(n10985), .B(n10986), .Z(n10982) );
  AND U10607 ( .A(n666), .B(n10981), .Z(n10986) );
  XNOR U10608 ( .A(n10985), .B(n10979), .Z(n10981) );
  XOR U10609 ( .A(n10987), .B(n10988), .Z(n10979) );
  AND U10610 ( .A(n681), .B(n10989), .Z(n10988) );
  XNOR U10611 ( .A(n10990), .B(n10991), .Z(n10985) );
  AND U10612 ( .A(n673), .B(n10992), .Z(n10991) );
  XOR U10613 ( .A(p_input[942]), .B(n10990), .Z(n10992) );
  XNOR U10614 ( .A(n10993), .B(n10994), .Z(n10990) );
  AND U10615 ( .A(n677), .B(n10989), .Z(n10994) );
  XNOR U10616 ( .A(n10993), .B(n10987), .Z(n10989) );
  XOR U10617 ( .A(n10995), .B(n10996), .Z(n10987) );
  AND U10618 ( .A(n692), .B(n10997), .Z(n10996) );
  XNOR U10619 ( .A(n10998), .B(n10999), .Z(n10993) );
  AND U10620 ( .A(n684), .B(n11000), .Z(n10999) );
  XOR U10621 ( .A(p_input[958]), .B(n10998), .Z(n11000) );
  XNOR U10622 ( .A(n11001), .B(n11002), .Z(n10998) );
  AND U10623 ( .A(n688), .B(n10997), .Z(n11002) );
  XNOR U10624 ( .A(n11001), .B(n10995), .Z(n10997) );
  XOR U10625 ( .A(n11003), .B(n11004), .Z(n10995) );
  AND U10626 ( .A(n703), .B(n11005), .Z(n11004) );
  XNOR U10627 ( .A(n11006), .B(n11007), .Z(n11001) );
  AND U10628 ( .A(n695), .B(n11008), .Z(n11007) );
  XOR U10629 ( .A(p_input[974]), .B(n11006), .Z(n11008) );
  XNOR U10630 ( .A(n11009), .B(n11010), .Z(n11006) );
  AND U10631 ( .A(n699), .B(n11005), .Z(n11010) );
  XNOR U10632 ( .A(n11009), .B(n11003), .Z(n11005) );
  XOR U10633 ( .A(n11011), .B(n11012), .Z(n11003) );
  AND U10634 ( .A(n714), .B(n11013), .Z(n11012) );
  XNOR U10635 ( .A(n11014), .B(n11015), .Z(n11009) );
  AND U10636 ( .A(n706), .B(n11016), .Z(n11015) );
  XOR U10637 ( .A(p_input[990]), .B(n11014), .Z(n11016) );
  XNOR U10638 ( .A(n11017), .B(n11018), .Z(n11014) );
  AND U10639 ( .A(n710), .B(n11013), .Z(n11018) );
  XNOR U10640 ( .A(n11017), .B(n11011), .Z(n11013) );
  XOR U10641 ( .A(n11019), .B(n11020), .Z(n11011) );
  AND U10642 ( .A(n725), .B(n11021), .Z(n11020) );
  XNOR U10643 ( .A(n11022), .B(n11023), .Z(n11017) );
  AND U10644 ( .A(n717), .B(n11024), .Z(n11023) );
  XOR U10645 ( .A(p_input[1006]), .B(n11022), .Z(n11024) );
  XNOR U10646 ( .A(n11025), .B(n11026), .Z(n11022) );
  AND U10647 ( .A(n721), .B(n11021), .Z(n11026) );
  XNOR U10648 ( .A(n11025), .B(n11019), .Z(n11021) );
  XOR U10649 ( .A(n11027), .B(n11028), .Z(n11019) );
  AND U10650 ( .A(n736), .B(n11029), .Z(n11028) );
  XNOR U10651 ( .A(n11030), .B(n11031), .Z(n11025) );
  AND U10652 ( .A(n728), .B(n11032), .Z(n11031) );
  XOR U10653 ( .A(p_input[1022]), .B(n11030), .Z(n11032) );
  XNOR U10654 ( .A(n11033), .B(n11034), .Z(n11030) );
  AND U10655 ( .A(n732), .B(n11029), .Z(n11034) );
  XNOR U10656 ( .A(n11033), .B(n11027), .Z(n11029) );
  XOR U10657 ( .A(n11035), .B(n11036), .Z(n11027) );
  AND U10658 ( .A(n747), .B(n11037), .Z(n11036) );
  XNOR U10659 ( .A(n11038), .B(n11039), .Z(n11033) );
  AND U10660 ( .A(n739), .B(n11040), .Z(n11039) );
  XOR U10661 ( .A(p_input[1038]), .B(n11038), .Z(n11040) );
  XNOR U10662 ( .A(n11041), .B(n11042), .Z(n11038) );
  AND U10663 ( .A(n743), .B(n11037), .Z(n11042) );
  XNOR U10664 ( .A(n11041), .B(n11035), .Z(n11037) );
  XOR U10665 ( .A(n11043), .B(n11044), .Z(n11035) );
  AND U10666 ( .A(n758), .B(n11045), .Z(n11044) );
  XNOR U10667 ( .A(n11046), .B(n11047), .Z(n11041) );
  AND U10668 ( .A(n750), .B(n11048), .Z(n11047) );
  XOR U10669 ( .A(p_input[1054]), .B(n11046), .Z(n11048) );
  XNOR U10670 ( .A(n11049), .B(n11050), .Z(n11046) );
  AND U10671 ( .A(n754), .B(n11045), .Z(n11050) );
  XNOR U10672 ( .A(n11049), .B(n11043), .Z(n11045) );
  XOR U10673 ( .A(n11051), .B(n11052), .Z(n11043) );
  AND U10674 ( .A(n769), .B(n11053), .Z(n11052) );
  XNOR U10675 ( .A(n11054), .B(n11055), .Z(n11049) );
  AND U10676 ( .A(n761), .B(n11056), .Z(n11055) );
  XOR U10677 ( .A(p_input[1070]), .B(n11054), .Z(n11056) );
  XNOR U10678 ( .A(n11057), .B(n11058), .Z(n11054) );
  AND U10679 ( .A(n765), .B(n11053), .Z(n11058) );
  XNOR U10680 ( .A(n11057), .B(n11051), .Z(n11053) );
  XOR U10681 ( .A(n11059), .B(n11060), .Z(n11051) );
  AND U10682 ( .A(n780), .B(n11061), .Z(n11060) );
  XNOR U10683 ( .A(n11062), .B(n11063), .Z(n11057) );
  AND U10684 ( .A(n772), .B(n11064), .Z(n11063) );
  XOR U10685 ( .A(p_input[1086]), .B(n11062), .Z(n11064) );
  XNOR U10686 ( .A(n11065), .B(n11066), .Z(n11062) );
  AND U10687 ( .A(n776), .B(n11061), .Z(n11066) );
  XNOR U10688 ( .A(n11065), .B(n11059), .Z(n11061) );
  XOR U10689 ( .A(n11067), .B(n11068), .Z(n11059) );
  AND U10690 ( .A(n791), .B(n11069), .Z(n11068) );
  XNOR U10691 ( .A(n11070), .B(n11071), .Z(n11065) );
  AND U10692 ( .A(n783), .B(n11072), .Z(n11071) );
  XOR U10693 ( .A(p_input[1102]), .B(n11070), .Z(n11072) );
  XNOR U10694 ( .A(n11073), .B(n11074), .Z(n11070) );
  AND U10695 ( .A(n787), .B(n11069), .Z(n11074) );
  XNOR U10696 ( .A(n11073), .B(n11067), .Z(n11069) );
  XOR U10697 ( .A(n11075), .B(n11076), .Z(n11067) );
  AND U10698 ( .A(n802), .B(n11077), .Z(n11076) );
  XNOR U10699 ( .A(n11078), .B(n11079), .Z(n11073) );
  AND U10700 ( .A(n794), .B(n11080), .Z(n11079) );
  XOR U10701 ( .A(p_input[1118]), .B(n11078), .Z(n11080) );
  XNOR U10702 ( .A(n11081), .B(n11082), .Z(n11078) );
  AND U10703 ( .A(n798), .B(n11077), .Z(n11082) );
  XNOR U10704 ( .A(n11081), .B(n11075), .Z(n11077) );
  XOR U10705 ( .A(n11083), .B(n11084), .Z(n11075) );
  AND U10706 ( .A(n813), .B(n11085), .Z(n11084) );
  XNOR U10707 ( .A(n11086), .B(n11087), .Z(n11081) );
  AND U10708 ( .A(n805), .B(n11088), .Z(n11087) );
  XOR U10709 ( .A(p_input[1134]), .B(n11086), .Z(n11088) );
  XNOR U10710 ( .A(n11089), .B(n11090), .Z(n11086) );
  AND U10711 ( .A(n809), .B(n11085), .Z(n11090) );
  XNOR U10712 ( .A(n11089), .B(n11083), .Z(n11085) );
  XOR U10713 ( .A(n11091), .B(n11092), .Z(n11083) );
  AND U10714 ( .A(n824), .B(n11093), .Z(n11092) );
  XNOR U10715 ( .A(n11094), .B(n11095), .Z(n11089) );
  AND U10716 ( .A(n816), .B(n11096), .Z(n11095) );
  XOR U10717 ( .A(p_input[1150]), .B(n11094), .Z(n11096) );
  XNOR U10718 ( .A(n11097), .B(n11098), .Z(n11094) );
  AND U10719 ( .A(n820), .B(n11093), .Z(n11098) );
  XNOR U10720 ( .A(n11097), .B(n11091), .Z(n11093) );
  XOR U10721 ( .A(n11099), .B(n11100), .Z(n11091) );
  AND U10722 ( .A(n835), .B(n11101), .Z(n11100) );
  XNOR U10723 ( .A(n11102), .B(n11103), .Z(n11097) );
  AND U10724 ( .A(n827), .B(n11104), .Z(n11103) );
  XOR U10725 ( .A(p_input[1166]), .B(n11102), .Z(n11104) );
  XNOR U10726 ( .A(n11105), .B(n11106), .Z(n11102) );
  AND U10727 ( .A(n831), .B(n11101), .Z(n11106) );
  XNOR U10728 ( .A(n11105), .B(n11099), .Z(n11101) );
  XOR U10729 ( .A(n11107), .B(n11108), .Z(n11099) );
  AND U10730 ( .A(n846), .B(n11109), .Z(n11108) );
  XNOR U10731 ( .A(n11110), .B(n11111), .Z(n11105) );
  AND U10732 ( .A(n838), .B(n11112), .Z(n11111) );
  XOR U10733 ( .A(p_input[1182]), .B(n11110), .Z(n11112) );
  XNOR U10734 ( .A(n11113), .B(n11114), .Z(n11110) );
  AND U10735 ( .A(n842), .B(n11109), .Z(n11114) );
  XNOR U10736 ( .A(n11113), .B(n11107), .Z(n11109) );
  XOR U10737 ( .A(n11115), .B(n11116), .Z(n11107) );
  AND U10738 ( .A(n857), .B(n11117), .Z(n11116) );
  XNOR U10739 ( .A(n11118), .B(n11119), .Z(n11113) );
  AND U10740 ( .A(n849), .B(n11120), .Z(n11119) );
  XOR U10741 ( .A(p_input[1198]), .B(n11118), .Z(n11120) );
  XNOR U10742 ( .A(n11121), .B(n11122), .Z(n11118) );
  AND U10743 ( .A(n853), .B(n11117), .Z(n11122) );
  XNOR U10744 ( .A(n11121), .B(n11115), .Z(n11117) );
  XOR U10745 ( .A(n11123), .B(n11124), .Z(n11115) );
  AND U10746 ( .A(n868), .B(n11125), .Z(n11124) );
  XNOR U10747 ( .A(n11126), .B(n11127), .Z(n11121) );
  AND U10748 ( .A(n860), .B(n11128), .Z(n11127) );
  XOR U10749 ( .A(p_input[1214]), .B(n11126), .Z(n11128) );
  XNOR U10750 ( .A(n11129), .B(n11130), .Z(n11126) );
  AND U10751 ( .A(n864), .B(n11125), .Z(n11130) );
  XNOR U10752 ( .A(n11129), .B(n11123), .Z(n11125) );
  XOR U10753 ( .A(n11131), .B(n11132), .Z(n11123) );
  AND U10754 ( .A(n879), .B(n11133), .Z(n11132) );
  XNOR U10755 ( .A(n11134), .B(n11135), .Z(n11129) );
  AND U10756 ( .A(n871), .B(n11136), .Z(n11135) );
  XOR U10757 ( .A(p_input[1230]), .B(n11134), .Z(n11136) );
  XNOR U10758 ( .A(n11137), .B(n11138), .Z(n11134) );
  AND U10759 ( .A(n875), .B(n11133), .Z(n11138) );
  XNOR U10760 ( .A(n11137), .B(n11131), .Z(n11133) );
  XOR U10761 ( .A(n11139), .B(n11140), .Z(n11131) );
  AND U10762 ( .A(n890), .B(n11141), .Z(n11140) );
  XNOR U10763 ( .A(n11142), .B(n11143), .Z(n11137) );
  AND U10764 ( .A(n882), .B(n11144), .Z(n11143) );
  XOR U10765 ( .A(p_input[1246]), .B(n11142), .Z(n11144) );
  XNOR U10766 ( .A(n11145), .B(n11146), .Z(n11142) );
  AND U10767 ( .A(n886), .B(n11141), .Z(n11146) );
  XNOR U10768 ( .A(n11145), .B(n11139), .Z(n11141) );
  XOR U10769 ( .A(n11147), .B(n11148), .Z(n11139) );
  AND U10770 ( .A(n901), .B(n11149), .Z(n11148) );
  XNOR U10771 ( .A(n11150), .B(n11151), .Z(n11145) );
  AND U10772 ( .A(n893), .B(n11152), .Z(n11151) );
  XOR U10773 ( .A(p_input[1262]), .B(n11150), .Z(n11152) );
  XNOR U10774 ( .A(n11153), .B(n11154), .Z(n11150) );
  AND U10775 ( .A(n897), .B(n11149), .Z(n11154) );
  XNOR U10776 ( .A(n11153), .B(n11147), .Z(n11149) );
  XOR U10777 ( .A(n11155), .B(n11156), .Z(n11147) );
  AND U10778 ( .A(n912), .B(n11157), .Z(n11156) );
  XNOR U10779 ( .A(n11158), .B(n11159), .Z(n11153) );
  AND U10780 ( .A(n904), .B(n11160), .Z(n11159) );
  XOR U10781 ( .A(p_input[1278]), .B(n11158), .Z(n11160) );
  XNOR U10782 ( .A(n11161), .B(n11162), .Z(n11158) );
  AND U10783 ( .A(n908), .B(n11157), .Z(n11162) );
  XNOR U10784 ( .A(n11161), .B(n11155), .Z(n11157) );
  XOR U10785 ( .A(n11163), .B(n11164), .Z(n11155) );
  AND U10786 ( .A(n923), .B(n11165), .Z(n11164) );
  XNOR U10787 ( .A(n11166), .B(n11167), .Z(n11161) );
  AND U10788 ( .A(n915), .B(n11168), .Z(n11167) );
  XOR U10789 ( .A(p_input[1294]), .B(n11166), .Z(n11168) );
  XNOR U10790 ( .A(n11169), .B(n11170), .Z(n11166) );
  AND U10791 ( .A(n919), .B(n11165), .Z(n11170) );
  XNOR U10792 ( .A(n11169), .B(n11163), .Z(n11165) );
  XOR U10793 ( .A(n11171), .B(n11172), .Z(n11163) );
  AND U10794 ( .A(n934), .B(n11173), .Z(n11172) );
  XNOR U10795 ( .A(n11174), .B(n11175), .Z(n11169) );
  AND U10796 ( .A(n926), .B(n11176), .Z(n11175) );
  XOR U10797 ( .A(p_input[1310]), .B(n11174), .Z(n11176) );
  XNOR U10798 ( .A(n11177), .B(n11178), .Z(n11174) );
  AND U10799 ( .A(n930), .B(n11173), .Z(n11178) );
  XNOR U10800 ( .A(n11177), .B(n11171), .Z(n11173) );
  XOR U10801 ( .A(n11179), .B(n11180), .Z(n11171) );
  AND U10802 ( .A(n945), .B(n11181), .Z(n11180) );
  XNOR U10803 ( .A(n11182), .B(n11183), .Z(n11177) );
  AND U10804 ( .A(n937), .B(n11184), .Z(n11183) );
  XOR U10805 ( .A(p_input[1326]), .B(n11182), .Z(n11184) );
  XNOR U10806 ( .A(n11185), .B(n11186), .Z(n11182) );
  AND U10807 ( .A(n941), .B(n11181), .Z(n11186) );
  XNOR U10808 ( .A(n11185), .B(n11179), .Z(n11181) );
  XOR U10809 ( .A(n11187), .B(n11188), .Z(n11179) );
  AND U10810 ( .A(n956), .B(n11189), .Z(n11188) );
  XNOR U10811 ( .A(n11190), .B(n11191), .Z(n11185) );
  AND U10812 ( .A(n948), .B(n11192), .Z(n11191) );
  XOR U10813 ( .A(p_input[1342]), .B(n11190), .Z(n11192) );
  XNOR U10814 ( .A(n11193), .B(n11194), .Z(n11190) );
  AND U10815 ( .A(n952), .B(n11189), .Z(n11194) );
  XNOR U10816 ( .A(n11193), .B(n11187), .Z(n11189) );
  XOR U10817 ( .A(n11195), .B(n11196), .Z(n11187) );
  AND U10818 ( .A(n967), .B(n11197), .Z(n11196) );
  XNOR U10819 ( .A(n11198), .B(n11199), .Z(n11193) );
  AND U10820 ( .A(n959), .B(n11200), .Z(n11199) );
  XOR U10821 ( .A(p_input[1358]), .B(n11198), .Z(n11200) );
  XNOR U10822 ( .A(n11201), .B(n11202), .Z(n11198) );
  AND U10823 ( .A(n963), .B(n11197), .Z(n11202) );
  XNOR U10824 ( .A(n11201), .B(n11195), .Z(n11197) );
  XOR U10825 ( .A(n11203), .B(n11204), .Z(n11195) );
  AND U10826 ( .A(n978), .B(n11205), .Z(n11204) );
  XNOR U10827 ( .A(n11206), .B(n11207), .Z(n11201) );
  AND U10828 ( .A(n970), .B(n11208), .Z(n11207) );
  XOR U10829 ( .A(p_input[1374]), .B(n11206), .Z(n11208) );
  XNOR U10830 ( .A(n11209), .B(n11210), .Z(n11206) );
  AND U10831 ( .A(n974), .B(n11205), .Z(n11210) );
  XNOR U10832 ( .A(n11209), .B(n11203), .Z(n11205) );
  XOR U10833 ( .A(n11211), .B(n11212), .Z(n11203) );
  AND U10834 ( .A(n989), .B(n11213), .Z(n11212) );
  XNOR U10835 ( .A(n11214), .B(n11215), .Z(n11209) );
  AND U10836 ( .A(n981), .B(n11216), .Z(n11215) );
  XOR U10837 ( .A(p_input[1390]), .B(n11214), .Z(n11216) );
  XNOR U10838 ( .A(n11217), .B(n11218), .Z(n11214) );
  AND U10839 ( .A(n985), .B(n11213), .Z(n11218) );
  XNOR U10840 ( .A(n11217), .B(n11211), .Z(n11213) );
  XOR U10841 ( .A(n11219), .B(n11220), .Z(n11211) );
  AND U10842 ( .A(n1000), .B(n11221), .Z(n11220) );
  XNOR U10843 ( .A(n11222), .B(n11223), .Z(n11217) );
  AND U10844 ( .A(n992), .B(n11224), .Z(n11223) );
  XOR U10845 ( .A(p_input[1406]), .B(n11222), .Z(n11224) );
  XNOR U10846 ( .A(n11225), .B(n11226), .Z(n11222) );
  AND U10847 ( .A(n996), .B(n11221), .Z(n11226) );
  XNOR U10848 ( .A(n11225), .B(n11219), .Z(n11221) );
  XOR U10849 ( .A(n11227), .B(n11228), .Z(n11219) );
  AND U10850 ( .A(n1011), .B(n11229), .Z(n11228) );
  XNOR U10851 ( .A(n11230), .B(n11231), .Z(n11225) );
  AND U10852 ( .A(n1003), .B(n11232), .Z(n11231) );
  XOR U10853 ( .A(p_input[1422]), .B(n11230), .Z(n11232) );
  XNOR U10854 ( .A(n11233), .B(n11234), .Z(n11230) );
  AND U10855 ( .A(n1007), .B(n11229), .Z(n11234) );
  XNOR U10856 ( .A(n11233), .B(n11227), .Z(n11229) );
  XOR U10857 ( .A(n11235), .B(n11236), .Z(n11227) );
  AND U10858 ( .A(n1022), .B(n11237), .Z(n11236) );
  XNOR U10859 ( .A(n11238), .B(n11239), .Z(n11233) );
  AND U10860 ( .A(n1014), .B(n11240), .Z(n11239) );
  XOR U10861 ( .A(p_input[1438]), .B(n11238), .Z(n11240) );
  XNOR U10862 ( .A(n11241), .B(n11242), .Z(n11238) );
  AND U10863 ( .A(n1018), .B(n11237), .Z(n11242) );
  XNOR U10864 ( .A(n11241), .B(n11235), .Z(n11237) );
  XOR U10865 ( .A(n11243), .B(n11244), .Z(n11235) );
  AND U10866 ( .A(n1033), .B(n11245), .Z(n11244) );
  XNOR U10867 ( .A(n11246), .B(n11247), .Z(n11241) );
  AND U10868 ( .A(n1025), .B(n11248), .Z(n11247) );
  XOR U10869 ( .A(p_input[1454]), .B(n11246), .Z(n11248) );
  XNOR U10870 ( .A(n11249), .B(n11250), .Z(n11246) );
  AND U10871 ( .A(n1029), .B(n11245), .Z(n11250) );
  XNOR U10872 ( .A(n11249), .B(n11243), .Z(n11245) );
  XOR U10873 ( .A(n11251), .B(n11252), .Z(n11243) );
  AND U10874 ( .A(n1044), .B(n11253), .Z(n11252) );
  XNOR U10875 ( .A(n11254), .B(n11255), .Z(n11249) );
  AND U10876 ( .A(n1036), .B(n11256), .Z(n11255) );
  XOR U10877 ( .A(p_input[1470]), .B(n11254), .Z(n11256) );
  XNOR U10878 ( .A(n11257), .B(n11258), .Z(n11254) );
  AND U10879 ( .A(n1040), .B(n11253), .Z(n11258) );
  XNOR U10880 ( .A(n11257), .B(n11251), .Z(n11253) );
  XOR U10881 ( .A(n11259), .B(n11260), .Z(n11251) );
  AND U10882 ( .A(n1055), .B(n11261), .Z(n11260) );
  XNOR U10883 ( .A(n11262), .B(n11263), .Z(n11257) );
  AND U10884 ( .A(n1047), .B(n11264), .Z(n11263) );
  XOR U10885 ( .A(p_input[1486]), .B(n11262), .Z(n11264) );
  XNOR U10886 ( .A(n11265), .B(n11266), .Z(n11262) );
  AND U10887 ( .A(n1051), .B(n11261), .Z(n11266) );
  XNOR U10888 ( .A(n11265), .B(n11259), .Z(n11261) );
  XOR U10889 ( .A(n11267), .B(n11268), .Z(n11259) );
  AND U10890 ( .A(n1066), .B(n11269), .Z(n11268) );
  XNOR U10891 ( .A(n11270), .B(n11271), .Z(n11265) );
  AND U10892 ( .A(n1058), .B(n11272), .Z(n11271) );
  XOR U10893 ( .A(p_input[1502]), .B(n11270), .Z(n11272) );
  XNOR U10894 ( .A(n11273), .B(n11274), .Z(n11270) );
  AND U10895 ( .A(n1062), .B(n11269), .Z(n11274) );
  XNOR U10896 ( .A(n11273), .B(n11267), .Z(n11269) );
  XOR U10897 ( .A(n11275), .B(n11276), .Z(n11267) );
  AND U10898 ( .A(n1077), .B(n11277), .Z(n11276) );
  XNOR U10899 ( .A(n11278), .B(n11279), .Z(n11273) );
  AND U10900 ( .A(n1069), .B(n11280), .Z(n11279) );
  XOR U10901 ( .A(p_input[1518]), .B(n11278), .Z(n11280) );
  XNOR U10902 ( .A(n11281), .B(n11282), .Z(n11278) );
  AND U10903 ( .A(n1073), .B(n11277), .Z(n11282) );
  XNOR U10904 ( .A(n11281), .B(n11275), .Z(n11277) );
  XOR U10905 ( .A(n11283), .B(n11284), .Z(n11275) );
  AND U10906 ( .A(n1088), .B(n11285), .Z(n11284) );
  XNOR U10907 ( .A(n11286), .B(n11287), .Z(n11281) );
  AND U10908 ( .A(n1080), .B(n11288), .Z(n11287) );
  XOR U10909 ( .A(p_input[1534]), .B(n11286), .Z(n11288) );
  XNOR U10910 ( .A(n11289), .B(n11290), .Z(n11286) );
  AND U10911 ( .A(n1084), .B(n11285), .Z(n11290) );
  XNOR U10912 ( .A(n11289), .B(n11283), .Z(n11285) );
  XOR U10913 ( .A(n11291), .B(n11292), .Z(n11283) );
  AND U10914 ( .A(n1099), .B(n11293), .Z(n11292) );
  XNOR U10915 ( .A(n11294), .B(n11295), .Z(n11289) );
  AND U10916 ( .A(n1091), .B(n11296), .Z(n11295) );
  XOR U10917 ( .A(p_input[1550]), .B(n11294), .Z(n11296) );
  XNOR U10918 ( .A(n11297), .B(n11298), .Z(n11294) );
  AND U10919 ( .A(n1095), .B(n11293), .Z(n11298) );
  XNOR U10920 ( .A(n11297), .B(n11291), .Z(n11293) );
  XOR U10921 ( .A(n11299), .B(n11300), .Z(n11291) );
  AND U10922 ( .A(n1110), .B(n11301), .Z(n11300) );
  XNOR U10923 ( .A(n11302), .B(n11303), .Z(n11297) );
  AND U10924 ( .A(n1102), .B(n11304), .Z(n11303) );
  XOR U10925 ( .A(p_input[1566]), .B(n11302), .Z(n11304) );
  XNOR U10926 ( .A(n11305), .B(n11306), .Z(n11302) );
  AND U10927 ( .A(n1106), .B(n11301), .Z(n11306) );
  XNOR U10928 ( .A(n11305), .B(n11299), .Z(n11301) );
  XOR U10929 ( .A(n11307), .B(n11308), .Z(n11299) );
  AND U10930 ( .A(n1121), .B(n11309), .Z(n11308) );
  XNOR U10931 ( .A(n11310), .B(n11311), .Z(n11305) );
  AND U10932 ( .A(n1113), .B(n11312), .Z(n11311) );
  XOR U10933 ( .A(p_input[1582]), .B(n11310), .Z(n11312) );
  XNOR U10934 ( .A(n11313), .B(n11314), .Z(n11310) );
  AND U10935 ( .A(n1117), .B(n11309), .Z(n11314) );
  XNOR U10936 ( .A(n11313), .B(n11307), .Z(n11309) );
  XOR U10937 ( .A(n11315), .B(n11316), .Z(n11307) );
  AND U10938 ( .A(n1132), .B(n11317), .Z(n11316) );
  XNOR U10939 ( .A(n11318), .B(n11319), .Z(n11313) );
  AND U10940 ( .A(n1124), .B(n11320), .Z(n11319) );
  XOR U10941 ( .A(p_input[1598]), .B(n11318), .Z(n11320) );
  XNOR U10942 ( .A(n11321), .B(n11322), .Z(n11318) );
  AND U10943 ( .A(n1128), .B(n11317), .Z(n11322) );
  XNOR U10944 ( .A(n11321), .B(n11315), .Z(n11317) );
  XOR U10945 ( .A(n11323), .B(n11324), .Z(n11315) );
  AND U10946 ( .A(n1143), .B(n11325), .Z(n11324) );
  XNOR U10947 ( .A(n11326), .B(n11327), .Z(n11321) );
  AND U10948 ( .A(n1135), .B(n11328), .Z(n11327) );
  XOR U10949 ( .A(p_input[1614]), .B(n11326), .Z(n11328) );
  XNOR U10950 ( .A(n11329), .B(n11330), .Z(n11326) );
  AND U10951 ( .A(n1139), .B(n11325), .Z(n11330) );
  XNOR U10952 ( .A(n11329), .B(n11323), .Z(n11325) );
  XOR U10953 ( .A(n11331), .B(n11332), .Z(n11323) );
  AND U10954 ( .A(n1154), .B(n11333), .Z(n11332) );
  XNOR U10955 ( .A(n11334), .B(n11335), .Z(n11329) );
  AND U10956 ( .A(n1146), .B(n11336), .Z(n11335) );
  XOR U10957 ( .A(p_input[1630]), .B(n11334), .Z(n11336) );
  XNOR U10958 ( .A(n11337), .B(n11338), .Z(n11334) );
  AND U10959 ( .A(n1150), .B(n11333), .Z(n11338) );
  XNOR U10960 ( .A(n11337), .B(n11331), .Z(n11333) );
  XOR U10961 ( .A(n11339), .B(n11340), .Z(n11331) );
  AND U10962 ( .A(n1165), .B(n11341), .Z(n11340) );
  XNOR U10963 ( .A(n11342), .B(n11343), .Z(n11337) );
  AND U10964 ( .A(n1157), .B(n11344), .Z(n11343) );
  XOR U10965 ( .A(p_input[1646]), .B(n11342), .Z(n11344) );
  XNOR U10966 ( .A(n11345), .B(n11346), .Z(n11342) );
  AND U10967 ( .A(n1161), .B(n11341), .Z(n11346) );
  XNOR U10968 ( .A(n11345), .B(n11339), .Z(n11341) );
  XOR U10969 ( .A(n11347), .B(n11348), .Z(n11339) );
  AND U10970 ( .A(n1176), .B(n11349), .Z(n11348) );
  XNOR U10971 ( .A(n11350), .B(n11351), .Z(n11345) );
  AND U10972 ( .A(n1168), .B(n11352), .Z(n11351) );
  XOR U10973 ( .A(p_input[1662]), .B(n11350), .Z(n11352) );
  XNOR U10974 ( .A(n11353), .B(n11354), .Z(n11350) );
  AND U10975 ( .A(n1172), .B(n11349), .Z(n11354) );
  XNOR U10976 ( .A(n11353), .B(n11347), .Z(n11349) );
  XOR U10977 ( .A(n11355), .B(n11356), .Z(n11347) );
  AND U10978 ( .A(n1187), .B(n11357), .Z(n11356) );
  XNOR U10979 ( .A(n11358), .B(n11359), .Z(n11353) );
  AND U10980 ( .A(n1179), .B(n11360), .Z(n11359) );
  XOR U10981 ( .A(p_input[1678]), .B(n11358), .Z(n11360) );
  XNOR U10982 ( .A(n11361), .B(n11362), .Z(n11358) );
  AND U10983 ( .A(n1183), .B(n11357), .Z(n11362) );
  XNOR U10984 ( .A(n11361), .B(n11355), .Z(n11357) );
  XOR U10985 ( .A(n11363), .B(n11364), .Z(n11355) );
  AND U10986 ( .A(n1198), .B(n11365), .Z(n11364) );
  XNOR U10987 ( .A(n11366), .B(n11367), .Z(n11361) );
  AND U10988 ( .A(n1190), .B(n11368), .Z(n11367) );
  XOR U10989 ( .A(p_input[1694]), .B(n11366), .Z(n11368) );
  XNOR U10990 ( .A(n11369), .B(n11370), .Z(n11366) );
  AND U10991 ( .A(n1194), .B(n11365), .Z(n11370) );
  XNOR U10992 ( .A(n11369), .B(n11363), .Z(n11365) );
  XOR U10993 ( .A(n11371), .B(n11372), .Z(n11363) );
  AND U10994 ( .A(n1209), .B(n11373), .Z(n11372) );
  XNOR U10995 ( .A(n11374), .B(n11375), .Z(n11369) );
  AND U10996 ( .A(n1201), .B(n11376), .Z(n11375) );
  XOR U10997 ( .A(p_input[1710]), .B(n11374), .Z(n11376) );
  XNOR U10998 ( .A(n11377), .B(n11378), .Z(n11374) );
  AND U10999 ( .A(n1205), .B(n11373), .Z(n11378) );
  XNOR U11000 ( .A(n11377), .B(n11371), .Z(n11373) );
  XOR U11001 ( .A(n11379), .B(n11380), .Z(n11371) );
  AND U11002 ( .A(n1220), .B(n11381), .Z(n11380) );
  XNOR U11003 ( .A(n11382), .B(n11383), .Z(n11377) );
  AND U11004 ( .A(n1212), .B(n11384), .Z(n11383) );
  XOR U11005 ( .A(p_input[1726]), .B(n11382), .Z(n11384) );
  XNOR U11006 ( .A(n11385), .B(n11386), .Z(n11382) );
  AND U11007 ( .A(n1216), .B(n11381), .Z(n11386) );
  XNOR U11008 ( .A(n11385), .B(n11379), .Z(n11381) );
  XOR U11009 ( .A(n11387), .B(n11388), .Z(n11379) );
  AND U11010 ( .A(n1231), .B(n11389), .Z(n11388) );
  XNOR U11011 ( .A(n11390), .B(n11391), .Z(n11385) );
  AND U11012 ( .A(n1223), .B(n11392), .Z(n11391) );
  XOR U11013 ( .A(p_input[1742]), .B(n11390), .Z(n11392) );
  XNOR U11014 ( .A(n11393), .B(n11394), .Z(n11390) );
  AND U11015 ( .A(n1227), .B(n11389), .Z(n11394) );
  XNOR U11016 ( .A(n11393), .B(n11387), .Z(n11389) );
  XOR U11017 ( .A(n11395), .B(n11396), .Z(n11387) );
  AND U11018 ( .A(n1242), .B(n11397), .Z(n11396) );
  XNOR U11019 ( .A(n11398), .B(n11399), .Z(n11393) );
  AND U11020 ( .A(n1234), .B(n11400), .Z(n11399) );
  XOR U11021 ( .A(p_input[1758]), .B(n11398), .Z(n11400) );
  XNOR U11022 ( .A(n11401), .B(n11402), .Z(n11398) );
  AND U11023 ( .A(n1238), .B(n11397), .Z(n11402) );
  XNOR U11024 ( .A(n11401), .B(n11395), .Z(n11397) );
  XOR U11025 ( .A(n11403), .B(n11404), .Z(n11395) );
  AND U11026 ( .A(n1253), .B(n11405), .Z(n11404) );
  XNOR U11027 ( .A(n11406), .B(n11407), .Z(n11401) );
  AND U11028 ( .A(n1245), .B(n11408), .Z(n11407) );
  XOR U11029 ( .A(p_input[1774]), .B(n11406), .Z(n11408) );
  XNOR U11030 ( .A(n11409), .B(n11410), .Z(n11406) );
  AND U11031 ( .A(n1249), .B(n11405), .Z(n11410) );
  XNOR U11032 ( .A(n11409), .B(n11403), .Z(n11405) );
  XOR U11033 ( .A(n11411), .B(n11412), .Z(n11403) );
  AND U11034 ( .A(n1264), .B(n11413), .Z(n11412) );
  XNOR U11035 ( .A(n11414), .B(n11415), .Z(n11409) );
  AND U11036 ( .A(n1256), .B(n11416), .Z(n11415) );
  XOR U11037 ( .A(p_input[1790]), .B(n11414), .Z(n11416) );
  XNOR U11038 ( .A(n11417), .B(n11418), .Z(n11414) );
  AND U11039 ( .A(n1260), .B(n11413), .Z(n11418) );
  XNOR U11040 ( .A(n11417), .B(n11411), .Z(n11413) );
  XOR U11041 ( .A(n11419), .B(n11420), .Z(n11411) );
  AND U11042 ( .A(n1275), .B(n11421), .Z(n11420) );
  XNOR U11043 ( .A(n11422), .B(n11423), .Z(n11417) );
  AND U11044 ( .A(n1267), .B(n11424), .Z(n11423) );
  XOR U11045 ( .A(p_input[1806]), .B(n11422), .Z(n11424) );
  XNOR U11046 ( .A(n11425), .B(n11426), .Z(n11422) );
  AND U11047 ( .A(n1271), .B(n11421), .Z(n11426) );
  XNOR U11048 ( .A(n11425), .B(n11419), .Z(n11421) );
  XOR U11049 ( .A(n11427), .B(n11428), .Z(n11419) );
  AND U11050 ( .A(n1286), .B(n11429), .Z(n11428) );
  XNOR U11051 ( .A(n11430), .B(n11431), .Z(n11425) );
  AND U11052 ( .A(n1278), .B(n11432), .Z(n11431) );
  XOR U11053 ( .A(p_input[1822]), .B(n11430), .Z(n11432) );
  XNOR U11054 ( .A(n11433), .B(n11434), .Z(n11430) );
  AND U11055 ( .A(n1282), .B(n11429), .Z(n11434) );
  XNOR U11056 ( .A(n11433), .B(n11427), .Z(n11429) );
  XOR U11057 ( .A(n11435), .B(n11436), .Z(n11427) );
  AND U11058 ( .A(n1297), .B(n11437), .Z(n11436) );
  XNOR U11059 ( .A(n11438), .B(n11439), .Z(n11433) );
  AND U11060 ( .A(n1289), .B(n11440), .Z(n11439) );
  XOR U11061 ( .A(p_input[1838]), .B(n11438), .Z(n11440) );
  XNOR U11062 ( .A(n11441), .B(n11442), .Z(n11438) );
  AND U11063 ( .A(n1293), .B(n11437), .Z(n11442) );
  XNOR U11064 ( .A(n11441), .B(n11435), .Z(n11437) );
  XOR U11065 ( .A(n11443), .B(n11444), .Z(n11435) );
  AND U11066 ( .A(n1308), .B(n11445), .Z(n11444) );
  XNOR U11067 ( .A(n11446), .B(n11447), .Z(n11441) );
  AND U11068 ( .A(n1300), .B(n11448), .Z(n11447) );
  XOR U11069 ( .A(p_input[1854]), .B(n11446), .Z(n11448) );
  XNOR U11070 ( .A(n11449), .B(n11450), .Z(n11446) );
  AND U11071 ( .A(n1304), .B(n11445), .Z(n11450) );
  XNOR U11072 ( .A(n11449), .B(n11443), .Z(n11445) );
  XOR U11073 ( .A(n11451), .B(n11452), .Z(n11443) );
  AND U11074 ( .A(n1319), .B(n11453), .Z(n11452) );
  XNOR U11075 ( .A(n11454), .B(n11455), .Z(n11449) );
  AND U11076 ( .A(n1311), .B(n11456), .Z(n11455) );
  XOR U11077 ( .A(p_input[1870]), .B(n11454), .Z(n11456) );
  XNOR U11078 ( .A(n11457), .B(n11458), .Z(n11454) );
  AND U11079 ( .A(n1315), .B(n11453), .Z(n11458) );
  XNOR U11080 ( .A(n11457), .B(n11451), .Z(n11453) );
  XOR U11081 ( .A(n11459), .B(n11460), .Z(n11451) );
  AND U11082 ( .A(n1330), .B(n11461), .Z(n11460) );
  XNOR U11083 ( .A(n11462), .B(n11463), .Z(n11457) );
  AND U11084 ( .A(n1322), .B(n11464), .Z(n11463) );
  XOR U11085 ( .A(p_input[1886]), .B(n11462), .Z(n11464) );
  XNOR U11086 ( .A(n11465), .B(n11466), .Z(n11462) );
  AND U11087 ( .A(n1326), .B(n11461), .Z(n11466) );
  XNOR U11088 ( .A(n11465), .B(n11459), .Z(n11461) );
  XOR U11089 ( .A(n11467), .B(n11468), .Z(n11459) );
  AND U11090 ( .A(n1341), .B(n11469), .Z(n11468) );
  XNOR U11091 ( .A(n11470), .B(n11471), .Z(n11465) );
  AND U11092 ( .A(n1333), .B(n11472), .Z(n11471) );
  XOR U11093 ( .A(p_input[1902]), .B(n11470), .Z(n11472) );
  XNOR U11094 ( .A(n11473), .B(n11474), .Z(n11470) );
  AND U11095 ( .A(n1337), .B(n11469), .Z(n11474) );
  XNOR U11096 ( .A(n11473), .B(n11467), .Z(n11469) );
  XOR U11097 ( .A(n11475), .B(n11476), .Z(n11467) );
  AND U11098 ( .A(n1352), .B(n11477), .Z(n11476) );
  XNOR U11099 ( .A(n11478), .B(n11479), .Z(n11473) );
  AND U11100 ( .A(n1344), .B(n11480), .Z(n11479) );
  XOR U11101 ( .A(p_input[1918]), .B(n11478), .Z(n11480) );
  XNOR U11102 ( .A(n11481), .B(n11482), .Z(n11478) );
  AND U11103 ( .A(n1348), .B(n11477), .Z(n11482) );
  XNOR U11104 ( .A(n11481), .B(n11475), .Z(n11477) );
  XOR U11105 ( .A(n11483), .B(n11484), .Z(n11475) );
  AND U11106 ( .A(n1363), .B(n11485), .Z(n11484) );
  XNOR U11107 ( .A(n11486), .B(n11487), .Z(n11481) );
  AND U11108 ( .A(n1355), .B(n11488), .Z(n11487) );
  XOR U11109 ( .A(p_input[1934]), .B(n11486), .Z(n11488) );
  XNOR U11110 ( .A(n11489), .B(n11490), .Z(n11486) );
  AND U11111 ( .A(n1359), .B(n11485), .Z(n11490) );
  XNOR U11112 ( .A(n11489), .B(n11483), .Z(n11485) );
  XOR U11113 ( .A(n11491), .B(n11492), .Z(n11483) );
  AND U11114 ( .A(n1374), .B(n11493), .Z(n11492) );
  XNOR U11115 ( .A(n11494), .B(n11495), .Z(n11489) );
  AND U11116 ( .A(n1366), .B(n11496), .Z(n11495) );
  XOR U11117 ( .A(p_input[1950]), .B(n11494), .Z(n11496) );
  XNOR U11118 ( .A(n11497), .B(n11498), .Z(n11494) );
  AND U11119 ( .A(n1370), .B(n11493), .Z(n11498) );
  XNOR U11120 ( .A(n11497), .B(n11491), .Z(n11493) );
  XOR U11121 ( .A(n11499), .B(n11500), .Z(n11491) );
  AND U11122 ( .A(n1385), .B(n11501), .Z(n11500) );
  XNOR U11123 ( .A(n11502), .B(n11503), .Z(n11497) );
  AND U11124 ( .A(n1377), .B(n11504), .Z(n11503) );
  XOR U11125 ( .A(p_input[1966]), .B(n11502), .Z(n11504) );
  XNOR U11126 ( .A(n11505), .B(n11506), .Z(n11502) );
  AND U11127 ( .A(n1381), .B(n11501), .Z(n11506) );
  XNOR U11128 ( .A(n11505), .B(n11499), .Z(n11501) );
  XOR U11129 ( .A(n11507), .B(n11508), .Z(n11499) );
  AND U11130 ( .A(n1396), .B(n11509), .Z(n11508) );
  XNOR U11131 ( .A(n11510), .B(n11511), .Z(n11505) );
  AND U11132 ( .A(n1388), .B(n11512), .Z(n11511) );
  XOR U11133 ( .A(p_input[1982]), .B(n11510), .Z(n11512) );
  XNOR U11134 ( .A(n11513), .B(n11514), .Z(n11510) );
  AND U11135 ( .A(n1392), .B(n11509), .Z(n11514) );
  XNOR U11136 ( .A(n11513), .B(n11507), .Z(n11509) );
  XOR U11137 ( .A(n11515), .B(n11516), .Z(n11507) );
  AND U11138 ( .A(n1407), .B(n11517), .Z(n11516) );
  XNOR U11139 ( .A(n11518), .B(n11519), .Z(n11513) );
  AND U11140 ( .A(n1399), .B(n11520), .Z(n11519) );
  XOR U11141 ( .A(p_input[1998]), .B(n11518), .Z(n11520) );
  XNOR U11142 ( .A(n11521), .B(n11522), .Z(n11518) );
  AND U11143 ( .A(n1403), .B(n11517), .Z(n11522) );
  XNOR U11144 ( .A(n11521), .B(n11515), .Z(n11517) );
  XOR U11145 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n11523), .Z(n11515) );
  AND U11146 ( .A(n1417), .B(n11524), .Z(n11523) );
  XNOR U11147 ( .A(n11525), .B(n11526), .Z(n11521) );
  AND U11148 ( .A(n1410), .B(n11527), .Z(n11526) );
  XOR U11149 ( .A(p_input[2014]), .B(n11525), .Z(n11527) );
  XNOR U11150 ( .A(n11528), .B(n11529), .Z(n11525) );
  AND U11151 ( .A(n1414), .B(n11524), .Z(n11529) );
  XOR U11152 ( .A(n11530), .B(n11528), .Z(n11524) );
  IV U11153 ( .A(\knn_comb_/min_val_out[0][14] ), .Z(n11530) );
  IV U11154 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n11528)
         );
  XOR U11155 ( .A(n21), .B(n11531), .Z(o[13]) );
  AND U11156 ( .A(n30), .B(n11532), .Z(n21) );
  XOR U11157 ( .A(n22), .B(n11531), .Z(n11532) );
  XOR U11158 ( .A(n11533), .B(n11534), .Z(n11531) );
  AND U11159 ( .A(n42), .B(n11535), .Z(n11534) );
  XOR U11160 ( .A(n11536), .B(n11537), .Z(n22) );
  AND U11161 ( .A(n34), .B(n11538), .Z(n11537) );
  XOR U11162 ( .A(p_input[13]), .B(n11536), .Z(n11538) );
  XNOR U11163 ( .A(n11539), .B(n11540), .Z(n11536) );
  AND U11164 ( .A(n38), .B(n11535), .Z(n11540) );
  XNOR U11165 ( .A(n11539), .B(n11533), .Z(n11535) );
  XOR U11166 ( .A(n11541), .B(n11542), .Z(n11533) );
  AND U11167 ( .A(n54), .B(n11543), .Z(n11542) );
  XNOR U11168 ( .A(n11544), .B(n11545), .Z(n11539) );
  AND U11169 ( .A(n46), .B(n11546), .Z(n11545) );
  XOR U11170 ( .A(p_input[29]), .B(n11544), .Z(n11546) );
  XNOR U11171 ( .A(n11547), .B(n11548), .Z(n11544) );
  AND U11172 ( .A(n50), .B(n11543), .Z(n11548) );
  XNOR U11173 ( .A(n11547), .B(n11541), .Z(n11543) );
  XOR U11174 ( .A(n11549), .B(n11550), .Z(n11541) );
  AND U11175 ( .A(n65), .B(n11551), .Z(n11550) );
  XNOR U11176 ( .A(n11552), .B(n11553), .Z(n11547) );
  AND U11177 ( .A(n57), .B(n11554), .Z(n11553) );
  XOR U11178 ( .A(p_input[45]), .B(n11552), .Z(n11554) );
  XNOR U11179 ( .A(n11555), .B(n11556), .Z(n11552) );
  AND U11180 ( .A(n61), .B(n11551), .Z(n11556) );
  XNOR U11181 ( .A(n11555), .B(n11549), .Z(n11551) );
  XOR U11182 ( .A(n11557), .B(n11558), .Z(n11549) );
  AND U11183 ( .A(n76), .B(n11559), .Z(n11558) );
  XNOR U11184 ( .A(n11560), .B(n11561), .Z(n11555) );
  AND U11185 ( .A(n68), .B(n11562), .Z(n11561) );
  XOR U11186 ( .A(p_input[61]), .B(n11560), .Z(n11562) );
  XNOR U11187 ( .A(n11563), .B(n11564), .Z(n11560) );
  AND U11188 ( .A(n72), .B(n11559), .Z(n11564) );
  XNOR U11189 ( .A(n11563), .B(n11557), .Z(n11559) );
  XOR U11190 ( .A(n11565), .B(n11566), .Z(n11557) );
  AND U11191 ( .A(n87), .B(n11567), .Z(n11566) );
  XNOR U11192 ( .A(n11568), .B(n11569), .Z(n11563) );
  AND U11193 ( .A(n79), .B(n11570), .Z(n11569) );
  XOR U11194 ( .A(p_input[77]), .B(n11568), .Z(n11570) );
  XNOR U11195 ( .A(n11571), .B(n11572), .Z(n11568) );
  AND U11196 ( .A(n83), .B(n11567), .Z(n11572) );
  XNOR U11197 ( .A(n11571), .B(n11565), .Z(n11567) );
  XOR U11198 ( .A(n11573), .B(n11574), .Z(n11565) );
  AND U11199 ( .A(n98), .B(n11575), .Z(n11574) );
  XNOR U11200 ( .A(n11576), .B(n11577), .Z(n11571) );
  AND U11201 ( .A(n90), .B(n11578), .Z(n11577) );
  XOR U11202 ( .A(p_input[93]), .B(n11576), .Z(n11578) );
  XNOR U11203 ( .A(n11579), .B(n11580), .Z(n11576) );
  AND U11204 ( .A(n94), .B(n11575), .Z(n11580) );
  XNOR U11205 ( .A(n11579), .B(n11573), .Z(n11575) );
  XOR U11206 ( .A(n11581), .B(n11582), .Z(n11573) );
  AND U11207 ( .A(n109), .B(n11583), .Z(n11582) );
  XNOR U11208 ( .A(n11584), .B(n11585), .Z(n11579) );
  AND U11209 ( .A(n101), .B(n11586), .Z(n11585) );
  XOR U11210 ( .A(p_input[109]), .B(n11584), .Z(n11586) );
  XNOR U11211 ( .A(n11587), .B(n11588), .Z(n11584) );
  AND U11212 ( .A(n105), .B(n11583), .Z(n11588) );
  XNOR U11213 ( .A(n11587), .B(n11581), .Z(n11583) );
  XOR U11214 ( .A(n11589), .B(n11590), .Z(n11581) );
  AND U11215 ( .A(n120), .B(n11591), .Z(n11590) );
  XNOR U11216 ( .A(n11592), .B(n11593), .Z(n11587) );
  AND U11217 ( .A(n112), .B(n11594), .Z(n11593) );
  XOR U11218 ( .A(p_input[125]), .B(n11592), .Z(n11594) );
  XNOR U11219 ( .A(n11595), .B(n11596), .Z(n11592) );
  AND U11220 ( .A(n116), .B(n11591), .Z(n11596) );
  XNOR U11221 ( .A(n11595), .B(n11589), .Z(n11591) );
  XOR U11222 ( .A(n11597), .B(n11598), .Z(n11589) );
  AND U11223 ( .A(n131), .B(n11599), .Z(n11598) );
  XNOR U11224 ( .A(n11600), .B(n11601), .Z(n11595) );
  AND U11225 ( .A(n123), .B(n11602), .Z(n11601) );
  XOR U11226 ( .A(p_input[141]), .B(n11600), .Z(n11602) );
  XNOR U11227 ( .A(n11603), .B(n11604), .Z(n11600) );
  AND U11228 ( .A(n127), .B(n11599), .Z(n11604) );
  XNOR U11229 ( .A(n11603), .B(n11597), .Z(n11599) );
  XOR U11230 ( .A(n11605), .B(n11606), .Z(n11597) );
  AND U11231 ( .A(n142), .B(n11607), .Z(n11606) );
  XNOR U11232 ( .A(n11608), .B(n11609), .Z(n11603) );
  AND U11233 ( .A(n134), .B(n11610), .Z(n11609) );
  XOR U11234 ( .A(p_input[157]), .B(n11608), .Z(n11610) );
  XNOR U11235 ( .A(n11611), .B(n11612), .Z(n11608) );
  AND U11236 ( .A(n138), .B(n11607), .Z(n11612) );
  XNOR U11237 ( .A(n11611), .B(n11605), .Z(n11607) );
  XOR U11238 ( .A(n11613), .B(n11614), .Z(n11605) );
  AND U11239 ( .A(n153), .B(n11615), .Z(n11614) );
  XNOR U11240 ( .A(n11616), .B(n11617), .Z(n11611) );
  AND U11241 ( .A(n145), .B(n11618), .Z(n11617) );
  XOR U11242 ( .A(p_input[173]), .B(n11616), .Z(n11618) );
  XNOR U11243 ( .A(n11619), .B(n11620), .Z(n11616) );
  AND U11244 ( .A(n149), .B(n11615), .Z(n11620) );
  XNOR U11245 ( .A(n11619), .B(n11613), .Z(n11615) );
  XOR U11246 ( .A(n11621), .B(n11622), .Z(n11613) );
  AND U11247 ( .A(n164), .B(n11623), .Z(n11622) );
  XNOR U11248 ( .A(n11624), .B(n11625), .Z(n11619) );
  AND U11249 ( .A(n156), .B(n11626), .Z(n11625) );
  XOR U11250 ( .A(p_input[189]), .B(n11624), .Z(n11626) );
  XNOR U11251 ( .A(n11627), .B(n11628), .Z(n11624) );
  AND U11252 ( .A(n160), .B(n11623), .Z(n11628) );
  XNOR U11253 ( .A(n11627), .B(n11621), .Z(n11623) );
  XOR U11254 ( .A(n11629), .B(n11630), .Z(n11621) );
  AND U11255 ( .A(n175), .B(n11631), .Z(n11630) );
  XNOR U11256 ( .A(n11632), .B(n11633), .Z(n11627) );
  AND U11257 ( .A(n167), .B(n11634), .Z(n11633) );
  XOR U11258 ( .A(p_input[205]), .B(n11632), .Z(n11634) );
  XNOR U11259 ( .A(n11635), .B(n11636), .Z(n11632) );
  AND U11260 ( .A(n171), .B(n11631), .Z(n11636) );
  XNOR U11261 ( .A(n11635), .B(n11629), .Z(n11631) );
  XOR U11262 ( .A(n11637), .B(n11638), .Z(n11629) );
  AND U11263 ( .A(n186), .B(n11639), .Z(n11638) );
  XNOR U11264 ( .A(n11640), .B(n11641), .Z(n11635) );
  AND U11265 ( .A(n178), .B(n11642), .Z(n11641) );
  XOR U11266 ( .A(p_input[221]), .B(n11640), .Z(n11642) );
  XNOR U11267 ( .A(n11643), .B(n11644), .Z(n11640) );
  AND U11268 ( .A(n182), .B(n11639), .Z(n11644) );
  XNOR U11269 ( .A(n11643), .B(n11637), .Z(n11639) );
  XOR U11270 ( .A(n11645), .B(n11646), .Z(n11637) );
  AND U11271 ( .A(n197), .B(n11647), .Z(n11646) );
  XNOR U11272 ( .A(n11648), .B(n11649), .Z(n11643) );
  AND U11273 ( .A(n189), .B(n11650), .Z(n11649) );
  XOR U11274 ( .A(p_input[237]), .B(n11648), .Z(n11650) );
  XNOR U11275 ( .A(n11651), .B(n11652), .Z(n11648) );
  AND U11276 ( .A(n193), .B(n11647), .Z(n11652) );
  XNOR U11277 ( .A(n11651), .B(n11645), .Z(n11647) );
  XOR U11278 ( .A(n11653), .B(n11654), .Z(n11645) );
  AND U11279 ( .A(n208), .B(n11655), .Z(n11654) );
  XNOR U11280 ( .A(n11656), .B(n11657), .Z(n11651) );
  AND U11281 ( .A(n200), .B(n11658), .Z(n11657) );
  XOR U11282 ( .A(p_input[253]), .B(n11656), .Z(n11658) );
  XNOR U11283 ( .A(n11659), .B(n11660), .Z(n11656) );
  AND U11284 ( .A(n204), .B(n11655), .Z(n11660) );
  XNOR U11285 ( .A(n11659), .B(n11653), .Z(n11655) );
  XOR U11286 ( .A(n11661), .B(n11662), .Z(n11653) );
  AND U11287 ( .A(n219), .B(n11663), .Z(n11662) );
  XNOR U11288 ( .A(n11664), .B(n11665), .Z(n11659) );
  AND U11289 ( .A(n211), .B(n11666), .Z(n11665) );
  XOR U11290 ( .A(p_input[269]), .B(n11664), .Z(n11666) );
  XNOR U11291 ( .A(n11667), .B(n11668), .Z(n11664) );
  AND U11292 ( .A(n215), .B(n11663), .Z(n11668) );
  XNOR U11293 ( .A(n11667), .B(n11661), .Z(n11663) );
  XOR U11294 ( .A(n11669), .B(n11670), .Z(n11661) );
  AND U11295 ( .A(n230), .B(n11671), .Z(n11670) );
  XNOR U11296 ( .A(n11672), .B(n11673), .Z(n11667) );
  AND U11297 ( .A(n222), .B(n11674), .Z(n11673) );
  XOR U11298 ( .A(p_input[285]), .B(n11672), .Z(n11674) );
  XNOR U11299 ( .A(n11675), .B(n11676), .Z(n11672) );
  AND U11300 ( .A(n226), .B(n11671), .Z(n11676) );
  XNOR U11301 ( .A(n11675), .B(n11669), .Z(n11671) );
  XOR U11302 ( .A(n11677), .B(n11678), .Z(n11669) );
  AND U11303 ( .A(n241), .B(n11679), .Z(n11678) );
  XNOR U11304 ( .A(n11680), .B(n11681), .Z(n11675) );
  AND U11305 ( .A(n233), .B(n11682), .Z(n11681) );
  XOR U11306 ( .A(p_input[301]), .B(n11680), .Z(n11682) );
  XNOR U11307 ( .A(n11683), .B(n11684), .Z(n11680) );
  AND U11308 ( .A(n237), .B(n11679), .Z(n11684) );
  XNOR U11309 ( .A(n11683), .B(n11677), .Z(n11679) );
  XOR U11310 ( .A(n11685), .B(n11686), .Z(n11677) );
  AND U11311 ( .A(n252), .B(n11687), .Z(n11686) );
  XNOR U11312 ( .A(n11688), .B(n11689), .Z(n11683) );
  AND U11313 ( .A(n244), .B(n11690), .Z(n11689) );
  XOR U11314 ( .A(p_input[317]), .B(n11688), .Z(n11690) );
  XNOR U11315 ( .A(n11691), .B(n11692), .Z(n11688) );
  AND U11316 ( .A(n248), .B(n11687), .Z(n11692) );
  XNOR U11317 ( .A(n11691), .B(n11685), .Z(n11687) );
  XOR U11318 ( .A(n11693), .B(n11694), .Z(n11685) );
  AND U11319 ( .A(n263), .B(n11695), .Z(n11694) );
  XNOR U11320 ( .A(n11696), .B(n11697), .Z(n11691) );
  AND U11321 ( .A(n255), .B(n11698), .Z(n11697) );
  XOR U11322 ( .A(p_input[333]), .B(n11696), .Z(n11698) );
  XNOR U11323 ( .A(n11699), .B(n11700), .Z(n11696) );
  AND U11324 ( .A(n259), .B(n11695), .Z(n11700) );
  XNOR U11325 ( .A(n11699), .B(n11693), .Z(n11695) );
  XOR U11326 ( .A(n11701), .B(n11702), .Z(n11693) );
  AND U11327 ( .A(n274), .B(n11703), .Z(n11702) );
  XNOR U11328 ( .A(n11704), .B(n11705), .Z(n11699) );
  AND U11329 ( .A(n266), .B(n11706), .Z(n11705) );
  XOR U11330 ( .A(p_input[349]), .B(n11704), .Z(n11706) );
  XNOR U11331 ( .A(n11707), .B(n11708), .Z(n11704) );
  AND U11332 ( .A(n270), .B(n11703), .Z(n11708) );
  XNOR U11333 ( .A(n11707), .B(n11701), .Z(n11703) );
  XOR U11334 ( .A(n11709), .B(n11710), .Z(n11701) );
  AND U11335 ( .A(n285), .B(n11711), .Z(n11710) );
  XNOR U11336 ( .A(n11712), .B(n11713), .Z(n11707) );
  AND U11337 ( .A(n277), .B(n11714), .Z(n11713) );
  XOR U11338 ( .A(p_input[365]), .B(n11712), .Z(n11714) );
  XNOR U11339 ( .A(n11715), .B(n11716), .Z(n11712) );
  AND U11340 ( .A(n281), .B(n11711), .Z(n11716) );
  XNOR U11341 ( .A(n11715), .B(n11709), .Z(n11711) );
  XOR U11342 ( .A(n11717), .B(n11718), .Z(n11709) );
  AND U11343 ( .A(n296), .B(n11719), .Z(n11718) );
  XNOR U11344 ( .A(n11720), .B(n11721), .Z(n11715) );
  AND U11345 ( .A(n288), .B(n11722), .Z(n11721) );
  XOR U11346 ( .A(p_input[381]), .B(n11720), .Z(n11722) );
  XNOR U11347 ( .A(n11723), .B(n11724), .Z(n11720) );
  AND U11348 ( .A(n292), .B(n11719), .Z(n11724) );
  XNOR U11349 ( .A(n11723), .B(n11717), .Z(n11719) );
  XOR U11350 ( .A(n11725), .B(n11726), .Z(n11717) );
  AND U11351 ( .A(n307), .B(n11727), .Z(n11726) );
  XNOR U11352 ( .A(n11728), .B(n11729), .Z(n11723) );
  AND U11353 ( .A(n299), .B(n11730), .Z(n11729) );
  XOR U11354 ( .A(p_input[397]), .B(n11728), .Z(n11730) );
  XNOR U11355 ( .A(n11731), .B(n11732), .Z(n11728) );
  AND U11356 ( .A(n303), .B(n11727), .Z(n11732) );
  XNOR U11357 ( .A(n11731), .B(n11725), .Z(n11727) );
  XOR U11358 ( .A(n11733), .B(n11734), .Z(n11725) );
  AND U11359 ( .A(n318), .B(n11735), .Z(n11734) );
  XNOR U11360 ( .A(n11736), .B(n11737), .Z(n11731) );
  AND U11361 ( .A(n310), .B(n11738), .Z(n11737) );
  XOR U11362 ( .A(p_input[413]), .B(n11736), .Z(n11738) );
  XNOR U11363 ( .A(n11739), .B(n11740), .Z(n11736) );
  AND U11364 ( .A(n314), .B(n11735), .Z(n11740) );
  XNOR U11365 ( .A(n11739), .B(n11733), .Z(n11735) );
  XOR U11366 ( .A(n11741), .B(n11742), .Z(n11733) );
  AND U11367 ( .A(n329), .B(n11743), .Z(n11742) );
  XNOR U11368 ( .A(n11744), .B(n11745), .Z(n11739) );
  AND U11369 ( .A(n321), .B(n11746), .Z(n11745) );
  XOR U11370 ( .A(p_input[429]), .B(n11744), .Z(n11746) );
  XNOR U11371 ( .A(n11747), .B(n11748), .Z(n11744) );
  AND U11372 ( .A(n325), .B(n11743), .Z(n11748) );
  XNOR U11373 ( .A(n11747), .B(n11741), .Z(n11743) );
  XOR U11374 ( .A(n11749), .B(n11750), .Z(n11741) );
  AND U11375 ( .A(n340), .B(n11751), .Z(n11750) );
  XNOR U11376 ( .A(n11752), .B(n11753), .Z(n11747) );
  AND U11377 ( .A(n332), .B(n11754), .Z(n11753) );
  XOR U11378 ( .A(p_input[445]), .B(n11752), .Z(n11754) );
  XNOR U11379 ( .A(n11755), .B(n11756), .Z(n11752) );
  AND U11380 ( .A(n336), .B(n11751), .Z(n11756) );
  XNOR U11381 ( .A(n11755), .B(n11749), .Z(n11751) );
  XOR U11382 ( .A(n11757), .B(n11758), .Z(n11749) );
  AND U11383 ( .A(n351), .B(n11759), .Z(n11758) );
  XNOR U11384 ( .A(n11760), .B(n11761), .Z(n11755) );
  AND U11385 ( .A(n343), .B(n11762), .Z(n11761) );
  XOR U11386 ( .A(p_input[461]), .B(n11760), .Z(n11762) );
  XNOR U11387 ( .A(n11763), .B(n11764), .Z(n11760) );
  AND U11388 ( .A(n347), .B(n11759), .Z(n11764) );
  XNOR U11389 ( .A(n11763), .B(n11757), .Z(n11759) );
  XOR U11390 ( .A(n11765), .B(n11766), .Z(n11757) );
  AND U11391 ( .A(n362), .B(n11767), .Z(n11766) );
  XNOR U11392 ( .A(n11768), .B(n11769), .Z(n11763) );
  AND U11393 ( .A(n354), .B(n11770), .Z(n11769) );
  XOR U11394 ( .A(p_input[477]), .B(n11768), .Z(n11770) );
  XNOR U11395 ( .A(n11771), .B(n11772), .Z(n11768) );
  AND U11396 ( .A(n358), .B(n11767), .Z(n11772) );
  XNOR U11397 ( .A(n11771), .B(n11765), .Z(n11767) );
  XOR U11398 ( .A(n11773), .B(n11774), .Z(n11765) );
  AND U11399 ( .A(n373), .B(n11775), .Z(n11774) );
  XNOR U11400 ( .A(n11776), .B(n11777), .Z(n11771) );
  AND U11401 ( .A(n365), .B(n11778), .Z(n11777) );
  XOR U11402 ( .A(p_input[493]), .B(n11776), .Z(n11778) );
  XNOR U11403 ( .A(n11779), .B(n11780), .Z(n11776) );
  AND U11404 ( .A(n369), .B(n11775), .Z(n11780) );
  XNOR U11405 ( .A(n11779), .B(n11773), .Z(n11775) );
  XOR U11406 ( .A(n11781), .B(n11782), .Z(n11773) );
  AND U11407 ( .A(n384), .B(n11783), .Z(n11782) );
  XNOR U11408 ( .A(n11784), .B(n11785), .Z(n11779) );
  AND U11409 ( .A(n376), .B(n11786), .Z(n11785) );
  XOR U11410 ( .A(p_input[509]), .B(n11784), .Z(n11786) );
  XNOR U11411 ( .A(n11787), .B(n11788), .Z(n11784) );
  AND U11412 ( .A(n380), .B(n11783), .Z(n11788) );
  XNOR U11413 ( .A(n11787), .B(n11781), .Z(n11783) );
  XOR U11414 ( .A(n11789), .B(n11790), .Z(n11781) );
  AND U11415 ( .A(n395), .B(n11791), .Z(n11790) );
  XNOR U11416 ( .A(n11792), .B(n11793), .Z(n11787) );
  AND U11417 ( .A(n387), .B(n11794), .Z(n11793) );
  XOR U11418 ( .A(p_input[525]), .B(n11792), .Z(n11794) );
  XNOR U11419 ( .A(n11795), .B(n11796), .Z(n11792) );
  AND U11420 ( .A(n391), .B(n11791), .Z(n11796) );
  XNOR U11421 ( .A(n11795), .B(n11789), .Z(n11791) );
  XOR U11422 ( .A(n11797), .B(n11798), .Z(n11789) );
  AND U11423 ( .A(n406), .B(n11799), .Z(n11798) );
  XNOR U11424 ( .A(n11800), .B(n11801), .Z(n11795) );
  AND U11425 ( .A(n398), .B(n11802), .Z(n11801) );
  XOR U11426 ( .A(p_input[541]), .B(n11800), .Z(n11802) );
  XNOR U11427 ( .A(n11803), .B(n11804), .Z(n11800) );
  AND U11428 ( .A(n402), .B(n11799), .Z(n11804) );
  XNOR U11429 ( .A(n11803), .B(n11797), .Z(n11799) );
  XOR U11430 ( .A(n11805), .B(n11806), .Z(n11797) );
  AND U11431 ( .A(n417), .B(n11807), .Z(n11806) );
  XNOR U11432 ( .A(n11808), .B(n11809), .Z(n11803) );
  AND U11433 ( .A(n409), .B(n11810), .Z(n11809) );
  XOR U11434 ( .A(p_input[557]), .B(n11808), .Z(n11810) );
  XNOR U11435 ( .A(n11811), .B(n11812), .Z(n11808) );
  AND U11436 ( .A(n413), .B(n11807), .Z(n11812) );
  XNOR U11437 ( .A(n11811), .B(n11805), .Z(n11807) );
  XOR U11438 ( .A(n11813), .B(n11814), .Z(n11805) );
  AND U11439 ( .A(n428), .B(n11815), .Z(n11814) );
  XNOR U11440 ( .A(n11816), .B(n11817), .Z(n11811) );
  AND U11441 ( .A(n420), .B(n11818), .Z(n11817) );
  XOR U11442 ( .A(p_input[573]), .B(n11816), .Z(n11818) );
  XNOR U11443 ( .A(n11819), .B(n11820), .Z(n11816) );
  AND U11444 ( .A(n424), .B(n11815), .Z(n11820) );
  XNOR U11445 ( .A(n11819), .B(n11813), .Z(n11815) );
  XOR U11446 ( .A(n11821), .B(n11822), .Z(n11813) );
  AND U11447 ( .A(n439), .B(n11823), .Z(n11822) );
  XNOR U11448 ( .A(n11824), .B(n11825), .Z(n11819) );
  AND U11449 ( .A(n431), .B(n11826), .Z(n11825) );
  XOR U11450 ( .A(p_input[589]), .B(n11824), .Z(n11826) );
  XNOR U11451 ( .A(n11827), .B(n11828), .Z(n11824) );
  AND U11452 ( .A(n435), .B(n11823), .Z(n11828) );
  XNOR U11453 ( .A(n11827), .B(n11821), .Z(n11823) );
  XOR U11454 ( .A(n11829), .B(n11830), .Z(n11821) );
  AND U11455 ( .A(n450), .B(n11831), .Z(n11830) );
  XNOR U11456 ( .A(n11832), .B(n11833), .Z(n11827) );
  AND U11457 ( .A(n442), .B(n11834), .Z(n11833) );
  XOR U11458 ( .A(p_input[605]), .B(n11832), .Z(n11834) );
  XNOR U11459 ( .A(n11835), .B(n11836), .Z(n11832) );
  AND U11460 ( .A(n446), .B(n11831), .Z(n11836) );
  XNOR U11461 ( .A(n11835), .B(n11829), .Z(n11831) );
  XOR U11462 ( .A(n11837), .B(n11838), .Z(n11829) );
  AND U11463 ( .A(n461), .B(n11839), .Z(n11838) );
  XNOR U11464 ( .A(n11840), .B(n11841), .Z(n11835) );
  AND U11465 ( .A(n453), .B(n11842), .Z(n11841) );
  XOR U11466 ( .A(p_input[621]), .B(n11840), .Z(n11842) );
  XNOR U11467 ( .A(n11843), .B(n11844), .Z(n11840) );
  AND U11468 ( .A(n457), .B(n11839), .Z(n11844) );
  XNOR U11469 ( .A(n11843), .B(n11837), .Z(n11839) );
  XOR U11470 ( .A(n11845), .B(n11846), .Z(n11837) );
  AND U11471 ( .A(n472), .B(n11847), .Z(n11846) );
  XNOR U11472 ( .A(n11848), .B(n11849), .Z(n11843) );
  AND U11473 ( .A(n464), .B(n11850), .Z(n11849) );
  XOR U11474 ( .A(p_input[637]), .B(n11848), .Z(n11850) );
  XNOR U11475 ( .A(n11851), .B(n11852), .Z(n11848) );
  AND U11476 ( .A(n468), .B(n11847), .Z(n11852) );
  XNOR U11477 ( .A(n11851), .B(n11845), .Z(n11847) );
  XOR U11478 ( .A(n11853), .B(n11854), .Z(n11845) );
  AND U11479 ( .A(n483), .B(n11855), .Z(n11854) );
  XNOR U11480 ( .A(n11856), .B(n11857), .Z(n11851) );
  AND U11481 ( .A(n475), .B(n11858), .Z(n11857) );
  XOR U11482 ( .A(p_input[653]), .B(n11856), .Z(n11858) );
  XNOR U11483 ( .A(n11859), .B(n11860), .Z(n11856) );
  AND U11484 ( .A(n479), .B(n11855), .Z(n11860) );
  XNOR U11485 ( .A(n11859), .B(n11853), .Z(n11855) );
  XOR U11486 ( .A(n11861), .B(n11862), .Z(n11853) );
  AND U11487 ( .A(n494), .B(n11863), .Z(n11862) );
  XNOR U11488 ( .A(n11864), .B(n11865), .Z(n11859) );
  AND U11489 ( .A(n486), .B(n11866), .Z(n11865) );
  XOR U11490 ( .A(p_input[669]), .B(n11864), .Z(n11866) );
  XNOR U11491 ( .A(n11867), .B(n11868), .Z(n11864) );
  AND U11492 ( .A(n490), .B(n11863), .Z(n11868) );
  XNOR U11493 ( .A(n11867), .B(n11861), .Z(n11863) );
  XOR U11494 ( .A(n11869), .B(n11870), .Z(n11861) );
  AND U11495 ( .A(n505), .B(n11871), .Z(n11870) );
  XNOR U11496 ( .A(n11872), .B(n11873), .Z(n11867) );
  AND U11497 ( .A(n497), .B(n11874), .Z(n11873) );
  XOR U11498 ( .A(p_input[685]), .B(n11872), .Z(n11874) );
  XNOR U11499 ( .A(n11875), .B(n11876), .Z(n11872) );
  AND U11500 ( .A(n501), .B(n11871), .Z(n11876) );
  XNOR U11501 ( .A(n11875), .B(n11869), .Z(n11871) );
  XOR U11502 ( .A(n11877), .B(n11878), .Z(n11869) );
  AND U11503 ( .A(n516), .B(n11879), .Z(n11878) );
  XNOR U11504 ( .A(n11880), .B(n11881), .Z(n11875) );
  AND U11505 ( .A(n508), .B(n11882), .Z(n11881) );
  XOR U11506 ( .A(p_input[701]), .B(n11880), .Z(n11882) );
  XNOR U11507 ( .A(n11883), .B(n11884), .Z(n11880) );
  AND U11508 ( .A(n512), .B(n11879), .Z(n11884) );
  XNOR U11509 ( .A(n11883), .B(n11877), .Z(n11879) );
  XOR U11510 ( .A(n11885), .B(n11886), .Z(n11877) );
  AND U11511 ( .A(n527), .B(n11887), .Z(n11886) );
  XNOR U11512 ( .A(n11888), .B(n11889), .Z(n11883) );
  AND U11513 ( .A(n519), .B(n11890), .Z(n11889) );
  XOR U11514 ( .A(p_input[717]), .B(n11888), .Z(n11890) );
  XNOR U11515 ( .A(n11891), .B(n11892), .Z(n11888) );
  AND U11516 ( .A(n523), .B(n11887), .Z(n11892) );
  XNOR U11517 ( .A(n11891), .B(n11885), .Z(n11887) );
  XOR U11518 ( .A(n11893), .B(n11894), .Z(n11885) );
  AND U11519 ( .A(n538), .B(n11895), .Z(n11894) );
  XNOR U11520 ( .A(n11896), .B(n11897), .Z(n11891) );
  AND U11521 ( .A(n530), .B(n11898), .Z(n11897) );
  XOR U11522 ( .A(p_input[733]), .B(n11896), .Z(n11898) );
  XNOR U11523 ( .A(n11899), .B(n11900), .Z(n11896) );
  AND U11524 ( .A(n534), .B(n11895), .Z(n11900) );
  XNOR U11525 ( .A(n11899), .B(n11893), .Z(n11895) );
  XOR U11526 ( .A(n11901), .B(n11902), .Z(n11893) );
  AND U11527 ( .A(n549), .B(n11903), .Z(n11902) );
  XNOR U11528 ( .A(n11904), .B(n11905), .Z(n11899) );
  AND U11529 ( .A(n541), .B(n11906), .Z(n11905) );
  XOR U11530 ( .A(p_input[749]), .B(n11904), .Z(n11906) );
  XNOR U11531 ( .A(n11907), .B(n11908), .Z(n11904) );
  AND U11532 ( .A(n545), .B(n11903), .Z(n11908) );
  XNOR U11533 ( .A(n11907), .B(n11901), .Z(n11903) );
  XOR U11534 ( .A(n11909), .B(n11910), .Z(n11901) );
  AND U11535 ( .A(n560), .B(n11911), .Z(n11910) );
  XNOR U11536 ( .A(n11912), .B(n11913), .Z(n11907) );
  AND U11537 ( .A(n552), .B(n11914), .Z(n11913) );
  XOR U11538 ( .A(p_input[765]), .B(n11912), .Z(n11914) );
  XNOR U11539 ( .A(n11915), .B(n11916), .Z(n11912) );
  AND U11540 ( .A(n556), .B(n11911), .Z(n11916) );
  XNOR U11541 ( .A(n11915), .B(n11909), .Z(n11911) );
  XOR U11542 ( .A(n11917), .B(n11918), .Z(n11909) );
  AND U11543 ( .A(n571), .B(n11919), .Z(n11918) );
  XNOR U11544 ( .A(n11920), .B(n11921), .Z(n11915) );
  AND U11545 ( .A(n563), .B(n11922), .Z(n11921) );
  XOR U11546 ( .A(p_input[781]), .B(n11920), .Z(n11922) );
  XNOR U11547 ( .A(n11923), .B(n11924), .Z(n11920) );
  AND U11548 ( .A(n567), .B(n11919), .Z(n11924) );
  XNOR U11549 ( .A(n11923), .B(n11917), .Z(n11919) );
  XOR U11550 ( .A(n11925), .B(n11926), .Z(n11917) );
  AND U11551 ( .A(n582), .B(n11927), .Z(n11926) );
  XNOR U11552 ( .A(n11928), .B(n11929), .Z(n11923) );
  AND U11553 ( .A(n574), .B(n11930), .Z(n11929) );
  XOR U11554 ( .A(p_input[797]), .B(n11928), .Z(n11930) );
  XNOR U11555 ( .A(n11931), .B(n11932), .Z(n11928) );
  AND U11556 ( .A(n578), .B(n11927), .Z(n11932) );
  XNOR U11557 ( .A(n11931), .B(n11925), .Z(n11927) );
  XOR U11558 ( .A(n11933), .B(n11934), .Z(n11925) );
  AND U11559 ( .A(n593), .B(n11935), .Z(n11934) );
  XNOR U11560 ( .A(n11936), .B(n11937), .Z(n11931) );
  AND U11561 ( .A(n585), .B(n11938), .Z(n11937) );
  XOR U11562 ( .A(p_input[813]), .B(n11936), .Z(n11938) );
  XNOR U11563 ( .A(n11939), .B(n11940), .Z(n11936) );
  AND U11564 ( .A(n589), .B(n11935), .Z(n11940) );
  XNOR U11565 ( .A(n11939), .B(n11933), .Z(n11935) );
  XOR U11566 ( .A(n11941), .B(n11942), .Z(n11933) );
  AND U11567 ( .A(n604), .B(n11943), .Z(n11942) );
  XNOR U11568 ( .A(n11944), .B(n11945), .Z(n11939) );
  AND U11569 ( .A(n596), .B(n11946), .Z(n11945) );
  XOR U11570 ( .A(p_input[829]), .B(n11944), .Z(n11946) );
  XNOR U11571 ( .A(n11947), .B(n11948), .Z(n11944) );
  AND U11572 ( .A(n600), .B(n11943), .Z(n11948) );
  XNOR U11573 ( .A(n11947), .B(n11941), .Z(n11943) );
  XOR U11574 ( .A(n11949), .B(n11950), .Z(n11941) );
  AND U11575 ( .A(n615), .B(n11951), .Z(n11950) );
  XNOR U11576 ( .A(n11952), .B(n11953), .Z(n11947) );
  AND U11577 ( .A(n607), .B(n11954), .Z(n11953) );
  XOR U11578 ( .A(p_input[845]), .B(n11952), .Z(n11954) );
  XNOR U11579 ( .A(n11955), .B(n11956), .Z(n11952) );
  AND U11580 ( .A(n611), .B(n11951), .Z(n11956) );
  XNOR U11581 ( .A(n11955), .B(n11949), .Z(n11951) );
  XOR U11582 ( .A(n11957), .B(n11958), .Z(n11949) );
  AND U11583 ( .A(n626), .B(n11959), .Z(n11958) );
  XNOR U11584 ( .A(n11960), .B(n11961), .Z(n11955) );
  AND U11585 ( .A(n618), .B(n11962), .Z(n11961) );
  XOR U11586 ( .A(p_input[861]), .B(n11960), .Z(n11962) );
  XNOR U11587 ( .A(n11963), .B(n11964), .Z(n11960) );
  AND U11588 ( .A(n622), .B(n11959), .Z(n11964) );
  XNOR U11589 ( .A(n11963), .B(n11957), .Z(n11959) );
  XOR U11590 ( .A(n11965), .B(n11966), .Z(n11957) );
  AND U11591 ( .A(n637), .B(n11967), .Z(n11966) );
  XNOR U11592 ( .A(n11968), .B(n11969), .Z(n11963) );
  AND U11593 ( .A(n629), .B(n11970), .Z(n11969) );
  XOR U11594 ( .A(p_input[877]), .B(n11968), .Z(n11970) );
  XNOR U11595 ( .A(n11971), .B(n11972), .Z(n11968) );
  AND U11596 ( .A(n633), .B(n11967), .Z(n11972) );
  XNOR U11597 ( .A(n11971), .B(n11965), .Z(n11967) );
  XOR U11598 ( .A(n11973), .B(n11974), .Z(n11965) );
  AND U11599 ( .A(n648), .B(n11975), .Z(n11974) );
  XNOR U11600 ( .A(n11976), .B(n11977), .Z(n11971) );
  AND U11601 ( .A(n640), .B(n11978), .Z(n11977) );
  XOR U11602 ( .A(p_input[893]), .B(n11976), .Z(n11978) );
  XNOR U11603 ( .A(n11979), .B(n11980), .Z(n11976) );
  AND U11604 ( .A(n644), .B(n11975), .Z(n11980) );
  XNOR U11605 ( .A(n11979), .B(n11973), .Z(n11975) );
  XOR U11606 ( .A(n11981), .B(n11982), .Z(n11973) );
  AND U11607 ( .A(n659), .B(n11983), .Z(n11982) );
  XNOR U11608 ( .A(n11984), .B(n11985), .Z(n11979) );
  AND U11609 ( .A(n651), .B(n11986), .Z(n11985) );
  XOR U11610 ( .A(p_input[909]), .B(n11984), .Z(n11986) );
  XNOR U11611 ( .A(n11987), .B(n11988), .Z(n11984) );
  AND U11612 ( .A(n655), .B(n11983), .Z(n11988) );
  XNOR U11613 ( .A(n11987), .B(n11981), .Z(n11983) );
  XOR U11614 ( .A(n11989), .B(n11990), .Z(n11981) );
  AND U11615 ( .A(n670), .B(n11991), .Z(n11990) );
  XNOR U11616 ( .A(n11992), .B(n11993), .Z(n11987) );
  AND U11617 ( .A(n662), .B(n11994), .Z(n11993) );
  XOR U11618 ( .A(p_input[925]), .B(n11992), .Z(n11994) );
  XNOR U11619 ( .A(n11995), .B(n11996), .Z(n11992) );
  AND U11620 ( .A(n666), .B(n11991), .Z(n11996) );
  XNOR U11621 ( .A(n11995), .B(n11989), .Z(n11991) );
  XOR U11622 ( .A(n11997), .B(n11998), .Z(n11989) );
  AND U11623 ( .A(n681), .B(n11999), .Z(n11998) );
  XNOR U11624 ( .A(n12000), .B(n12001), .Z(n11995) );
  AND U11625 ( .A(n673), .B(n12002), .Z(n12001) );
  XOR U11626 ( .A(p_input[941]), .B(n12000), .Z(n12002) );
  XNOR U11627 ( .A(n12003), .B(n12004), .Z(n12000) );
  AND U11628 ( .A(n677), .B(n11999), .Z(n12004) );
  XNOR U11629 ( .A(n12003), .B(n11997), .Z(n11999) );
  XOR U11630 ( .A(n12005), .B(n12006), .Z(n11997) );
  AND U11631 ( .A(n692), .B(n12007), .Z(n12006) );
  XNOR U11632 ( .A(n12008), .B(n12009), .Z(n12003) );
  AND U11633 ( .A(n684), .B(n12010), .Z(n12009) );
  XOR U11634 ( .A(p_input[957]), .B(n12008), .Z(n12010) );
  XNOR U11635 ( .A(n12011), .B(n12012), .Z(n12008) );
  AND U11636 ( .A(n688), .B(n12007), .Z(n12012) );
  XNOR U11637 ( .A(n12011), .B(n12005), .Z(n12007) );
  XOR U11638 ( .A(n12013), .B(n12014), .Z(n12005) );
  AND U11639 ( .A(n703), .B(n12015), .Z(n12014) );
  XNOR U11640 ( .A(n12016), .B(n12017), .Z(n12011) );
  AND U11641 ( .A(n695), .B(n12018), .Z(n12017) );
  XOR U11642 ( .A(p_input[973]), .B(n12016), .Z(n12018) );
  XNOR U11643 ( .A(n12019), .B(n12020), .Z(n12016) );
  AND U11644 ( .A(n699), .B(n12015), .Z(n12020) );
  XNOR U11645 ( .A(n12019), .B(n12013), .Z(n12015) );
  XOR U11646 ( .A(n12021), .B(n12022), .Z(n12013) );
  AND U11647 ( .A(n714), .B(n12023), .Z(n12022) );
  XNOR U11648 ( .A(n12024), .B(n12025), .Z(n12019) );
  AND U11649 ( .A(n706), .B(n12026), .Z(n12025) );
  XOR U11650 ( .A(p_input[989]), .B(n12024), .Z(n12026) );
  XNOR U11651 ( .A(n12027), .B(n12028), .Z(n12024) );
  AND U11652 ( .A(n710), .B(n12023), .Z(n12028) );
  XNOR U11653 ( .A(n12027), .B(n12021), .Z(n12023) );
  XOR U11654 ( .A(n12029), .B(n12030), .Z(n12021) );
  AND U11655 ( .A(n725), .B(n12031), .Z(n12030) );
  XNOR U11656 ( .A(n12032), .B(n12033), .Z(n12027) );
  AND U11657 ( .A(n717), .B(n12034), .Z(n12033) );
  XOR U11658 ( .A(p_input[1005]), .B(n12032), .Z(n12034) );
  XNOR U11659 ( .A(n12035), .B(n12036), .Z(n12032) );
  AND U11660 ( .A(n721), .B(n12031), .Z(n12036) );
  XNOR U11661 ( .A(n12035), .B(n12029), .Z(n12031) );
  XOR U11662 ( .A(n12037), .B(n12038), .Z(n12029) );
  AND U11663 ( .A(n736), .B(n12039), .Z(n12038) );
  XNOR U11664 ( .A(n12040), .B(n12041), .Z(n12035) );
  AND U11665 ( .A(n728), .B(n12042), .Z(n12041) );
  XOR U11666 ( .A(p_input[1021]), .B(n12040), .Z(n12042) );
  XNOR U11667 ( .A(n12043), .B(n12044), .Z(n12040) );
  AND U11668 ( .A(n732), .B(n12039), .Z(n12044) );
  XNOR U11669 ( .A(n12043), .B(n12037), .Z(n12039) );
  XOR U11670 ( .A(n12045), .B(n12046), .Z(n12037) );
  AND U11671 ( .A(n747), .B(n12047), .Z(n12046) );
  XNOR U11672 ( .A(n12048), .B(n12049), .Z(n12043) );
  AND U11673 ( .A(n739), .B(n12050), .Z(n12049) );
  XOR U11674 ( .A(p_input[1037]), .B(n12048), .Z(n12050) );
  XNOR U11675 ( .A(n12051), .B(n12052), .Z(n12048) );
  AND U11676 ( .A(n743), .B(n12047), .Z(n12052) );
  XNOR U11677 ( .A(n12051), .B(n12045), .Z(n12047) );
  XOR U11678 ( .A(n12053), .B(n12054), .Z(n12045) );
  AND U11679 ( .A(n758), .B(n12055), .Z(n12054) );
  XNOR U11680 ( .A(n12056), .B(n12057), .Z(n12051) );
  AND U11681 ( .A(n750), .B(n12058), .Z(n12057) );
  XOR U11682 ( .A(p_input[1053]), .B(n12056), .Z(n12058) );
  XNOR U11683 ( .A(n12059), .B(n12060), .Z(n12056) );
  AND U11684 ( .A(n754), .B(n12055), .Z(n12060) );
  XNOR U11685 ( .A(n12059), .B(n12053), .Z(n12055) );
  XOR U11686 ( .A(n12061), .B(n12062), .Z(n12053) );
  AND U11687 ( .A(n769), .B(n12063), .Z(n12062) );
  XNOR U11688 ( .A(n12064), .B(n12065), .Z(n12059) );
  AND U11689 ( .A(n761), .B(n12066), .Z(n12065) );
  XOR U11690 ( .A(p_input[1069]), .B(n12064), .Z(n12066) );
  XNOR U11691 ( .A(n12067), .B(n12068), .Z(n12064) );
  AND U11692 ( .A(n765), .B(n12063), .Z(n12068) );
  XNOR U11693 ( .A(n12067), .B(n12061), .Z(n12063) );
  XOR U11694 ( .A(n12069), .B(n12070), .Z(n12061) );
  AND U11695 ( .A(n780), .B(n12071), .Z(n12070) );
  XNOR U11696 ( .A(n12072), .B(n12073), .Z(n12067) );
  AND U11697 ( .A(n772), .B(n12074), .Z(n12073) );
  XOR U11698 ( .A(p_input[1085]), .B(n12072), .Z(n12074) );
  XNOR U11699 ( .A(n12075), .B(n12076), .Z(n12072) );
  AND U11700 ( .A(n776), .B(n12071), .Z(n12076) );
  XNOR U11701 ( .A(n12075), .B(n12069), .Z(n12071) );
  XOR U11702 ( .A(n12077), .B(n12078), .Z(n12069) );
  AND U11703 ( .A(n791), .B(n12079), .Z(n12078) );
  XNOR U11704 ( .A(n12080), .B(n12081), .Z(n12075) );
  AND U11705 ( .A(n783), .B(n12082), .Z(n12081) );
  XOR U11706 ( .A(p_input[1101]), .B(n12080), .Z(n12082) );
  XNOR U11707 ( .A(n12083), .B(n12084), .Z(n12080) );
  AND U11708 ( .A(n787), .B(n12079), .Z(n12084) );
  XNOR U11709 ( .A(n12083), .B(n12077), .Z(n12079) );
  XOR U11710 ( .A(n12085), .B(n12086), .Z(n12077) );
  AND U11711 ( .A(n802), .B(n12087), .Z(n12086) );
  XNOR U11712 ( .A(n12088), .B(n12089), .Z(n12083) );
  AND U11713 ( .A(n794), .B(n12090), .Z(n12089) );
  XOR U11714 ( .A(p_input[1117]), .B(n12088), .Z(n12090) );
  XNOR U11715 ( .A(n12091), .B(n12092), .Z(n12088) );
  AND U11716 ( .A(n798), .B(n12087), .Z(n12092) );
  XNOR U11717 ( .A(n12091), .B(n12085), .Z(n12087) );
  XOR U11718 ( .A(n12093), .B(n12094), .Z(n12085) );
  AND U11719 ( .A(n813), .B(n12095), .Z(n12094) );
  XNOR U11720 ( .A(n12096), .B(n12097), .Z(n12091) );
  AND U11721 ( .A(n805), .B(n12098), .Z(n12097) );
  XOR U11722 ( .A(p_input[1133]), .B(n12096), .Z(n12098) );
  XNOR U11723 ( .A(n12099), .B(n12100), .Z(n12096) );
  AND U11724 ( .A(n809), .B(n12095), .Z(n12100) );
  XNOR U11725 ( .A(n12099), .B(n12093), .Z(n12095) );
  XOR U11726 ( .A(n12101), .B(n12102), .Z(n12093) );
  AND U11727 ( .A(n824), .B(n12103), .Z(n12102) );
  XNOR U11728 ( .A(n12104), .B(n12105), .Z(n12099) );
  AND U11729 ( .A(n816), .B(n12106), .Z(n12105) );
  XOR U11730 ( .A(p_input[1149]), .B(n12104), .Z(n12106) );
  XNOR U11731 ( .A(n12107), .B(n12108), .Z(n12104) );
  AND U11732 ( .A(n820), .B(n12103), .Z(n12108) );
  XNOR U11733 ( .A(n12107), .B(n12101), .Z(n12103) );
  XOR U11734 ( .A(n12109), .B(n12110), .Z(n12101) );
  AND U11735 ( .A(n835), .B(n12111), .Z(n12110) );
  XNOR U11736 ( .A(n12112), .B(n12113), .Z(n12107) );
  AND U11737 ( .A(n827), .B(n12114), .Z(n12113) );
  XOR U11738 ( .A(p_input[1165]), .B(n12112), .Z(n12114) );
  XNOR U11739 ( .A(n12115), .B(n12116), .Z(n12112) );
  AND U11740 ( .A(n831), .B(n12111), .Z(n12116) );
  XNOR U11741 ( .A(n12115), .B(n12109), .Z(n12111) );
  XOR U11742 ( .A(n12117), .B(n12118), .Z(n12109) );
  AND U11743 ( .A(n846), .B(n12119), .Z(n12118) );
  XNOR U11744 ( .A(n12120), .B(n12121), .Z(n12115) );
  AND U11745 ( .A(n838), .B(n12122), .Z(n12121) );
  XOR U11746 ( .A(p_input[1181]), .B(n12120), .Z(n12122) );
  XNOR U11747 ( .A(n12123), .B(n12124), .Z(n12120) );
  AND U11748 ( .A(n842), .B(n12119), .Z(n12124) );
  XNOR U11749 ( .A(n12123), .B(n12117), .Z(n12119) );
  XOR U11750 ( .A(n12125), .B(n12126), .Z(n12117) );
  AND U11751 ( .A(n857), .B(n12127), .Z(n12126) );
  XNOR U11752 ( .A(n12128), .B(n12129), .Z(n12123) );
  AND U11753 ( .A(n849), .B(n12130), .Z(n12129) );
  XOR U11754 ( .A(p_input[1197]), .B(n12128), .Z(n12130) );
  XNOR U11755 ( .A(n12131), .B(n12132), .Z(n12128) );
  AND U11756 ( .A(n853), .B(n12127), .Z(n12132) );
  XNOR U11757 ( .A(n12131), .B(n12125), .Z(n12127) );
  XOR U11758 ( .A(n12133), .B(n12134), .Z(n12125) );
  AND U11759 ( .A(n868), .B(n12135), .Z(n12134) );
  XNOR U11760 ( .A(n12136), .B(n12137), .Z(n12131) );
  AND U11761 ( .A(n860), .B(n12138), .Z(n12137) );
  XOR U11762 ( .A(p_input[1213]), .B(n12136), .Z(n12138) );
  XNOR U11763 ( .A(n12139), .B(n12140), .Z(n12136) );
  AND U11764 ( .A(n864), .B(n12135), .Z(n12140) );
  XNOR U11765 ( .A(n12139), .B(n12133), .Z(n12135) );
  XOR U11766 ( .A(n12141), .B(n12142), .Z(n12133) );
  AND U11767 ( .A(n879), .B(n12143), .Z(n12142) );
  XNOR U11768 ( .A(n12144), .B(n12145), .Z(n12139) );
  AND U11769 ( .A(n871), .B(n12146), .Z(n12145) );
  XOR U11770 ( .A(p_input[1229]), .B(n12144), .Z(n12146) );
  XNOR U11771 ( .A(n12147), .B(n12148), .Z(n12144) );
  AND U11772 ( .A(n875), .B(n12143), .Z(n12148) );
  XNOR U11773 ( .A(n12147), .B(n12141), .Z(n12143) );
  XOR U11774 ( .A(n12149), .B(n12150), .Z(n12141) );
  AND U11775 ( .A(n890), .B(n12151), .Z(n12150) );
  XNOR U11776 ( .A(n12152), .B(n12153), .Z(n12147) );
  AND U11777 ( .A(n882), .B(n12154), .Z(n12153) );
  XOR U11778 ( .A(p_input[1245]), .B(n12152), .Z(n12154) );
  XNOR U11779 ( .A(n12155), .B(n12156), .Z(n12152) );
  AND U11780 ( .A(n886), .B(n12151), .Z(n12156) );
  XNOR U11781 ( .A(n12155), .B(n12149), .Z(n12151) );
  XOR U11782 ( .A(n12157), .B(n12158), .Z(n12149) );
  AND U11783 ( .A(n901), .B(n12159), .Z(n12158) );
  XNOR U11784 ( .A(n12160), .B(n12161), .Z(n12155) );
  AND U11785 ( .A(n893), .B(n12162), .Z(n12161) );
  XOR U11786 ( .A(p_input[1261]), .B(n12160), .Z(n12162) );
  XNOR U11787 ( .A(n12163), .B(n12164), .Z(n12160) );
  AND U11788 ( .A(n897), .B(n12159), .Z(n12164) );
  XNOR U11789 ( .A(n12163), .B(n12157), .Z(n12159) );
  XOR U11790 ( .A(n12165), .B(n12166), .Z(n12157) );
  AND U11791 ( .A(n912), .B(n12167), .Z(n12166) );
  XNOR U11792 ( .A(n12168), .B(n12169), .Z(n12163) );
  AND U11793 ( .A(n904), .B(n12170), .Z(n12169) );
  XOR U11794 ( .A(p_input[1277]), .B(n12168), .Z(n12170) );
  XNOR U11795 ( .A(n12171), .B(n12172), .Z(n12168) );
  AND U11796 ( .A(n908), .B(n12167), .Z(n12172) );
  XNOR U11797 ( .A(n12171), .B(n12165), .Z(n12167) );
  XOR U11798 ( .A(n12173), .B(n12174), .Z(n12165) );
  AND U11799 ( .A(n923), .B(n12175), .Z(n12174) );
  XNOR U11800 ( .A(n12176), .B(n12177), .Z(n12171) );
  AND U11801 ( .A(n915), .B(n12178), .Z(n12177) );
  XOR U11802 ( .A(p_input[1293]), .B(n12176), .Z(n12178) );
  XNOR U11803 ( .A(n12179), .B(n12180), .Z(n12176) );
  AND U11804 ( .A(n919), .B(n12175), .Z(n12180) );
  XNOR U11805 ( .A(n12179), .B(n12173), .Z(n12175) );
  XOR U11806 ( .A(n12181), .B(n12182), .Z(n12173) );
  AND U11807 ( .A(n934), .B(n12183), .Z(n12182) );
  XNOR U11808 ( .A(n12184), .B(n12185), .Z(n12179) );
  AND U11809 ( .A(n926), .B(n12186), .Z(n12185) );
  XOR U11810 ( .A(p_input[1309]), .B(n12184), .Z(n12186) );
  XNOR U11811 ( .A(n12187), .B(n12188), .Z(n12184) );
  AND U11812 ( .A(n930), .B(n12183), .Z(n12188) );
  XNOR U11813 ( .A(n12187), .B(n12181), .Z(n12183) );
  XOR U11814 ( .A(n12189), .B(n12190), .Z(n12181) );
  AND U11815 ( .A(n945), .B(n12191), .Z(n12190) );
  XNOR U11816 ( .A(n12192), .B(n12193), .Z(n12187) );
  AND U11817 ( .A(n937), .B(n12194), .Z(n12193) );
  XOR U11818 ( .A(p_input[1325]), .B(n12192), .Z(n12194) );
  XNOR U11819 ( .A(n12195), .B(n12196), .Z(n12192) );
  AND U11820 ( .A(n941), .B(n12191), .Z(n12196) );
  XNOR U11821 ( .A(n12195), .B(n12189), .Z(n12191) );
  XOR U11822 ( .A(n12197), .B(n12198), .Z(n12189) );
  AND U11823 ( .A(n956), .B(n12199), .Z(n12198) );
  XNOR U11824 ( .A(n12200), .B(n12201), .Z(n12195) );
  AND U11825 ( .A(n948), .B(n12202), .Z(n12201) );
  XOR U11826 ( .A(p_input[1341]), .B(n12200), .Z(n12202) );
  XNOR U11827 ( .A(n12203), .B(n12204), .Z(n12200) );
  AND U11828 ( .A(n952), .B(n12199), .Z(n12204) );
  XNOR U11829 ( .A(n12203), .B(n12197), .Z(n12199) );
  XOR U11830 ( .A(n12205), .B(n12206), .Z(n12197) );
  AND U11831 ( .A(n967), .B(n12207), .Z(n12206) );
  XNOR U11832 ( .A(n12208), .B(n12209), .Z(n12203) );
  AND U11833 ( .A(n959), .B(n12210), .Z(n12209) );
  XOR U11834 ( .A(p_input[1357]), .B(n12208), .Z(n12210) );
  XNOR U11835 ( .A(n12211), .B(n12212), .Z(n12208) );
  AND U11836 ( .A(n963), .B(n12207), .Z(n12212) );
  XNOR U11837 ( .A(n12211), .B(n12205), .Z(n12207) );
  XOR U11838 ( .A(n12213), .B(n12214), .Z(n12205) );
  AND U11839 ( .A(n978), .B(n12215), .Z(n12214) );
  XNOR U11840 ( .A(n12216), .B(n12217), .Z(n12211) );
  AND U11841 ( .A(n970), .B(n12218), .Z(n12217) );
  XOR U11842 ( .A(p_input[1373]), .B(n12216), .Z(n12218) );
  XNOR U11843 ( .A(n12219), .B(n12220), .Z(n12216) );
  AND U11844 ( .A(n974), .B(n12215), .Z(n12220) );
  XNOR U11845 ( .A(n12219), .B(n12213), .Z(n12215) );
  XOR U11846 ( .A(n12221), .B(n12222), .Z(n12213) );
  AND U11847 ( .A(n989), .B(n12223), .Z(n12222) );
  XNOR U11848 ( .A(n12224), .B(n12225), .Z(n12219) );
  AND U11849 ( .A(n981), .B(n12226), .Z(n12225) );
  XOR U11850 ( .A(p_input[1389]), .B(n12224), .Z(n12226) );
  XNOR U11851 ( .A(n12227), .B(n12228), .Z(n12224) );
  AND U11852 ( .A(n985), .B(n12223), .Z(n12228) );
  XNOR U11853 ( .A(n12227), .B(n12221), .Z(n12223) );
  XOR U11854 ( .A(n12229), .B(n12230), .Z(n12221) );
  AND U11855 ( .A(n1000), .B(n12231), .Z(n12230) );
  XNOR U11856 ( .A(n12232), .B(n12233), .Z(n12227) );
  AND U11857 ( .A(n992), .B(n12234), .Z(n12233) );
  XOR U11858 ( .A(p_input[1405]), .B(n12232), .Z(n12234) );
  XNOR U11859 ( .A(n12235), .B(n12236), .Z(n12232) );
  AND U11860 ( .A(n996), .B(n12231), .Z(n12236) );
  XNOR U11861 ( .A(n12235), .B(n12229), .Z(n12231) );
  XOR U11862 ( .A(n12237), .B(n12238), .Z(n12229) );
  AND U11863 ( .A(n1011), .B(n12239), .Z(n12238) );
  XNOR U11864 ( .A(n12240), .B(n12241), .Z(n12235) );
  AND U11865 ( .A(n1003), .B(n12242), .Z(n12241) );
  XOR U11866 ( .A(p_input[1421]), .B(n12240), .Z(n12242) );
  XNOR U11867 ( .A(n12243), .B(n12244), .Z(n12240) );
  AND U11868 ( .A(n1007), .B(n12239), .Z(n12244) );
  XNOR U11869 ( .A(n12243), .B(n12237), .Z(n12239) );
  XOR U11870 ( .A(n12245), .B(n12246), .Z(n12237) );
  AND U11871 ( .A(n1022), .B(n12247), .Z(n12246) );
  XNOR U11872 ( .A(n12248), .B(n12249), .Z(n12243) );
  AND U11873 ( .A(n1014), .B(n12250), .Z(n12249) );
  XOR U11874 ( .A(p_input[1437]), .B(n12248), .Z(n12250) );
  XNOR U11875 ( .A(n12251), .B(n12252), .Z(n12248) );
  AND U11876 ( .A(n1018), .B(n12247), .Z(n12252) );
  XNOR U11877 ( .A(n12251), .B(n12245), .Z(n12247) );
  XOR U11878 ( .A(n12253), .B(n12254), .Z(n12245) );
  AND U11879 ( .A(n1033), .B(n12255), .Z(n12254) );
  XNOR U11880 ( .A(n12256), .B(n12257), .Z(n12251) );
  AND U11881 ( .A(n1025), .B(n12258), .Z(n12257) );
  XOR U11882 ( .A(p_input[1453]), .B(n12256), .Z(n12258) );
  XNOR U11883 ( .A(n12259), .B(n12260), .Z(n12256) );
  AND U11884 ( .A(n1029), .B(n12255), .Z(n12260) );
  XNOR U11885 ( .A(n12259), .B(n12253), .Z(n12255) );
  XOR U11886 ( .A(n12261), .B(n12262), .Z(n12253) );
  AND U11887 ( .A(n1044), .B(n12263), .Z(n12262) );
  XNOR U11888 ( .A(n12264), .B(n12265), .Z(n12259) );
  AND U11889 ( .A(n1036), .B(n12266), .Z(n12265) );
  XOR U11890 ( .A(p_input[1469]), .B(n12264), .Z(n12266) );
  XNOR U11891 ( .A(n12267), .B(n12268), .Z(n12264) );
  AND U11892 ( .A(n1040), .B(n12263), .Z(n12268) );
  XNOR U11893 ( .A(n12267), .B(n12261), .Z(n12263) );
  XOR U11894 ( .A(n12269), .B(n12270), .Z(n12261) );
  AND U11895 ( .A(n1055), .B(n12271), .Z(n12270) );
  XNOR U11896 ( .A(n12272), .B(n12273), .Z(n12267) );
  AND U11897 ( .A(n1047), .B(n12274), .Z(n12273) );
  XOR U11898 ( .A(p_input[1485]), .B(n12272), .Z(n12274) );
  XNOR U11899 ( .A(n12275), .B(n12276), .Z(n12272) );
  AND U11900 ( .A(n1051), .B(n12271), .Z(n12276) );
  XNOR U11901 ( .A(n12275), .B(n12269), .Z(n12271) );
  XOR U11902 ( .A(n12277), .B(n12278), .Z(n12269) );
  AND U11903 ( .A(n1066), .B(n12279), .Z(n12278) );
  XNOR U11904 ( .A(n12280), .B(n12281), .Z(n12275) );
  AND U11905 ( .A(n1058), .B(n12282), .Z(n12281) );
  XOR U11906 ( .A(p_input[1501]), .B(n12280), .Z(n12282) );
  XNOR U11907 ( .A(n12283), .B(n12284), .Z(n12280) );
  AND U11908 ( .A(n1062), .B(n12279), .Z(n12284) );
  XNOR U11909 ( .A(n12283), .B(n12277), .Z(n12279) );
  XOR U11910 ( .A(n12285), .B(n12286), .Z(n12277) );
  AND U11911 ( .A(n1077), .B(n12287), .Z(n12286) );
  XNOR U11912 ( .A(n12288), .B(n12289), .Z(n12283) );
  AND U11913 ( .A(n1069), .B(n12290), .Z(n12289) );
  XOR U11914 ( .A(p_input[1517]), .B(n12288), .Z(n12290) );
  XNOR U11915 ( .A(n12291), .B(n12292), .Z(n12288) );
  AND U11916 ( .A(n1073), .B(n12287), .Z(n12292) );
  XNOR U11917 ( .A(n12291), .B(n12285), .Z(n12287) );
  XOR U11918 ( .A(n12293), .B(n12294), .Z(n12285) );
  AND U11919 ( .A(n1088), .B(n12295), .Z(n12294) );
  XNOR U11920 ( .A(n12296), .B(n12297), .Z(n12291) );
  AND U11921 ( .A(n1080), .B(n12298), .Z(n12297) );
  XOR U11922 ( .A(p_input[1533]), .B(n12296), .Z(n12298) );
  XNOR U11923 ( .A(n12299), .B(n12300), .Z(n12296) );
  AND U11924 ( .A(n1084), .B(n12295), .Z(n12300) );
  XNOR U11925 ( .A(n12299), .B(n12293), .Z(n12295) );
  XOR U11926 ( .A(n12301), .B(n12302), .Z(n12293) );
  AND U11927 ( .A(n1099), .B(n12303), .Z(n12302) );
  XNOR U11928 ( .A(n12304), .B(n12305), .Z(n12299) );
  AND U11929 ( .A(n1091), .B(n12306), .Z(n12305) );
  XOR U11930 ( .A(p_input[1549]), .B(n12304), .Z(n12306) );
  XNOR U11931 ( .A(n12307), .B(n12308), .Z(n12304) );
  AND U11932 ( .A(n1095), .B(n12303), .Z(n12308) );
  XNOR U11933 ( .A(n12307), .B(n12301), .Z(n12303) );
  XOR U11934 ( .A(n12309), .B(n12310), .Z(n12301) );
  AND U11935 ( .A(n1110), .B(n12311), .Z(n12310) );
  XNOR U11936 ( .A(n12312), .B(n12313), .Z(n12307) );
  AND U11937 ( .A(n1102), .B(n12314), .Z(n12313) );
  XOR U11938 ( .A(p_input[1565]), .B(n12312), .Z(n12314) );
  XNOR U11939 ( .A(n12315), .B(n12316), .Z(n12312) );
  AND U11940 ( .A(n1106), .B(n12311), .Z(n12316) );
  XNOR U11941 ( .A(n12315), .B(n12309), .Z(n12311) );
  XOR U11942 ( .A(n12317), .B(n12318), .Z(n12309) );
  AND U11943 ( .A(n1121), .B(n12319), .Z(n12318) );
  XNOR U11944 ( .A(n12320), .B(n12321), .Z(n12315) );
  AND U11945 ( .A(n1113), .B(n12322), .Z(n12321) );
  XOR U11946 ( .A(p_input[1581]), .B(n12320), .Z(n12322) );
  XNOR U11947 ( .A(n12323), .B(n12324), .Z(n12320) );
  AND U11948 ( .A(n1117), .B(n12319), .Z(n12324) );
  XNOR U11949 ( .A(n12323), .B(n12317), .Z(n12319) );
  XOR U11950 ( .A(n12325), .B(n12326), .Z(n12317) );
  AND U11951 ( .A(n1132), .B(n12327), .Z(n12326) );
  XNOR U11952 ( .A(n12328), .B(n12329), .Z(n12323) );
  AND U11953 ( .A(n1124), .B(n12330), .Z(n12329) );
  XOR U11954 ( .A(p_input[1597]), .B(n12328), .Z(n12330) );
  XNOR U11955 ( .A(n12331), .B(n12332), .Z(n12328) );
  AND U11956 ( .A(n1128), .B(n12327), .Z(n12332) );
  XNOR U11957 ( .A(n12331), .B(n12325), .Z(n12327) );
  XOR U11958 ( .A(n12333), .B(n12334), .Z(n12325) );
  AND U11959 ( .A(n1143), .B(n12335), .Z(n12334) );
  XNOR U11960 ( .A(n12336), .B(n12337), .Z(n12331) );
  AND U11961 ( .A(n1135), .B(n12338), .Z(n12337) );
  XOR U11962 ( .A(p_input[1613]), .B(n12336), .Z(n12338) );
  XNOR U11963 ( .A(n12339), .B(n12340), .Z(n12336) );
  AND U11964 ( .A(n1139), .B(n12335), .Z(n12340) );
  XNOR U11965 ( .A(n12339), .B(n12333), .Z(n12335) );
  XOR U11966 ( .A(n12341), .B(n12342), .Z(n12333) );
  AND U11967 ( .A(n1154), .B(n12343), .Z(n12342) );
  XNOR U11968 ( .A(n12344), .B(n12345), .Z(n12339) );
  AND U11969 ( .A(n1146), .B(n12346), .Z(n12345) );
  XOR U11970 ( .A(p_input[1629]), .B(n12344), .Z(n12346) );
  XNOR U11971 ( .A(n12347), .B(n12348), .Z(n12344) );
  AND U11972 ( .A(n1150), .B(n12343), .Z(n12348) );
  XNOR U11973 ( .A(n12347), .B(n12341), .Z(n12343) );
  XOR U11974 ( .A(n12349), .B(n12350), .Z(n12341) );
  AND U11975 ( .A(n1165), .B(n12351), .Z(n12350) );
  XNOR U11976 ( .A(n12352), .B(n12353), .Z(n12347) );
  AND U11977 ( .A(n1157), .B(n12354), .Z(n12353) );
  XOR U11978 ( .A(p_input[1645]), .B(n12352), .Z(n12354) );
  XNOR U11979 ( .A(n12355), .B(n12356), .Z(n12352) );
  AND U11980 ( .A(n1161), .B(n12351), .Z(n12356) );
  XNOR U11981 ( .A(n12355), .B(n12349), .Z(n12351) );
  XOR U11982 ( .A(n12357), .B(n12358), .Z(n12349) );
  AND U11983 ( .A(n1176), .B(n12359), .Z(n12358) );
  XNOR U11984 ( .A(n12360), .B(n12361), .Z(n12355) );
  AND U11985 ( .A(n1168), .B(n12362), .Z(n12361) );
  XOR U11986 ( .A(p_input[1661]), .B(n12360), .Z(n12362) );
  XNOR U11987 ( .A(n12363), .B(n12364), .Z(n12360) );
  AND U11988 ( .A(n1172), .B(n12359), .Z(n12364) );
  XNOR U11989 ( .A(n12363), .B(n12357), .Z(n12359) );
  XOR U11990 ( .A(n12365), .B(n12366), .Z(n12357) );
  AND U11991 ( .A(n1187), .B(n12367), .Z(n12366) );
  XNOR U11992 ( .A(n12368), .B(n12369), .Z(n12363) );
  AND U11993 ( .A(n1179), .B(n12370), .Z(n12369) );
  XOR U11994 ( .A(p_input[1677]), .B(n12368), .Z(n12370) );
  XNOR U11995 ( .A(n12371), .B(n12372), .Z(n12368) );
  AND U11996 ( .A(n1183), .B(n12367), .Z(n12372) );
  XNOR U11997 ( .A(n12371), .B(n12365), .Z(n12367) );
  XOR U11998 ( .A(n12373), .B(n12374), .Z(n12365) );
  AND U11999 ( .A(n1198), .B(n12375), .Z(n12374) );
  XNOR U12000 ( .A(n12376), .B(n12377), .Z(n12371) );
  AND U12001 ( .A(n1190), .B(n12378), .Z(n12377) );
  XOR U12002 ( .A(p_input[1693]), .B(n12376), .Z(n12378) );
  XNOR U12003 ( .A(n12379), .B(n12380), .Z(n12376) );
  AND U12004 ( .A(n1194), .B(n12375), .Z(n12380) );
  XNOR U12005 ( .A(n12379), .B(n12373), .Z(n12375) );
  XOR U12006 ( .A(n12381), .B(n12382), .Z(n12373) );
  AND U12007 ( .A(n1209), .B(n12383), .Z(n12382) );
  XNOR U12008 ( .A(n12384), .B(n12385), .Z(n12379) );
  AND U12009 ( .A(n1201), .B(n12386), .Z(n12385) );
  XOR U12010 ( .A(p_input[1709]), .B(n12384), .Z(n12386) );
  XNOR U12011 ( .A(n12387), .B(n12388), .Z(n12384) );
  AND U12012 ( .A(n1205), .B(n12383), .Z(n12388) );
  XNOR U12013 ( .A(n12387), .B(n12381), .Z(n12383) );
  XOR U12014 ( .A(n12389), .B(n12390), .Z(n12381) );
  AND U12015 ( .A(n1220), .B(n12391), .Z(n12390) );
  XNOR U12016 ( .A(n12392), .B(n12393), .Z(n12387) );
  AND U12017 ( .A(n1212), .B(n12394), .Z(n12393) );
  XOR U12018 ( .A(p_input[1725]), .B(n12392), .Z(n12394) );
  XNOR U12019 ( .A(n12395), .B(n12396), .Z(n12392) );
  AND U12020 ( .A(n1216), .B(n12391), .Z(n12396) );
  XNOR U12021 ( .A(n12395), .B(n12389), .Z(n12391) );
  XOR U12022 ( .A(n12397), .B(n12398), .Z(n12389) );
  AND U12023 ( .A(n1231), .B(n12399), .Z(n12398) );
  XNOR U12024 ( .A(n12400), .B(n12401), .Z(n12395) );
  AND U12025 ( .A(n1223), .B(n12402), .Z(n12401) );
  XOR U12026 ( .A(p_input[1741]), .B(n12400), .Z(n12402) );
  XNOR U12027 ( .A(n12403), .B(n12404), .Z(n12400) );
  AND U12028 ( .A(n1227), .B(n12399), .Z(n12404) );
  XNOR U12029 ( .A(n12403), .B(n12397), .Z(n12399) );
  XOR U12030 ( .A(n12405), .B(n12406), .Z(n12397) );
  AND U12031 ( .A(n1242), .B(n12407), .Z(n12406) );
  XNOR U12032 ( .A(n12408), .B(n12409), .Z(n12403) );
  AND U12033 ( .A(n1234), .B(n12410), .Z(n12409) );
  XOR U12034 ( .A(p_input[1757]), .B(n12408), .Z(n12410) );
  XNOR U12035 ( .A(n12411), .B(n12412), .Z(n12408) );
  AND U12036 ( .A(n1238), .B(n12407), .Z(n12412) );
  XNOR U12037 ( .A(n12411), .B(n12405), .Z(n12407) );
  XOR U12038 ( .A(n12413), .B(n12414), .Z(n12405) );
  AND U12039 ( .A(n1253), .B(n12415), .Z(n12414) );
  XNOR U12040 ( .A(n12416), .B(n12417), .Z(n12411) );
  AND U12041 ( .A(n1245), .B(n12418), .Z(n12417) );
  XOR U12042 ( .A(p_input[1773]), .B(n12416), .Z(n12418) );
  XNOR U12043 ( .A(n12419), .B(n12420), .Z(n12416) );
  AND U12044 ( .A(n1249), .B(n12415), .Z(n12420) );
  XNOR U12045 ( .A(n12419), .B(n12413), .Z(n12415) );
  XOR U12046 ( .A(n12421), .B(n12422), .Z(n12413) );
  AND U12047 ( .A(n1264), .B(n12423), .Z(n12422) );
  XNOR U12048 ( .A(n12424), .B(n12425), .Z(n12419) );
  AND U12049 ( .A(n1256), .B(n12426), .Z(n12425) );
  XOR U12050 ( .A(p_input[1789]), .B(n12424), .Z(n12426) );
  XNOR U12051 ( .A(n12427), .B(n12428), .Z(n12424) );
  AND U12052 ( .A(n1260), .B(n12423), .Z(n12428) );
  XNOR U12053 ( .A(n12427), .B(n12421), .Z(n12423) );
  XOR U12054 ( .A(n12429), .B(n12430), .Z(n12421) );
  AND U12055 ( .A(n1275), .B(n12431), .Z(n12430) );
  XNOR U12056 ( .A(n12432), .B(n12433), .Z(n12427) );
  AND U12057 ( .A(n1267), .B(n12434), .Z(n12433) );
  XOR U12058 ( .A(p_input[1805]), .B(n12432), .Z(n12434) );
  XNOR U12059 ( .A(n12435), .B(n12436), .Z(n12432) );
  AND U12060 ( .A(n1271), .B(n12431), .Z(n12436) );
  XNOR U12061 ( .A(n12435), .B(n12429), .Z(n12431) );
  XOR U12062 ( .A(n12437), .B(n12438), .Z(n12429) );
  AND U12063 ( .A(n1286), .B(n12439), .Z(n12438) );
  XNOR U12064 ( .A(n12440), .B(n12441), .Z(n12435) );
  AND U12065 ( .A(n1278), .B(n12442), .Z(n12441) );
  XOR U12066 ( .A(p_input[1821]), .B(n12440), .Z(n12442) );
  XNOR U12067 ( .A(n12443), .B(n12444), .Z(n12440) );
  AND U12068 ( .A(n1282), .B(n12439), .Z(n12444) );
  XNOR U12069 ( .A(n12443), .B(n12437), .Z(n12439) );
  XOR U12070 ( .A(n12445), .B(n12446), .Z(n12437) );
  AND U12071 ( .A(n1297), .B(n12447), .Z(n12446) );
  XNOR U12072 ( .A(n12448), .B(n12449), .Z(n12443) );
  AND U12073 ( .A(n1289), .B(n12450), .Z(n12449) );
  XOR U12074 ( .A(p_input[1837]), .B(n12448), .Z(n12450) );
  XNOR U12075 ( .A(n12451), .B(n12452), .Z(n12448) );
  AND U12076 ( .A(n1293), .B(n12447), .Z(n12452) );
  XNOR U12077 ( .A(n12451), .B(n12445), .Z(n12447) );
  XOR U12078 ( .A(n12453), .B(n12454), .Z(n12445) );
  AND U12079 ( .A(n1308), .B(n12455), .Z(n12454) );
  XNOR U12080 ( .A(n12456), .B(n12457), .Z(n12451) );
  AND U12081 ( .A(n1300), .B(n12458), .Z(n12457) );
  XOR U12082 ( .A(p_input[1853]), .B(n12456), .Z(n12458) );
  XNOR U12083 ( .A(n12459), .B(n12460), .Z(n12456) );
  AND U12084 ( .A(n1304), .B(n12455), .Z(n12460) );
  XNOR U12085 ( .A(n12459), .B(n12453), .Z(n12455) );
  XOR U12086 ( .A(n12461), .B(n12462), .Z(n12453) );
  AND U12087 ( .A(n1319), .B(n12463), .Z(n12462) );
  XNOR U12088 ( .A(n12464), .B(n12465), .Z(n12459) );
  AND U12089 ( .A(n1311), .B(n12466), .Z(n12465) );
  XOR U12090 ( .A(p_input[1869]), .B(n12464), .Z(n12466) );
  XNOR U12091 ( .A(n12467), .B(n12468), .Z(n12464) );
  AND U12092 ( .A(n1315), .B(n12463), .Z(n12468) );
  XNOR U12093 ( .A(n12467), .B(n12461), .Z(n12463) );
  XOR U12094 ( .A(n12469), .B(n12470), .Z(n12461) );
  AND U12095 ( .A(n1330), .B(n12471), .Z(n12470) );
  XNOR U12096 ( .A(n12472), .B(n12473), .Z(n12467) );
  AND U12097 ( .A(n1322), .B(n12474), .Z(n12473) );
  XOR U12098 ( .A(p_input[1885]), .B(n12472), .Z(n12474) );
  XNOR U12099 ( .A(n12475), .B(n12476), .Z(n12472) );
  AND U12100 ( .A(n1326), .B(n12471), .Z(n12476) );
  XNOR U12101 ( .A(n12475), .B(n12469), .Z(n12471) );
  XOR U12102 ( .A(n12477), .B(n12478), .Z(n12469) );
  AND U12103 ( .A(n1341), .B(n12479), .Z(n12478) );
  XNOR U12104 ( .A(n12480), .B(n12481), .Z(n12475) );
  AND U12105 ( .A(n1333), .B(n12482), .Z(n12481) );
  XOR U12106 ( .A(p_input[1901]), .B(n12480), .Z(n12482) );
  XNOR U12107 ( .A(n12483), .B(n12484), .Z(n12480) );
  AND U12108 ( .A(n1337), .B(n12479), .Z(n12484) );
  XNOR U12109 ( .A(n12483), .B(n12477), .Z(n12479) );
  XOR U12110 ( .A(n12485), .B(n12486), .Z(n12477) );
  AND U12111 ( .A(n1352), .B(n12487), .Z(n12486) );
  XNOR U12112 ( .A(n12488), .B(n12489), .Z(n12483) );
  AND U12113 ( .A(n1344), .B(n12490), .Z(n12489) );
  XOR U12114 ( .A(p_input[1917]), .B(n12488), .Z(n12490) );
  XNOR U12115 ( .A(n12491), .B(n12492), .Z(n12488) );
  AND U12116 ( .A(n1348), .B(n12487), .Z(n12492) );
  XNOR U12117 ( .A(n12491), .B(n12485), .Z(n12487) );
  XOR U12118 ( .A(n12493), .B(n12494), .Z(n12485) );
  AND U12119 ( .A(n1363), .B(n12495), .Z(n12494) );
  XNOR U12120 ( .A(n12496), .B(n12497), .Z(n12491) );
  AND U12121 ( .A(n1355), .B(n12498), .Z(n12497) );
  XOR U12122 ( .A(p_input[1933]), .B(n12496), .Z(n12498) );
  XNOR U12123 ( .A(n12499), .B(n12500), .Z(n12496) );
  AND U12124 ( .A(n1359), .B(n12495), .Z(n12500) );
  XNOR U12125 ( .A(n12499), .B(n12493), .Z(n12495) );
  XOR U12126 ( .A(n12501), .B(n12502), .Z(n12493) );
  AND U12127 ( .A(n1374), .B(n12503), .Z(n12502) );
  XNOR U12128 ( .A(n12504), .B(n12505), .Z(n12499) );
  AND U12129 ( .A(n1366), .B(n12506), .Z(n12505) );
  XOR U12130 ( .A(p_input[1949]), .B(n12504), .Z(n12506) );
  XNOR U12131 ( .A(n12507), .B(n12508), .Z(n12504) );
  AND U12132 ( .A(n1370), .B(n12503), .Z(n12508) );
  XNOR U12133 ( .A(n12507), .B(n12501), .Z(n12503) );
  XOR U12134 ( .A(n12509), .B(n12510), .Z(n12501) );
  AND U12135 ( .A(n1385), .B(n12511), .Z(n12510) );
  XNOR U12136 ( .A(n12512), .B(n12513), .Z(n12507) );
  AND U12137 ( .A(n1377), .B(n12514), .Z(n12513) );
  XOR U12138 ( .A(p_input[1965]), .B(n12512), .Z(n12514) );
  XNOR U12139 ( .A(n12515), .B(n12516), .Z(n12512) );
  AND U12140 ( .A(n1381), .B(n12511), .Z(n12516) );
  XNOR U12141 ( .A(n12515), .B(n12509), .Z(n12511) );
  XOR U12142 ( .A(n12517), .B(n12518), .Z(n12509) );
  AND U12143 ( .A(n1396), .B(n12519), .Z(n12518) );
  XNOR U12144 ( .A(n12520), .B(n12521), .Z(n12515) );
  AND U12145 ( .A(n1388), .B(n12522), .Z(n12521) );
  XOR U12146 ( .A(p_input[1981]), .B(n12520), .Z(n12522) );
  XNOR U12147 ( .A(n12523), .B(n12524), .Z(n12520) );
  AND U12148 ( .A(n1392), .B(n12519), .Z(n12524) );
  XNOR U12149 ( .A(n12523), .B(n12517), .Z(n12519) );
  XOR U12150 ( .A(n12525), .B(n12526), .Z(n12517) );
  AND U12151 ( .A(n1407), .B(n12527), .Z(n12526) );
  XNOR U12152 ( .A(n12528), .B(n12529), .Z(n12523) );
  AND U12153 ( .A(n1399), .B(n12530), .Z(n12529) );
  XOR U12154 ( .A(p_input[1997]), .B(n12528), .Z(n12530) );
  XNOR U12155 ( .A(n12531), .B(n12532), .Z(n12528) );
  AND U12156 ( .A(n1403), .B(n12527), .Z(n12532) );
  XNOR U12157 ( .A(n12531), .B(n12525), .Z(n12527) );
  XOR U12158 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n12533), .Z(n12525) );
  AND U12159 ( .A(n1417), .B(n12534), .Z(n12533) );
  XNOR U12160 ( .A(n12535), .B(n12536), .Z(n12531) );
  AND U12161 ( .A(n1410), .B(n12537), .Z(n12536) );
  XOR U12162 ( .A(p_input[2013]), .B(n12535), .Z(n12537) );
  XNOR U12163 ( .A(n12538), .B(n12539), .Z(n12535) );
  AND U12164 ( .A(n1414), .B(n12534), .Z(n12539) );
  XOR U12165 ( .A(\knn_comb_/min_val_out[0][13] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n12534) );
  XOR U12166 ( .A(n23), .B(n12540), .Z(o[12]) );
  AND U12167 ( .A(n30), .B(n12541), .Z(n23) );
  XOR U12168 ( .A(n24), .B(n12540), .Z(n12541) );
  XOR U12169 ( .A(n12542), .B(n12543), .Z(n12540) );
  AND U12170 ( .A(n42), .B(n12544), .Z(n12543) );
  XOR U12171 ( .A(n12545), .B(n12546), .Z(n24) );
  AND U12172 ( .A(n34), .B(n12547), .Z(n12546) );
  XOR U12173 ( .A(p_input[12]), .B(n12545), .Z(n12547) );
  XNOR U12174 ( .A(n12548), .B(n12549), .Z(n12545) );
  AND U12175 ( .A(n38), .B(n12544), .Z(n12549) );
  XNOR U12176 ( .A(n12548), .B(n12542), .Z(n12544) );
  XOR U12177 ( .A(n12550), .B(n12551), .Z(n12542) );
  AND U12178 ( .A(n54), .B(n12552), .Z(n12551) );
  XNOR U12179 ( .A(n12553), .B(n12554), .Z(n12548) );
  AND U12180 ( .A(n46), .B(n12555), .Z(n12554) );
  XOR U12181 ( .A(p_input[28]), .B(n12553), .Z(n12555) );
  XNOR U12182 ( .A(n12556), .B(n12557), .Z(n12553) );
  AND U12183 ( .A(n50), .B(n12552), .Z(n12557) );
  XNOR U12184 ( .A(n12556), .B(n12550), .Z(n12552) );
  XOR U12185 ( .A(n12558), .B(n12559), .Z(n12550) );
  AND U12186 ( .A(n65), .B(n12560), .Z(n12559) );
  XNOR U12187 ( .A(n12561), .B(n12562), .Z(n12556) );
  AND U12188 ( .A(n57), .B(n12563), .Z(n12562) );
  XOR U12189 ( .A(p_input[44]), .B(n12561), .Z(n12563) );
  XNOR U12190 ( .A(n12564), .B(n12565), .Z(n12561) );
  AND U12191 ( .A(n61), .B(n12560), .Z(n12565) );
  XNOR U12192 ( .A(n12564), .B(n12558), .Z(n12560) );
  XOR U12193 ( .A(n12566), .B(n12567), .Z(n12558) );
  AND U12194 ( .A(n76), .B(n12568), .Z(n12567) );
  XNOR U12195 ( .A(n12569), .B(n12570), .Z(n12564) );
  AND U12196 ( .A(n68), .B(n12571), .Z(n12570) );
  XOR U12197 ( .A(p_input[60]), .B(n12569), .Z(n12571) );
  XNOR U12198 ( .A(n12572), .B(n12573), .Z(n12569) );
  AND U12199 ( .A(n72), .B(n12568), .Z(n12573) );
  XNOR U12200 ( .A(n12572), .B(n12566), .Z(n12568) );
  XOR U12201 ( .A(n12574), .B(n12575), .Z(n12566) );
  AND U12202 ( .A(n87), .B(n12576), .Z(n12575) );
  XNOR U12203 ( .A(n12577), .B(n12578), .Z(n12572) );
  AND U12204 ( .A(n79), .B(n12579), .Z(n12578) );
  XOR U12205 ( .A(p_input[76]), .B(n12577), .Z(n12579) );
  XNOR U12206 ( .A(n12580), .B(n12581), .Z(n12577) );
  AND U12207 ( .A(n83), .B(n12576), .Z(n12581) );
  XNOR U12208 ( .A(n12580), .B(n12574), .Z(n12576) );
  XOR U12209 ( .A(n12582), .B(n12583), .Z(n12574) );
  AND U12210 ( .A(n98), .B(n12584), .Z(n12583) );
  XNOR U12211 ( .A(n12585), .B(n12586), .Z(n12580) );
  AND U12212 ( .A(n90), .B(n12587), .Z(n12586) );
  XOR U12213 ( .A(p_input[92]), .B(n12585), .Z(n12587) );
  XNOR U12214 ( .A(n12588), .B(n12589), .Z(n12585) );
  AND U12215 ( .A(n94), .B(n12584), .Z(n12589) );
  XNOR U12216 ( .A(n12588), .B(n12582), .Z(n12584) );
  XOR U12217 ( .A(n12590), .B(n12591), .Z(n12582) );
  AND U12218 ( .A(n109), .B(n12592), .Z(n12591) );
  XNOR U12219 ( .A(n12593), .B(n12594), .Z(n12588) );
  AND U12220 ( .A(n101), .B(n12595), .Z(n12594) );
  XOR U12221 ( .A(p_input[108]), .B(n12593), .Z(n12595) );
  XNOR U12222 ( .A(n12596), .B(n12597), .Z(n12593) );
  AND U12223 ( .A(n105), .B(n12592), .Z(n12597) );
  XNOR U12224 ( .A(n12596), .B(n12590), .Z(n12592) );
  XOR U12225 ( .A(n12598), .B(n12599), .Z(n12590) );
  AND U12226 ( .A(n120), .B(n12600), .Z(n12599) );
  XNOR U12227 ( .A(n12601), .B(n12602), .Z(n12596) );
  AND U12228 ( .A(n112), .B(n12603), .Z(n12602) );
  XOR U12229 ( .A(p_input[124]), .B(n12601), .Z(n12603) );
  XNOR U12230 ( .A(n12604), .B(n12605), .Z(n12601) );
  AND U12231 ( .A(n116), .B(n12600), .Z(n12605) );
  XNOR U12232 ( .A(n12604), .B(n12598), .Z(n12600) );
  XOR U12233 ( .A(n12606), .B(n12607), .Z(n12598) );
  AND U12234 ( .A(n131), .B(n12608), .Z(n12607) );
  XNOR U12235 ( .A(n12609), .B(n12610), .Z(n12604) );
  AND U12236 ( .A(n123), .B(n12611), .Z(n12610) );
  XOR U12237 ( .A(p_input[140]), .B(n12609), .Z(n12611) );
  XNOR U12238 ( .A(n12612), .B(n12613), .Z(n12609) );
  AND U12239 ( .A(n127), .B(n12608), .Z(n12613) );
  XNOR U12240 ( .A(n12612), .B(n12606), .Z(n12608) );
  XOR U12241 ( .A(n12614), .B(n12615), .Z(n12606) );
  AND U12242 ( .A(n142), .B(n12616), .Z(n12615) );
  XNOR U12243 ( .A(n12617), .B(n12618), .Z(n12612) );
  AND U12244 ( .A(n134), .B(n12619), .Z(n12618) );
  XOR U12245 ( .A(p_input[156]), .B(n12617), .Z(n12619) );
  XNOR U12246 ( .A(n12620), .B(n12621), .Z(n12617) );
  AND U12247 ( .A(n138), .B(n12616), .Z(n12621) );
  XNOR U12248 ( .A(n12620), .B(n12614), .Z(n12616) );
  XOR U12249 ( .A(n12622), .B(n12623), .Z(n12614) );
  AND U12250 ( .A(n153), .B(n12624), .Z(n12623) );
  XNOR U12251 ( .A(n12625), .B(n12626), .Z(n12620) );
  AND U12252 ( .A(n145), .B(n12627), .Z(n12626) );
  XOR U12253 ( .A(p_input[172]), .B(n12625), .Z(n12627) );
  XNOR U12254 ( .A(n12628), .B(n12629), .Z(n12625) );
  AND U12255 ( .A(n149), .B(n12624), .Z(n12629) );
  XNOR U12256 ( .A(n12628), .B(n12622), .Z(n12624) );
  XOR U12257 ( .A(n12630), .B(n12631), .Z(n12622) );
  AND U12258 ( .A(n164), .B(n12632), .Z(n12631) );
  XNOR U12259 ( .A(n12633), .B(n12634), .Z(n12628) );
  AND U12260 ( .A(n156), .B(n12635), .Z(n12634) );
  XOR U12261 ( .A(p_input[188]), .B(n12633), .Z(n12635) );
  XNOR U12262 ( .A(n12636), .B(n12637), .Z(n12633) );
  AND U12263 ( .A(n160), .B(n12632), .Z(n12637) );
  XNOR U12264 ( .A(n12636), .B(n12630), .Z(n12632) );
  XOR U12265 ( .A(n12638), .B(n12639), .Z(n12630) );
  AND U12266 ( .A(n175), .B(n12640), .Z(n12639) );
  XNOR U12267 ( .A(n12641), .B(n12642), .Z(n12636) );
  AND U12268 ( .A(n167), .B(n12643), .Z(n12642) );
  XOR U12269 ( .A(p_input[204]), .B(n12641), .Z(n12643) );
  XNOR U12270 ( .A(n12644), .B(n12645), .Z(n12641) );
  AND U12271 ( .A(n171), .B(n12640), .Z(n12645) );
  XNOR U12272 ( .A(n12644), .B(n12638), .Z(n12640) );
  XOR U12273 ( .A(n12646), .B(n12647), .Z(n12638) );
  AND U12274 ( .A(n186), .B(n12648), .Z(n12647) );
  XNOR U12275 ( .A(n12649), .B(n12650), .Z(n12644) );
  AND U12276 ( .A(n178), .B(n12651), .Z(n12650) );
  XOR U12277 ( .A(p_input[220]), .B(n12649), .Z(n12651) );
  XNOR U12278 ( .A(n12652), .B(n12653), .Z(n12649) );
  AND U12279 ( .A(n182), .B(n12648), .Z(n12653) );
  XNOR U12280 ( .A(n12652), .B(n12646), .Z(n12648) );
  XOR U12281 ( .A(n12654), .B(n12655), .Z(n12646) );
  AND U12282 ( .A(n197), .B(n12656), .Z(n12655) );
  XNOR U12283 ( .A(n12657), .B(n12658), .Z(n12652) );
  AND U12284 ( .A(n189), .B(n12659), .Z(n12658) );
  XOR U12285 ( .A(p_input[236]), .B(n12657), .Z(n12659) );
  XNOR U12286 ( .A(n12660), .B(n12661), .Z(n12657) );
  AND U12287 ( .A(n193), .B(n12656), .Z(n12661) );
  XNOR U12288 ( .A(n12660), .B(n12654), .Z(n12656) );
  XOR U12289 ( .A(n12662), .B(n12663), .Z(n12654) );
  AND U12290 ( .A(n208), .B(n12664), .Z(n12663) );
  XNOR U12291 ( .A(n12665), .B(n12666), .Z(n12660) );
  AND U12292 ( .A(n200), .B(n12667), .Z(n12666) );
  XOR U12293 ( .A(p_input[252]), .B(n12665), .Z(n12667) );
  XNOR U12294 ( .A(n12668), .B(n12669), .Z(n12665) );
  AND U12295 ( .A(n204), .B(n12664), .Z(n12669) );
  XNOR U12296 ( .A(n12668), .B(n12662), .Z(n12664) );
  XOR U12297 ( .A(n12670), .B(n12671), .Z(n12662) );
  AND U12298 ( .A(n219), .B(n12672), .Z(n12671) );
  XNOR U12299 ( .A(n12673), .B(n12674), .Z(n12668) );
  AND U12300 ( .A(n211), .B(n12675), .Z(n12674) );
  XOR U12301 ( .A(p_input[268]), .B(n12673), .Z(n12675) );
  XNOR U12302 ( .A(n12676), .B(n12677), .Z(n12673) );
  AND U12303 ( .A(n215), .B(n12672), .Z(n12677) );
  XNOR U12304 ( .A(n12676), .B(n12670), .Z(n12672) );
  XOR U12305 ( .A(n12678), .B(n12679), .Z(n12670) );
  AND U12306 ( .A(n230), .B(n12680), .Z(n12679) );
  XNOR U12307 ( .A(n12681), .B(n12682), .Z(n12676) );
  AND U12308 ( .A(n222), .B(n12683), .Z(n12682) );
  XOR U12309 ( .A(p_input[284]), .B(n12681), .Z(n12683) );
  XNOR U12310 ( .A(n12684), .B(n12685), .Z(n12681) );
  AND U12311 ( .A(n226), .B(n12680), .Z(n12685) );
  XNOR U12312 ( .A(n12684), .B(n12678), .Z(n12680) );
  XOR U12313 ( .A(n12686), .B(n12687), .Z(n12678) );
  AND U12314 ( .A(n241), .B(n12688), .Z(n12687) );
  XNOR U12315 ( .A(n12689), .B(n12690), .Z(n12684) );
  AND U12316 ( .A(n233), .B(n12691), .Z(n12690) );
  XOR U12317 ( .A(p_input[300]), .B(n12689), .Z(n12691) );
  XNOR U12318 ( .A(n12692), .B(n12693), .Z(n12689) );
  AND U12319 ( .A(n237), .B(n12688), .Z(n12693) );
  XNOR U12320 ( .A(n12692), .B(n12686), .Z(n12688) );
  XOR U12321 ( .A(n12694), .B(n12695), .Z(n12686) );
  AND U12322 ( .A(n252), .B(n12696), .Z(n12695) );
  XNOR U12323 ( .A(n12697), .B(n12698), .Z(n12692) );
  AND U12324 ( .A(n244), .B(n12699), .Z(n12698) );
  XOR U12325 ( .A(p_input[316]), .B(n12697), .Z(n12699) );
  XNOR U12326 ( .A(n12700), .B(n12701), .Z(n12697) );
  AND U12327 ( .A(n248), .B(n12696), .Z(n12701) );
  XNOR U12328 ( .A(n12700), .B(n12694), .Z(n12696) );
  XOR U12329 ( .A(n12702), .B(n12703), .Z(n12694) );
  AND U12330 ( .A(n263), .B(n12704), .Z(n12703) );
  XNOR U12331 ( .A(n12705), .B(n12706), .Z(n12700) );
  AND U12332 ( .A(n255), .B(n12707), .Z(n12706) );
  XOR U12333 ( .A(p_input[332]), .B(n12705), .Z(n12707) );
  XNOR U12334 ( .A(n12708), .B(n12709), .Z(n12705) );
  AND U12335 ( .A(n259), .B(n12704), .Z(n12709) );
  XNOR U12336 ( .A(n12708), .B(n12702), .Z(n12704) );
  XOR U12337 ( .A(n12710), .B(n12711), .Z(n12702) );
  AND U12338 ( .A(n274), .B(n12712), .Z(n12711) );
  XNOR U12339 ( .A(n12713), .B(n12714), .Z(n12708) );
  AND U12340 ( .A(n266), .B(n12715), .Z(n12714) );
  XOR U12341 ( .A(p_input[348]), .B(n12713), .Z(n12715) );
  XNOR U12342 ( .A(n12716), .B(n12717), .Z(n12713) );
  AND U12343 ( .A(n270), .B(n12712), .Z(n12717) );
  XNOR U12344 ( .A(n12716), .B(n12710), .Z(n12712) );
  XOR U12345 ( .A(n12718), .B(n12719), .Z(n12710) );
  AND U12346 ( .A(n285), .B(n12720), .Z(n12719) );
  XNOR U12347 ( .A(n12721), .B(n12722), .Z(n12716) );
  AND U12348 ( .A(n277), .B(n12723), .Z(n12722) );
  XOR U12349 ( .A(p_input[364]), .B(n12721), .Z(n12723) );
  XNOR U12350 ( .A(n12724), .B(n12725), .Z(n12721) );
  AND U12351 ( .A(n281), .B(n12720), .Z(n12725) );
  XNOR U12352 ( .A(n12724), .B(n12718), .Z(n12720) );
  XOR U12353 ( .A(n12726), .B(n12727), .Z(n12718) );
  AND U12354 ( .A(n296), .B(n12728), .Z(n12727) );
  XNOR U12355 ( .A(n12729), .B(n12730), .Z(n12724) );
  AND U12356 ( .A(n288), .B(n12731), .Z(n12730) );
  XOR U12357 ( .A(p_input[380]), .B(n12729), .Z(n12731) );
  XNOR U12358 ( .A(n12732), .B(n12733), .Z(n12729) );
  AND U12359 ( .A(n292), .B(n12728), .Z(n12733) );
  XNOR U12360 ( .A(n12732), .B(n12726), .Z(n12728) );
  XOR U12361 ( .A(n12734), .B(n12735), .Z(n12726) );
  AND U12362 ( .A(n307), .B(n12736), .Z(n12735) );
  XNOR U12363 ( .A(n12737), .B(n12738), .Z(n12732) );
  AND U12364 ( .A(n299), .B(n12739), .Z(n12738) );
  XOR U12365 ( .A(p_input[396]), .B(n12737), .Z(n12739) );
  XNOR U12366 ( .A(n12740), .B(n12741), .Z(n12737) );
  AND U12367 ( .A(n303), .B(n12736), .Z(n12741) );
  XNOR U12368 ( .A(n12740), .B(n12734), .Z(n12736) );
  XOR U12369 ( .A(n12742), .B(n12743), .Z(n12734) );
  AND U12370 ( .A(n318), .B(n12744), .Z(n12743) );
  XNOR U12371 ( .A(n12745), .B(n12746), .Z(n12740) );
  AND U12372 ( .A(n310), .B(n12747), .Z(n12746) );
  XOR U12373 ( .A(p_input[412]), .B(n12745), .Z(n12747) );
  XNOR U12374 ( .A(n12748), .B(n12749), .Z(n12745) );
  AND U12375 ( .A(n314), .B(n12744), .Z(n12749) );
  XNOR U12376 ( .A(n12748), .B(n12742), .Z(n12744) );
  XOR U12377 ( .A(n12750), .B(n12751), .Z(n12742) );
  AND U12378 ( .A(n329), .B(n12752), .Z(n12751) );
  XNOR U12379 ( .A(n12753), .B(n12754), .Z(n12748) );
  AND U12380 ( .A(n321), .B(n12755), .Z(n12754) );
  XOR U12381 ( .A(p_input[428]), .B(n12753), .Z(n12755) );
  XNOR U12382 ( .A(n12756), .B(n12757), .Z(n12753) );
  AND U12383 ( .A(n325), .B(n12752), .Z(n12757) );
  XNOR U12384 ( .A(n12756), .B(n12750), .Z(n12752) );
  XOR U12385 ( .A(n12758), .B(n12759), .Z(n12750) );
  AND U12386 ( .A(n340), .B(n12760), .Z(n12759) );
  XNOR U12387 ( .A(n12761), .B(n12762), .Z(n12756) );
  AND U12388 ( .A(n332), .B(n12763), .Z(n12762) );
  XOR U12389 ( .A(p_input[444]), .B(n12761), .Z(n12763) );
  XNOR U12390 ( .A(n12764), .B(n12765), .Z(n12761) );
  AND U12391 ( .A(n336), .B(n12760), .Z(n12765) );
  XNOR U12392 ( .A(n12764), .B(n12758), .Z(n12760) );
  XOR U12393 ( .A(n12766), .B(n12767), .Z(n12758) );
  AND U12394 ( .A(n351), .B(n12768), .Z(n12767) );
  XNOR U12395 ( .A(n12769), .B(n12770), .Z(n12764) );
  AND U12396 ( .A(n343), .B(n12771), .Z(n12770) );
  XOR U12397 ( .A(p_input[460]), .B(n12769), .Z(n12771) );
  XNOR U12398 ( .A(n12772), .B(n12773), .Z(n12769) );
  AND U12399 ( .A(n347), .B(n12768), .Z(n12773) );
  XNOR U12400 ( .A(n12772), .B(n12766), .Z(n12768) );
  XOR U12401 ( .A(n12774), .B(n12775), .Z(n12766) );
  AND U12402 ( .A(n362), .B(n12776), .Z(n12775) );
  XNOR U12403 ( .A(n12777), .B(n12778), .Z(n12772) );
  AND U12404 ( .A(n354), .B(n12779), .Z(n12778) );
  XOR U12405 ( .A(p_input[476]), .B(n12777), .Z(n12779) );
  XNOR U12406 ( .A(n12780), .B(n12781), .Z(n12777) );
  AND U12407 ( .A(n358), .B(n12776), .Z(n12781) );
  XNOR U12408 ( .A(n12780), .B(n12774), .Z(n12776) );
  XOR U12409 ( .A(n12782), .B(n12783), .Z(n12774) );
  AND U12410 ( .A(n373), .B(n12784), .Z(n12783) );
  XNOR U12411 ( .A(n12785), .B(n12786), .Z(n12780) );
  AND U12412 ( .A(n365), .B(n12787), .Z(n12786) );
  XOR U12413 ( .A(p_input[492]), .B(n12785), .Z(n12787) );
  XNOR U12414 ( .A(n12788), .B(n12789), .Z(n12785) );
  AND U12415 ( .A(n369), .B(n12784), .Z(n12789) );
  XNOR U12416 ( .A(n12788), .B(n12782), .Z(n12784) );
  XOR U12417 ( .A(n12790), .B(n12791), .Z(n12782) );
  AND U12418 ( .A(n384), .B(n12792), .Z(n12791) );
  XNOR U12419 ( .A(n12793), .B(n12794), .Z(n12788) );
  AND U12420 ( .A(n376), .B(n12795), .Z(n12794) );
  XOR U12421 ( .A(p_input[508]), .B(n12793), .Z(n12795) );
  XNOR U12422 ( .A(n12796), .B(n12797), .Z(n12793) );
  AND U12423 ( .A(n380), .B(n12792), .Z(n12797) );
  XNOR U12424 ( .A(n12796), .B(n12790), .Z(n12792) );
  XOR U12425 ( .A(n12798), .B(n12799), .Z(n12790) );
  AND U12426 ( .A(n395), .B(n12800), .Z(n12799) );
  XNOR U12427 ( .A(n12801), .B(n12802), .Z(n12796) );
  AND U12428 ( .A(n387), .B(n12803), .Z(n12802) );
  XOR U12429 ( .A(p_input[524]), .B(n12801), .Z(n12803) );
  XNOR U12430 ( .A(n12804), .B(n12805), .Z(n12801) );
  AND U12431 ( .A(n391), .B(n12800), .Z(n12805) );
  XNOR U12432 ( .A(n12804), .B(n12798), .Z(n12800) );
  XOR U12433 ( .A(n12806), .B(n12807), .Z(n12798) );
  AND U12434 ( .A(n406), .B(n12808), .Z(n12807) );
  XNOR U12435 ( .A(n12809), .B(n12810), .Z(n12804) );
  AND U12436 ( .A(n398), .B(n12811), .Z(n12810) );
  XOR U12437 ( .A(p_input[540]), .B(n12809), .Z(n12811) );
  XNOR U12438 ( .A(n12812), .B(n12813), .Z(n12809) );
  AND U12439 ( .A(n402), .B(n12808), .Z(n12813) );
  XNOR U12440 ( .A(n12812), .B(n12806), .Z(n12808) );
  XOR U12441 ( .A(n12814), .B(n12815), .Z(n12806) );
  AND U12442 ( .A(n417), .B(n12816), .Z(n12815) );
  XNOR U12443 ( .A(n12817), .B(n12818), .Z(n12812) );
  AND U12444 ( .A(n409), .B(n12819), .Z(n12818) );
  XOR U12445 ( .A(p_input[556]), .B(n12817), .Z(n12819) );
  XNOR U12446 ( .A(n12820), .B(n12821), .Z(n12817) );
  AND U12447 ( .A(n413), .B(n12816), .Z(n12821) );
  XNOR U12448 ( .A(n12820), .B(n12814), .Z(n12816) );
  XOR U12449 ( .A(n12822), .B(n12823), .Z(n12814) );
  AND U12450 ( .A(n428), .B(n12824), .Z(n12823) );
  XNOR U12451 ( .A(n12825), .B(n12826), .Z(n12820) );
  AND U12452 ( .A(n420), .B(n12827), .Z(n12826) );
  XOR U12453 ( .A(p_input[572]), .B(n12825), .Z(n12827) );
  XNOR U12454 ( .A(n12828), .B(n12829), .Z(n12825) );
  AND U12455 ( .A(n424), .B(n12824), .Z(n12829) );
  XNOR U12456 ( .A(n12828), .B(n12822), .Z(n12824) );
  XOR U12457 ( .A(n12830), .B(n12831), .Z(n12822) );
  AND U12458 ( .A(n439), .B(n12832), .Z(n12831) );
  XNOR U12459 ( .A(n12833), .B(n12834), .Z(n12828) );
  AND U12460 ( .A(n431), .B(n12835), .Z(n12834) );
  XOR U12461 ( .A(p_input[588]), .B(n12833), .Z(n12835) );
  XNOR U12462 ( .A(n12836), .B(n12837), .Z(n12833) );
  AND U12463 ( .A(n435), .B(n12832), .Z(n12837) );
  XNOR U12464 ( .A(n12836), .B(n12830), .Z(n12832) );
  XOR U12465 ( .A(n12838), .B(n12839), .Z(n12830) );
  AND U12466 ( .A(n450), .B(n12840), .Z(n12839) );
  XNOR U12467 ( .A(n12841), .B(n12842), .Z(n12836) );
  AND U12468 ( .A(n442), .B(n12843), .Z(n12842) );
  XOR U12469 ( .A(p_input[604]), .B(n12841), .Z(n12843) );
  XNOR U12470 ( .A(n12844), .B(n12845), .Z(n12841) );
  AND U12471 ( .A(n446), .B(n12840), .Z(n12845) );
  XNOR U12472 ( .A(n12844), .B(n12838), .Z(n12840) );
  XOR U12473 ( .A(n12846), .B(n12847), .Z(n12838) );
  AND U12474 ( .A(n461), .B(n12848), .Z(n12847) );
  XNOR U12475 ( .A(n12849), .B(n12850), .Z(n12844) );
  AND U12476 ( .A(n453), .B(n12851), .Z(n12850) );
  XOR U12477 ( .A(p_input[620]), .B(n12849), .Z(n12851) );
  XNOR U12478 ( .A(n12852), .B(n12853), .Z(n12849) );
  AND U12479 ( .A(n457), .B(n12848), .Z(n12853) );
  XNOR U12480 ( .A(n12852), .B(n12846), .Z(n12848) );
  XOR U12481 ( .A(n12854), .B(n12855), .Z(n12846) );
  AND U12482 ( .A(n472), .B(n12856), .Z(n12855) );
  XNOR U12483 ( .A(n12857), .B(n12858), .Z(n12852) );
  AND U12484 ( .A(n464), .B(n12859), .Z(n12858) );
  XOR U12485 ( .A(p_input[636]), .B(n12857), .Z(n12859) );
  XNOR U12486 ( .A(n12860), .B(n12861), .Z(n12857) );
  AND U12487 ( .A(n468), .B(n12856), .Z(n12861) );
  XNOR U12488 ( .A(n12860), .B(n12854), .Z(n12856) );
  XOR U12489 ( .A(n12862), .B(n12863), .Z(n12854) );
  AND U12490 ( .A(n483), .B(n12864), .Z(n12863) );
  XNOR U12491 ( .A(n12865), .B(n12866), .Z(n12860) );
  AND U12492 ( .A(n475), .B(n12867), .Z(n12866) );
  XOR U12493 ( .A(p_input[652]), .B(n12865), .Z(n12867) );
  XNOR U12494 ( .A(n12868), .B(n12869), .Z(n12865) );
  AND U12495 ( .A(n479), .B(n12864), .Z(n12869) );
  XNOR U12496 ( .A(n12868), .B(n12862), .Z(n12864) );
  XOR U12497 ( .A(n12870), .B(n12871), .Z(n12862) );
  AND U12498 ( .A(n494), .B(n12872), .Z(n12871) );
  XNOR U12499 ( .A(n12873), .B(n12874), .Z(n12868) );
  AND U12500 ( .A(n486), .B(n12875), .Z(n12874) );
  XOR U12501 ( .A(p_input[668]), .B(n12873), .Z(n12875) );
  XNOR U12502 ( .A(n12876), .B(n12877), .Z(n12873) );
  AND U12503 ( .A(n490), .B(n12872), .Z(n12877) );
  XNOR U12504 ( .A(n12876), .B(n12870), .Z(n12872) );
  XOR U12505 ( .A(n12878), .B(n12879), .Z(n12870) );
  AND U12506 ( .A(n505), .B(n12880), .Z(n12879) );
  XNOR U12507 ( .A(n12881), .B(n12882), .Z(n12876) );
  AND U12508 ( .A(n497), .B(n12883), .Z(n12882) );
  XOR U12509 ( .A(p_input[684]), .B(n12881), .Z(n12883) );
  XNOR U12510 ( .A(n12884), .B(n12885), .Z(n12881) );
  AND U12511 ( .A(n501), .B(n12880), .Z(n12885) );
  XNOR U12512 ( .A(n12884), .B(n12878), .Z(n12880) );
  XOR U12513 ( .A(n12886), .B(n12887), .Z(n12878) );
  AND U12514 ( .A(n516), .B(n12888), .Z(n12887) );
  XNOR U12515 ( .A(n12889), .B(n12890), .Z(n12884) );
  AND U12516 ( .A(n508), .B(n12891), .Z(n12890) );
  XOR U12517 ( .A(p_input[700]), .B(n12889), .Z(n12891) );
  XNOR U12518 ( .A(n12892), .B(n12893), .Z(n12889) );
  AND U12519 ( .A(n512), .B(n12888), .Z(n12893) );
  XNOR U12520 ( .A(n12892), .B(n12886), .Z(n12888) );
  XOR U12521 ( .A(n12894), .B(n12895), .Z(n12886) );
  AND U12522 ( .A(n527), .B(n12896), .Z(n12895) );
  XNOR U12523 ( .A(n12897), .B(n12898), .Z(n12892) );
  AND U12524 ( .A(n519), .B(n12899), .Z(n12898) );
  XOR U12525 ( .A(p_input[716]), .B(n12897), .Z(n12899) );
  XNOR U12526 ( .A(n12900), .B(n12901), .Z(n12897) );
  AND U12527 ( .A(n523), .B(n12896), .Z(n12901) );
  XNOR U12528 ( .A(n12900), .B(n12894), .Z(n12896) );
  XOR U12529 ( .A(n12902), .B(n12903), .Z(n12894) );
  AND U12530 ( .A(n538), .B(n12904), .Z(n12903) );
  XNOR U12531 ( .A(n12905), .B(n12906), .Z(n12900) );
  AND U12532 ( .A(n530), .B(n12907), .Z(n12906) );
  XOR U12533 ( .A(p_input[732]), .B(n12905), .Z(n12907) );
  XNOR U12534 ( .A(n12908), .B(n12909), .Z(n12905) );
  AND U12535 ( .A(n534), .B(n12904), .Z(n12909) );
  XNOR U12536 ( .A(n12908), .B(n12902), .Z(n12904) );
  XOR U12537 ( .A(n12910), .B(n12911), .Z(n12902) );
  AND U12538 ( .A(n549), .B(n12912), .Z(n12911) );
  XNOR U12539 ( .A(n12913), .B(n12914), .Z(n12908) );
  AND U12540 ( .A(n541), .B(n12915), .Z(n12914) );
  XOR U12541 ( .A(p_input[748]), .B(n12913), .Z(n12915) );
  XNOR U12542 ( .A(n12916), .B(n12917), .Z(n12913) );
  AND U12543 ( .A(n545), .B(n12912), .Z(n12917) );
  XNOR U12544 ( .A(n12916), .B(n12910), .Z(n12912) );
  XOR U12545 ( .A(n12918), .B(n12919), .Z(n12910) );
  AND U12546 ( .A(n560), .B(n12920), .Z(n12919) );
  XNOR U12547 ( .A(n12921), .B(n12922), .Z(n12916) );
  AND U12548 ( .A(n552), .B(n12923), .Z(n12922) );
  XOR U12549 ( .A(p_input[764]), .B(n12921), .Z(n12923) );
  XNOR U12550 ( .A(n12924), .B(n12925), .Z(n12921) );
  AND U12551 ( .A(n556), .B(n12920), .Z(n12925) );
  XNOR U12552 ( .A(n12924), .B(n12918), .Z(n12920) );
  XOR U12553 ( .A(n12926), .B(n12927), .Z(n12918) );
  AND U12554 ( .A(n571), .B(n12928), .Z(n12927) );
  XNOR U12555 ( .A(n12929), .B(n12930), .Z(n12924) );
  AND U12556 ( .A(n563), .B(n12931), .Z(n12930) );
  XOR U12557 ( .A(p_input[780]), .B(n12929), .Z(n12931) );
  XNOR U12558 ( .A(n12932), .B(n12933), .Z(n12929) );
  AND U12559 ( .A(n567), .B(n12928), .Z(n12933) );
  XNOR U12560 ( .A(n12932), .B(n12926), .Z(n12928) );
  XOR U12561 ( .A(n12934), .B(n12935), .Z(n12926) );
  AND U12562 ( .A(n582), .B(n12936), .Z(n12935) );
  XNOR U12563 ( .A(n12937), .B(n12938), .Z(n12932) );
  AND U12564 ( .A(n574), .B(n12939), .Z(n12938) );
  XOR U12565 ( .A(p_input[796]), .B(n12937), .Z(n12939) );
  XNOR U12566 ( .A(n12940), .B(n12941), .Z(n12937) );
  AND U12567 ( .A(n578), .B(n12936), .Z(n12941) );
  XNOR U12568 ( .A(n12940), .B(n12934), .Z(n12936) );
  XOR U12569 ( .A(n12942), .B(n12943), .Z(n12934) );
  AND U12570 ( .A(n593), .B(n12944), .Z(n12943) );
  XNOR U12571 ( .A(n12945), .B(n12946), .Z(n12940) );
  AND U12572 ( .A(n585), .B(n12947), .Z(n12946) );
  XOR U12573 ( .A(p_input[812]), .B(n12945), .Z(n12947) );
  XNOR U12574 ( .A(n12948), .B(n12949), .Z(n12945) );
  AND U12575 ( .A(n589), .B(n12944), .Z(n12949) );
  XNOR U12576 ( .A(n12948), .B(n12942), .Z(n12944) );
  XOR U12577 ( .A(n12950), .B(n12951), .Z(n12942) );
  AND U12578 ( .A(n604), .B(n12952), .Z(n12951) );
  XNOR U12579 ( .A(n12953), .B(n12954), .Z(n12948) );
  AND U12580 ( .A(n596), .B(n12955), .Z(n12954) );
  XOR U12581 ( .A(p_input[828]), .B(n12953), .Z(n12955) );
  XNOR U12582 ( .A(n12956), .B(n12957), .Z(n12953) );
  AND U12583 ( .A(n600), .B(n12952), .Z(n12957) );
  XNOR U12584 ( .A(n12956), .B(n12950), .Z(n12952) );
  XOR U12585 ( .A(n12958), .B(n12959), .Z(n12950) );
  AND U12586 ( .A(n615), .B(n12960), .Z(n12959) );
  XNOR U12587 ( .A(n12961), .B(n12962), .Z(n12956) );
  AND U12588 ( .A(n607), .B(n12963), .Z(n12962) );
  XOR U12589 ( .A(p_input[844]), .B(n12961), .Z(n12963) );
  XNOR U12590 ( .A(n12964), .B(n12965), .Z(n12961) );
  AND U12591 ( .A(n611), .B(n12960), .Z(n12965) );
  XNOR U12592 ( .A(n12964), .B(n12958), .Z(n12960) );
  XOR U12593 ( .A(n12966), .B(n12967), .Z(n12958) );
  AND U12594 ( .A(n626), .B(n12968), .Z(n12967) );
  XNOR U12595 ( .A(n12969), .B(n12970), .Z(n12964) );
  AND U12596 ( .A(n618), .B(n12971), .Z(n12970) );
  XOR U12597 ( .A(p_input[860]), .B(n12969), .Z(n12971) );
  XNOR U12598 ( .A(n12972), .B(n12973), .Z(n12969) );
  AND U12599 ( .A(n622), .B(n12968), .Z(n12973) );
  XNOR U12600 ( .A(n12972), .B(n12966), .Z(n12968) );
  XOR U12601 ( .A(n12974), .B(n12975), .Z(n12966) );
  AND U12602 ( .A(n637), .B(n12976), .Z(n12975) );
  XNOR U12603 ( .A(n12977), .B(n12978), .Z(n12972) );
  AND U12604 ( .A(n629), .B(n12979), .Z(n12978) );
  XOR U12605 ( .A(p_input[876]), .B(n12977), .Z(n12979) );
  XNOR U12606 ( .A(n12980), .B(n12981), .Z(n12977) );
  AND U12607 ( .A(n633), .B(n12976), .Z(n12981) );
  XNOR U12608 ( .A(n12980), .B(n12974), .Z(n12976) );
  XOR U12609 ( .A(n12982), .B(n12983), .Z(n12974) );
  AND U12610 ( .A(n648), .B(n12984), .Z(n12983) );
  XNOR U12611 ( .A(n12985), .B(n12986), .Z(n12980) );
  AND U12612 ( .A(n640), .B(n12987), .Z(n12986) );
  XOR U12613 ( .A(p_input[892]), .B(n12985), .Z(n12987) );
  XNOR U12614 ( .A(n12988), .B(n12989), .Z(n12985) );
  AND U12615 ( .A(n644), .B(n12984), .Z(n12989) );
  XNOR U12616 ( .A(n12988), .B(n12982), .Z(n12984) );
  XOR U12617 ( .A(n12990), .B(n12991), .Z(n12982) );
  AND U12618 ( .A(n659), .B(n12992), .Z(n12991) );
  XNOR U12619 ( .A(n12993), .B(n12994), .Z(n12988) );
  AND U12620 ( .A(n651), .B(n12995), .Z(n12994) );
  XOR U12621 ( .A(p_input[908]), .B(n12993), .Z(n12995) );
  XNOR U12622 ( .A(n12996), .B(n12997), .Z(n12993) );
  AND U12623 ( .A(n655), .B(n12992), .Z(n12997) );
  XNOR U12624 ( .A(n12996), .B(n12990), .Z(n12992) );
  XOR U12625 ( .A(n12998), .B(n12999), .Z(n12990) );
  AND U12626 ( .A(n670), .B(n13000), .Z(n12999) );
  XNOR U12627 ( .A(n13001), .B(n13002), .Z(n12996) );
  AND U12628 ( .A(n662), .B(n13003), .Z(n13002) );
  XOR U12629 ( .A(p_input[924]), .B(n13001), .Z(n13003) );
  XNOR U12630 ( .A(n13004), .B(n13005), .Z(n13001) );
  AND U12631 ( .A(n666), .B(n13000), .Z(n13005) );
  XNOR U12632 ( .A(n13004), .B(n12998), .Z(n13000) );
  XOR U12633 ( .A(n13006), .B(n13007), .Z(n12998) );
  AND U12634 ( .A(n681), .B(n13008), .Z(n13007) );
  XNOR U12635 ( .A(n13009), .B(n13010), .Z(n13004) );
  AND U12636 ( .A(n673), .B(n13011), .Z(n13010) );
  XOR U12637 ( .A(p_input[940]), .B(n13009), .Z(n13011) );
  XNOR U12638 ( .A(n13012), .B(n13013), .Z(n13009) );
  AND U12639 ( .A(n677), .B(n13008), .Z(n13013) );
  XNOR U12640 ( .A(n13012), .B(n13006), .Z(n13008) );
  XOR U12641 ( .A(n13014), .B(n13015), .Z(n13006) );
  AND U12642 ( .A(n692), .B(n13016), .Z(n13015) );
  XNOR U12643 ( .A(n13017), .B(n13018), .Z(n13012) );
  AND U12644 ( .A(n684), .B(n13019), .Z(n13018) );
  XOR U12645 ( .A(p_input[956]), .B(n13017), .Z(n13019) );
  XNOR U12646 ( .A(n13020), .B(n13021), .Z(n13017) );
  AND U12647 ( .A(n688), .B(n13016), .Z(n13021) );
  XNOR U12648 ( .A(n13020), .B(n13014), .Z(n13016) );
  XOR U12649 ( .A(n13022), .B(n13023), .Z(n13014) );
  AND U12650 ( .A(n703), .B(n13024), .Z(n13023) );
  XNOR U12651 ( .A(n13025), .B(n13026), .Z(n13020) );
  AND U12652 ( .A(n695), .B(n13027), .Z(n13026) );
  XOR U12653 ( .A(p_input[972]), .B(n13025), .Z(n13027) );
  XNOR U12654 ( .A(n13028), .B(n13029), .Z(n13025) );
  AND U12655 ( .A(n699), .B(n13024), .Z(n13029) );
  XNOR U12656 ( .A(n13028), .B(n13022), .Z(n13024) );
  XOR U12657 ( .A(n13030), .B(n13031), .Z(n13022) );
  AND U12658 ( .A(n714), .B(n13032), .Z(n13031) );
  XNOR U12659 ( .A(n13033), .B(n13034), .Z(n13028) );
  AND U12660 ( .A(n706), .B(n13035), .Z(n13034) );
  XOR U12661 ( .A(p_input[988]), .B(n13033), .Z(n13035) );
  XNOR U12662 ( .A(n13036), .B(n13037), .Z(n13033) );
  AND U12663 ( .A(n710), .B(n13032), .Z(n13037) );
  XNOR U12664 ( .A(n13036), .B(n13030), .Z(n13032) );
  XOR U12665 ( .A(n13038), .B(n13039), .Z(n13030) );
  AND U12666 ( .A(n725), .B(n13040), .Z(n13039) );
  XNOR U12667 ( .A(n13041), .B(n13042), .Z(n13036) );
  AND U12668 ( .A(n717), .B(n13043), .Z(n13042) );
  XOR U12669 ( .A(p_input[1004]), .B(n13041), .Z(n13043) );
  XNOR U12670 ( .A(n13044), .B(n13045), .Z(n13041) );
  AND U12671 ( .A(n721), .B(n13040), .Z(n13045) );
  XNOR U12672 ( .A(n13044), .B(n13038), .Z(n13040) );
  XOR U12673 ( .A(n13046), .B(n13047), .Z(n13038) );
  AND U12674 ( .A(n736), .B(n13048), .Z(n13047) );
  XNOR U12675 ( .A(n13049), .B(n13050), .Z(n13044) );
  AND U12676 ( .A(n728), .B(n13051), .Z(n13050) );
  XOR U12677 ( .A(p_input[1020]), .B(n13049), .Z(n13051) );
  XNOR U12678 ( .A(n13052), .B(n13053), .Z(n13049) );
  AND U12679 ( .A(n732), .B(n13048), .Z(n13053) );
  XNOR U12680 ( .A(n13052), .B(n13046), .Z(n13048) );
  XOR U12681 ( .A(n13054), .B(n13055), .Z(n13046) );
  AND U12682 ( .A(n747), .B(n13056), .Z(n13055) );
  XNOR U12683 ( .A(n13057), .B(n13058), .Z(n13052) );
  AND U12684 ( .A(n739), .B(n13059), .Z(n13058) );
  XOR U12685 ( .A(p_input[1036]), .B(n13057), .Z(n13059) );
  XNOR U12686 ( .A(n13060), .B(n13061), .Z(n13057) );
  AND U12687 ( .A(n743), .B(n13056), .Z(n13061) );
  XNOR U12688 ( .A(n13060), .B(n13054), .Z(n13056) );
  XOR U12689 ( .A(n13062), .B(n13063), .Z(n13054) );
  AND U12690 ( .A(n758), .B(n13064), .Z(n13063) );
  XNOR U12691 ( .A(n13065), .B(n13066), .Z(n13060) );
  AND U12692 ( .A(n750), .B(n13067), .Z(n13066) );
  XOR U12693 ( .A(p_input[1052]), .B(n13065), .Z(n13067) );
  XNOR U12694 ( .A(n13068), .B(n13069), .Z(n13065) );
  AND U12695 ( .A(n754), .B(n13064), .Z(n13069) );
  XNOR U12696 ( .A(n13068), .B(n13062), .Z(n13064) );
  XOR U12697 ( .A(n13070), .B(n13071), .Z(n13062) );
  AND U12698 ( .A(n769), .B(n13072), .Z(n13071) );
  XNOR U12699 ( .A(n13073), .B(n13074), .Z(n13068) );
  AND U12700 ( .A(n761), .B(n13075), .Z(n13074) );
  XOR U12701 ( .A(p_input[1068]), .B(n13073), .Z(n13075) );
  XNOR U12702 ( .A(n13076), .B(n13077), .Z(n13073) );
  AND U12703 ( .A(n765), .B(n13072), .Z(n13077) );
  XNOR U12704 ( .A(n13076), .B(n13070), .Z(n13072) );
  XOR U12705 ( .A(n13078), .B(n13079), .Z(n13070) );
  AND U12706 ( .A(n780), .B(n13080), .Z(n13079) );
  XNOR U12707 ( .A(n13081), .B(n13082), .Z(n13076) );
  AND U12708 ( .A(n772), .B(n13083), .Z(n13082) );
  XOR U12709 ( .A(p_input[1084]), .B(n13081), .Z(n13083) );
  XNOR U12710 ( .A(n13084), .B(n13085), .Z(n13081) );
  AND U12711 ( .A(n776), .B(n13080), .Z(n13085) );
  XNOR U12712 ( .A(n13084), .B(n13078), .Z(n13080) );
  XOR U12713 ( .A(n13086), .B(n13087), .Z(n13078) );
  AND U12714 ( .A(n791), .B(n13088), .Z(n13087) );
  XNOR U12715 ( .A(n13089), .B(n13090), .Z(n13084) );
  AND U12716 ( .A(n783), .B(n13091), .Z(n13090) );
  XOR U12717 ( .A(p_input[1100]), .B(n13089), .Z(n13091) );
  XNOR U12718 ( .A(n13092), .B(n13093), .Z(n13089) );
  AND U12719 ( .A(n787), .B(n13088), .Z(n13093) );
  XNOR U12720 ( .A(n13092), .B(n13086), .Z(n13088) );
  XOR U12721 ( .A(n13094), .B(n13095), .Z(n13086) );
  AND U12722 ( .A(n802), .B(n13096), .Z(n13095) );
  XNOR U12723 ( .A(n13097), .B(n13098), .Z(n13092) );
  AND U12724 ( .A(n794), .B(n13099), .Z(n13098) );
  XOR U12725 ( .A(p_input[1116]), .B(n13097), .Z(n13099) );
  XNOR U12726 ( .A(n13100), .B(n13101), .Z(n13097) );
  AND U12727 ( .A(n798), .B(n13096), .Z(n13101) );
  XNOR U12728 ( .A(n13100), .B(n13094), .Z(n13096) );
  XOR U12729 ( .A(n13102), .B(n13103), .Z(n13094) );
  AND U12730 ( .A(n813), .B(n13104), .Z(n13103) );
  XNOR U12731 ( .A(n13105), .B(n13106), .Z(n13100) );
  AND U12732 ( .A(n805), .B(n13107), .Z(n13106) );
  XOR U12733 ( .A(p_input[1132]), .B(n13105), .Z(n13107) );
  XNOR U12734 ( .A(n13108), .B(n13109), .Z(n13105) );
  AND U12735 ( .A(n809), .B(n13104), .Z(n13109) );
  XNOR U12736 ( .A(n13108), .B(n13102), .Z(n13104) );
  XOR U12737 ( .A(n13110), .B(n13111), .Z(n13102) );
  AND U12738 ( .A(n824), .B(n13112), .Z(n13111) );
  XNOR U12739 ( .A(n13113), .B(n13114), .Z(n13108) );
  AND U12740 ( .A(n816), .B(n13115), .Z(n13114) );
  XOR U12741 ( .A(p_input[1148]), .B(n13113), .Z(n13115) );
  XNOR U12742 ( .A(n13116), .B(n13117), .Z(n13113) );
  AND U12743 ( .A(n820), .B(n13112), .Z(n13117) );
  XNOR U12744 ( .A(n13116), .B(n13110), .Z(n13112) );
  XOR U12745 ( .A(n13118), .B(n13119), .Z(n13110) );
  AND U12746 ( .A(n835), .B(n13120), .Z(n13119) );
  XNOR U12747 ( .A(n13121), .B(n13122), .Z(n13116) );
  AND U12748 ( .A(n827), .B(n13123), .Z(n13122) );
  XOR U12749 ( .A(p_input[1164]), .B(n13121), .Z(n13123) );
  XNOR U12750 ( .A(n13124), .B(n13125), .Z(n13121) );
  AND U12751 ( .A(n831), .B(n13120), .Z(n13125) );
  XNOR U12752 ( .A(n13124), .B(n13118), .Z(n13120) );
  XOR U12753 ( .A(n13126), .B(n13127), .Z(n13118) );
  AND U12754 ( .A(n846), .B(n13128), .Z(n13127) );
  XNOR U12755 ( .A(n13129), .B(n13130), .Z(n13124) );
  AND U12756 ( .A(n838), .B(n13131), .Z(n13130) );
  XOR U12757 ( .A(p_input[1180]), .B(n13129), .Z(n13131) );
  XNOR U12758 ( .A(n13132), .B(n13133), .Z(n13129) );
  AND U12759 ( .A(n842), .B(n13128), .Z(n13133) );
  XNOR U12760 ( .A(n13132), .B(n13126), .Z(n13128) );
  XOR U12761 ( .A(n13134), .B(n13135), .Z(n13126) );
  AND U12762 ( .A(n857), .B(n13136), .Z(n13135) );
  XNOR U12763 ( .A(n13137), .B(n13138), .Z(n13132) );
  AND U12764 ( .A(n849), .B(n13139), .Z(n13138) );
  XOR U12765 ( .A(p_input[1196]), .B(n13137), .Z(n13139) );
  XNOR U12766 ( .A(n13140), .B(n13141), .Z(n13137) );
  AND U12767 ( .A(n853), .B(n13136), .Z(n13141) );
  XNOR U12768 ( .A(n13140), .B(n13134), .Z(n13136) );
  XOR U12769 ( .A(n13142), .B(n13143), .Z(n13134) );
  AND U12770 ( .A(n868), .B(n13144), .Z(n13143) );
  XNOR U12771 ( .A(n13145), .B(n13146), .Z(n13140) );
  AND U12772 ( .A(n860), .B(n13147), .Z(n13146) );
  XOR U12773 ( .A(p_input[1212]), .B(n13145), .Z(n13147) );
  XNOR U12774 ( .A(n13148), .B(n13149), .Z(n13145) );
  AND U12775 ( .A(n864), .B(n13144), .Z(n13149) );
  XNOR U12776 ( .A(n13148), .B(n13142), .Z(n13144) );
  XOR U12777 ( .A(n13150), .B(n13151), .Z(n13142) );
  AND U12778 ( .A(n879), .B(n13152), .Z(n13151) );
  XNOR U12779 ( .A(n13153), .B(n13154), .Z(n13148) );
  AND U12780 ( .A(n871), .B(n13155), .Z(n13154) );
  XOR U12781 ( .A(p_input[1228]), .B(n13153), .Z(n13155) );
  XNOR U12782 ( .A(n13156), .B(n13157), .Z(n13153) );
  AND U12783 ( .A(n875), .B(n13152), .Z(n13157) );
  XNOR U12784 ( .A(n13156), .B(n13150), .Z(n13152) );
  XOR U12785 ( .A(n13158), .B(n13159), .Z(n13150) );
  AND U12786 ( .A(n890), .B(n13160), .Z(n13159) );
  XNOR U12787 ( .A(n13161), .B(n13162), .Z(n13156) );
  AND U12788 ( .A(n882), .B(n13163), .Z(n13162) );
  XOR U12789 ( .A(p_input[1244]), .B(n13161), .Z(n13163) );
  XNOR U12790 ( .A(n13164), .B(n13165), .Z(n13161) );
  AND U12791 ( .A(n886), .B(n13160), .Z(n13165) );
  XNOR U12792 ( .A(n13164), .B(n13158), .Z(n13160) );
  XOR U12793 ( .A(n13166), .B(n13167), .Z(n13158) );
  AND U12794 ( .A(n901), .B(n13168), .Z(n13167) );
  XNOR U12795 ( .A(n13169), .B(n13170), .Z(n13164) );
  AND U12796 ( .A(n893), .B(n13171), .Z(n13170) );
  XOR U12797 ( .A(p_input[1260]), .B(n13169), .Z(n13171) );
  XNOR U12798 ( .A(n13172), .B(n13173), .Z(n13169) );
  AND U12799 ( .A(n897), .B(n13168), .Z(n13173) );
  XNOR U12800 ( .A(n13172), .B(n13166), .Z(n13168) );
  XOR U12801 ( .A(n13174), .B(n13175), .Z(n13166) );
  AND U12802 ( .A(n912), .B(n13176), .Z(n13175) );
  XNOR U12803 ( .A(n13177), .B(n13178), .Z(n13172) );
  AND U12804 ( .A(n904), .B(n13179), .Z(n13178) );
  XOR U12805 ( .A(p_input[1276]), .B(n13177), .Z(n13179) );
  XNOR U12806 ( .A(n13180), .B(n13181), .Z(n13177) );
  AND U12807 ( .A(n908), .B(n13176), .Z(n13181) );
  XNOR U12808 ( .A(n13180), .B(n13174), .Z(n13176) );
  XOR U12809 ( .A(n13182), .B(n13183), .Z(n13174) );
  AND U12810 ( .A(n923), .B(n13184), .Z(n13183) );
  XNOR U12811 ( .A(n13185), .B(n13186), .Z(n13180) );
  AND U12812 ( .A(n915), .B(n13187), .Z(n13186) );
  XOR U12813 ( .A(p_input[1292]), .B(n13185), .Z(n13187) );
  XNOR U12814 ( .A(n13188), .B(n13189), .Z(n13185) );
  AND U12815 ( .A(n919), .B(n13184), .Z(n13189) );
  XNOR U12816 ( .A(n13188), .B(n13182), .Z(n13184) );
  XOR U12817 ( .A(n13190), .B(n13191), .Z(n13182) );
  AND U12818 ( .A(n934), .B(n13192), .Z(n13191) );
  XNOR U12819 ( .A(n13193), .B(n13194), .Z(n13188) );
  AND U12820 ( .A(n926), .B(n13195), .Z(n13194) );
  XOR U12821 ( .A(p_input[1308]), .B(n13193), .Z(n13195) );
  XNOR U12822 ( .A(n13196), .B(n13197), .Z(n13193) );
  AND U12823 ( .A(n930), .B(n13192), .Z(n13197) );
  XNOR U12824 ( .A(n13196), .B(n13190), .Z(n13192) );
  XOR U12825 ( .A(n13198), .B(n13199), .Z(n13190) );
  AND U12826 ( .A(n945), .B(n13200), .Z(n13199) );
  XNOR U12827 ( .A(n13201), .B(n13202), .Z(n13196) );
  AND U12828 ( .A(n937), .B(n13203), .Z(n13202) );
  XOR U12829 ( .A(p_input[1324]), .B(n13201), .Z(n13203) );
  XNOR U12830 ( .A(n13204), .B(n13205), .Z(n13201) );
  AND U12831 ( .A(n941), .B(n13200), .Z(n13205) );
  XNOR U12832 ( .A(n13204), .B(n13198), .Z(n13200) );
  XOR U12833 ( .A(n13206), .B(n13207), .Z(n13198) );
  AND U12834 ( .A(n956), .B(n13208), .Z(n13207) );
  XNOR U12835 ( .A(n13209), .B(n13210), .Z(n13204) );
  AND U12836 ( .A(n948), .B(n13211), .Z(n13210) );
  XOR U12837 ( .A(p_input[1340]), .B(n13209), .Z(n13211) );
  XNOR U12838 ( .A(n13212), .B(n13213), .Z(n13209) );
  AND U12839 ( .A(n952), .B(n13208), .Z(n13213) );
  XNOR U12840 ( .A(n13212), .B(n13206), .Z(n13208) );
  XOR U12841 ( .A(n13214), .B(n13215), .Z(n13206) );
  AND U12842 ( .A(n967), .B(n13216), .Z(n13215) );
  XNOR U12843 ( .A(n13217), .B(n13218), .Z(n13212) );
  AND U12844 ( .A(n959), .B(n13219), .Z(n13218) );
  XOR U12845 ( .A(p_input[1356]), .B(n13217), .Z(n13219) );
  XNOR U12846 ( .A(n13220), .B(n13221), .Z(n13217) );
  AND U12847 ( .A(n963), .B(n13216), .Z(n13221) );
  XNOR U12848 ( .A(n13220), .B(n13214), .Z(n13216) );
  XOR U12849 ( .A(n13222), .B(n13223), .Z(n13214) );
  AND U12850 ( .A(n978), .B(n13224), .Z(n13223) );
  XNOR U12851 ( .A(n13225), .B(n13226), .Z(n13220) );
  AND U12852 ( .A(n970), .B(n13227), .Z(n13226) );
  XOR U12853 ( .A(p_input[1372]), .B(n13225), .Z(n13227) );
  XNOR U12854 ( .A(n13228), .B(n13229), .Z(n13225) );
  AND U12855 ( .A(n974), .B(n13224), .Z(n13229) );
  XNOR U12856 ( .A(n13228), .B(n13222), .Z(n13224) );
  XOR U12857 ( .A(n13230), .B(n13231), .Z(n13222) );
  AND U12858 ( .A(n989), .B(n13232), .Z(n13231) );
  XNOR U12859 ( .A(n13233), .B(n13234), .Z(n13228) );
  AND U12860 ( .A(n981), .B(n13235), .Z(n13234) );
  XOR U12861 ( .A(p_input[1388]), .B(n13233), .Z(n13235) );
  XNOR U12862 ( .A(n13236), .B(n13237), .Z(n13233) );
  AND U12863 ( .A(n985), .B(n13232), .Z(n13237) );
  XNOR U12864 ( .A(n13236), .B(n13230), .Z(n13232) );
  XOR U12865 ( .A(n13238), .B(n13239), .Z(n13230) );
  AND U12866 ( .A(n1000), .B(n13240), .Z(n13239) );
  XNOR U12867 ( .A(n13241), .B(n13242), .Z(n13236) );
  AND U12868 ( .A(n992), .B(n13243), .Z(n13242) );
  XOR U12869 ( .A(p_input[1404]), .B(n13241), .Z(n13243) );
  XNOR U12870 ( .A(n13244), .B(n13245), .Z(n13241) );
  AND U12871 ( .A(n996), .B(n13240), .Z(n13245) );
  XNOR U12872 ( .A(n13244), .B(n13238), .Z(n13240) );
  XOR U12873 ( .A(n13246), .B(n13247), .Z(n13238) );
  AND U12874 ( .A(n1011), .B(n13248), .Z(n13247) );
  XNOR U12875 ( .A(n13249), .B(n13250), .Z(n13244) );
  AND U12876 ( .A(n1003), .B(n13251), .Z(n13250) );
  XOR U12877 ( .A(p_input[1420]), .B(n13249), .Z(n13251) );
  XNOR U12878 ( .A(n13252), .B(n13253), .Z(n13249) );
  AND U12879 ( .A(n1007), .B(n13248), .Z(n13253) );
  XNOR U12880 ( .A(n13252), .B(n13246), .Z(n13248) );
  XOR U12881 ( .A(n13254), .B(n13255), .Z(n13246) );
  AND U12882 ( .A(n1022), .B(n13256), .Z(n13255) );
  XNOR U12883 ( .A(n13257), .B(n13258), .Z(n13252) );
  AND U12884 ( .A(n1014), .B(n13259), .Z(n13258) );
  XOR U12885 ( .A(p_input[1436]), .B(n13257), .Z(n13259) );
  XNOR U12886 ( .A(n13260), .B(n13261), .Z(n13257) );
  AND U12887 ( .A(n1018), .B(n13256), .Z(n13261) );
  XNOR U12888 ( .A(n13260), .B(n13254), .Z(n13256) );
  XOR U12889 ( .A(n13262), .B(n13263), .Z(n13254) );
  AND U12890 ( .A(n1033), .B(n13264), .Z(n13263) );
  XNOR U12891 ( .A(n13265), .B(n13266), .Z(n13260) );
  AND U12892 ( .A(n1025), .B(n13267), .Z(n13266) );
  XOR U12893 ( .A(p_input[1452]), .B(n13265), .Z(n13267) );
  XNOR U12894 ( .A(n13268), .B(n13269), .Z(n13265) );
  AND U12895 ( .A(n1029), .B(n13264), .Z(n13269) );
  XNOR U12896 ( .A(n13268), .B(n13262), .Z(n13264) );
  XOR U12897 ( .A(n13270), .B(n13271), .Z(n13262) );
  AND U12898 ( .A(n1044), .B(n13272), .Z(n13271) );
  XNOR U12899 ( .A(n13273), .B(n13274), .Z(n13268) );
  AND U12900 ( .A(n1036), .B(n13275), .Z(n13274) );
  XOR U12901 ( .A(p_input[1468]), .B(n13273), .Z(n13275) );
  XNOR U12902 ( .A(n13276), .B(n13277), .Z(n13273) );
  AND U12903 ( .A(n1040), .B(n13272), .Z(n13277) );
  XNOR U12904 ( .A(n13276), .B(n13270), .Z(n13272) );
  XOR U12905 ( .A(n13278), .B(n13279), .Z(n13270) );
  AND U12906 ( .A(n1055), .B(n13280), .Z(n13279) );
  XNOR U12907 ( .A(n13281), .B(n13282), .Z(n13276) );
  AND U12908 ( .A(n1047), .B(n13283), .Z(n13282) );
  XOR U12909 ( .A(p_input[1484]), .B(n13281), .Z(n13283) );
  XNOR U12910 ( .A(n13284), .B(n13285), .Z(n13281) );
  AND U12911 ( .A(n1051), .B(n13280), .Z(n13285) );
  XNOR U12912 ( .A(n13284), .B(n13278), .Z(n13280) );
  XOR U12913 ( .A(n13286), .B(n13287), .Z(n13278) );
  AND U12914 ( .A(n1066), .B(n13288), .Z(n13287) );
  XNOR U12915 ( .A(n13289), .B(n13290), .Z(n13284) );
  AND U12916 ( .A(n1058), .B(n13291), .Z(n13290) );
  XOR U12917 ( .A(p_input[1500]), .B(n13289), .Z(n13291) );
  XNOR U12918 ( .A(n13292), .B(n13293), .Z(n13289) );
  AND U12919 ( .A(n1062), .B(n13288), .Z(n13293) );
  XNOR U12920 ( .A(n13292), .B(n13286), .Z(n13288) );
  XOR U12921 ( .A(n13294), .B(n13295), .Z(n13286) );
  AND U12922 ( .A(n1077), .B(n13296), .Z(n13295) );
  XNOR U12923 ( .A(n13297), .B(n13298), .Z(n13292) );
  AND U12924 ( .A(n1069), .B(n13299), .Z(n13298) );
  XOR U12925 ( .A(p_input[1516]), .B(n13297), .Z(n13299) );
  XNOR U12926 ( .A(n13300), .B(n13301), .Z(n13297) );
  AND U12927 ( .A(n1073), .B(n13296), .Z(n13301) );
  XNOR U12928 ( .A(n13300), .B(n13294), .Z(n13296) );
  XOR U12929 ( .A(n13302), .B(n13303), .Z(n13294) );
  AND U12930 ( .A(n1088), .B(n13304), .Z(n13303) );
  XNOR U12931 ( .A(n13305), .B(n13306), .Z(n13300) );
  AND U12932 ( .A(n1080), .B(n13307), .Z(n13306) );
  XOR U12933 ( .A(p_input[1532]), .B(n13305), .Z(n13307) );
  XNOR U12934 ( .A(n13308), .B(n13309), .Z(n13305) );
  AND U12935 ( .A(n1084), .B(n13304), .Z(n13309) );
  XNOR U12936 ( .A(n13308), .B(n13302), .Z(n13304) );
  XOR U12937 ( .A(n13310), .B(n13311), .Z(n13302) );
  AND U12938 ( .A(n1099), .B(n13312), .Z(n13311) );
  XNOR U12939 ( .A(n13313), .B(n13314), .Z(n13308) );
  AND U12940 ( .A(n1091), .B(n13315), .Z(n13314) );
  XOR U12941 ( .A(p_input[1548]), .B(n13313), .Z(n13315) );
  XNOR U12942 ( .A(n13316), .B(n13317), .Z(n13313) );
  AND U12943 ( .A(n1095), .B(n13312), .Z(n13317) );
  XNOR U12944 ( .A(n13316), .B(n13310), .Z(n13312) );
  XOR U12945 ( .A(n13318), .B(n13319), .Z(n13310) );
  AND U12946 ( .A(n1110), .B(n13320), .Z(n13319) );
  XNOR U12947 ( .A(n13321), .B(n13322), .Z(n13316) );
  AND U12948 ( .A(n1102), .B(n13323), .Z(n13322) );
  XOR U12949 ( .A(p_input[1564]), .B(n13321), .Z(n13323) );
  XNOR U12950 ( .A(n13324), .B(n13325), .Z(n13321) );
  AND U12951 ( .A(n1106), .B(n13320), .Z(n13325) );
  XNOR U12952 ( .A(n13324), .B(n13318), .Z(n13320) );
  XOR U12953 ( .A(n13326), .B(n13327), .Z(n13318) );
  AND U12954 ( .A(n1121), .B(n13328), .Z(n13327) );
  XNOR U12955 ( .A(n13329), .B(n13330), .Z(n13324) );
  AND U12956 ( .A(n1113), .B(n13331), .Z(n13330) );
  XOR U12957 ( .A(p_input[1580]), .B(n13329), .Z(n13331) );
  XNOR U12958 ( .A(n13332), .B(n13333), .Z(n13329) );
  AND U12959 ( .A(n1117), .B(n13328), .Z(n13333) );
  XNOR U12960 ( .A(n13332), .B(n13326), .Z(n13328) );
  XOR U12961 ( .A(n13334), .B(n13335), .Z(n13326) );
  AND U12962 ( .A(n1132), .B(n13336), .Z(n13335) );
  XNOR U12963 ( .A(n13337), .B(n13338), .Z(n13332) );
  AND U12964 ( .A(n1124), .B(n13339), .Z(n13338) );
  XOR U12965 ( .A(p_input[1596]), .B(n13337), .Z(n13339) );
  XNOR U12966 ( .A(n13340), .B(n13341), .Z(n13337) );
  AND U12967 ( .A(n1128), .B(n13336), .Z(n13341) );
  XNOR U12968 ( .A(n13340), .B(n13334), .Z(n13336) );
  XOR U12969 ( .A(n13342), .B(n13343), .Z(n13334) );
  AND U12970 ( .A(n1143), .B(n13344), .Z(n13343) );
  XNOR U12971 ( .A(n13345), .B(n13346), .Z(n13340) );
  AND U12972 ( .A(n1135), .B(n13347), .Z(n13346) );
  XOR U12973 ( .A(p_input[1612]), .B(n13345), .Z(n13347) );
  XNOR U12974 ( .A(n13348), .B(n13349), .Z(n13345) );
  AND U12975 ( .A(n1139), .B(n13344), .Z(n13349) );
  XNOR U12976 ( .A(n13348), .B(n13342), .Z(n13344) );
  XOR U12977 ( .A(n13350), .B(n13351), .Z(n13342) );
  AND U12978 ( .A(n1154), .B(n13352), .Z(n13351) );
  XNOR U12979 ( .A(n13353), .B(n13354), .Z(n13348) );
  AND U12980 ( .A(n1146), .B(n13355), .Z(n13354) );
  XOR U12981 ( .A(p_input[1628]), .B(n13353), .Z(n13355) );
  XNOR U12982 ( .A(n13356), .B(n13357), .Z(n13353) );
  AND U12983 ( .A(n1150), .B(n13352), .Z(n13357) );
  XNOR U12984 ( .A(n13356), .B(n13350), .Z(n13352) );
  XOR U12985 ( .A(n13358), .B(n13359), .Z(n13350) );
  AND U12986 ( .A(n1165), .B(n13360), .Z(n13359) );
  XNOR U12987 ( .A(n13361), .B(n13362), .Z(n13356) );
  AND U12988 ( .A(n1157), .B(n13363), .Z(n13362) );
  XOR U12989 ( .A(p_input[1644]), .B(n13361), .Z(n13363) );
  XNOR U12990 ( .A(n13364), .B(n13365), .Z(n13361) );
  AND U12991 ( .A(n1161), .B(n13360), .Z(n13365) );
  XNOR U12992 ( .A(n13364), .B(n13358), .Z(n13360) );
  XOR U12993 ( .A(n13366), .B(n13367), .Z(n13358) );
  AND U12994 ( .A(n1176), .B(n13368), .Z(n13367) );
  XNOR U12995 ( .A(n13369), .B(n13370), .Z(n13364) );
  AND U12996 ( .A(n1168), .B(n13371), .Z(n13370) );
  XOR U12997 ( .A(p_input[1660]), .B(n13369), .Z(n13371) );
  XNOR U12998 ( .A(n13372), .B(n13373), .Z(n13369) );
  AND U12999 ( .A(n1172), .B(n13368), .Z(n13373) );
  XNOR U13000 ( .A(n13372), .B(n13366), .Z(n13368) );
  XOR U13001 ( .A(n13374), .B(n13375), .Z(n13366) );
  AND U13002 ( .A(n1187), .B(n13376), .Z(n13375) );
  XNOR U13003 ( .A(n13377), .B(n13378), .Z(n13372) );
  AND U13004 ( .A(n1179), .B(n13379), .Z(n13378) );
  XOR U13005 ( .A(p_input[1676]), .B(n13377), .Z(n13379) );
  XNOR U13006 ( .A(n13380), .B(n13381), .Z(n13377) );
  AND U13007 ( .A(n1183), .B(n13376), .Z(n13381) );
  XNOR U13008 ( .A(n13380), .B(n13374), .Z(n13376) );
  XOR U13009 ( .A(n13382), .B(n13383), .Z(n13374) );
  AND U13010 ( .A(n1198), .B(n13384), .Z(n13383) );
  XNOR U13011 ( .A(n13385), .B(n13386), .Z(n13380) );
  AND U13012 ( .A(n1190), .B(n13387), .Z(n13386) );
  XOR U13013 ( .A(p_input[1692]), .B(n13385), .Z(n13387) );
  XNOR U13014 ( .A(n13388), .B(n13389), .Z(n13385) );
  AND U13015 ( .A(n1194), .B(n13384), .Z(n13389) );
  XNOR U13016 ( .A(n13388), .B(n13382), .Z(n13384) );
  XOR U13017 ( .A(n13390), .B(n13391), .Z(n13382) );
  AND U13018 ( .A(n1209), .B(n13392), .Z(n13391) );
  XNOR U13019 ( .A(n13393), .B(n13394), .Z(n13388) );
  AND U13020 ( .A(n1201), .B(n13395), .Z(n13394) );
  XOR U13021 ( .A(p_input[1708]), .B(n13393), .Z(n13395) );
  XNOR U13022 ( .A(n13396), .B(n13397), .Z(n13393) );
  AND U13023 ( .A(n1205), .B(n13392), .Z(n13397) );
  XNOR U13024 ( .A(n13396), .B(n13390), .Z(n13392) );
  XOR U13025 ( .A(n13398), .B(n13399), .Z(n13390) );
  AND U13026 ( .A(n1220), .B(n13400), .Z(n13399) );
  XNOR U13027 ( .A(n13401), .B(n13402), .Z(n13396) );
  AND U13028 ( .A(n1212), .B(n13403), .Z(n13402) );
  XOR U13029 ( .A(p_input[1724]), .B(n13401), .Z(n13403) );
  XNOR U13030 ( .A(n13404), .B(n13405), .Z(n13401) );
  AND U13031 ( .A(n1216), .B(n13400), .Z(n13405) );
  XNOR U13032 ( .A(n13404), .B(n13398), .Z(n13400) );
  XOR U13033 ( .A(n13406), .B(n13407), .Z(n13398) );
  AND U13034 ( .A(n1231), .B(n13408), .Z(n13407) );
  XNOR U13035 ( .A(n13409), .B(n13410), .Z(n13404) );
  AND U13036 ( .A(n1223), .B(n13411), .Z(n13410) );
  XOR U13037 ( .A(p_input[1740]), .B(n13409), .Z(n13411) );
  XNOR U13038 ( .A(n13412), .B(n13413), .Z(n13409) );
  AND U13039 ( .A(n1227), .B(n13408), .Z(n13413) );
  XNOR U13040 ( .A(n13412), .B(n13406), .Z(n13408) );
  XOR U13041 ( .A(n13414), .B(n13415), .Z(n13406) );
  AND U13042 ( .A(n1242), .B(n13416), .Z(n13415) );
  XNOR U13043 ( .A(n13417), .B(n13418), .Z(n13412) );
  AND U13044 ( .A(n1234), .B(n13419), .Z(n13418) );
  XOR U13045 ( .A(p_input[1756]), .B(n13417), .Z(n13419) );
  XNOR U13046 ( .A(n13420), .B(n13421), .Z(n13417) );
  AND U13047 ( .A(n1238), .B(n13416), .Z(n13421) );
  XNOR U13048 ( .A(n13420), .B(n13414), .Z(n13416) );
  XOR U13049 ( .A(n13422), .B(n13423), .Z(n13414) );
  AND U13050 ( .A(n1253), .B(n13424), .Z(n13423) );
  XNOR U13051 ( .A(n13425), .B(n13426), .Z(n13420) );
  AND U13052 ( .A(n1245), .B(n13427), .Z(n13426) );
  XOR U13053 ( .A(p_input[1772]), .B(n13425), .Z(n13427) );
  XNOR U13054 ( .A(n13428), .B(n13429), .Z(n13425) );
  AND U13055 ( .A(n1249), .B(n13424), .Z(n13429) );
  XNOR U13056 ( .A(n13428), .B(n13422), .Z(n13424) );
  XOR U13057 ( .A(n13430), .B(n13431), .Z(n13422) );
  AND U13058 ( .A(n1264), .B(n13432), .Z(n13431) );
  XNOR U13059 ( .A(n13433), .B(n13434), .Z(n13428) );
  AND U13060 ( .A(n1256), .B(n13435), .Z(n13434) );
  XOR U13061 ( .A(p_input[1788]), .B(n13433), .Z(n13435) );
  XNOR U13062 ( .A(n13436), .B(n13437), .Z(n13433) );
  AND U13063 ( .A(n1260), .B(n13432), .Z(n13437) );
  XNOR U13064 ( .A(n13436), .B(n13430), .Z(n13432) );
  XOR U13065 ( .A(n13438), .B(n13439), .Z(n13430) );
  AND U13066 ( .A(n1275), .B(n13440), .Z(n13439) );
  XNOR U13067 ( .A(n13441), .B(n13442), .Z(n13436) );
  AND U13068 ( .A(n1267), .B(n13443), .Z(n13442) );
  XOR U13069 ( .A(p_input[1804]), .B(n13441), .Z(n13443) );
  XNOR U13070 ( .A(n13444), .B(n13445), .Z(n13441) );
  AND U13071 ( .A(n1271), .B(n13440), .Z(n13445) );
  XNOR U13072 ( .A(n13444), .B(n13438), .Z(n13440) );
  XOR U13073 ( .A(n13446), .B(n13447), .Z(n13438) );
  AND U13074 ( .A(n1286), .B(n13448), .Z(n13447) );
  XNOR U13075 ( .A(n13449), .B(n13450), .Z(n13444) );
  AND U13076 ( .A(n1278), .B(n13451), .Z(n13450) );
  XOR U13077 ( .A(p_input[1820]), .B(n13449), .Z(n13451) );
  XNOR U13078 ( .A(n13452), .B(n13453), .Z(n13449) );
  AND U13079 ( .A(n1282), .B(n13448), .Z(n13453) );
  XNOR U13080 ( .A(n13452), .B(n13446), .Z(n13448) );
  XOR U13081 ( .A(n13454), .B(n13455), .Z(n13446) );
  AND U13082 ( .A(n1297), .B(n13456), .Z(n13455) );
  XNOR U13083 ( .A(n13457), .B(n13458), .Z(n13452) );
  AND U13084 ( .A(n1289), .B(n13459), .Z(n13458) );
  XOR U13085 ( .A(p_input[1836]), .B(n13457), .Z(n13459) );
  XNOR U13086 ( .A(n13460), .B(n13461), .Z(n13457) );
  AND U13087 ( .A(n1293), .B(n13456), .Z(n13461) );
  XNOR U13088 ( .A(n13460), .B(n13454), .Z(n13456) );
  XOR U13089 ( .A(n13462), .B(n13463), .Z(n13454) );
  AND U13090 ( .A(n1308), .B(n13464), .Z(n13463) );
  XNOR U13091 ( .A(n13465), .B(n13466), .Z(n13460) );
  AND U13092 ( .A(n1300), .B(n13467), .Z(n13466) );
  XOR U13093 ( .A(p_input[1852]), .B(n13465), .Z(n13467) );
  XNOR U13094 ( .A(n13468), .B(n13469), .Z(n13465) );
  AND U13095 ( .A(n1304), .B(n13464), .Z(n13469) );
  XNOR U13096 ( .A(n13468), .B(n13462), .Z(n13464) );
  XOR U13097 ( .A(n13470), .B(n13471), .Z(n13462) );
  AND U13098 ( .A(n1319), .B(n13472), .Z(n13471) );
  XNOR U13099 ( .A(n13473), .B(n13474), .Z(n13468) );
  AND U13100 ( .A(n1311), .B(n13475), .Z(n13474) );
  XOR U13101 ( .A(p_input[1868]), .B(n13473), .Z(n13475) );
  XNOR U13102 ( .A(n13476), .B(n13477), .Z(n13473) );
  AND U13103 ( .A(n1315), .B(n13472), .Z(n13477) );
  XNOR U13104 ( .A(n13476), .B(n13470), .Z(n13472) );
  XOR U13105 ( .A(n13478), .B(n13479), .Z(n13470) );
  AND U13106 ( .A(n1330), .B(n13480), .Z(n13479) );
  XNOR U13107 ( .A(n13481), .B(n13482), .Z(n13476) );
  AND U13108 ( .A(n1322), .B(n13483), .Z(n13482) );
  XOR U13109 ( .A(p_input[1884]), .B(n13481), .Z(n13483) );
  XNOR U13110 ( .A(n13484), .B(n13485), .Z(n13481) );
  AND U13111 ( .A(n1326), .B(n13480), .Z(n13485) );
  XNOR U13112 ( .A(n13484), .B(n13478), .Z(n13480) );
  XOR U13113 ( .A(n13486), .B(n13487), .Z(n13478) );
  AND U13114 ( .A(n1341), .B(n13488), .Z(n13487) );
  XNOR U13115 ( .A(n13489), .B(n13490), .Z(n13484) );
  AND U13116 ( .A(n1333), .B(n13491), .Z(n13490) );
  XOR U13117 ( .A(p_input[1900]), .B(n13489), .Z(n13491) );
  XNOR U13118 ( .A(n13492), .B(n13493), .Z(n13489) );
  AND U13119 ( .A(n1337), .B(n13488), .Z(n13493) );
  XNOR U13120 ( .A(n13492), .B(n13486), .Z(n13488) );
  XOR U13121 ( .A(n13494), .B(n13495), .Z(n13486) );
  AND U13122 ( .A(n1352), .B(n13496), .Z(n13495) );
  XNOR U13123 ( .A(n13497), .B(n13498), .Z(n13492) );
  AND U13124 ( .A(n1344), .B(n13499), .Z(n13498) );
  XOR U13125 ( .A(p_input[1916]), .B(n13497), .Z(n13499) );
  XNOR U13126 ( .A(n13500), .B(n13501), .Z(n13497) );
  AND U13127 ( .A(n1348), .B(n13496), .Z(n13501) );
  XNOR U13128 ( .A(n13500), .B(n13494), .Z(n13496) );
  XOR U13129 ( .A(n13502), .B(n13503), .Z(n13494) );
  AND U13130 ( .A(n1363), .B(n13504), .Z(n13503) );
  XNOR U13131 ( .A(n13505), .B(n13506), .Z(n13500) );
  AND U13132 ( .A(n1355), .B(n13507), .Z(n13506) );
  XOR U13133 ( .A(p_input[1932]), .B(n13505), .Z(n13507) );
  XNOR U13134 ( .A(n13508), .B(n13509), .Z(n13505) );
  AND U13135 ( .A(n1359), .B(n13504), .Z(n13509) );
  XNOR U13136 ( .A(n13508), .B(n13502), .Z(n13504) );
  XOR U13137 ( .A(n13510), .B(n13511), .Z(n13502) );
  AND U13138 ( .A(n1374), .B(n13512), .Z(n13511) );
  XNOR U13139 ( .A(n13513), .B(n13514), .Z(n13508) );
  AND U13140 ( .A(n1366), .B(n13515), .Z(n13514) );
  XOR U13141 ( .A(p_input[1948]), .B(n13513), .Z(n13515) );
  XNOR U13142 ( .A(n13516), .B(n13517), .Z(n13513) );
  AND U13143 ( .A(n1370), .B(n13512), .Z(n13517) );
  XNOR U13144 ( .A(n13516), .B(n13510), .Z(n13512) );
  XOR U13145 ( .A(n13518), .B(n13519), .Z(n13510) );
  AND U13146 ( .A(n1385), .B(n13520), .Z(n13519) );
  XNOR U13147 ( .A(n13521), .B(n13522), .Z(n13516) );
  AND U13148 ( .A(n1377), .B(n13523), .Z(n13522) );
  XOR U13149 ( .A(p_input[1964]), .B(n13521), .Z(n13523) );
  XNOR U13150 ( .A(n13524), .B(n13525), .Z(n13521) );
  AND U13151 ( .A(n1381), .B(n13520), .Z(n13525) );
  XNOR U13152 ( .A(n13524), .B(n13518), .Z(n13520) );
  XOR U13153 ( .A(n13526), .B(n13527), .Z(n13518) );
  AND U13154 ( .A(n1396), .B(n13528), .Z(n13527) );
  XNOR U13155 ( .A(n13529), .B(n13530), .Z(n13524) );
  AND U13156 ( .A(n1388), .B(n13531), .Z(n13530) );
  XOR U13157 ( .A(p_input[1980]), .B(n13529), .Z(n13531) );
  XNOR U13158 ( .A(n13532), .B(n13533), .Z(n13529) );
  AND U13159 ( .A(n1392), .B(n13528), .Z(n13533) );
  XNOR U13160 ( .A(n13532), .B(n13526), .Z(n13528) );
  XOR U13161 ( .A(n13534), .B(n13535), .Z(n13526) );
  AND U13162 ( .A(n1407), .B(n13536), .Z(n13535) );
  XNOR U13163 ( .A(n13537), .B(n13538), .Z(n13532) );
  AND U13164 ( .A(n1399), .B(n13539), .Z(n13538) );
  XOR U13165 ( .A(p_input[1996]), .B(n13537), .Z(n13539) );
  XNOR U13166 ( .A(n13540), .B(n13541), .Z(n13537) );
  AND U13167 ( .A(n1403), .B(n13536), .Z(n13541) );
  XNOR U13168 ( .A(n13540), .B(n13534), .Z(n13536) );
  XOR U13169 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n13542), .Z(n13534) );
  AND U13170 ( .A(n1417), .B(n13543), .Z(n13542) );
  XNOR U13171 ( .A(n13544), .B(n13545), .Z(n13540) );
  AND U13172 ( .A(n1410), .B(n13546), .Z(n13545) );
  XOR U13173 ( .A(p_input[2012]), .B(n13544), .Z(n13546) );
  XNOR U13174 ( .A(n13547), .B(n13548), .Z(n13544) );
  AND U13175 ( .A(n1414), .B(n13543), .Z(n13548) );
  XOR U13176 ( .A(\knn_comb_/min_val_out[0][12] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n13543) );
  XOR U13177 ( .A(n25), .B(n13549), .Z(o[11]) );
  AND U13178 ( .A(n30), .B(n13550), .Z(n25) );
  XOR U13179 ( .A(n26), .B(n13549), .Z(n13550) );
  XOR U13180 ( .A(n13551), .B(n13552), .Z(n13549) );
  AND U13181 ( .A(n42), .B(n13553), .Z(n13552) );
  XOR U13182 ( .A(n13554), .B(n13555), .Z(n26) );
  AND U13183 ( .A(n34), .B(n13556), .Z(n13555) );
  XOR U13184 ( .A(p_input[11]), .B(n13554), .Z(n13556) );
  XNOR U13185 ( .A(n13557), .B(n13558), .Z(n13554) );
  AND U13186 ( .A(n38), .B(n13553), .Z(n13558) );
  XNOR U13187 ( .A(n13557), .B(n13551), .Z(n13553) );
  XOR U13188 ( .A(n13559), .B(n13560), .Z(n13551) );
  AND U13189 ( .A(n54), .B(n13561), .Z(n13560) );
  XNOR U13190 ( .A(n13562), .B(n13563), .Z(n13557) );
  AND U13191 ( .A(n46), .B(n13564), .Z(n13563) );
  XOR U13192 ( .A(p_input[27]), .B(n13562), .Z(n13564) );
  XNOR U13193 ( .A(n13565), .B(n13566), .Z(n13562) );
  AND U13194 ( .A(n50), .B(n13561), .Z(n13566) );
  XNOR U13195 ( .A(n13565), .B(n13559), .Z(n13561) );
  XOR U13196 ( .A(n13567), .B(n13568), .Z(n13559) );
  AND U13197 ( .A(n65), .B(n13569), .Z(n13568) );
  XNOR U13198 ( .A(n13570), .B(n13571), .Z(n13565) );
  AND U13199 ( .A(n57), .B(n13572), .Z(n13571) );
  XOR U13200 ( .A(p_input[43]), .B(n13570), .Z(n13572) );
  XNOR U13201 ( .A(n13573), .B(n13574), .Z(n13570) );
  AND U13202 ( .A(n61), .B(n13569), .Z(n13574) );
  XNOR U13203 ( .A(n13573), .B(n13567), .Z(n13569) );
  XOR U13204 ( .A(n13575), .B(n13576), .Z(n13567) );
  AND U13205 ( .A(n76), .B(n13577), .Z(n13576) );
  XNOR U13206 ( .A(n13578), .B(n13579), .Z(n13573) );
  AND U13207 ( .A(n68), .B(n13580), .Z(n13579) );
  XOR U13208 ( .A(p_input[59]), .B(n13578), .Z(n13580) );
  XNOR U13209 ( .A(n13581), .B(n13582), .Z(n13578) );
  AND U13210 ( .A(n72), .B(n13577), .Z(n13582) );
  XNOR U13211 ( .A(n13581), .B(n13575), .Z(n13577) );
  XOR U13212 ( .A(n13583), .B(n13584), .Z(n13575) );
  AND U13213 ( .A(n87), .B(n13585), .Z(n13584) );
  XNOR U13214 ( .A(n13586), .B(n13587), .Z(n13581) );
  AND U13215 ( .A(n79), .B(n13588), .Z(n13587) );
  XOR U13216 ( .A(p_input[75]), .B(n13586), .Z(n13588) );
  XNOR U13217 ( .A(n13589), .B(n13590), .Z(n13586) );
  AND U13218 ( .A(n83), .B(n13585), .Z(n13590) );
  XNOR U13219 ( .A(n13589), .B(n13583), .Z(n13585) );
  XOR U13220 ( .A(n13591), .B(n13592), .Z(n13583) );
  AND U13221 ( .A(n98), .B(n13593), .Z(n13592) );
  XNOR U13222 ( .A(n13594), .B(n13595), .Z(n13589) );
  AND U13223 ( .A(n90), .B(n13596), .Z(n13595) );
  XOR U13224 ( .A(p_input[91]), .B(n13594), .Z(n13596) );
  XNOR U13225 ( .A(n13597), .B(n13598), .Z(n13594) );
  AND U13226 ( .A(n94), .B(n13593), .Z(n13598) );
  XNOR U13227 ( .A(n13597), .B(n13591), .Z(n13593) );
  XOR U13228 ( .A(n13599), .B(n13600), .Z(n13591) );
  AND U13229 ( .A(n109), .B(n13601), .Z(n13600) );
  XNOR U13230 ( .A(n13602), .B(n13603), .Z(n13597) );
  AND U13231 ( .A(n101), .B(n13604), .Z(n13603) );
  XOR U13232 ( .A(p_input[107]), .B(n13602), .Z(n13604) );
  XNOR U13233 ( .A(n13605), .B(n13606), .Z(n13602) );
  AND U13234 ( .A(n105), .B(n13601), .Z(n13606) );
  XNOR U13235 ( .A(n13605), .B(n13599), .Z(n13601) );
  XOR U13236 ( .A(n13607), .B(n13608), .Z(n13599) );
  AND U13237 ( .A(n120), .B(n13609), .Z(n13608) );
  XNOR U13238 ( .A(n13610), .B(n13611), .Z(n13605) );
  AND U13239 ( .A(n112), .B(n13612), .Z(n13611) );
  XOR U13240 ( .A(p_input[123]), .B(n13610), .Z(n13612) );
  XNOR U13241 ( .A(n13613), .B(n13614), .Z(n13610) );
  AND U13242 ( .A(n116), .B(n13609), .Z(n13614) );
  XNOR U13243 ( .A(n13613), .B(n13607), .Z(n13609) );
  XOR U13244 ( .A(n13615), .B(n13616), .Z(n13607) );
  AND U13245 ( .A(n131), .B(n13617), .Z(n13616) );
  XNOR U13246 ( .A(n13618), .B(n13619), .Z(n13613) );
  AND U13247 ( .A(n123), .B(n13620), .Z(n13619) );
  XOR U13248 ( .A(p_input[139]), .B(n13618), .Z(n13620) );
  XNOR U13249 ( .A(n13621), .B(n13622), .Z(n13618) );
  AND U13250 ( .A(n127), .B(n13617), .Z(n13622) );
  XNOR U13251 ( .A(n13621), .B(n13615), .Z(n13617) );
  XOR U13252 ( .A(n13623), .B(n13624), .Z(n13615) );
  AND U13253 ( .A(n142), .B(n13625), .Z(n13624) );
  XNOR U13254 ( .A(n13626), .B(n13627), .Z(n13621) );
  AND U13255 ( .A(n134), .B(n13628), .Z(n13627) );
  XOR U13256 ( .A(p_input[155]), .B(n13626), .Z(n13628) );
  XNOR U13257 ( .A(n13629), .B(n13630), .Z(n13626) );
  AND U13258 ( .A(n138), .B(n13625), .Z(n13630) );
  XNOR U13259 ( .A(n13629), .B(n13623), .Z(n13625) );
  XOR U13260 ( .A(n13631), .B(n13632), .Z(n13623) );
  AND U13261 ( .A(n153), .B(n13633), .Z(n13632) );
  XNOR U13262 ( .A(n13634), .B(n13635), .Z(n13629) );
  AND U13263 ( .A(n145), .B(n13636), .Z(n13635) );
  XOR U13264 ( .A(p_input[171]), .B(n13634), .Z(n13636) );
  XNOR U13265 ( .A(n13637), .B(n13638), .Z(n13634) );
  AND U13266 ( .A(n149), .B(n13633), .Z(n13638) );
  XNOR U13267 ( .A(n13637), .B(n13631), .Z(n13633) );
  XOR U13268 ( .A(n13639), .B(n13640), .Z(n13631) );
  AND U13269 ( .A(n164), .B(n13641), .Z(n13640) );
  XNOR U13270 ( .A(n13642), .B(n13643), .Z(n13637) );
  AND U13271 ( .A(n156), .B(n13644), .Z(n13643) );
  XOR U13272 ( .A(p_input[187]), .B(n13642), .Z(n13644) );
  XNOR U13273 ( .A(n13645), .B(n13646), .Z(n13642) );
  AND U13274 ( .A(n160), .B(n13641), .Z(n13646) );
  XNOR U13275 ( .A(n13645), .B(n13639), .Z(n13641) );
  XOR U13276 ( .A(n13647), .B(n13648), .Z(n13639) );
  AND U13277 ( .A(n175), .B(n13649), .Z(n13648) );
  XNOR U13278 ( .A(n13650), .B(n13651), .Z(n13645) );
  AND U13279 ( .A(n167), .B(n13652), .Z(n13651) );
  XOR U13280 ( .A(p_input[203]), .B(n13650), .Z(n13652) );
  XNOR U13281 ( .A(n13653), .B(n13654), .Z(n13650) );
  AND U13282 ( .A(n171), .B(n13649), .Z(n13654) );
  XNOR U13283 ( .A(n13653), .B(n13647), .Z(n13649) );
  XOR U13284 ( .A(n13655), .B(n13656), .Z(n13647) );
  AND U13285 ( .A(n186), .B(n13657), .Z(n13656) );
  XNOR U13286 ( .A(n13658), .B(n13659), .Z(n13653) );
  AND U13287 ( .A(n178), .B(n13660), .Z(n13659) );
  XOR U13288 ( .A(p_input[219]), .B(n13658), .Z(n13660) );
  XNOR U13289 ( .A(n13661), .B(n13662), .Z(n13658) );
  AND U13290 ( .A(n182), .B(n13657), .Z(n13662) );
  XNOR U13291 ( .A(n13661), .B(n13655), .Z(n13657) );
  XOR U13292 ( .A(n13663), .B(n13664), .Z(n13655) );
  AND U13293 ( .A(n197), .B(n13665), .Z(n13664) );
  XNOR U13294 ( .A(n13666), .B(n13667), .Z(n13661) );
  AND U13295 ( .A(n189), .B(n13668), .Z(n13667) );
  XOR U13296 ( .A(p_input[235]), .B(n13666), .Z(n13668) );
  XNOR U13297 ( .A(n13669), .B(n13670), .Z(n13666) );
  AND U13298 ( .A(n193), .B(n13665), .Z(n13670) );
  XNOR U13299 ( .A(n13669), .B(n13663), .Z(n13665) );
  XOR U13300 ( .A(n13671), .B(n13672), .Z(n13663) );
  AND U13301 ( .A(n208), .B(n13673), .Z(n13672) );
  XNOR U13302 ( .A(n13674), .B(n13675), .Z(n13669) );
  AND U13303 ( .A(n200), .B(n13676), .Z(n13675) );
  XOR U13304 ( .A(p_input[251]), .B(n13674), .Z(n13676) );
  XNOR U13305 ( .A(n13677), .B(n13678), .Z(n13674) );
  AND U13306 ( .A(n204), .B(n13673), .Z(n13678) );
  XNOR U13307 ( .A(n13677), .B(n13671), .Z(n13673) );
  XOR U13308 ( .A(n13679), .B(n13680), .Z(n13671) );
  AND U13309 ( .A(n219), .B(n13681), .Z(n13680) );
  XNOR U13310 ( .A(n13682), .B(n13683), .Z(n13677) );
  AND U13311 ( .A(n211), .B(n13684), .Z(n13683) );
  XOR U13312 ( .A(p_input[267]), .B(n13682), .Z(n13684) );
  XNOR U13313 ( .A(n13685), .B(n13686), .Z(n13682) );
  AND U13314 ( .A(n215), .B(n13681), .Z(n13686) );
  XNOR U13315 ( .A(n13685), .B(n13679), .Z(n13681) );
  XOR U13316 ( .A(n13687), .B(n13688), .Z(n13679) );
  AND U13317 ( .A(n230), .B(n13689), .Z(n13688) );
  XNOR U13318 ( .A(n13690), .B(n13691), .Z(n13685) );
  AND U13319 ( .A(n222), .B(n13692), .Z(n13691) );
  XOR U13320 ( .A(p_input[283]), .B(n13690), .Z(n13692) );
  XNOR U13321 ( .A(n13693), .B(n13694), .Z(n13690) );
  AND U13322 ( .A(n226), .B(n13689), .Z(n13694) );
  XNOR U13323 ( .A(n13693), .B(n13687), .Z(n13689) );
  XOR U13324 ( .A(n13695), .B(n13696), .Z(n13687) );
  AND U13325 ( .A(n241), .B(n13697), .Z(n13696) );
  XNOR U13326 ( .A(n13698), .B(n13699), .Z(n13693) );
  AND U13327 ( .A(n233), .B(n13700), .Z(n13699) );
  XOR U13328 ( .A(p_input[299]), .B(n13698), .Z(n13700) );
  XNOR U13329 ( .A(n13701), .B(n13702), .Z(n13698) );
  AND U13330 ( .A(n237), .B(n13697), .Z(n13702) );
  XNOR U13331 ( .A(n13701), .B(n13695), .Z(n13697) );
  XOR U13332 ( .A(n13703), .B(n13704), .Z(n13695) );
  AND U13333 ( .A(n252), .B(n13705), .Z(n13704) );
  XNOR U13334 ( .A(n13706), .B(n13707), .Z(n13701) );
  AND U13335 ( .A(n244), .B(n13708), .Z(n13707) );
  XOR U13336 ( .A(p_input[315]), .B(n13706), .Z(n13708) );
  XNOR U13337 ( .A(n13709), .B(n13710), .Z(n13706) );
  AND U13338 ( .A(n248), .B(n13705), .Z(n13710) );
  XNOR U13339 ( .A(n13709), .B(n13703), .Z(n13705) );
  XOR U13340 ( .A(n13711), .B(n13712), .Z(n13703) );
  AND U13341 ( .A(n263), .B(n13713), .Z(n13712) );
  XNOR U13342 ( .A(n13714), .B(n13715), .Z(n13709) );
  AND U13343 ( .A(n255), .B(n13716), .Z(n13715) );
  XOR U13344 ( .A(p_input[331]), .B(n13714), .Z(n13716) );
  XNOR U13345 ( .A(n13717), .B(n13718), .Z(n13714) );
  AND U13346 ( .A(n259), .B(n13713), .Z(n13718) );
  XNOR U13347 ( .A(n13717), .B(n13711), .Z(n13713) );
  XOR U13348 ( .A(n13719), .B(n13720), .Z(n13711) );
  AND U13349 ( .A(n274), .B(n13721), .Z(n13720) );
  XNOR U13350 ( .A(n13722), .B(n13723), .Z(n13717) );
  AND U13351 ( .A(n266), .B(n13724), .Z(n13723) );
  XOR U13352 ( .A(p_input[347]), .B(n13722), .Z(n13724) );
  XNOR U13353 ( .A(n13725), .B(n13726), .Z(n13722) );
  AND U13354 ( .A(n270), .B(n13721), .Z(n13726) );
  XNOR U13355 ( .A(n13725), .B(n13719), .Z(n13721) );
  XOR U13356 ( .A(n13727), .B(n13728), .Z(n13719) );
  AND U13357 ( .A(n285), .B(n13729), .Z(n13728) );
  XNOR U13358 ( .A(n13730), .B(n13731), .Z(n13725) );
  AND U13359 ( .A(n277), .B(n13732), .Z(n13731) );
  XOR U13360 ( .A(p_input[363]), .B(n13730), .Z(n13732) );
  XNOR U13361 ( .A(n13733), .B(n13734), .Z(n13730) );
  AND U13362 ( .A(n281), .B(n13729), .Z(n13734) );
  XNOR U13363 ( .A(n13733), .B(n13727), .Z(n13729) );
  XOR U13364 ( .A(n13735), .B(n13736), .Z(n13727) );
  AND U13365 ( .A(n296), .B(n13737), .Z(n13736) );
  XNOR U13366 ( .A(n13738), .B(n13739), .Z(n13733) );
  AND U13367 ( .A(n288), .B(n13740), .Z(n13739) );
  XOR U13368 ( .A(p_input[379]), .B(n13738), .Z(n13740) );
  XNOR U13369 ( .A(n13741), .B(n13742), .Z(n13738) );
  AND U13370 ( .A(n292), .B(n13737), .Z(n13742) );
  XNOR U13371 ( .A(n13741), .B(n13735), .Z(n13737) );
  XOR U13372 ( .A(n13743), .B(n13744), .Z(n13735) );
  AND U13373 ( .A(n307), .B(n13745), .Z(n13744) );
  XNOR U13374 ( .A(n13746), .B(n13747), .Z(n13741) );
  AND U13375 ( .A(n299), .B(n13748), .Z(n13747) );
  XOR U13376 ( .A(p_input[395]), .B(n13746), .Z(n13748) );
  XNOR U13377 ( .A(n13749), .B(n13750), .Z(n13746) );
  AND U13378 ( .A(n303), .B(n13745), .Z(n13750) );
  XNOR U13379 ( .A(n13749), .B(n13743), .Z(n13745) );
  XOR U13380 ( .A(n13751), .B(n13752), .Z(n13743) );
  AND U13381 ( .A(n318), .B(n13753), .Z(n13752) );
  XNOR U13382 ( .A(n13754), .B(n13755), .Z(n13749) );
  AND U13383 ( .A(n310), .B(n13756), .Z(n13755) );
  XOR U13384 ( .A(p_input[411]), .B(n13754), .Z(n13756) );
  XNOR U13385 ( .A(n13757), .B(n13758), .Z(n13754) );
  AND U13386 ( .A(n314), .B(n13753), .Z(n13758) );
  XNOR U13387 ( .A(n13757), .B(n13751), .Z(n13753) );
  XOR U13388 ( .A(n13759), .B(n13760), .Z(n13751) );
  AND U13389 ( .A(n329), .B(n13761), .Z(n13760) );
  XNOR U13390 ( .A(n13762), .B(n13763), .Z(n13757) );
  AND U13391 ( .A(n321), .B(n13764), .Z(n13763) );
  XOR U13392 ( .A(p_input[427]), .B(n13762), .Z(n13764) );
  XNOR U13393 ( .A(n13765), .B(n13766), .Z(n13762) );
  AND U13394 ( .A(n325), .B(n13761), .Z(n13766) );
  XNOR U13395 ( .A(n13765), .B(n13759), .Z(n13761) );
  XOR U13396 ( .A(n13767), .B(n13768), .Z(n13759) );
  AND U13397 ( .A(n340), .B(n13769), .Z(n13768) );
  XNOR U13398 ( .A(n13770), .B(n13771), .Z(n13765) );
  AND U13399 ( .A(n332), .B(n13772), .Z(n13771) );
  XOR U13400 ( .A(p_input[443]), .B(n13770), .Z(n13772) );
  XNOR U13401 ( .A(n13773), .B(n13774), .Z(n13770) );
  AND U13402 ( .A(n336), .B(n13769), .Z(n13774) );
  XNOR U13403 ( .A(n13773), .B(n13767), .Z(n13769) );
  XOR U13404 ( .A(n13775), .B(n13776), .Z(n13767) );
  AND U13405 ( .A(n351), .B(n13777), .Z(n13776) );
  XNOR U13406 ( .A(n13778), .B(n13779), .Z(n13773) );
  AND U13407 ( .A(n343), .B(n13780), .Z(n13779) );
  XOR U13408 ( .A(p_input[459]), .B(n13778), .Z(n13780) );
  XNOR U13409 ( .A(n13781), .B(n13782), .Z(n13778) );
  AND U13410 ( .A(n347), .B(n13777), .Z(n13782) );
  XNOR U13411 ( .A(n13781), .B(n13775), .Z(n13777) );
  XOR U13412 ( .A(n13783), .B(n13784), .Z(n13775) );
  AND U13413 ( .A(n362), .B(n13785), .Z(n13784) );
  XNOR U13414 ( .A(n13786), .B(n13787), .Z(n13781) );
  AND U13415 ( .A(n354), .B(n13788), .Z(n13787) );
  XOR U13416 ( .A(p_input[475]), .B(n13786), .Z(n13788) );
  XNOR U13417 ( .A(n13789), .B(n13790), .Z(n13786) );
  AND U13418 ( .A(n358), .B(n13785), .Z(n13790) );
  XNOR U13419 ( .A(n13789), .B(n13783), .Z(n13785) );
  XOR U13420 ( .A(n13791), .B(n13792), .Z(n13783) );
  AND U13421 ( .A(n373), .B(n13793), .Z(n13792) );
  XNOR U13422 ( .A(n13794), .B(n13795), .Z(n13789) );
  AND U13423 ( .A(n365), .B(n13796), .Z(n13795) );
  XOR U13424 ( .A(p_input[491]), .B(n13794), .Z(n13796) );
  XNOR U13425 ( .A(n13797), .B(n13798), .Z(n13794) );
  AND U13426 ( .A(n369), .B(n13793), .Z(n13798) );
  XNOR U13427 ( .A(n13797), .B(n13791), .Z(n13793) );
  XOR U13428 ( .A(n13799), .B(n13800), .Z(n13791) );
  AND U13429 ( .A(n384), .B(n13801), .Z(n13800) );
  XNOR U13430 ( .A(n13802), .B(n13803), .Z(n13797) );
  AND U13431 ( .A(n376), .B(n13804), .Z(n13803) );
  XOR U13432 ( .A(p_input[507]), .B(n13802), .Z(n13804) );
  XNOR U13433 ( .A(n13805), .B(n13806), .Z(n13802) );
  AND U13434 ( .A(n380), .B(n13801), .Z(n13806) );
  XNOR U13435 ( .A(n13805), .B(n13799), .Z(n13801) );
  XOR U13436 ( .A(n13807), .B(n13808), .Z(n13799) );
  AND U13437 ( .A(n395), .B(n13809), .Z(n13808) );
  XNOR U13438 ( .A(n13810), .B(n13811), .Z(n13805) );
  AND U13439 ( .A(n387), .B(n13812), .Z(n13811) );
  XOR U13440 ( .A(p_input[523]), .B(n13810), .Z(n13812) );
  XNOR U13441 ( .A(n13813), .B(n13814), .Z(n13810) );
  AND U13442 ( .A(n391), .B(n13809), .Z(n13814) );
  XNOR U13443 ( .A(n13813), .B(n13807), .Z(n13809) );
  XOR U13444 ( .A(n13815), .B(n13816), .Z(n13807) );
  AND U13445 ( .A(n406), .B(n13817), .Z(n13816) );
  XNOR U13446 ( .A(n13818), .B(n13819), .Z(n13813) );
  AND U13447 ( .A(n398), .B(n13820), .Z(n13819) );
  XOR U13448 ( .A(p_input[539]), .B(n13818), .Z(n13820) );
  XNOR U13449 ( .A(n13821), .B(n13822), .Z(n13818) );
  AND U13450 ( .A(n402), .B(n13817), .Z(n13822) );
  XNOR U13451 ( .A(n13821), .B(n13815), .Z(n13817) );
  XOR U13452 ( .A(n13823), .B(n13824), .Z(n13815) );
  AND U13453 ( .A(n417), .B(n13825), .Z(n13824) );
  XNOR U13454 ( .A(n13826), .B(n13827), .Z(n13821) );
  AND U13455 ( .A(n409), .B(n13828), .Z(n13827) );
  XOR U13456 ( .A(p_input[555]), .B(n13826), .Z(n13828) );
  XNOR U13457 ( .A(n13829), .B(n13830), .Z(n13826) );
  AND U13458 ( .A(n413), .B(n13825), .Z(n13830) );
  XNOR U13459 ( .A(n13829), .B(n13823), .Z(n13825) );
  XOR U13460 ( .A(n13831), .B(n13832), .Z(n13823) );
  AND U13461 ( .A(n428), .B(n13833), .Z(n13832) );
  XNOR U13462 ( .A(n13834), .B(n13835), .Z(n13829) );
  AND U13463 ( .A(n420), .B(n13836), .Z(n13835) );
  XOR U13464 ( .A(p_input[571]), .B(n13834), .Z(n13836) );
  XNOR U13465 ( .A(n13837), .B(n13838), .Z(n13834) );
  AND U13466 ( .A(n424), .B(n13833), .Z(n13838) );
  XNOR U13467 ( .A(n13837), .B(n13831), .Z(n13833) );
  XOR U13468 ( .A(n13839), .B(n13840), .Z(n13831) );
  AND U13469 ( .A(n439), .B(n13841), .Z(n13840) );
  XNOR U13470 ( .A(n13842), .B(n13843), .Z(n13837) );
  AND U13471 ( .A(n431), .B(n13844), .Z(n13843) );
  XOR U13472 ( .A(p_input[587]), .B(n13842), .Z(n13844) );
  XNOR U13473 ( .A(n13845), .B(n13846), .Z(n13842) );
  AND U13474 ( .A(n435), .B(n13841), .Z(n13846) );
  XNOR U13475 ( .A(n13845), .B(n13839), .Z(n13841) );
  XOR U13476 ( .A(n13847), .B(n13848), .Z(n13839) );
  AND U13477 ( .A(n450), .B(n13849), .Z(n13848) );
  XNOR U13478 ( .A(n13850), .B(n13851), .Z(n13845) );
  AND U13479 ( .A(n442), .B(n13852), .Z(n13851) );
  XOR U13480 ( .A(p_input[603]), .B(n13850), .Z(n13852) );
  XNOR U13481 ( .A(n13853), .B(n13854), .Z(n13850) );
  AND U13482 ( .A(n446), .B(n13849), .Z(n13854) );
  XNOR U13483 ( .A(n13853), .B(n13847), .Z(n13849) );
  XOR U13484 ( .A(n13855), .B(n13856), .Z(n13847) );
  AND U13485 ( .A(n461), .B(n13857), .Z(n13856) );
  XNOR U13486 ( .A(n13858), .B(n13859), .Z(n13853) );
  AND U13487 ( .A(n453), .B(n13860), .Z(n13859) );
  XOR U13488 ( .A(p_input[619]), .B(n13858), .Z(n13860) );
  XNOR U13489 ( .A(n13861), .B(n13862), .Z(n13858) );
  AND U13490 ( .A(n457), .B(n13857), .Z(n13862) );
  XNOR U13491 ( .A(n13861), .B(n13855), .Z(n13857) );
  XOR U13492 ( .A(n13863), .B(n13864), .Z(n13855) );
  AND U13493 ( .A(n472), .B(n13865), .Z(n13864) );
  XNOR U13494 ( .A(n13866), .B(n13867), .Z(n13861) );
  AND U13495 ( .A(n464), .B(n13868), .Z(n13867) );
  XOR U13496 ( .A(p_input[635]), .B(n13866), .Z(n13868) );
  XNOR U13497 ( .A(n13869), .B(n13870), .Z(n13866) );
  AND U13498 ( .A(n468), .B(n13865), .Z(n13870) );
  XNOR U13499 ( .A(n13869), .B(n13863), .Z(n13865) );
  XOR U13500 ( .A(n13871), .B(n13872), .Z(n13863) );
  AND U13501 ( .A(n483), .B(n13873), .Z(n13872) );
  XNOR U13502 ( .A(n13874), .B(n13875), .Z(n13869) );
  AND U13503 ( .A(n475), .B(n13876), .Z(n13875) );
  XOR U13504 ( .A(p_input[651]), .B(n13874), .Z(n13876) );
  XNOR U13505 ( .A(n13877), .B(n13878), .Z(n13874) );
  AND U13506 ( .A(n479), .B(n13873), .Z(n13878) );
  XNOR U13507 ( .A(n13877), .B(n13871), .Z(n13873) );
  XOR U13508 ( .A(n13879), .B(n13880), .Z(n13871) );
  AND U13509 ( .A(n494), .B(n13881), .Z(n13880) );
  XNOR U13510 ( .A(n13882), .B(n13883), .Z(n13877) );
  AND U13511 ( .A(n486), .B(n13884), .Z(n13883) );
  XOR U13512 ( .A(p_input[667]), .B(n13882), .Z(n13884) );
  XNOR U13513 ( .A(n13885), .B(n13886), .Z(n13882) );
  AND U13514 ( .A(n490), .B(n13881), .Z(n13886) );
  XNOR U13515 ( .A(n13885), .B(n13879), .Z(n13881) );
  XOR U13516 ( .A(n13887), .B(n13888), .Z(n13879) );
  AND U13517 ( .A(n505), .B(n13889), .Z(n13888) );
  XNOR U13518 ( .A(n13890), .B(n13891), .Z(n13885) );
  AND U13519 ( .A(n497), .B(n13892), .Z(n13891) );
  XOR U13520 ( .A(p_input[683]), .B(n13890), .Z(n13892) );
  XNOR U13521 ( .A(n13893), .B(n13894), .Z(n13890) );
  AND U13522 ( .A(n501), .B(n13889), .Z(n13894) );
  XNOR U13523 ( .A(n13893), .B(n13887), .Z(n13889) );
  XOR U13524 ( .A(n13895), .B(n13896), .Z(n13887) );
  AND U13525 ( .A(n516), .B(n13897), .Z(n13896) );
  XNOR U13526 ( .A(n13898), .B(n13899), .Z(n13893) );
  AND U13527 ( .A(n508), .B(n13900), .Z(n13899) );
  XOR U13528 ( .A(p_input[699]), .B(n13898), .Z(n13900) );
  XNOR U13529 ( .A(n13901), .B(n13902), .Z(n13898) );
  AND U13530 ( .A(n512), .B(n13897), .Z(n13902) );
  XNOR U13531 ( .A(n13901), .B(n13895), .Z(n13897) );
  XOR U13532 ( .A(n13903), .B(n13904), .Z(n13895) );
  AND U13533 ( .A(n527), .B(n13905), .Z(n13904) );
  XNOR U13534 ( .A(n13906), .B(n13907), .Z(n13901) );
  AND U13535 ( .A(n519), .B(n13908), .Z(n13907) );
  XOR U13536 ( .A(p_input[715]), .B(n13906), .Z(n13908) );
  XNOR U13537 ( .A(n13909), .B(n13910), .Z(n13906) );
  AND U13538 ( .A(n523), .B(n13905), .Z(n13910) );
  XNOR U13539 ( .A(n13909), .B(n13903), .Z(n13905) );
  XOR U13540 ( .A(n13911), .B(n13912), .Z(n13903) );
  AND U13541 ( .A(n538), .B(n13913), .Z(n13912) );
  XNOR U13542 ( .A(n13914), .B(n13915), .Z(n13909) );
  AND U13543 ( .A(n530), .B(n13916), .Z(n13915) );
  XOR U13544 ( .A(p_input[731]), .B(n13914), .Z(n13916) );
  XNOR U13545 ( .A(n13917), .B(n13918), .Z(n13914) );
  AND U13546 ( .A(n534), .B(n13913), .Z(n13918) );
  XNOR U13547 ( .A(n13917), .B(n13911), .Z(n13913) );
  XOR U13548 ( .A(n13919), .B(n13920), .Z(n13911) );
  AND U13549 ( .A(n549), .B(n13921), .Z(n13920) );
  XNOR U13550 ( .A(n13922), .B(n13923), .Z(n13917) );
  AND U13551 ( .A(n541), .B(n13924), .Z(n13923) );
  XOR U13552 ( .A(p_input[747]), .B(n13922), .Z(n13924) );
  XNOR U13553 ( .A(n13925), .B(n13926), .Z(n13922) );
  AND U13554 ( .A(n545), .B(n13921), .Z(n13926) );
  XNOR U13555 ( .A(n13925), .B(n13919), .Z(n13921) );
  XOR U13556 ( .A(n13927), .B(n13928), .Z(n13919) );
  AND U13557 ( .A(n560), .B(n13929), .Z(n13928) );
  XNOR U13558 ( .A(n13930), .B(n13931), .Z(n13925) );
  AND U13559 ( .A(n552), .B(n13932), .Z(n13931) );
  XOR U13560 ( .A(p_input[763]), .B(n13930), .Z(n13932) );
  XNOR U13561 ( .A(n13933), .B(n13934), .Z(n13930) );
  AND U13562 ( .A(n556), .B(n13929), .Z(n13934) );
  XNOR U13563 ( .A(n13933), .B(n13927), .Z(n13929) );
  XOR U13564 ( .A(n13935), .B(n13936), .Z(n13927) );
  AND U13565 ( .A(n571), .B(n13937), .Z(n13936) );
  XNOR U13566 ( .A(n13938), .B(n13939), .Z(n13933) );
  AND U13567 ( .A(n563), .B(n13940), .Z(n13939) );
  XOR U13568 ( .A(p_input[779]), .B(n13938), .Z(n13940) );
  XNOR U13569 ( .A(n13941), .B(n13942), .Z(n13938) );
  AND U13570 ( .A(n567), .B(n13937), .Z(n13942) );
  XNOR U13571 ( .A(n13941), .B(n13935), .Z(n13937) );
  XOR U13572 ( .A(n13943), .B(n13944), .Z(n13935) );
  AND U13573 ( .A(n582), .B(n13945), .Z(n13944) );
  XNOR U13574 ( .A(n13946), .B(n13947), .Z(n13941) );
  AND U13575 ( .A(n574), .B(n13948), .Z(n13947) );
  XOR U13576 ( .A(p_input[795]), .B(n13946), .Z(n13948) );
  XNOR U13577 ( .A(n13949), .B(n13950), .Z(n13946) );
  AND U13578 ( .A(n578), .B(n13945), .Z(n13950) );
  XNOR U13579 ( .A(n13949), .B(n13943), .Z(n13945) );
  XOR U13580 ( .A(n13951), .B(n13952), .Z(n13943) );
  AND U13581 ( .A(n593), .B(n13953), .Z(n13952) );
  XNOR U13582 ( .A(n13954), .B(n13955), .Z(n13949) );
  AND U13583 ( .A(n585), .B(n13956), .Z(n13955) );
  XOR U13584 ( .A(p_input[811]), .B(n13954), .Z(n13956) );
  XNOR U13585 ( .A(n13957), .B(n13958), .Z(n13954) );
  AND U13586 ( .A(n589), .B(n13953), .Z(n13958) );
  XNOR U13587 ( .A(n13957), .B(n13951), .Z(n13953) );
  XOR U13588 ( .A(n13959), .B(n13960), .Z(n13951) );
  AND U13589 ( .A(n604), .B(n13961), .Z(n13960) );
  XNOR U13590 ( .A(n13962), .B(n13963), .Z(n13957) );
  AND U13591 ( .A(n596), .B(n13964), .Z(n13963) );
  XOR U13592 ( .A(p_input[827]), .B(n13962), .Z(n13964) );
  XNOR U13593 ( .A(n13965), .B(n13966), .Z(n13962) );
  AND U13594 ( .A(n600), .B(n13961), .Z(n13966) );
  XNOR U13595 ( .A(n13965), .B(n13959), .Z(n13961) );
  XOR U13596 ( .A(n13967), .B(n13968), .Z(n13959) );
  AND U13597 ( .A(n615), .B(n13969), .Z(n13968) );
  XNOR U13598 ( .A(n13970), .B(n13971), .Z(n13965) );
  AND U13599 ( .A(n607), .B(n13972), .Z(n13971) );
  XOR U13600 ( .A(p_input[843]), .B(n13970), .Z(n13972) );
  XNOR U13601 ( .A(n13973), .B(n13974), .Z(n13970) );
  AND U13602 ( .A(n611), .B(n13969), .Z(n13974) );
  XNOR U13603 ( .A(n13973), .B(n13967), .Z(n13969) );
  XOR U13604 ( .A(n13975), .B(n13976), .Z(n13967) );
  AND U13605 ( .A(n626), .B(n13977), .Z(n13976) );
  XNOR U13606 ( .A(n13978), .B(n13979), .Z(n13973) );
  AND U13607 ( .A(n618), .B(n13980), .Z(n13979) );
  XOR U13608 ( .A(p_input[859]), .B(n13978), .Z(n13980) );
  XNOR U13609 ( .A(n13981), .B(n13982), .Z(n13978) );
  AND U13610 ( .A(n622), .B(n13977), .Z(n13982) );
  XNOR U13611 ( .A(n13981), .B(n13975), .Z(n13977) );
  XOR U13612 ( .A(n13983), .B(n13984), .Z(n13975) );
  AND U13613 ( .A(n637), .B(n13985), .Z(n13984) );
  XNOR U13614 ( .A(n13986), .B(n13987), .Z(n13981) );
  AND U13615 ( .A(n629), .B(n13988), .Z(n13987) );
  XOR U13616 ( .A(p_input[875]), .B(n13986), .Z(n13988) );
  XNOR U13617 ( .A(n13989), .B(n13990), .Z(n13986) );
  AND U13618 ( .A(n633), .B(n13985), .Z(n13990) );
  XNOR U13619 ( .A(n13989), .B(n13983), .Z(n13985) );
  XOR U13620 ( .A(n13991), .B(n13992), .Z(n13983) );
  AND U13621 ( .A(n648), .B(n13993), .Z(n13992) );
  XNOR U13622 ( .A(n13994), .B(n13995), .Z(n13989) );
  AND U13623 ( .A(n640), .B(n13996), .Z(n13995) );
  XOR U13624 ( .A(p_input[891]), .B(n13994), .Z(n13996) );
  XNOR U13625 ( .A(n13997), .B(n13998), .Z(n13994) );
  AND U13626 ( .A(n644), .B(n13993), .Z(n13998) );
  XNOR U13627 ( .A(n13997), .B(n13991), .Z(n13993) );
  XOR U13628 ( .A(n13999), .B(n14000), .Z(n13991) );
  AND U13629 ( .A(n659), .B(n14001), .Z(n14000) );
  XNOR U13630 ( .A(n14002), .B(n14003), .Z(n13997) );
  AND U13631 ( .A(n651), .B(n14004), .Z(n14003) );
  XOR U13632 ( .A(p_input[907]), .B(n14002), .Z(n14004) );
  XNOR U13633 ( .A(n14005), .B(n14006), .Z(n14002) );
  AND U13634 ( .A(n655), .B(n14001), .Z(n14006) );
  XNOR U13635 ( .A(n14005), .B(n13999), .Z(n14001) );
  XOR U13636 ( .A(n14007), .B(n14008), .Z(n13999) );
  AND U13637 ( .A(n670), .B(n14009), .Z(n14008) );
  XNOR U13638 ( .A(n14010), .B(n14011), .Z(n14005) );
  AND U13639 ( .A(n662), .B(n14012), .Z(n14011) );
  XOR U13640 ( .A(p_input[923]), .B(n14010), .Z(n14012) );
  XNOR U13641 ( .A(n14013), .B(n14014), .Z(n14010) );
  AND U13642 ( .A(n666), .B(n14009), .Z(n14014) );
  XNOR U13643 ( .A(n14013), .B(n14007), .Z(n14009) );
  XOR U13644 ( .A(n14015), .B(n14016), .Z(n14007) );
  AND U13645 ( .A(n681), .B(n14017), .Z(n14016) );
  XNOR U13646 ( .A(n14018), .B(n14019), .Z(n14013) );
  AND U13647 ( .A(n673), .B(n14020), .Z(n14019) );
  XOR U13648 ( .A(p_input[939]), .B(n14018), .Z(n14020) );
  XNOR U13649 ( .A(n14021), .B(n14022), .Z(n14018) );
  AND U13650 ( .A(n677), .B(n14017), .Z(n14022) );
  XNOR U13651 ( .A(n14021), .B(n14015), .Z(n14017) );
  XOR U13652 ( .A(n14023), .B(n14024), .Z(n14015) );
  AND U13653 ( .A(n692), .B(n14025), .Z(n14024) );
  XNOR U13654 ( .A(n14026), .B(n14027), .Z(n14021) );
  AND U13655 ( .A(n684), .B(n14028), .Z(n14027) );
  XOR U13656 ( .A(p_input[955]), .B(n14026), .Z(n14028) );
  XNOR U13657 ( .A(n14029), .B(n14030), .Z(n14026) );
  AND U13658 ( .A(n688), .B(n14025), .Z(n14030) );
  XNOR U13659 ( .A(n14029), .B(n14023), .Z(n14025) );
  XOR U13660 ( .A(n14031), .B(n14032), .Z(n14023) );
  AND U13661 ( .A(n703), .B(n14033), .Z(n14032) );
  XNOR U13662 ( .A(n14034), .B(n14035), .Z(n14029) );
  AND U13663 ( .A(n695), .B(n14036), .Z(n14035) );
  XOR U13664 ( .A(p_input[971]), .B(n14034), .Z(n14036) );
  XNOR U13665 ( .A(n14037), .B(n14038), .Z(n14034) );
  AND U13666 ( .A(n699), .B(n14033), .Z(n14038) );
  XNOR U13667 ( .A(n14037), .B(n14031), .Z(n14033) );
  XOR U13668 ( .A(n14039), .B(n14040), .Z(n14031) );
  AND U13669 ( .A(n714), .B(n14041), .Z(n14040) );
  XNOR U13670 ( .A(n14042), .B(n14043), .Z(n14037) );
  AND U13671 ( .A(n706), .B(n14044), .Z(n14043) );
  XOR U13672 ( .A(p_input[987]), .B(n14042), .Z(n14044) );
  XNOR U13673 ( .A(n14045), .B(n14046), .Z(n14042) );
  AND U13674 ( .A(n710), .B(n14041), .Z(n14046) );
  XNOR U13675 ( .A(n14045), .B(n14039), .Z(n14041) );
  XOR U13676 ( .A(n14047), .B(n14048), .Z(n14039) );
  AND U13677 ( .A(n725), .B(n14049), .Z(n14048) );
  XNOR U13678 ( .A(n14050), .B(n14051), .Z(n14045) );
  AND U13679 ( .A(n717), .B(n14052), .Z(n14051) );
  XOR U13680 ( .A(p_input[1003]), .B(n14050), .Z(n14052) );
  XNOR U13681 ( .A(n14053), .B(n14054), .Z(n14050) );
  AND U13682 ( .A(n721), .B(n14049), .Z(n14054) );
  XNOR U13683 ( .A(n14053), .B(n14047), .Z(n14049) );
  XOR U13684 ( .A(n14055), .B(n14056), .Z(n14047) );
  AND U13685 ( .A(n736), .B(n14057), .Z(n14056) );
  XNOR U13686 ( .A(n14058), .B(n14059), .Z(n14053) );
  AND U13687 ( .A(n728), .B(n14060), .Z(n14059) );
  XOR U13688 ( .A(p_input[1019]), .B(n14058), .Z(n14060) );
  XNOR U13689 ( .A(n14061), .B(n14062), .Z(n14058) );
  AND U13690 ( .A(n732), .B(n14057), .Z(n14062) );
  XNOR U13691 ( .A(n14061), .B(n14055), .Z(n14057) );
  XOR U13692 ( .A(n14063), .B(n14064), .Z(n14055) );
  AND U13693 ( .A(n747), .B(n14065), .Z(n14064) );
  XNOR U13694 ( .A(n14066), .B(n14067), .Z(n14061) );
  AND U13695 ( .A(n739), .B(n14068), .Z(n14067) );
  XOR U13696 ( .A(p_input[1035]), .B(n14066), .Z(n14068) );
  XNOR U13697 ( .A(n14069), .B(n14070), .Z(n14066) );
  AND U13698 ( .A(n743), .B(n14065), .Z(n14070) );
  XNOR U13699 ( .A(n14069), .B(n14063), .Z(n14065) );
  XOR U13700 ( .A(n14071), .B(n14072), .Z(n14063) );
  AND U13701 ( .A(n758), .B(n14073), .Z(n14072) );
  XNOR U13702 ( .A(n14074), .B(n14075), .Z(n14069) );
  AND U13703 ( .A(n750), .B(n14076), .Z(n14075) );
  XOR U13704 ( .A(p_input[1051]), .B(n14074), .Z(n14076) );
  XNOR U13705 ( .A(n14077), .B(n14078), .Z(n14074) );
  AND U13706 ( .A(n754), .B(n14073), .Z(n14078) );
  XNOR U13707 ( .A(n14077), .B(n14071), .Z(n14073) );
  XOR U13708 ( .A(n14079), .B(n14080), .Z(n14071) );
  AND U13709 ( .A(n769), .B(n14081), .Z(n14080) );
  XNOR U13710 ( .A(n14082), .B(n14083), .Z(n14077) );
  AND U13711 ( .A(n761), .B(n14084), .Z(n14083) );
  XOR U13712 ( .A(p_input[1067]), .B(n14082), .Z(n14084) );
  XNOR U13713 ( .A(n14085), .B(n14086), .Z(n14082) );
  AND U13714 ( .A(n765), .B(n14081), .Z(n14086) );
  XNOR U13715 ( .A(n14085), .B(n14079), .Z(n14081) );
  XOR U13716 ( .A(n14087), .B(n14088), .Z(n14079) );
  AND U13717 ( .A(n780), .B(n14089), .Z(n14088) );
  XNOR U13718 ( .A(n14090), .B(n14091), .Z(n14085) );
  AND U13719 ( .A(n772), .B(n14092), .Z(n14091) );
  XOR U13720 ( .A(p_input[1083]), .B(n14090), .Z(n14092) );
  XNOR U13721 ( .A(n14093), .B(n14094), .Z(n14090) );
  AND U13722 ( .A(n776), .B(n14089), .Z(n14094) );
  XNOR U13723 ( .A(n14093), .B(n14087), .Z(n14089) );
  XOR U13724 ( .A(n14095), .B(n14096), .Z(n14087) );
  AND U13725 ( .A(n791), .B(n14097), .Z(n14096) );
  XNOR U13726 ( .A(n14098), .B(n14099), .Z(n14093) );
  AND U13727 ( .A(n783), .B(n14100), .Z(n14099) );
  XOR U13728 ( .A(p_input[1099]), .B(n14098), .Z(n14100) );
  XNOR U13729 ( .A(n14101), .B(n14102), .Z(n14098) );
  AND U13730 ( .A(n787), .B(n14097), .Z(n14102) );
  XNOR U13731 ( .A(n14101), .B(n14095), .Z(n14097) );
  XOR U13732 ( .A(n14103), .B(n14104), .Z(n14095) );
  AND U13733 ( .A(n802), .B(n14105), .Z(n14104) );
  XNOR U13734 ( .A(n14106), .B(n14107), .Z(n14101) );
  AND U13735 ( .A(n794), .B(n14108), .Z(n14107) );
  XOR U13736 ( .A(p_input[1115]), .B(n14106), .Z(n14108) );
  XNOR U13737 ( .A(n14109), .B(n14110), .Z(n14106) );
  AND U13738 ( .A(n798), .B(n14105), .Z(n14110) );
  XNOR U13739 ( .A(n14109), .B(n14103), .Z(n14105) );
  XOR U13740 ( .A(n14111), .B(n14112), .Z(n14103) );
  AND U13741 ( .A(n813), .B(n14113), .Z(n14112) );
  XNOR U13742 ( .A(n14114), .B(n14115), .Z(n14109) );
  AND U13743 ( .A(n805), .B(n14116), .Z(n14115) );
  XOR U13744 ( .A(p_input[1131]), .B(n14114), .Z(n14116) );
  XNOR U13745 ( .A(n14117), .B(n14118), .Z(n14114) );
  AND U13746 ( .A(n809), .B(n14113), .Z(n14118) );
  XNOR U13747 ( .A(n14117), .B(n14111), .Z(n14113) );
  XOR U13748 ( .A(n14119), .B(n14120), .Z(n14111) );
  AND U13749 ( .A(n824), .B(n14121), .Z(n14120) );
  XNOR U13750 ( .A(n14122), .B(n14123), .Z(n14117) );
  AND U13751 ( .A(n816), .B(n14124), .Z(n14123) );
  XOR U13752 ( .A(p_input[1147]), .B(n14122), .Z(n14124) );
  XNOR U13753 ( .A(n14125), .B(n14126), .Z(n14122) );
  AND U13754 ( .A(n820), .B(n14121), .Z(n14126) );
  XNOR U13755 ( .A(n14125), .B(n14119), .Z(n14121) );
  XOR U13756 ( .A(n14127), .B(n14128), .Z(n14119) );
  AND U13757 ( .A(n835), .B(n14129), .Z(n14128) );
  XNOR U13758 ( .A(n14130), .B(n14131), .Z(n14125) );
  AND U13759 ( .A(n827), .B(n14132), .Z(n14131) );
  XOR U13760 ( .A(p_input[1163]), .B(n14130), .Z(n14132) );
  XNOR U13761 ( .A(n14133), .B(n14134), .Z(n14130) );
  AND U13762 ( .A(n831), .B(n14129), .Z(n14134) );
  XNOR U13763 ( .A(n14133), .B(n14127), .Z(n14129) );
  XOR U13764 ( .A(n14135), .B(n14136), .Z(n14127) );
  AND U13765 ( .A(n846), .B(n14137), .Z(n14136) );
  XNOR U13766 ( .A(n14138), .B(n14139), .Z(n14133) );
  AND U13767 ( .A(n838), .B(n14140), .Z(n14139) );
  XOR U13768 ( .A(p_input[1179]), .B(n14138), .Z(n14140) );
  XNOR U13769 ( .A(n14141), .B(n14142), .Z(n14138) );
  AND U13770 ( .A(n842), .B(n14137), .Z(n14142) );
  XNOR U13771 ( .A(n14141), .B(n14135), .Z(n14137) );
  XOR U13772 ( .A(n14143), .B(n14144), .Z(n14135) );
  AND U13773 ( .A(n857), .B(n14145), .Z(n14144) );
  XNOR U13774 ( .A(n14146), .B(n14147), .Z(n14141) );
  AND U13775 ( .A(n849), .B(n14148), .Z(n14147) );
  XOR U13776 ( .A(p_input[1195]), .B(n14146), .Z(n14148) );
  XNOR U13777 ( .A(n14149), .B(n14150), .Z(n14146) );
  AND U13778 ( .A(n853), .B(n14145), .Z(n14150) );
  XNOR U13779 ( .A(n14149), .B(n14143), .Z(n14145) );
  XOR U13780 ( .A(n14151), .B(n14152), .Z(n14143) );
  AND U13781 ( .A(n868), .B(n14153), .Z(n14152) );
  XNOR U13782 ( .A(n14154), .B(n14155), .Z(n14149) );
  AND U13783 ( .A(n860), .B(n14156), .Z(n14155) );
  XOR U13784 ( .A(p_input[1211]), .B(n14154), .Z(n14156) );
  XNOR U13785 ( .A(n14157), .B(n14158), .Z(n14154) );
  AND U13786 ( .A(n864), .B(n14153), .Z(n14158) );
  XNOR U13787 ( .A(n14157), .B(n14151), .Z(n14153) );
  XOR U13788 ( .A(n14159), .B(n14160), .Z(n14151) );
  AND U13789 ( .A(n879), .B(n14161), .Z(n14160) );
  XNOR U13790 ( .A(n14162), .B(n14163), .Z(n14157) );
  AND U13791 ( .A(n871), .B(n14164), .Z(n14163) );
  XOR U13792 ( .A(p_input[1227]), .B(n14162), .Z(n14164) );
  XNOR U13793 ( .A(n14165), .B(n14166), .Z(n14162) );
  AND U13794 ( .A(n875), .B(n14161), .Z(n14166) );
  XNOR U13795 ( .A(n14165), .B(n14159), .Z(n14161) );
  XOR U13796 ( .A(n14167), .B(n14168), .Z(n14159) );
  AND U13797 ( .A(n890), .B(n14169), .Z(n14168) );
  XNOR U13798 ( .A(n14170), .B(n14171), .Z(n14165) );
  AND U13799 ( .A(n882), .B(n14172), .Z(n14171) );
  XOR U13800 ( .A(p_input[1243]), .B(n14170), .Z(n14172) );
  XNOR U13801 ( .A(n14173), .B(n14174), .Z(n14170) );
  AND U13802 ( .A(n886), .B(n14169), .Z(n14174) );
  XNOR U13803 ( .A(n14173), .B(n14167), .Z(n14169) );
  XOR U13804 ( .A(n14175), .B(n14176), .Z(n14167) );
  AND U13805 ( .A(n901), .B(n14177), .Z(n14176) );
  XNOR U13806 ( .A(n14178), .B(n14179), .Z(n14173) );
  AND U13807 ( .A(n893), .B(n14180), .Z(n14179) );
  XOR U13808 ( .A(p_input[1259]), .B(n14178), .Z(n14180) );
  XNOR U13809 ( .A(n14181), .B(n14182), .Z(n14178) );
  AND U13810 ( .A(n897), .B(n14177), .Z(n14182) );
  XNOR U13811 ( .A(n14181), .B(n14175), .Z(n14177) );
  XOR U13812 ( .A(n14183), .B(n14184), .Z(n14175) );
  AND U13813 ( .A(n912), .B(n14185), .Z(n14184) );
  XNOR U13814 ( .A(n14186), .B(n14187), .Z(n14181) );
  AND U13815 ( .A(n904), .B(n14188), .Z(n14187) );
  XOR U13816 ( .A(p_input[1275]), .B(n14186), .Z(n14188) );
  XNOR U13817 ( .A(n14189), .B(n14190), .Z(n14186) );
  AND U13818 ( .A(n908), .B(n14185), .Z(n14190) );
  XNOR U13819 ( .A(n14189), .B(n14183), .Z(n14185) );
  XOR U13820 ( .A(n14191), .B(n14192), .Z(n14183) );
  AND U13821 ( .A(n923), .B(n14193), .Z(n14192) );
  XNOR U13822 ( .A(n14194), .B(n14195), .Z(n14189) );
  AND U13823 ( .A(n915), .B(n14196), .Z(n14195) );
  XOR U13824 ( .A(p_input[1291]), .B(n14194), .Z(n14196) );
  XNOR U13825 ( .A(n14197), .B(n14198), .Z(n14194) );
  AND U13826 ( .A(n919), .B(n14193), .Z(n14198) );
  XNOR U13827 ( .A(n14197), .B(n14191), .Z(n14193) );
  XOR U13828 ( .A(n14199), .B(n14200), .Z(n14191) );
  AND U13829 ( .A(n934), .B(n14201), .Z(n14200) );
  XNOR U13830 ( .A(n14202), .B(n14203), .Z(n14197) );
  AND U13831 ( .A(n926), .B(n14204), .Z(n14203) );
  XOR U13832 ( .A(p_input[1307]), .B(n14202), .Z(n14204) );
  XNOR U13833 ( .A(n14205), .B(n14206), .Z(n14202) );
  AND U13834 ( .A(n930), .B(n14201), .Z(n14206) );
  XNOR U13835 ( .A(n14205), .B(n14199), .Z(n14201) );
  XOR U13836 ( .A(n14207), .B(n14208), .Z(n14199) );
  AND U13837 ( .A(n945), .B(n14209), .Z(n14208) );
  XNOR U13838 ( .A(n14210), .B(n14211), .Z(n14205) );
  AND U13839 ( .A(n937), .B(n14212), .Z(n14211) );
  XOR U13840 ( .A(p_input[1323]), .B(n14210), .Z(n14212) );
  XNOR U13841 ( .A(n14213), .B(n14214), .Z(n14210) );
  AND U13842 ( .A(n941), .B(n14209), .Z(n14214) );
  XNOR U13843 ( .A(n14213), .B(n14207), .Z(n14209) );
  XOR U13844 ( .A(n14215), .B(n14216), .Z(n14207) );
  AND U13845 ( .A(n956), .B(n14217), .Z(n14216) );
  XNOR U13846 ( .A(n14218), .B(n14219), .Z(n14213) );
  AND U13847 ( .A(n948), .B(n14220), .Z(n14219) );
  XOR U13848 ( .A(p_input[1339]), .B(n14218), .Z(n14220) );
  XNOR U13849 ( .A(n14221), .B(n14222), .Z(n14218) );
  AND U13850 ( .A(n952), .B(n14217), .Z(n14222) );
  XNOR U13851 ( .A(n14221), .B(n14215), .Z(n14217) );
  XOR U13852 ( .A(n14223), .B(n14224), .Z(n14215) );
  AND U13853 ( .A(n967), .B(n14225), .Z(n14224) );
  XNOR U13854 ( .A(n14226), .B(n14227), .Z(n14221) );
  AND U13855 ( .A(n959), .B(n14228), .Z(n14227) );
  XOR U13856 ( .A(p_input[1355]), .B(n14226), .Z(n14228) );
  XNOR U13857 ( .A(n14229), .B(n14230), .Z(n14226) );
  AND U13858 ( .A(n963), .B(n14225), .Z(n14230) );
  XNOR U13859 ( .A(n14229), .B(n14223), .Z(n14225) );
  XOR U13860 ( .A(n14231), .B(n14232), .Z(n14223) );
  AND U13861 ( .A(n978), .B(n14233), .Z(n14232) );
  XNOR U13862 ( .A(n14234), .B(n14235), .Z(n14229) );
  AND U13863 ( .A(n970), .B(n14236), .Z(n14235) );
  XOR U13864 ( .A(p_input[1371]), .B(n14234), .Z(n14236) );
  XNOR U13865 ( .A(n14237), .B(n14238), .Z(n14234) );
  AND U13866 ( .A(n974), .B(n14233), .Z(n14238) );
  XNOR U13867 ( .A(n14237), .B(n14231), .Z(n14233) );
  XOR U13868 ( .A(n14239), .B(n14240), .Z(n14231) );
  AND U13869 ( .A(n989), .B(n14241), .Z(n14240) );
  XNOR U13870 ( .A(n14242), .B(n14243), .Z(n14237) );
  AND U13871 ( .A(n981), .B(n14244), .Z(n14243) );
  XOR U13872 ( .A(p_input[1387]), .B(n14242), .Z(n14244) );
  XNOR U13873 ( .A(n14245), .B(n14246), .Z(n14242) );
  AND U13874 ( .A(n985), .B(n14241), .Z(n14246) );
  XNOR U13875 ( .A(n14245), .B(n14239), .Z(n14241) );
  XOR U13876 ( .A(n14247), .B(n14248), .Z(n14239) );
  AND U13877 ( .A(n1000), .B(n14249), .Z(n14248) );
  XNOR U13878 ( .A(n14250), .B(n14251), .Z(n14245) );
  AND U13879 ( .A(n992), .B(n14252), .Z(n14251) );
  XOR U13880 ( .A(p_input[1403]), .B(n14250), .Z(n14252) );
  XNOR U13881 ( .A(n14253), .B(n14254), .Z(n14250) );
  AND U13882 ( .A(n996), .B(n14249), .Z(n14254) );
  XNOR U13883 ( .A(n14253), .B(n14247), .Z(n14249) );
  XOR U13884 ( .A(n14255), .B(n14256), .Z(n14247) );
  AND U13885 ( .A(n1011), .B(n14257), .Z(n14256) );
  XNOR U13886 ( .A(n14258), .B(n14259), .Z(n14253) );
  AND U13887 ( .A(n1003), .B(n14260), .Z(n14259) );
  XOR U13888 ( .A(p_input[1419]), .B(n14258), .Z(n14260) );
  XNOR U13889 ( .A(n14261), .B(n14262), .Z(n14258) );
  AND U13890 ( .A(n1007), .B(n14257), .Z(n14262) );
  XNOR U13891 ( .A(n14261), .B(n14255), .Z(n14257) );
  XOR U13892 ( .A(n14263), .B(n14264), .Z(n14255) );
  AND U13893 ( .A(n1022), .B(n14265), .Z(n14264) );
  XNOR U13894 ( .A(n14266), .B(n14267), .Z(n14261) );
  AND U13895 ( .A(n1014), .B(n14268), .Z(n14267) );
  XOR U13896 ( .A(p_input[1435]), .B(n14266), .Z(n14268) );
  XNOR U13897 ( .A(n14269), .B(n14270), .Z(n14266) );
  AND U13898 ( .A(n1018), .B(n14265), .Z(n14270) );
  XNOR U13899 ( .A(n14269), .B(n14263), .Z(n14265) );
  XOR U13900 ( .A(n14271), .B(n14272), .Z(n14263) );
  AND U13901 ( .A(n1033), .B(n14273), .Z(n14272) );
  XNOR U13902 ( .A(n14274), .B(n14275), .Z(n14269) );
  AND U13903 ( .A(n1025), .B(n14276), .Z(n14275) );
  XOR U13904 ( .A(p_input[1451]), .B(n14274), .Z(n14276) );
  XNOR U13905 ( .A(n14277), .B(n14278), .Z(n14274) );
  AND U13906 ( .A(n1029), .B(n14273), .Z(n14278) );
  XNOR U13907 ( .A(n14277), .B(n14271), .Z(n14273) );
  XOR U13908 ( .A(n14279), .B(n14280), .Z(n14271) );
  AND U13909 ( .A(n1044), .B(n14281), .Z(n14280) );
  XNOR U13910 ( .A(n14282), .B(n14283), .Z(n14277) );
  AND U13911 ( .A(n1036), .B(n14284), .Z(n14283) );
  XOR U13912 ( .A(p_input[1467]), .B(n14282), .Z(n14284) );
  XNOR U13913 ( .A(n14285), .B(n14286), .Z(n14282) );
  AND U13914 ( .A(n1040), .B(n14281), .Z(n14286) );
  XNOR U13915 ( .A(n14285), .B(n14279), .Z(n14281) );
  XOR U13916 ( .A(n14287), .B(n14288), .Z(n14279) );
  AND U13917 ( .A(n1055), .B(n14289), .Z(n14288) );
  XNOR U13918 ( .A(n14290), .B(n14291), .Z(n14285) );
  AND U13919 ( .A(n1047), .B(n14292), .Z(n14291) );
  XOR U13920 ( .A(p_input[1483]), .B(n14290), .Z(n14292) );
  XNOR U13921 ( .A(n14293), .B(n14294), .Z(n14290) );
  AND U13922 ( .A(n1051), .B(n14289), .Z(n14294) );
  XNOR U13923 ( .A(n14293), .B(n14287), .Z(n14289) );
  XOR U13924 ( .A(n14295), .B(n14296), .Z(n14287) );
  AND U13925 ( .A(n1066), .B(n14297), .Z(n14296) );
  XNOR U13926 ( .A(n14298), .B(n14299), .Z(n14293) );
  AND U13927 ( .A(n1058), .B(n14300), .Z(n14299) );
  XOR U13928 ( .A(p_input[1499]), .B(n14298), .Z(n14300) );
  XNOR U13929 ( .A(n14301), .B(n14302), .Z(n14298) );
  AND U13930 ( .A(n1062), .B(n14297), .Z(n14302) );
  XNOR U13931 ( .A(n14301), .B(n14295), .Z(n14297) );
  XOR U13932 ( .A(n14303), .B(n14304), .Z(n14295) );
  AND U13933 ( .A(n1077), .B(n14305), .Z(n14304) );
  XNOR U13934 ( .A(n14306), .B(n14307), .Z(n14301) );
  AND U13935 ( .A(n1069), .B(n14308), .Z(n14307) );
  XOR U13936 ( .A(p_input[1515]), .B(n14306), .Z(n14308) );
  XNOR U13937 ( .A(n14309), .B(n14310), .Z(n14306) );
  AND U13938 ( .A(n1073), .B(n14305), .Z(n14310) );
  XNOR U13939 ( .A(n14309), .B(n14303), .Z(n14305) );
  XOR U13940 ( .A(n14311), .B(n14312), .Z(n14303) );
  AND U13941 ( .A(n1088), .B(n14313), .Z(n14312) );
  XNOR U13942 ( .A(n14314), .B(n14315), .Z(n14309) );
  AND U13943 ( .A(n1080), .B(n14316), .Z(n14315) );
  XOR U13944 ( .A(p_input[1531]), .B(n14314), .Z(n14316) );
  XNOR U13945 ( .A(n14317), .B(n14318), .Z(n14314) );
  AND U13946 ( .A(n1084), .B(n14313), .Z(n14318) );
  XNOR U13947 ( .A(n14317), .B(n14311), .Z(n14313) );
  XOR U13948 ( .A(n14319), .B(n14320), .Z(n14311) );
  AND U13949 ( .A(n1099), .B(n14321), .Z(n14320) );
  XNOR U13950 ( .A(n14322), .B(n14323), .Z(n14317) );
  AND U13951 ( .A(n1091), .B(n14324), .Z(n14323) );
  XOR U13952 ( .A(p_input[1547]), .B(n14322), .Z(n14324) );
  XNOR U13953 ( .A(n14325), .B(n14326), .Z(n14322) );
  AND U13954 ( .A(n1095), .B(n14321), .Z(n14326) );
  XNOR U13955 ( .A(n14325), .B(n14319), .Z(n14321) );
  XOR U13956 ( .A(n14327), .B(n14328), .Z(n14319) );
  AND U13957 ( .A(n1110), .B(n14329), .Z(n14328) );
  XNOR U13958 ( .A(n14330), .B(n14331), .Z(n14325) );
  AND U13959 ( .A(n1102), .B(n14332), .Z(n14331) );
  XOR U13960 ( .A(p_input[1563]), .B(n14330), .Z(n14332) );
  XNOR U13961 ( .A(n14333), .B(n14334), .Z(n14330) );
  AND U13962 ( .A(n1106), .B(n14329), .Z(n14334) );
  XNOR U13963 ( .A(n14333), .B(n14327), .Z(n14329) );
  XOR U13964 ( .A(n14335), .B(n14336), .Z(n14327) );
  AND U13965 ( .A(n1121), .B(n14337), .Z(n14336) );
  XNOR U13966 ( .A(n14338), .B(n14339), .Z(n14333) );
  AND U13967 ( .A(n1113), .B(n14340), .Z(n14339) );
  XOR U13968 ( .A(p_input[1579]), .B(n14338), .Z(n14340) );
  XNOR U13969 ( .A(n14341), .B(n14342), .Z(n14338) );
  AND U13970 ( .A(n1117), .B(n14337), .Z(n14342) );
  XNOR U13971 ( .A(n14341), .B(n14335), .Z(n14337) );
  XOR U13972 ( .A(n14343), .B(n14344), .Z(n14335) );
  AND U13973 ( .A(n1132), .B(n14345), .Z(n14344) );
  XNOR U13974 ( .A(n14346), .B(n14347), .Z(n14341) );
  AND U13975 ( .A(n1124), .B(n14348), .Z(n14347) );
  XOR U13976 ( .A(p_input[1595]), .B(n14346), .Z(n14348) );
  XNOR U13977 ( .A(n14349), .B(n14350), .Z(n14346) );
  AND U13978 ( .A(n1128), .B(n14345), .Z(n14350) );
  XNOR U13979 ( .A(n14349), .B(n14343), .Z(n14345) );
  XOR U13980 ( .A(n14351), .B(n14352), .Z(n14343) );
  AND U13981 ( .A(n1143), .B(n14353), .Z(n14352) );
  XNOR U13982 ( .A(n14354), .B(n14355), .Z(n14349) );
  AND U13983 ( .A(n1135), .B(n14356), .Z(n14355) );
  XOR U13984 ( .A(p_input[1611]), .B(n14354), .Z(n14356) );
  XNOR U13985 ( .A(n14357), .B(n14358), .Z(n14354) );
  AND U13986 ( .A(n1139), .B(n14353), .Z(n14358) );
  XNOR U13987 ( .A(n14357), .B(n14351), .Z(n14353) );
  XOR U13988 ( .A(n14359), .B(n14360), .Z(n14351) );
  AND U13989 ( .A(n1154), .B(n14361), .Z(n14360) );
  XNOR U13990 ( .A(n14362), .B(n14363), .Z(n14357) );
  AND U13991 ( .A(n1146), .B(n14364), .Z(n14363) );
  XOR U13992 ( .A(p_input[1627]), .B(n14362), .Z(n14364) );
  XNOR U13993 ( .A(n14365), .B(n14366), .Z(n14362) );
  AND U13994 ( .A(n1150), .B(n14361), .Z(n14366) );
  XNOR U13995 ( .A(n14365), .B(n14359), .Z(n14361) );
  XOR U13996 ( .A(n14367), .B(n14368), .Z(n14359) );
  AND U13997 ( .A(n1165), .B(n14369), .Z(n14368) );
  XNOR U13998 ( .A(n14370), .B(n14371), .Z(n14365) );
  AND U13999 ( .A(n1157), .B(n14372), .Z(n14371) );
  XOR U14000 ( .A(p_input[1643]), .B(n14370), .Z(n14372) );
  XNOR U14001 ( .A(n14373), .B(n14374), .Z(n14370) );
  AND U14002 ( .A(n1161), .B(n14369), .Z(n14374) );
  XNOR U14003 ( .A(n14373), .B(n14367), .Z(n14369) );
  XOR U14004 ( .A(n14375), .B(n14376), .Z(n14367) );
  AND U14005 ( .A(n1176), .B(n14377), .Z(n14376) );
  XNOR U14006 ( .A(n14378), .B(n14379), .Z(n14373) );
  AND U14007 ( .A(n1168), .B(n14380), .Z(n14379) );
  XOR U14008 ( .A(p_input[1659]), .B(n14378), .Z(n14380) );
  XNOR U14009 ( .A(n14381), .B(n14382), .Z(n14378) );
  AND U14010 ( .A(n1172), .B(n14377), .Z(n14382) );
  XNOR U14011 ( .A(n14381), .B(n14375), .Z(n14377) );
  XOR U14012 ( .A(n14383), .B(n14384), .Z(n14375) );
  AND U14013 ( .A(n1187), .B(n14385), .Z(n14384) );
  XNOR U14014 ( .A(n14386), .B(n14387), .Z(n14381) );
  AND U14015 ( .A(n1179), .B(n14388), .Z(n14387) );
  XOR U14016 ( .A(p_input[1675]), .B(n14386), .Z(n14388) );
  XNOR U14017 ( .A(n14389), .B(n14390), .Z(n14386) );
  AND U14018 ( .A(n1183), .B(n14385), .Z(n14390) );
  XNOR U14019 ( .A(n14389), .B(n14383), .Z(n14385) );
  XOR U14020 ( .A(n14391), .B(n14392), .Z(n14383) );
  AND U14021 ( .A(n1198), .B(n14393), .Z(n14392) );
  XNOR U14022 ( .A(n14394), .B(n14395), .Z(n14389) );
  AND U14023 ( .A(n1190), .B(n14396), .Z(n14395) );
  XOR U14024 ( .A(p_input[1691]), .B(n14394), .Z(n14396) );
  XNOR U14025 ( .A(n14397), .B(n14398), .Z(n14394) );
  AND U14026 ( .A(n1194), .B(n14393), .Z(n14398) );
  XNOR U14027 ( .A(n14397), .B(n14391), .Z(n14393) );
  XOR U14028 ( .A(n14399), .B(n14400), .Z(n14391) );
  AND U14029 ( .A(n1209), .B(n14401), .Z(n14400) );
  XNOR U14030 ( .A(n14402), .B(n14403), .Z(n14397) );
  AND U14031 ( .A(n1201), .B(n14404), .Z(n14403) );
  XOR U14032 ( .A(p_input[1707]), .B(n14402), .Z(n14404) );
  XNOR U14033 ( .A(n14405), .B(n14406), .Z(n14402) );
  AND U14034 ( .A(n1205), .B(n14401), .Z(n14406) );
  XNOR U14035 ( .A(n14405), .B(n14399), .Z(n14401) );
  XOR U14036 ( .A(n14407), .B(n14408), .Z(n14399) );
  AND U14037 ( .A(n1220), .B(n14409), .Z(n14408) );
  XNOR U14038 ( .A(n14410), .B(n14411), .Z(n14405) );
  AND U14039 ( .A(n1212), .B(n14412), .Z(n14411) );
  XOR U14040 ( .A(p_input[1723]), .B(n14410), .Z(n14412) );
  XNOR U14041 ( .A(n14413), .B(n14414), .Z(n14410) );
  AND U14042 ( .A(n1216), .B(n14409), .Z(n14414) );
  XNOR U14043 ( .A(n14413), .B(n14407), .Z(n14409) );
  XOR U14044 ( .A(n14415), .B(n14416), .Z(n14407) );
  AND U14045 ( .A(n1231), .B(n14417), .Z(n14416) );
  XNOR U14046 ( .A(n14418), .B(n14419), .Z(n14413) );
  AND U14047 ( .A(n1223), .B(n14420), .Z(n14419) );
  XOR U14048 ( .A(p_input[1739]), .B(n14418), .Z(n14420) );
  XNOR U14049 ( .A(n14421), .B(n14422), .Z(n14418) );
  AND U14050 ( .A(n1227), .B(n14417), .Z(n14422) );
  XNOR U14051 ( .A(n14421), .B(n14415), .Z(n14417) );
  XOR U14052 ( .A(n14423), .B(n14424), .Z(n14415) );
  AND U14053 ( .A(n1242), .B(n14425), .Z(n14424) );
  XNOR U14054 ( .A(n14426), .B(n14427), .Z(n14421) );
  AND U14055 ( .A(n1234), .B(n14428), .Z(n14427) );
  XOR U14056 ( .A(p_input[1755]), .B(n14426), .Z(n14428) );
  XNOR U14057 ( .A(n14429), .B(n14430), .Z(n14426) );
  AND U14058 ( .A(n1238), .B(n14425), .Z(n14430) );
  XNOR U14059 ( .A(n14429), .B(n14423), .Z(n14425) );
  XOR U14060 ( .A(n14431), .B(n14432), .Z(n14423) );
  AND U14061 ( .A(n1253), .B(n14433), .Z(n14432) );
  XNOR U14062 ( .A(n14434), .B(n14435), .Z(n14429) );
  AND U14063 ( .A(n1245), .B(n14436), .Z(n14435) );
  XOR U14064 ( .A(p_input[1771]), .B(n14434), .Z(n14436) );
  XNOR U14065 ( .A(n14437), .B(n14438), .Z(n14434) );
  AND U14066 ( .A(n1249), .B(n14433), .Z(n14438) );
  XNOR U14067 ( .A(n14437), .B(n14431), .Z(n14433) );
  XOR U14068 ( .A(n14439), .B(n14440), .Z(n14431) );
  AND U14069 ( .A(n1264), .B(n14441), .Z(n14440) );
  XNOR U14070 ( .A(n14442), .B(n14443), .Z(n14437) );
  AND U14071 ( .A(n1256), .B(n14444), .Z(n14443) );
  XOR U14072 ( .A(p_input[1787]), .B(n14442), .Z(n14444) );
  XNOR U14073 ( .A(n14445), .B(n14446), .Z(n14442) );
  AND U14074 ( .A(n1260), .B(n14441), .Z(n14446) );
  XNOR U14075 ( .A(n14445), .B(n14439), .Z(n14441) );
  XOR U14076 ( .A(n14447), .B(n14448), .Z(n14439) );
  AND U14077 ( .A(n1275), .B(n14449), .Z(n14448) );
  XNOR U14078 ( .A(n14450), .B(n14451), .Z(n14445) );
  AND U14079 ( .A(n1267), .B(n14452), .Z(n14451) );
  XOR U14080 ( .A(p_input[1803]), .B(n14450), .Z(n14452) );
  XNOR U14081 ( .A(n14453), .B(n14454), .Z(n14450) );
  AND U14082 ( .A(n1271), .B(n14449), .Z(n14454) );
  XNOR U14083 ( .A(n14453), .B(n14447), .Z(n14449) );
  XOR U14084 ( .A(n14455), .B(n14456), .Z(n14447) );
  AND U14085 ( .A(n1286), .B(n14457), .Z(n14456) );
  XNOR U14086 ( .A(n14458), .B(n14459), .Z(n14453) );
  AND U14087 ( .A(n1278), .B(n14460), .Z(n14459) );
  XOR U14088 ( .A(p_input[1819]), .B(n14458), .Z(n14460) );
  XNOR U14089 ( .A(n14461), .B(n14462), .Z(n14458) );
  AND U14090 ( .A(n1282), .B(n14457), .Z(n14462) );
  XNOR U14091 ( .A(n14461), .B(n14455), .Z(n14457) );
  XOR U14092 ( .A(n14463), .B(n14464), .Z(n14455) );
  AND U14093 ( .A(n1297), .B(n14465), .Z(n14464) );
  XNOR U14094 ( .A(n14466), .B(n14467), .Z(n14461) );
  AND U14095 ( .A(n1289), .B(n14468), .Z(n14467) );
  XOR U14096 ( .A(p_input[1835]), .B(n14466), .Z(n14468) );
  XNOR U14097 ( .A(n14469), .B(n14470), .Z(n14466) );
  AND U14098 ( .A(n1293), .B(n14465), .Z(n14470) );
  XNOR U14099 ( .A(n14469), .B(n14463), .Z(n14465) );
  XOR U14100 ( .A(n14471), .B(n14472), .Z(n14463) );
  AND U14101 ( .A(n1308), .B(n14473), .Z(n14472) );
  XNOR U14102 ( .A(n14474), .B(n14475), .Z(n14469) );
  AND U14103 ( .A(n1300), .B(n14476), .Z(n14475) );
  XOR U14104 ( .A(p_input[1851]), .B(n14474), .Z(n14476) );
  XNOR U14105 ( .A(n14477), .B(n14478), .Z(n14474) );
  AND U14106 ( .A(n1304), .B(n14473), .Z(n14478) );
  XNOR U14107 ( .A(n14477), .B(n14471), .Z(n14473) );
  XOR U14108 ( .A(n14479), .B(n14480), .Z(n14471) );
  AND U14109 ( .A(n1319), .B(n14481), .Z(n14480) );
  XNOR U14110 ( .A(n14482), .B(n14483), .Z(n14477) );
  AND U14111 ( .A(n1311), .B(n14484), .Z(n14483) );
  XOR U14112 ( .A(p_input[1867]), .B(n14482), .Z(n14484) );
  XNOR U14113 ( .A(n14485), .B(n14486), .Z(n14482) );
  AND U14114 ( .A(n1315), .B(n14481), .Z(n14486) );
  XNOR U14115 ( .A(n14485), .B(n14479), .Z(n14481) );
  XOR U14116 ( .A(n14487), .B(n14488), .Z(n14479) );
  AND U14117 ( .A(n1330), .B(n14489), .Z(n14488) );
  XNOR U14118 ( .A(n14490), .B(n14491), .Z(n14485) );
  AND U14119 ( .A(n1322), .B(n14492), .Z(n14491) );
  XOR U14120 ( .A(p_input[1883]), .B(n14490), .Z(n14492) );
  XNOR U14121 ( .A(n14493), .B(n14494), .Z(n14490) );
  AND U14122 ( .A(n1326), .B(n14489), .Z(n14494) );
  XNOR U14123 ( .A(n14493), .B(n14487), .Z(n14489) );
  XOR U14124 ( .A(n14495), .B(n14496), .Z(n14487) );
  AND U14125 ( .A(n1341), .B(n14497), .Z(n14496) );
  XNOR U14126 ( .A(n14498), .B(n14499), .Z(n14493) );
  AND U14127 ( .A(n1333), .B(n14500), .Z(n14499) );
  XOR U14128 ( .A(p_input[1899]), .B(n14498), .Z(n14500) );
  XNOR U14129 ( .A(n14501), .B(n14502), .Z(n14498) );
  AND U14130 ( .A(n1337), .B(n14497), .Z(n14502) );
  XNOR U14131 ( .A(n14501), .B(n14495), .Z(n14497) );
  XOR U14132 ( .A(n14503), .B(n14504), .Z(n14495) );
  AND U14133 ( .A(n1352), .B(n14505), .Z(n14504) );
  XNOR U14134 ( .A(n14506), .B(n14507), .Z(n14501) );
  AND U14135 ( .A(n1344), .B(n14508), .Z(n14507) );
  XOR U14136 ( .A(p_input[1915]), .B(n14506), .Z(n14508) );
  XNOR U14137 ( .A(n14509), .B(n14510), .Z(n14506) );
  AND U14138 ( .A(n1348), .B(n14505), .Z(n14510) );
  XNOR U14139 ( .A(n14509), .B(n14503), .Z(n14505) );
  XOR U14140 ( .A(n14511), .B(n14512), .Z(n14503) );
  AND U14141 ( .A(n1363), .B(n14513), .Z(n14512) );
  XNOR U14142 ( .A(n14514), .B(n14515), .Z(n14509) );
  AND U14143 ( .A(n1355), .B(n14516), .Z(n14515) );
  XOR U14144 ( .A(p_input[1931]), .B(n14514), .Z(n14516) );
  XNOR U14145 ( .A(n14517), .B(n14518), .Z(n14514) );
  AND U14146 ( .A(n1359), .B(n14513), .Z(n14518) );
  XNOR U14147 ( .A(n14517), .B(n14511), .Z(n14513) );
  XOR U14148 ( .A(n14519), .B(n14520), .Z(n14511) );
  AND U14149 ( .A(n1374), .B(n14521), .Z(n14520) );
  XNOR U14150 ( .A(n14522), .B(n14523), .Z(n14517) );
  AND U14151 ( .A(n1366), .B(n14524), .Z(n14523) );
  XOR U14152 ( .A(p_input[1947]), .B(n14522), .Z(n14524) );
  XNOR U14153 ( .A(n14525), .B(n14526), .Z(n14522) );
  AND U14154 ( .A(n1370), .B(n14521), .Z(n14526) );
  XNOR U14155 ( .A(n14525), .B(n14519), .Z(n14521) );
  XOR U14156 ( .A(n14527), .B(n14528), .Z(n14519) );
  AND U14157 ( .A(n1385), .B(n14529), .Z(n14528) );
  XNOR U14158 ( .A(n14530), .B(n14531), .Z(n14525) );
  AND U14159 ( .A(n1377), .B(n14532), .Z(n14531) );
  XOR U14160 ( .A(p_input[1963]), .B(n14530), .Z(n14532) );
  XNOR U14161 ( .A(n14533), .B(n14534), .Z(n14530) );
  AND U14162 ( .A(n1381), .B(n14529), .Z(n14534) );
  XNOR U14163 ( .A(n14533), .B(n14527), .Z(n14529) );
  XOR U14164 ( .A(n14535), .B(n14536), .Z(n14527) );
  AND U14165 ( .A(n1396), .B(n14537), .Z(n14536) );
  XNOR U14166 ( .A(n14538), .B(n14539), .Z(n14533) );
  AND U14167 ( .A(n1388), .B(n14540), .Z(n14539) );
  XOR U14168 ( .A(p_input[1979]), .B(n14538), .Z(n14540) );
  XNOR U14169 ( .A(n14541), .B(n14542), .Z(n14538) );
  AND U14170 ( .A(n1392), .B(n14537), .Z(n14542) );
  XNOR U14171 ( .A(n14541), .B(n14535), .Z(n14537) );
  XOR U14172 ( .A(n14543), .B(n14544), .Z(n14535) );
  AND U14173 ( .A(n1407), .B(n14545), .Z(n14544) );
  XNOR U14174 ( .A(n14546), .B(n14547), .Z(n14541) );
  AND U14175 ( .A(n1399), .B(n14548), .Z(n14547) );
  XOR U14176 ( .A(p_input[1995]), .B(n14546), .Z(n14548) );
  XNOR U14177 ( .A(n14549), .B(n14550), .Z(n14546) );
  AND U14178 ( .A(n1403), .B(n14545), .Z(n14550) );
  XNOR U14179 ( .A(n14549), .B(n14543), .Z(n14545) );
  XOR U14180 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n14551), .Z(n14543) );
  AND U14181 ( .A(n1417), .B(n14552), .Z(n14551) );
  XNOR U14182 ( .A(n14553), .B(n14554), .Z(n14549) );
  AND U14183 ( .A(n1410), .B(n14555), .Z(n14554) );
  XOR U14184 ( .A(p_input[2011]), .B(n14553), .Z(n14555) );
  XNOR U14185 ( .A(n14556), .B(n14557), .Z(n14553) );
  AND U14186 ( .A(n1414), .B(n14552), .Z(n14557) );
  XOR U14187 ( .A(n14558), .B(n14556), .Z(n14552) );
  IV U14188 ( .A(\knn_comb_/min_val_out[0][11] ), .Z(n14558) );
  IV U14189 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n14556)
         );
  XOR U14190 ( .A(n27), .B(n14559), .Z(o[10]) );
  AND U14191 ( .A(n30), .B(n14560), .Z(n27) );
  XOR U14192 ( .A(n28), .B(n14559), .Z(n14560) );
  XOR U14193 ( .A(n14561), .B(n14562), .Z(n14559) );
  AND U14194 ( .A(n42), .B(n14563), .Z(n14562) );
  XOR U14195 ( .A(n14564), .B(n14565), .Z(n28) );
  AND U14196 ( .A(n34), .B(n14566), .Z(n14565) );
  XOR U14197 ( .A(p_input[10]), .B(n14564), .Z(n14566) );
  XNOR U14198 ( .A(n14567), .B(n14568), .Z(n14564) );
  AND U14199 ( .A(n38), .B(n14563), .Z(n14568) );
  XNOR U14200 ( .A(n14567), .B(n14561), .Z(n14563) );
  XOR U14201 ( .A(n14569), .B(n14570), .Z(n14561) );
  AND U14202 ( .A(n54), .B(n14571), .Z(n14570) );
  XNOR U14203 ( .A(n14572), .B(n14573), .Z(n14567) );
  AND U14204 ( .A(n46), .B(n14574), .Z(n14573) );
  XOR U14205 ( .A(p_input[26]), .B(n14572), .Z(n14574) );
  XNOR U14206 ( .A(n14575), .B(n14576), .Z(n14572) );
  AND U14207 ( .A(n50), .B(n14571), .Z(n14576) );
  XNOR U14208 ( .A(n14575), .B(n14569), .Z(n14571) );
  XOR U14209 ( .A(n14577), .B(n14578), .Z(n14569) );
  AND U14210 ( .A(n65), .B(n14579), .Z(n14578) );
  XNOR U14211 ( .A(n14580), .B(n14581), .Z(n14575) );
  AND U14212 ( .A(n57), .B(n14582), .Z(n14581) );
  XOR U14213 ( .A(p_input[42]), .B(n14580), .Z(n14582) );
  XNOR U14214 ( .A(n14583), .B(n14584), .Z(n14580) );
  AND U14215 ( .A(n61), .B(n14579), .Z(n14584) );
  XNOR U14216 ( .A(n14583), .B(n14577), .Z(n14579) );
  XOR U14217 ( .A(n14585), .B(n14586), .Z(n14577) );
  AND U14218 ( .A(n76), .B(n14587), .Z(n14586) );
  XNOR U14219 ( .A(n14588), .B(n14589), .Z(n14583) );
  AND U14220 ( .A(n68), .B(n14590), .Z(n14589) );
  XOR U14221 ( .A(p_input[58]), .B(n14588), .Z(n14590) );
  XNOR U14222 ( .A(n14591), .B(n14592), .Z(n14588) );
  AND U14223 ( .A(n72), .B(n14587), .Z(n14592) );
  XNOR U14224 ( .A(n14591), .B(n14585), .Z(n14587) );
  XOR U14225 ( .A(n14593), .B(n14594), .Z(n14585) );
  AND U14226 ( .A(n87), .B(n14595), .Z(n14594) );
  XNOR U14227 ( .A(n14596), .B(n14597), .Z(n14591) );
  AND U14228 ( .A(n79), .B(n14598), .Z(n14597) );
  XOR U14229 ( .A(p_input[74]), .B(n14596), .Z(n14598) );
  XNOR U14230 ( .A(n14599), .B(n14600), .Z(n14596) );
  AND U14231 ( .A(n83), .B(n14595), .Z(n14600) );
  XNOR U14232 ( .A(n14599), .B(n14593), .Z(n14595) );
  XOR U14233 ( .A(n14601), .B(n14602), .Z(n14593) );
  AND U14234 ( .A(n98), .B(n14603), .Z(n14602) );
  XNOR U14235 ( .A(n14604), .B(n14605), .Z(n14599) );
  AND U14236 ( .A(n90), .B(n14606), .Z(n14605) );
  XOR U14237 ( .A(p_input[90]), .B(n14604), .Z(n14606) );
  XNOR U14238 ( .A(n14607), .B(n14608), .Z(n14604) );
  AND U14239 ( .A(n94), .B(n14603), .Z(n14608) );
  XNOR U14240 ( .A(n14607), .B(n14601), .Z(n14603) );
  XOR U14241 ( .A(n14609), .B(n14610), .Z(n14601) );
  AND U14242 ( .A(n109), .B(n14611), .Z(n14610) );
  XNOR U14243 ( .A(n14612), .B(n14613), .Z(n14607) );
  AND U14244 ( .A(n101), .B(n14614), .Z(n14613) );
  XOR U14245 ( .A(p_input[106]), .B(n14612), .Z(n14614) );
  XNOR U14246 ( .A(n14615), .B(n14616), .Z(n14612) );
  AND U14247 ( .A(n105), .B(n14611), .Z(n14616) );
  XNOR U14248 ( .A(n14615), .B(n14609), .Z(n14611) );
  XOR U14249 ( .A(n14617), .B(n14618), .Z(n14609) );
  AND U14250 ( .A(n120), .B(n14619), .Z(n14618) );
  XNOR U14251 ( .A(n14620), .B(n14621), .Z(n14615) );
  AND U14252 ( .A(n112), .B(n14622), .Z(n14621) );
  XOR U14253 ( .A(p_input[122]), .B(n14620), .Z(n14622) );
  XNOR U14254 ( .A(n14623), .B(n14624), .Z(n14620) );
  AND U14255 ( .A(n116), .B(n14619), .Z(n14624) );
  XNOR U14256 ( .A(n14623), .B(n14617), .Z(n14619) );
  XOR U14257 ( .A(n14625), .B(n14626), .Z(n14617) );
  AND U14258 ( .A(n131), .B(n14627), .Z(n14626) );
  XNOR U14259 ( .A(n14628), .B(n14629), .Z(n14623) );
  AND U14260 ( .A(n123), .B(n14630), .Z(n14629) );
  XOR U14261 ( .A(p_input[138]), .B(n14628), .Z(n14630) );
  XNOR U14262 ( .A(n14631), .B(n14632), .Z(n14628) );
  AND U14263 ( .A(n127), .B(n14627), .Z(n14632) );
  XNOR U14264 ( .A(n14631), .B(n14625), .Z(n14627) );
  XOR U14265 ( .A(n14633), .B(n14634), .Z(n14625) );
  AND U14266 ( .A(n142), .B(n14635), .Z(n14634) );
  XNOR U14267 ( .A(n14636), .B(n14637), .Z(n14631) );
  AND U14268 ( .A(n134), .B(n14638), .Z(n14637) );
  XOR U14269 ( .A(p_input[154]), .B(n14636), .Z(n14638) );
  XNOR U14270 ( .A(n14639), .B(n14640), .Z(n14636) );
  AND U14271 ( .A(n138), .B(n14635), .Z(n14640) );
  XNOR U14272 ( .A(n14639), .B(n14633), .Z(n14635) );
  XOR U14273 ( .A(n14641), .B(n14642), .Z(n14633) );
  AND U14274 ( .A(n153), .B(n14643), .Z(n14642) );
  XNOR U14275 ( .A(n14644), .B(n14645), .Z(n14639) );
  AND U14276 ( .A(n145), .B(n14646), .Z(n14645) );
  XOR U14277 ( .A(p_input[170]), .B(n14644), .Z(n14646) );
  XNOR U14278 ( .A(n14647), .B(n14648), .Z(n14644) );
  AND U14279 ( .A(n149), .B(n14643), .Z(n14648) );
  XNOR U14280 ( .A(n14647), .B(n14641), .Z(n14643) );
  XOR U14281 ( .A(n14649), .B(n14650), .Z(n14641) );
  AND U14282 ( .A(n164), .B(n14651), .Z(n14650) );
  XNOR U14283 ( .A(n14652), .B(n14653), .Z(n14647) );
  AND U14284 ( .A(n156), .B(n14654), .Z(n14653) );
  XOR U14285 ( .A(p_input[186]), .B(n14652), .Z(n14654) );
  XNOR U14286 ( .A(n14655), .B(n14656), .Z(n14652) );
  AND U14287 ( .A(n160), .B(n14651), .Z(n14656) );
  XNOR U14288 ( .A(n14655), .B(n14649), .Z(n14651) );
  XOR U14289 ( .A(n14657), .B(n14658), .Z(n14649) );
  AND U14290 ( .A(n175), .B(n14659), .Z(n14658) );
  XNOR U14291 ( .A(n14660), .B(n14661), .Z(n14655) );
  AND U14292 ( .A(n167), .B(n14662), .Z(n14661) );
  XOR U14293 ( .A(p_input[202]), .B(n14660), .Z(n14662) );
  XNOR U14294 ( .A(n14663), .B(n14664), .Z(n14660) );
  AND U14295 ( .A(n171), .B(n14659), .Z(n14664) );
  XNOR U14296 ( .A(n14663), .B(n14657), .Z(n14659) );
  XOR U14297 ( .A(n14665), .B(n14666), .Z(n14657) );
  AND U14298 ( .A(n186), .B(n14667), .Z(n14666) );
  XNOR U14299 ( .A(n14668), .B(n14669), .Z(n14663) );
  AND U14300 ( .A(n178), .B(n14670), .Z(n14669) );
  XOR U14301 ( .A(p_input[218]), .B(n14668), .Z(n14670) );
  XNOR U14302 ( .A(n14671), .B(n14672), .Z(n14668) );
  AND U14303 ( .A(n182), .B(n14667), .Z(n14672) );
  XNOR U14304 ( .A(n14671), .B(n14665), .Z(n14667) );
  XOR U14305 ( .A(n14673), .B(n14674), .Z(n14665) );
  AND U14306 ( .A(n197), .B(n14675), .Z(n14674) );
  XNOR U14307 ( .A(n14676), .B(n14677), .Z(n14671) );
  AND U14308 ( .A(n189), .B(n14678), .Z(n14677) );
  XOR U14309 ( .A(p_input[234]), .B(n14676), .Z(n14678) );
  XNOR U14310 ( .A(n14679), .B(n14680), .Z(n14676) );
  AND U14311 ( .A(n193), .B(n14675), .Z(n14680) );
  XNOR U14312 ( .A(n14679), .B(n14673), .Z(n14675) );
  XOR U14313 ( .A(n14681), .B(n14682), .Z(n14673) );
  AND U14314 ( .A(n208), .B(n14683), .Z(n14682) );
  XNOR U14315 ( .A(n14684), .B(n14685), .Z(n14679) );
  AND U14316 ( .A(n200), .B(n14686), .Z(n14685) );
  XOR U14317 ( .A(p_input[250]), .B(n14684), .Z(n14686) );
  XNOR U14318 ( .A(n14687), .B(n14688), .Z(n14684) );
  AND U14319 ( .A(n204), .B(n14683), .Z(n14688) );
  XNOR U14320 ( .A(n14687), .B(n14681), .Z(n14683) );
  XOR U14321 ( .A(n14689), .B(n14690), .Z(n14681) );
  AND U14322 ( .A(n219), .B(n14691), .Z(n14690) );
  XNOR U14323 ( .A(n14692), .B(n14693), .Z(n14687) );
  AND U14324 ( .A(n211), .B(n14694), .Z(n14693) );
  XOR U14325 ( .A(p_input[266]), .B(n14692), .Z(n14694) );
  XNOR U14326 ( .A(n14695), .B(n14696), .Z(n14692) );
  AND U14327 ( .A(n215), .B(n14691), .Z(n14696) );
  XNOR U14328 ( .A(n14695), .B(n14689), .Z(n14691) );
  XOR U14329 ( .A(n14697), .B(n14698), .Z(n14689) );
  AND U14330 ( .A(n230), .B(n14699), .Z(n14698) );
  XNOR U14331 ( .A(n14700), .B(n14701), .Z(n14695) );
  AND U14332 ( .A(n222), .B(n14702), .Z(n14701) );
  XOR U14333 ( .A(p_input[282]), .B(n14700), .Z(n14702) );
  XNOR U14334 ( .A(n14703), .B(n14704), .Z(n14700) );
  AND U14335 ( .A(n226), .B(n14699), .Z(n14704) );
  XNOR U14336 ( .A(n14703), .B(n14697), .Z(n14699) );
  XOR U14337 ( .A(n14705), .B(n14706), .Z(n14697) );
  AND U14338 ( .A(n241), .B(n14707), .Z(n14706) );
  XNOR U14339 ( .A(n14708), .B(n14709), .Z(n14703) );
  AND U14340 ( .A(n233), .B(n14710), .Z(n14709) );
  XOR U14341 ( .A(p_input[298]), .B(n14708), .Z(n14710) );
  XNOR U14342 ( .A(n14711), .B(n14712), .Z(n14708) );
  AND U14343 ( .A(n237), .B(n14707), .Z(n14712) );
  XNOR U14344 ( .A(n14711), .B(n14705), .Z(n14707) );
  XOR U14345 ( .A(n14713), .B(n14714), .Z(n14705) );
  AND U14346 ( .A(n252), .B(n14715), .Z(n14714) );
  XNOR U14347 ( .A(n14716), .B(n14717), .Z(n14711) );
  AND U14348 ( .A(n244), .B(n14718), .Z(n14717) );
  XOR U14349 ( .A(p_input[314]), .B(n14716), .Z(n14718) );
  XNOR U14350 ( .A(n14719), .B(n14720), .Z(n14716) );
  AND U14351 ( .A(n248), .B(n14715), .Z(n14720) );
  XNOR U14352 ( .A(n14719), .B(n14713), .Z(n14715) );
  XOR U14353 ( .A(n14721), .B(n14722), .Z(n14713) );
  AND U14354 ( .A(n263), .B(n14723), .Z(n14722) );
  XNOR U14355 ( .A(n14724), .B(n14725), .Z(n14719) );
  AND U14356 ( .A(n255), .B(n14726), .Z(n14725) );
  XOR U14357 ( .A(p_input[330]), .B(n14724), .Z(n14726) );
  XNOR U14358 ( .A(n14727), .B(n14728), .Z(n14724) );
  AND U14359 ( .A(n259), .B(n14723), .Z(n14728) );
  XNOR U14360 ( .A(n14727), .B(n14721), .Z(n14723) );
  XOR U14361 ( .A(n14729), .B(n14730), .Z(n14721) );
  AND U14362 ( .A(n274), .B(n14731), .Z(n14730) );
  XNOR U14363 ( .A(n14732), .B(n14733), .Z(n14727) );
  AND U14364 ( .A(n266), .B(n14734), .Z(n14733) );
  XOR U14365 ( .A(p_input[346]), .B(n14732), .Z(n14734) );
  XNOR U14366 ( .A(n14735), .B(n14736), .Z(n14732) );
  AND U14367 ( .A(n270), .B(n14731), .Z(n14736) );
  XNOR U14368 ( .A(n14735), .B(n14729), .Z(n14731) );
  XOR U14369 ( .A(n14737), .B(n14738), .Z(n14729) );
  AND U14370 ( .A(n285), .B(n14739), .Z(n14738) );
  XNOR U14371 ( .A(n14740), .B(n14741), .Z(n14735) );
  AND U14372 ( .A(n277), .B(n14742), .Z(n14741) );
  XOR U14373 ( .A(p_input[362]), .B(n14740), .Z(n14742) );
  XNOR U14374 ( .A(n14743), .B(n14744), .Z(n14740) );
  AND U14375 ( .A(n281), .B(n14739), .Z(n14744) );
  XNOR U14376 ( .A(n14743), .B(n14737), .Z(n14739) );
  XOR U14377 ( .A(n14745), .B(n14746), .Z(n14737) );
  AND U14378 ( .A(n296), .B(n14747), .Z(n14746) );
  XNOR U14379 ( .A(n14748), .B(n14749), .Z(n14743) );
  AND U14380 ( .A(n288), .B(n14750), .Z(n14749) );
  XOR U14381 ( .A(p_input[378]), .B(n14748), .Z(n14750) );
  XNOR U14382 ( .A(n14751), .B(n14752), .Z(n14748) );
  AND U14383 ( .A(n292), .B(n14747), .Z(n14752) );
  XNOR U14384 ( .A(n14751), .B(n14745), .Z(n14747) );
  XOR U14385 ( .A(n14753), .B(n14754), .Z(n14745) );
  AND U14386 ( .A(n307), .B(n14755), .Z(n14754) );
  XNOR U14387 ( .A(n14756), .B(n14757), .Z(n14751) );
  AND U14388 ( .A(n299), .B(n14758), .Z(n14757) );
  XOR U14389 ( .A(p_input[394]), .B(n14756), .Z(n14758) );
  XNOR U14390 ( .A(n14759), .B(n14760), .Z(n14756) );
  AND U14391 ( .A(n303), .B(n14755), .Z(n14760) );
  XNOR U14392 ( .A(n14759), .B(n14753), .Z(n14755) );
  XOR U14393 ( .A(n14761), .B(n14762), .Z(n14753) );
  AND U14394 ( .A(n318), .B(n14763), .Z(n14762) );
  XNOR U14395 ( .A(n14764), .B(n14765), .Z(n14759) );
  AND U14396 ( .A(n310), .B(n14766), .Z(n14765) );
  XOR U14397 ( .A(p_input[410]), .B(n14764), .Z(n14766) );
  XNOR U14398 ( .A(n14767), .B(n14768), .Z(n14764) );
  AND U14399 ( .A(n314), .B(n14763), .Z(n14768) );
  XNOR U14400 ( .A(n14767), .B(n14761), .Z(n14763) );
  XOR U14401 ( .A(n14769), .B(n14770), .Z(n14761) );
  AND U14402 ( .A(n329), .B(n14771), .Z(n14770) );
  XNOR U14403 ( .A(n14772), .B(n14773), .Z(n14767) );
  AND U14404 ( .A(n321), .B(n14774), .Z(n14773) );
  XOR U14405 ( .A(p_input[426]), .B(n14772), .Z(n14774) );
  XNOR U14406 ( .A(n14775), .B(n14776), .Z(n14772) );
  AND U14407 ( .A(n325), .B(n14771), .Z(n14776) );
  XNOR U14408 ( .A(n14775), .B(n14769), .Z(n14771) );
  XOR U14409 ( .A(n14777), .B(n14778), .Z(n14769) );
  AND U14410 ( .A(n340), .B(n14779), .Z(n14778) );
  XNOR U14411 ( .A(n14780), .B(n14781), .Z(n14775) );
  AND U14412 ( .A(n332), .B(n14782), .Z(n14781) );
  XOR U14413 ( .A(p_input[442]), .B(n14780), .Z(n14782) );
  XNOR U14414 ( .A(n14783), .B(n14784), .Z(n14780) );
  AND U14415 ( .A(n336), .B(n14779), .Z(n14784) );
  XNOR U14416 ( .A(n14783), .B(n14777), .Z(n14779) );
  XOR U14417 ( .A(n14785), .B(n14786), .Z(n14777) );
  AND U14418 ( .A(n351), .B(n14787), .Z(n14786) );
  XNOR U14419 ( .A(n14788), .B(n14789), .Z(n14783) );
  AND U14420 ( .A(n343), .B(n14790), .Z(n14789) );
  XOR U14421 ( .A(p_input[458]), .B(n14788), .Z(n14790) );
  XNOR U14422 ( .A(n14791), .B(n14792), .Z(n14788) );
  AND U14423 ( .A(n347), .B(n14787), .Z(n14792) );
  XNOR U14424 ( .A(n14791), .B(n14785), .Z(n14787) );
  XOR U14425 ( .A(n14793), .B(n14794), .Z(n14785) );
  AND U14426 ( .A(n362), .B(n14795), .Z(n14794) );
  XNOR U14427 ( .A(n14796), .B(n14797), .Z(n14791) );
  AND U14428 ( .A(n354), .B(n14798), .Z(n14797) );
  XOR U14429 ( .A(p_input[474]), .B(n14796), .Z(n14798) );
  XNOR U14430 ( .A(n14799), .B(n14800), .Z(n14796) );
  AND U14431 ( .A(n358), .B(n14795), .Z(n14800) );
  XNOR U14432 ( .A(n14799), .B(n14793), .Z(n14795) );
  XOR U14433 ( .A(n14801), .B(n14802), .Z(n14793) );
  AND U14434 ( .A(n373), .B(n14803), .Z(n14802) );
  XNOR U14435 ( .A(n14804), .B(n14805), .Z(n14799) );
  AND U14436 ( .A(n365), .B(n14806), .Z(n14805) );
  XOR U14437 ( .A(p_input[490]), .B(n14804), .Z(n14806) );
  XNOR U14438 ( .A(n14807), .B(n14808), .Z(n14804) );
  AND U14439 ( .A(n369), .B(n14803), .Z(n14808) );
  XNOR U14440 ( .A(n14807), .B(n14801), .Z(n14803) );
  XOR U14441 ( .A(n14809), .B(n14810), .Z(n14801) );
  AND U14442 ( .A(n384), .B(n14811), .Z(n14810) );
  XNOR U14443 ( .A(n14812), .B(n14813), .Z(n14807) );
  AND U14444 ( .A(n376), .B(n14814), .Z(n14813) );
  XOR U14445 ( .A(p_input[506]), .B(n14812), .Z(n14814) );
  XNOR U14446 ( .A(n14815), .B(n14816), .Z(n14812) );
  AND U14447 ( .A(n380), .B(n14811), .Z(n14816) );
  XNOR U14448 ( .A(n14815), .B(n14809), .Z(n14811) );
  XOR U14449 ( .A(n14817), .B(n14818), .Z(n14809) );
  AND U14450 ( .A(n395), .B(n14819), .Z(n14818) );
  XNOR U14451 ( .A(n14820), .B(n14821), .Z(n14815) );
  AND U14452 ( .A(n387), .B(n14822), .Z(n14821) );
  XOR U14453 ( .A(p_input[522]), .B(n14820), .Z(n14822) );
  XNOR U14454 ( .A(n14823), .B(n14824), .Z(n14820) );
  AND U14455 ( .A(n391), .B(n14819), .Z(n14824) );
  XNOR U14456 ( .A(n14823), .B(n14817), .Z(n14819) );
  XOR U14457 ( .A(n14825), .B(n14826), .Z(n14817) );
  AND U14458 ( .A(n406), .B(n14827), .Z(n14826) );
  XNOR U14459 ( .A(n14828), .B(n14829), .Z(n14823) );
  AND U14460 ( .A(n398), .B(n14830), .Z(n14829) );
  XOR U14461 ( .A(p_input[538]), .B(n14828), .Z(n14830) );
  XNOR U14462 ( .A(n14831), .B(n14832), .Z(n14828) );
  AND U14463 ( .A(n402), .B(n14827), .Z(n14832) );
  XNOR U14464 ( .A(n14831), .B(n14825), .Z(n14827) );
  XOR U14465 ( .A(n14833), .B(n14834), .Z(n14825) );
  AND U14466 ( .A(n417), .B(n14835), .Z(n14834) );
  XNOR U14467 ( .A(n14836), .B(n14837), .Z(n14831) );
  AND U14468 ( .A(n409), .B(n14838), .Z(n14837) );
  XOR U14469 ( .A(p_input[554]), .B(n14836), .Z(n14838) );
  XNOR U14470 ( .A(n14839), .B(n14840), .Z(n14836) );
  AND U14471 ( .A(n413), .B(n14835), .Z(n14840) );
  XNOR U14472 ( .A(n14839), .B(n14833), .Z(n14835) );
  XOR U14473 ( .A(n14841), .B(n14842), .Z(n14833) );
  AND U14474 ( .A(n428), .B(n14843), .Z(n14842) );
  XNOR U14475 ( .A(n14844), .B(n14845), .Z(n14839) );
  AND U14476 ( .A(n420), .B(n14846), .Z(n14845) );
  XOR U14477 ( .A(p_input[570]), .B(n14844), .Z(n14846) );
  XNOR U14478 ( .A(n14847), .B(n14848), .Z(n14844) );
  AND U14479 ( .A(n424), .B(n14843), .Z(n14848) );
  XNOR U14480 ( .A(n14847), .B(n14841), .Z(n14843) );
  XOR U14481 ( .A(n14849), .B(n14850), .Z(n14841) );
  AND U14482 ( .A(n439), .B(n14851), .Z(n14850) );
  XNOR U14483 ( .A(n14852), .B(n14853), .Z(n14847) );
  AND U14484 ( .A(n431), .B(n14854), .Z(n14853) );
  XOR U14485 ( .A(p_input[586]), .B(n14852), .Z(n14854) );
  XNOR U14486 ( .A(n14855), .B(n14856), .Z(n14852) );
  AND U14487 ( .A(n435), .B(n14851), .Z(n14856) );
  XNOR U14488 ( .A(n14855), .B(n14849), .Z(n14851) );
  XOR U14489 ( .A(n14857), .B(n14858), .Z(n14849) );
  AND U14490 ( .A(n450), .B(n14859), .Z(n14858) );
  XNOR U14491 ( .A(n14860), .B(n14861), .Z(n14855) );
  AND U14492 ( .A(n442), .B(n14862), .Z(n14861) );
  XOR U14493 ( .A(p_input[602]), .B(n14860), .Z(n14862) );
  XNOR U14494 ( .A(n14863), .B(n14864), .Z(n14860) );
  AND U14495 ( .A(n446), .B(n14859), .Z(n14864) );
  XNOR U14496 ( .A(n14863), .B(n14857), .Z(n14859) );
  XOR U14497 ( .A(n14865), .B(n14866), .Z(n14857) );
  AND U14498 ( .A(n461), .B(n14867), .Z(n14866) );
  XNOR U14499 ( .A(n14868), .B(n14869), .Z(n14863) );
  AND U14500 ( .A(n453), .B(n14870), .Z(n14869) );
  XOR U14501 ( .A(p_input[618]), .B(n14868), .Z(n14870) );
  XNOR U14502 ( .A(n14871), .B(n14872), .Z(n14868) );
  AND U14503 ( .A(n457), .B(n14867), .Z(n14872) );
  XNOR U14504 ( .A(n14871), .B(n14865), .Z(n14867) );
  XOR U14505 ( .A(n14873), .B(n14874), .Z(n14865) );
  AND U14506 ( .A(n472), .B(n14875), .Z(n14874) );
  XNOR U14507 ( .A(n14876), .B(n14877), .Z(n14871) );
  AND U14508 ( .A(n464), .B(n14878), .Z(n14877) );
  XOR U14509 ( .A(p_input[634]), .B(n14876), .Z(n14878) );
  XNOR U14510 ( .A(n14879), .B(n14880), .Z(n14876) );
  AND U14511 ( .A(n468), .B(n14875), .Z(n14880) );
  XNOR U14512 ( .A(n14879), .B(n14873), .Z(n14875) );
  XOR U14513 ( .A(n14881), .B(n14882), .Z(n14873) );
  AND U14514 ( .A(n483), .B(n14883), .Z(n14882) );
  XNOR U14515 ( .A(n14884), .B(n14885), .Z(n14879) );
  AND U14516 ( .A(n475), .B(n14886), .Z(n14885) );
  XOR U14517 ( .A(p_input[650]), .B(n14884), .Z(n14886) );
  XNOR U14518 ( .A(n14887), .B(n14888), .Z(n14884) );
  AND U14519 ( .A(n479), .B(n14883), .Z(n14888) );
  XNOR U14520 ( .A(n14887), .B(n14881), .Z(n14883) );
  XOR U14521 ( .A(n14889), .B(n14890), .Z(n14881) );
  AND U14522 ( .A(n494), .B(n14891), .Z(n14890) );
  XNOR U14523 ( .A(n14892), .B(n14893), .Z(n14887) );
  AND U14524 ( .A(n486), .B(n14894), .Z(n14893) );
  XOR U14525 ( .A(p_input[666]), .B(n14892), .Z(n14894) );
  XNOR U14526 ( .A(n14895), .B(n14896), .Z(n14892) );
  AND U14527 ( .A(n490), .B(n14891), .Z(n14896) );
  XNOR U14528 ( .A(n14895), .B(n14889), .Z(n14891) );
  XOR U14529 ( .A(n14897), .B(n14898), .Z(n14889) );
  AND U14530 ( .A(n505), .B(n14899), .Z(n14898) );
  XNOR U14531 ( .A(n14900), .B(n14901), .Z(n14895) );
  AND U14532 ( .A(n497), .B(n14902), .Z(n14901) );
  XOR U14533 ( .A(p_input[682]), .B(n14900), .Z(n14902) );
  XNOR U14534 ( .A(n14903), .B(n14904), .Z(n14900) );
  AND U14535 ( .A(n501), .B(n14899), .Z(n14904) );
  XNOR U14536 ( .A(n14903), .B(n14897), .Z(n14899) );
  XOR U14537 ( .A(n14905), .B(n14906), .Z(n14897) );
  AND U14538 ( .A(n516), .B(n14907), .Z(n14906) );
  XNOR U14539 ( .A(n14908), .B(n14909), .Z(n14903) );
  AND U14540 ( .A(n508), .B(n14910), .Z(n14909) );
  XOR U14541 ( .A(p_input[698]), .B(n14908), .Z(n14910) );
  XNOR U14542 ( .A(n14911), .B(n14912), .Z(n14908) );
  AND U14543 ( .A(n512), .B(n14907), .Z(n14912) );
  XNOR U14544 ( .A(n14911), .B(n14905), .Z(n14907) );
  XOR U14545 ( .A(n14913), .B(n14914), .Z(n14905) );
  AND U14546 ( .A(n527), .B(n14915), .Z(n14914) );
  XNOR U14547 ( .A(n14916), .B(n14917), .Z(n14911) );
  AND U14548 ( .A(n519), .B(n14918), .Z(n14917) );
  XOR U14549 ( .A(p_input[714]), .B(n14916), .Z(n14918) );
  XNOR U14550 ( .A(n14919), .B(n14920), .Z(n14916) );
  AND U14551 ( .A(n523), .B(n14915), .Z(n14920) );
  XNOR U14552 ( .A(n14919), .B(n14913), .Z(n14915) );
  XOR U14553 ( .A(n14921), .B(n14922), .Z(n14913) );
  AND U14554 ( .A(n538), .B(n14923), .Z(n14922) );
  XNOR U14555 ( .A(n14924), .B(n14925), .Z(n14919) );
  AND U14556 ( .A(n530), .B(n14926), .Z(n14925) );
  XOR U14557 ( .A(p_input[730]), .B(n14924), .Z(n14926) );
  XNOR U14558 ( .A(n14927), .B(n14928), .Z(n14924) );
  AND U14559 ( .A(n534), .B(n14923), .Z(n14928) );
  XNOR U14560 ( .A(n14927), .B(n14921), .Z(n14923) );
  XOR U14561 ( .A(n14929), .B(n14930), .Z(n14921) );
  AND U14562 ( .A(n549), .B(n14931), .Z(n14930) );
  XNOR U14563 ( .A(n14932), .B(n14933), .Z(n14927) );
  AND U14564 ( .A(n541), .B(n14934), .Z(n14933) );
  XOR U14565 ( .A(p_input[746]), .B(n14932), .Z(n14934) );
  XNOR U14566 ( .A(n14935), .B(n14936), .Z(n14932) );
  AND U14567 ( .A(n545), .B(n14931), .Z(n14936) );
  XNOR U14568 ( .A(n14935), .B(n14929), .Z(n14931) );
  XOR U14569 ( .A(n14937), .B(n14938), .Z(n14929) );
  AND U14570 ( .A(n560), .B(n14939), .Z(n14938) );
  XNOR U14571 ( .A(n14940), .B(n14941), .Z(n14935) );
  AND U14572 ( .A(n552), .B(n14942), .Z(n14941) );
  XOR U14573 ( .A(p_input[762]), .B(n14940), .Z(n14942) );
  XNOR U14574 ( .A(n14943), .B(n14944), .Z(n14940) );
  AND U14575 ( .A(n556), .B(n14939), .Z(n14944) );
  XNOR U14576 ( .A(n14943), .B(n14937), .Z(n14939) );
  XOR U14577 ( .A(n14945), .B(n14946), .Z(n14937) );
  AND U14578 ( .A(n571), .B(n14947), .Z(n14946) );
  XNOR U14579 ( .A(n14948), .B(n14949), .Z(n14943) );
  AND U14580 ( .A(n563), .B(n14950), .Z(n14949) );
  XOR U14581 ( .A(p_input[778]), .B(n14948), .Z(n14950) );
  XNOR U14582 ( .A(n14951), .B(n14952), .Z(n14948) );
  AND U14583 ( .A(n567), .B(n14947), .Z(n14952) );
  XNOR U14584 ( .A(n14951), .B(n14945), .Z(n14947) );
  XOR U14585 ( .A(n14953), .B(n14954), .Z(n14945) );
  AND U14586 ( .A(n582), .B(n14955), .Z(n14954) );
  XNOR U14587 ( .A(n14956), .B(n14957), .Z(n14951) );
  AND U14588 ( .A(n574), .B(n14958), .Z(n14957) );
  XOR U14589 ( .A(p_input[794]), .B(n14956), .Z(n14958) );
  XNOR U14590 ( .A(n14959), .B(n14960), .Z(n14956) );
  AND U14591 ( .A(n578), .B(n14955), .Z(n14960) );
  XNOR U14592 ( .A(n14959), .B(n14953), .Z(n14955) );
  XOR U14593 ( .A(n14961), .B(n14962), .Z(n14953) );
  AND U14594 ( .A(n593), .B(n14963), .Z(n14962) );
  XNOR U14595 ( .A(n14964), .B(n14965), .Z(n14959) );
  AND U14596 ( .A(n585), .B(n14966), .Z(n14965) );
  XOR U14597 ( .A(p_input[810]), .B(n14964), .Z(n14966) );
  XNOR U14598 ( .A(n14967), .B(n14968), .Z(n14964) );
  AND U14599 ( .A(n589), .B(n14963), .Z(n14968) );
  XNOR U14600 ( .A(n14967), .B(n14961), .Z(n14963) );
  XOR U14601 ( .A(n14969), .B(n14970), .Z(n14961) );
  AND U14602 ( .A(n604), .B(n14971), .Z(n14970) );
  XNOR U14603 ( .A(n14972), .B(n14973), .Z(n14967) );
  AND U14604 ( .A(n596), .B(n14974), .Z(n14973) );
  XOR U14605 ( .A(p_input[826]), .B(n14972), .Z(n14974) );
  XNOR U14606 ( .A(n14975), .B(n14976), .Z(n14972) );
  AND U14607 ( .A(n600), .B(n14971), .Z(n14976) );
  XNOR U14608 ( .A(n14975), .B(n14969), .Z(n14971) );
  XOR U14609 ( .A(n14977), .B(n14978), .Z(n14969) );
  AND U14610 ( .A(n615), .B(n14979), .Z(n14978) );
  XNOR U14611 ( .A(n14980), .B(n14981), .Z(n14975) );
  AND U14612 ( .A(n607), .B(n14982), .Z(n14981) );
  XOR U14613 ( .A(p_input[842]), .B(n14980), .Z(n14982) );
  XNOR U14614 ( .A(n14983), .B(n14984), .Z(n14980) );
  AND U14615 ( .A(n611), .B(n14979), .Z(n14984) );
  XNOR U14616 ( .A(n14983), .B(n14977), .Z(n14979) );
  XOR U14617 ( .A(n14985), .B(n14986), .Z(n14977) );
  AND U14618 ( .A(n626), .B(n14987), .Z(n14986) );
  XNOR U14619 ( .A(n14988), .B(n14989), .Z(n14983) );
  AND U14620 ( .A(n618), .B(n14990), .Z(n14989) );
  XOR U14621 ( .A(p_input[858]), .B(n14988), .Z(n14990) );
  XNOR U14622 ( .A(n14991), .B(n14992), .Z(n14988) );
  AND U14623 ( .A(n622), .B(n14987), .Z(n14992) );
  XNOR U14624 ( .A(n14991), .B(n14985), .Z(n14987) );
  XOR U14625 ( .A(n14993), .B(n14994), .Z(n14985) );
  AND U14626 ( .A(n637), .B(n14995), .Z(n14994) );
  XNOR U14627 ( .A(n14996), .B(n14997), .Z(n14991) );
  AND U14628 ( .A(n629), .B(n14998), .Z(n14997) );
  XOR U14629 ( .A(p_input[874]), .B(n14996), .Z(n14998) );
  XNOR U14630 ( .A(n14999), .B(n15000), .Z(n14996) );
  AND U14631 ( .A(n633), .B(n14995), .Z(n15000) );
  XNOR U14632 ( .A(n14999), .B(n14993), .Z(n14995) );
  XOR U14633 ( .A(n15001), .B(n15002), .Z(n14993) );
  AND U14634 ( .A(n648), .B(n15003), .Z(n15002) );
  XNOR U14635 ( .A(n15004), .B(n15005), .Z(n14999) );
  AND U14636 ( .A(n640), .B(n15006), .Z(n15005) );
  XOR U14637 ( .A(p_input[890]), .B(n15004), .Z(n15006) );
  XNOR U14638 ( .A(n15007), .B(n15008), .Z(n15004) );
  AND U14639 ( .A(n644), .B(n15003), .Z(n15008) );
  XNOR U14640 ( .A(n15007), .B(n15001), .Z(n15003) );
  XOR U14641 ( .A(n15009), .B(n15010), .Z(n15001) );
  AND U14642 ( .A(n659), .B(n15011), .Z(n15010) );
  XNOR U14643 ( .A(n15012), .B(n15013), .Z(n15007) );
  AND U14644 ( .A(n651), .B(n15014), .Z(n15013) );
  XOR U14645 ( .A(p_input[906]), .B(n15012), .Z(n15014) );
  XNOR U14646 ( .A(n15015), .B(n15016), .Z(n15012) );
  AND U14647 ( .A(n655), .B(n15011), .Z(n15016) );
  XNOR U14648 ( .A(n15015), .B(n15009), .Z(n15011) );
  XOR U14649 ( .A(n15017), .B(n15018), .Z(n15009) );
  AND U14650 ( .A(n670), .B(n15019), .Z(n15018) );
  XNOR U14651 ( .A(n15020), .B(n15021), .Z(n15015) );
  AND U14652 ( .A(n662), .B(n15022), .Z(n15021) );
  XOR U14653 ( .A(p_input[922]), .B(n15020), .Z(n15022) );
  XNOR U14654 ( .A(n15023), .B(n15024), .Z(n15020) );
  AND U14655 ( .A(n666), .B(n15019), .Z(n15024) );
  XNOR U14656 ( .A(n15023), .B(n15017), .Z(n15019) );
  XOR U14657 ( .A(n15025), .B(n15026), .Z(n15017) );
  AND U14658 ( .A(n681), .B(n15027), .Z(n15026) );
  XNOR U14659 ( .A(n15028), .B(n15029), .Z(n15023) );
  AND U14660 ( .A(n673), .B(n15030), .Z(n15029) );
  XOR U14661 ( .A(p_input[938]), .B(n15028), .Z(n15030) );
  XNOR U14662 ( .A(n15031), .B(n15032), .Z(n15028) );
  AND U14663 ( .A(n677), .B(n15027), .Z(n15032) );
  XNOR U14664 ( .A(n15031), .B(n15025), .Z(n15027) );
  XOR U14665 ( .A(n15033), .B(n15034), .Z(n15025) );
  AND U14666 ( .A(n692), .B(n15035), .Z(n15034) );
  XNOR U14667 ( .A(n15036), .B(n15037), .Z(n15031) );
  AND U14668 ( .A(n684), .B(n15038), .Z(n15037) );
  XOR U14669 ( .A(p_input[954]), .B(n15036), .Z(n15038) );
  XNOR U14670 ( .A(n15039), .B(n15040), .Z(n15036) );
  AND U14671 ( .A(n688), .B(n15035), .Z(n15040) );
  XNOR U14672 ( .A(n15039), .B(n15033), .Z(n15035) );
  XOR U14673 ( .A(n15041), .B(n15042), .Z(n15033) );
  AND U14674 ( .A(n703), .B(n15043), .Z(n15042) );
  XNOR U14675 ( .A(n15044), .B(n15045), .Z(n15039) );
  AND U14676 ( .A(n695), .B(n15046), .Z(n15045) );
  XOR U14677 ( .A(p_input[970]), .B(n15044), .Z(n15046) );
  XNOR U14678 ( .A(n15047), .B(n15048), .Z(n15044) );
  AND U14679 ( .A(n699), .B(n15043), .Z(n15048) );
  XNOR U14680 ( .A(n15047), .B(n15041), .Z(n15043) );
  XOR U14681 ( .A(n15049), .B(n15050), .Z(n15041) );
  AND U14682 ( .A(n714), .B(n15051), .Z(n15050) );
  XNOR U14683 ( .A(n15052), .B(n15053), .Z(n15047) );
  AND U14684 ( .A(n706), .B(n15054), .Z(n15053) );
  XOR U14685 ( .A(p_input[986]), .B(n15052), .Z(n15054) );
  XNOR U14686 ( .A(n15055), .B(n15056), .Z(n15052) );
  AND U14687 ( .A(n710), .B(n15051), .Z(n15056) );
  XNOR U14688 ( .A(n15055), .B(n15049), .Z(n15051) );
  XOR U14689 ( .A(n15057), .B(n15058), .Z(n15049) );
  AND U14690 ( .A(n725), .B(n15059), .Z(n15058) );
  XNOR U14691 ( .A(n15060), .B(n15061), .Z(n15055) );
  AND U14692 ( .A(n717), .B(n15062), .Z(n15061) );
  XOR U14693 ( .A(p_input[1002]), .B(n15060), .Z(n15062) );
  XNOR U14694 ( .A(n15063), .B(n15064), .Z(n15060) );
  AND U14695 ( .A(n721), .B(n15059), .Z(n15064) );
  XNOR U14696 ( .A(n15063), .B(n15057), .Z(n15059) );
  XOR U14697 ( .A(n15065), .B(n15066), .Z(n15057) );
  AND U14698 ( .A(n736), .B(n15067), .Z(n15066) );
  XNOR U14699 ( .A(n15068), .B(n15069), .Z(n15063) );
  AND U14700 ( .A(n728), .B(n15070), .Z(n15069) );
  XOR U14701 ( .A(p_input[1018]), .B(n15068), .Z(n15070) );
  XNOR U14702 ( .A(n15071), .B(n15072), .Z(n15068) );
  AND U14703 ( .A(n732), .B(n15067), .Z(n15072) );
  XNOR U14704 ( .A(n15071), .B(n15065), .Z(n15067) );
  XOR U14705 ( .A(n15073), .B(n15074), .Z(n15065) );
  AND U14706 ( .A(n747), .B(n15075), .Z(n15074) );
  XNOR U14707 ( .A(n15076), .B(n15077), .Z(n15071) );
  AND U14708 ( .A(n739), .B(n15078), .Z(n15077) );
  XOR U14709 ( .A(p_input[1034]), .B(n15076), .Z(n15078) );
  XNOR U14710 ( .A(n15079), .B(n15080), .Z(n15076) );
  AND U14711 ( .A(n743), .B(n15075), .Z(n15080) );
  XNOR U14712 ( .A(n15079), .B(n15073), .Z(n15075) );
  XOR U14713 ( .A(n15081), .B(n15082), .Z(n15073) );
  AND U14714 ( .A(n758), .B(n15083), .Z(n15082) );
  XNOR U14715 ( .A(n15084), .B(n15085), .Z(n15079) );
  AND U14716 ( .A(n750), .B(n15086), .Z(n15085) );
  XOR U14717 ( .A(p_input[1050]), .B(n15084), .Z(n15086) );
  XNOR U14718 ( .A(n15087), .B(n15088), .Z(n15084) );
  AND U14719 ( .A(n754), .B(n15083), .Z(n15088) );
  XNOR U14720 ( .A(n15087), .B(n15081), .Z(n15083) );
  XOR U14721 ( .A(n15089), .B(n15090), .Z(n15081) );
  AND U14722 ( .A(n769), .B(n15091), .Z(n15090) );
  XNOR U14723 ( .A(n15092), .B(n15093), .Z(n15087) );
  AND U14724 ( .A(n761), .B(n15094), .Z(n15093) );
  XOR U14725 ( .A(p_input[1066]), .B(n15092), .Z(n15094) );
  XNOR U14726 ( .A(n15095), .B(n15096), .Z(n15092) );
  AND U14727 ( .A(n765), .B(n15091), .Z(n15096) );
  XNOR U14728 ( .A(n15095), .B(n15089), .Z(n15091) );
  XOR U14729 ( .A(n15097), .B(n15098), .Z(n15089) );
  AND U14730 ( .A(n780), .B(n15099), .Z(n15098) );
  XNOR U14731 ( .A(n15100), .B(n15101), .Z(n15095) );
  AND U14732 ( .A(n772), .B(n15102), .Z(n15101) );
  XOR U14733 ( .A(p_input[1082]), .B(n15100), .Z(n15102) );
  XNOR U14734 ( .A(n15103), .B(n15104), .Z(n15100) );
  AND U14735 ( .A(n776), .B(n15099), .Z(n15104) );
  XNOR U14736 ( .A(n15103), .B(n15097), .Z(n15099) );
  XOR U14737 ( .A(n15105), .B(n15106), .Z(n15097) );
  AND U14738 ( .A(n791), .B(n15107), .Z(n15106) );
  XNOR U14739 ( .A(n15108), .B(n15109), .Z(n15103) );
  AND U14740 ( .A(n783), .B(n15110), .Z(n15109) );
  XOR U14741 ( .A(p_input[1098]), .B(n15108), .Z(n15110) );
  XNOR U14742 ( .A(n15111), .B(n15112), .Z(n15108) );
  AND U14743 ( .A(n787), .B(n15107), .Z(n15112) );
  XNOR U14744 ( .A(n15111), .B(n15105), .Z(n15107) );
  XOR U14745 ( .A(n15113), .B(n15114), .Z(n15105) );
  AND U14746 ( .A(n802), .B(n15115), .Z(n15114) );
  XNOR U14747 ( .A(n15116), .B(n15117), .Z(n15111) );
  AND U14748 ( .A(n794), .B(n15118), .Z(n15117) );
  XOR U14749 ( .A(p_input[1114]), .B(n15116), .Z(n15118) );
  XNOR U14750 ( .A(n15119), .B(n15120), .Z(n15116) );
  AND U14751 ( .A(n798), .B(n15115), .Z(n15120) );
  XNOR U14752 ( .A(n15119), .B(n15113), .Z(n15115) );
  XOR U14753 ( .A(n15121), .B(n15122), .Z(n15113) );
  AND U14754 ( .A(n813), .B(n15123), .Z(n15122) );
  XNOR U14755 ( .A(n15124), .B(n15125), .Z(n15119) );
  AND U14756 ( .A(n805), .B(n15126), .Z(n15125) );
  XOR U14757 ( .A(p_input[1130]), .B(n15124), .Z(n15126) );
  XNOR U14758 ( .A(n15127), .B(n15128), .Z(n15124) );
  AND U14759 ( .A(n809), .B(n15123), .Z(n15128) );
  XNOR U14760 ( .A(n15127), .B(n15121), .Z(n15123) );
  XOR U14761 ( .A(n15129), .B(n15130), .Z(n15121) );
  AND U14762 ( .A(n824), .B(n15131), .Z(n15130) );
  XNOR U14763 ( .A(n15132), .B(n15133), .Z(n15127) );
  AND U14764 ( .A(n816), .B(n15134), .Z(n15133) );
  XOR U14765 ( .A(p_input[1146]), .B(n15132), .Z(n15134) );
  XNOR U14766 ( .A(n15135), .B(n15136), .Z(n15132) );
  AND U14767 ( .A(n820), .B(n15131), .Z(n15136) );
  XNOR U14768 ( .A(n15135), .B(n15129), .Z(n15131) );
  XOR U14769 ( .A(n15137), .B(n15138), .Z(n15129) );
  AND U14770 ( .A(n835), .B(n15139), .Z(n15138) );
  XNOR U14771 ( .A(n15140), .B(n15141), .Z(n15135) );
  AND U14772 ( .A(n827), .B(n15142), .Z(n15141) );
  XOR U14773 ( .A(p_input[1162]), .B(n15140), .Z(n15142) );
  XNOR U14774 ( .A(n15143), .B(n15144), .Z(n15140) );
  AND U14775 ( .A(n831), .B(n15139), .Z(n15144) );
  XNOR U14776 ( .A(n15143), .B(n15137), .Z(n15139) );
  XOR U14777 ( .A(n15145), .B(n15146), .Z(n15137) );
  AND U14778 ( .A(n846), .B(n15147), .Z(n15146) );
  XNOR U14779 ( .A(n15148), .B(n15149), .Z(n15143) );
  AND U14780 ( .A(n838), .B(n15150), .Z(n15149) );
  XOR U14781 ( .A(p_input[1178]), .B(n15148), .Z(n15150) );
  XNOR U14782 ( .A(n15151), .B(n15152), .Z(n15148) );
  AND U14783 ( .A(n842), .B(n15147), .Z(n15152) );
  XNOR U14784 ( .A(n15151), .B(n15145), .Z(n15147) );
  XOR U14785 ( .A(n15153), .B(n15154), .Z(n15145) );
  AND U14786 ( .A(n857), .B(n15155), .Z(n15154) );
  XNOR U14787 ( .A(n15156), .B(n15157), .Z(n15151) );
  AND U14788 ( .A(n849), .B(n15158), .Z(n15157) );
  XOR U14789 ( .A(p_input[1194]), .B(n15156), .Z(n15158) );
  XNOR U14790 ( .A(n15159), .B(n15160), .Z(n15156) );
  AND U14791 ( .A(n853), .B(n15155), .Z(n15160) );
  XNOR U14792 ( .A(n15159), .B(n15153), .Z(n15155) );
  XOR U14793 ( .A(n15161), .B(n15162), .Z(n15153) );
  AND U14794 ( .A(n868), .B(n15163), .Z(n15162) );
  XNOR U14795 ( .A(n15164), .B(n15165), .Z(n15159) );
  AND U14796 ( .A(n860), .B(n15166), .Z(n15165) );
  XOR U14797 ( .A(p_input[1210]), .B(n15164), .Z(n15166) );
  XNOR U14798 ( .A(n15167), .B(n15168), .Z(n15164) );
  AND U14799 ( .A(n864), .B(n15163), .Z(n15168) );
  XNOR U14800 ( .A(n15167), .B(n15161), .Z(n15163) );
  XOR U14801 ( .A(n15169), .B(n15170), .Z(n15161) );
  AND U14802 ( .A(n879), .B(n15171), .Z(n15170) );
  XNOR U14803 ( .A(n15172), .B(n15173), .Z(n15167) );
  AND U14804 ( .A(n871), .B(n15174), .Z(n15173) );
  XOR U14805 ( .A(p_input[1226]), .B(n15172), .Z(n15174) );
  XNOR U14806 ( .A(n15175), .B(n15176), .Z(n15172) );
  AND U14807 ( .A(n875), .B(n15171), .Z(n15176) );
  XNOR U14808 ( .A(n15175), .B(n15169), .Z(n15171) );
  XOR U14809 ( .A(n15177), .B(n15178), .Z(n15169) );
  AND U14810 ( .A(n890), .B(n15179), .Z(n15178) );
  XNOR U14811 ( .A(n15180), .B(n15181), .Z(n15175) );
  AND U14812 ( .A(n882), .B(n15182), .Z(n15181) );
  XOR U14813 ( .A(p_input[1242]), .B(n15180), .Z(n15182) );
  XNOR U14814 ( .A(n15183), .B(n15184), .Z(n15180) );
  AND U14815 ( .A(n886), .B(n15179), .Z(n15184) );
  XNOR U14816 ( .A(n15183), .B(n15177), .Z(n15179) );
  XOR U14817 ( .A(n15185), .B(n15186), .Z(n15177) );
  AND U14818 ( .A(n901), .B(n15187), .Z(n15186) );
  XNOR U14819 ( .A(n15188), .B(n15189), .Z(n15183) );
  AND U14820 ( .A(n893), .B(n15190), .Z(n15189) );
  XOR U14821 ( .A(p_input[1258]), .B(n15188), .Z(n15190) );
  XNOR U14822 ( .A(n15191), .B(n15192), .Z(n15188) );
  AND U14823 ( .A(n897), .B(n15187), .Z(n15192) );
  XNOR U14824 ( .A(n15191), .B(n15185), .Z(n15187) );
  XOR U14825 ( .A(n15193), .B(n15194), .Z(n15185) );
  AND U14826 ( .A(n912), .B(n15195), .Z(n15194) );
  XNOR U14827 ( .A(n15196), .B(n15197), .Z(n15191) );
  AND U14828 ( .A(n904), .B(n15198), .Z(n15197) );
  XOR U14829 ( .A(p_input[1274]), .B(n15196), .Z(n15198) );
  XNOR U14830 ( .A(n15199), .B(n15200), .Z(n15196) );
  AND U14831 ( .A(n908), .B(n15195), .Z(n15200) );
  XNOR U14832 ( .A(n15199), .B(n15193), .Z(n15195) );
  XOR U14833 ( .A(n15201), .B(n15202), .Z(n15193) );
  AND U14834 ( .A(n923), .B(n15203), .Z(n15202) );
  XNOR U14835 ( .A(n15204), .B(n15205), .Z(n15199) );
  AND U14836 ( .A(n915), .B(n15206), .Z(n15205) );
  XOR U14837 ( .A(p_input[1290]), .B(n15204), .Z(n15206) );
  XNOR U14838 ( .A(n15207), .B(n15208), .Z(n15204) );
  AND U14839 ( .A(n919), .B(n15203), .Z(n15208) );
  XNOR U14840 ( .A(n15207), .B(n15201), .Z(n15203) );
  XOR U14841 ( .A(n15209), .B(n15210), .Z(n15201) );
  AND U14842 ( .A(n934), .B(n15211), .Z(n15210) );
  XNOR U14843 ( .A(n15212), .B(n15213), .Z(n15207) );
  AND U14844 ( .A(n926), .B(n15214), .Z(n15213) );
  XOR U14845 ( .A(p_input[1306]), .B(n15212), .Z(n15214) );
  XNOR U14846 ( .A(n15215), .B(n15216), .Z(n15212) );
  AND U14847 ( .A(n930), .B(n15211), .Z(n15216) );
  XNOR U14848 ( .A(n15215), .B(n15209), .Z(n15211) );
  XOR U14849 ( .A(n15217), .B(n15218), .Z(n15209) );
  AND U14850 ( .A(n945), .B(n15219), .Z(n15218) );
  XNOR U14851 ( .A(n15220), .B(n15221), .Z(n15215) );
  AND U14852 ( .A(n937), .B(n15222), .Z(n15221) );
  XOR U14853 ( .A(p_input[1322]), .B(n15220), .Z(n15222) );
  XNOR U14854 ( .A(n15223), .B(n15224), .Z(n15220) );
  AND U14855 ( .A(n941), .B(n15219), .Z(n15224) );
  XNOR U14856 ( .A(n15223), .B(n15217), .Z(n15219) );
  XOR U14857 ( .A(n15225), .B(n15226), .Z(n15217) );
  AND U14858 ( .A(n956), .B(n15227), .Z(n15226) );
  XNOR U14859 ( .A(n15228), .B(n15229), .Z(n15223) );
  AND U14860 ( .A(n948), .B(n15230), .Z(n15229) );
  XOR U14861 ( .A(p_input[1338]), .B(n15228), .Z(n15230) );
  XNOR U14862 ( .A(n15231), .B(n15232), .Z(n15228) );
  AND U14863 ( .A(n952), .B(n15227), .Z(n15232) );
  XNOR U14864 ( .A(n15231), .B(n15225), .Z(n15227) );
  XOR U14865 ( .A(n15233), .B(n15234), .Z(n15225) );
  AND U14866 ( .A(n967), .B(n15235), .Z(n15234) );
  XNOR U14867 ( .A(n15236), .B(n15237), .Z(n15231) );
  AND U14868 ( .A(n959), .B(n15238), .Z(n15237) );
  XOR U14869 ( .A(p_input[1354]), .B(n15236), .Z(n15238) );
  XNOR U14870 ( .A(n15239), .B(n15240), .Z(n15236) );
  AND U14871 ( .A(n963), .B(n15235), .Z(n15240) );
  XNOR U14872 ( .A(n15239), .B(n15233), .Z(n15235) );
  XOR U14873 ( .A(n15241), .B(n15242), .Z(n15233) );
  AND U14874 ( .A(n978), .B(n15243), .Z(n15242) );
  XNOR U14875 ( .A(n15244), .B(n15245), .Z(n15239) );
  AND U14876 ( .A(n970), .B(n15246), .Z(n15245) );
  XOR U14877 ( .A(p_input[1370]), .B(n15244), .Z(n15246) );
  XNOR U14878 ( .A(n15247), .B(n15248), .Z(n15244) );
  AND U14879 ( .A(n974), .B(n15243), .Z(n15248) );
  XNOR U14880 ( .A(n15247), .B(n15241), .Z(n15243) );
  XOR U14881 ( .A(n15249), .B(n15250), .Z(n15241) );
  AND U14882 ( .A(n989), .B(n15251), .Z(n15250) );
  XNOR U14883 ( .A(n15252), .B(n15253), .Z(n15247) );
  AND U14884 ( .A(n981), .B(n15254), .Z(n15253) );
  XOR U14885 ( .A(p_input[1386]), .B(n15252), .Z(n15254) );
  XNOR U14886 ( .A(n15255), .B(n15256), .Z(n15252) );
  AND U14887 ( .A(n985), .B(n15251), .Z(n15256) );
  XNOR U14888 ( .A(n15255), .B(n15249), .Z(n15251) );
  XOR U14889 ( .A(n15257), .B(n15258), .Z(n15249) );
  AND U14890 ( .A(n1000), .B(n15259), .Z(n15258) );
  XNOR U14891 ( .A(n15260), .B(n15261), .Z(n15255) );
  AND U14892 ( .A(n992), .B(n15262), .Z(n15261) );
  XOR U14893 ( .A(p_input[1402]), .B(n15260), .Z(n15262) );
  XNOR U14894 ( .A(n15263), .B(n15264), .Z(n15260) );
  AND U14895 ( .A(n996), .B(n15259), .Z(n15264) );
  XNOR U14896 ( .A(n15263), .B(n15257), .Z(n15259) );
  XOR U14897 ( .A(n15265), .B(n15266), .Z(n15257) );
  AND U14898 ( .A(n1011), .B(n15267), .Z(n15266) );
  XNOR U14899 ( .A(n15268), .B(n15269), .Z(n15263) );
  AND U14900 ( .A(n1003), .B(n15270), .Z(n15269) );
  XOR U14901 ( .A(p_input[1418]), .B(n15268), .Z(n15270) );
  XNOR U14902 ( .A(n15271), .B(n15272), .Z(n15268) );
  AND U14903 ( .A(n1007), .B(n15267), .Z(n15272) );
  XNOR U14904 ( .A(n15271), .B(n15265), .Z(n15267) );
  XOR U14905 ( .A(n15273), .B(n15274), .Z(n15265) );
  AND U14906 ( .A(n1022), .B(n15275), .Z(n15274) );
  XNOR U14907 ( .A(n15276), .B(n15277), .Z(n15271) );
  AND U14908 ( .A(n1014), .B(n15278), .Z(n15277) );
  XOR U14909 ( .A(p_input[1434]), .B(n15276), .Z(n15278) );
  XNOR U14910 ( .A(n15279), .B(n15280), .Z(n15276) );
  AND U14911 ( .A(n1018), .B(n15275), .Z(n15280) );
  XNOR U14912 ( .A(n15279), .B(n15273), .Z(n15275) );
  XOR U14913 ( .A(n15281), .B(n15282), .Z(n15273) );
  AND U14914 ( .A(n1033), .B(n15283), .Z(n15282) );
  XNOR U14915 ( .A(n15284), .B(n15285), .Z(n15279) );
  AND U14916 ( .A(n1025), .B(n15286), .Z(n15285) );
  XOR U14917 ( .A(p_input[1450]), .B(n15284), .Z(n15286) );
  XNOR U14918 ( .A(n15287), .B(n15288), .Z(n15284) );
  AND U14919 ( .A(n1029), .B(n15283), .Z(n15288) );
  XNOR U14920 ( .A(n15287), .B(n15281), .Z(n15283) );
  XOR U14921 ( .A(n15289), .B(n15290), .Z(n15281) );
  AND U14922 ( .A(n1044), .B(n15291), .Z(n15290) );
  XNOR U14923 ( .A(n15292), .B(n15293), .Z(n15287) );
  AND U14924 ( .A(n1036), .B(n15294), .Z(n15293) );
  XOR U14925 ( .A(p_input[1466]), .B(n15292), .Z(n15294) );
  XNOR U14926 ( .A(n15295), .B(n15296), .Z(n15292) );
  AND U14927 ( .A(n1040), .B(n15291), .Z(n15296) );
  XNOR U14928 ( .A(n15295), .B(n15289), .Z(n15291) );
  XOR U14929 ( .A(n15297), .B(n15298), .Z(n15289) );
  AND U14930 ( .A(n1055), .B(n15299), .Z(n15298) );
  XNOR U14931 ( .A(n15300), .B(n15301), .Z(n15295) );
  AND U14932 ( .A(n1047), .B(n15302), .Z(n15301) );
  XOR U14933 ( .A(p_input[1482]), .B(n15300), .Z(n15302) );
  XNOR U14934 ( .A(n15303), .B(n15304), .Z(n15300) );
  AND U14935 ( .A(n1051), .B(n15299), .Z(n15304) );
  XNOR U14936 ( .A(n15303), .B(n15297), .Z(n15299) );
  XOR U14937 ( .A(n15305), .B(n15306), .Z(n15297) );
  AND U14938 ( .A(n1066), .B(n15307), .Z(n15306) );
  XNOR U14939 ( .A(n15308), .B(n15309), .Z(n15303) );
  AND U14940 ( .A(n1058), .B(n15310), .Z(n15309) );
  XOR U14941 ( .A(p_input[1498]), .B(n15308), .Z(n15310) );
  XNOR U14942 ( .A(n15311), .B(n15312), .Z(n15308) );
  AND U14943 ( .A(n1062), .B(n15307), .Z(n15312) );
  XNOR U14944 ( .A(n15311), .B(n15305), .Z(n15307) );
  XOR U14945 ( .A(n15313), .B(n15314), .Z(n15305) );
  AND U14946 ( .A(n1077), .B(n15315), .Z(n15314) );
  XNOR U14947 ( .A(n15316), .B(n15317), .Z(n15311) );
  AND U14948 ( .A(n1069), .B(n15318), .Z(n15317) );
  XOR U14949 ( .A(p_input[1514]), .B(n15316), .Z(n15318) );
  XNOR U14950 ( .A(n15319), .B(n15320), .Z(n15316) );
  AND U14951 ( .A(n1073), .B(n15315), .Z(n15320) );
  XNOR U14952 ( .A(n15319), .B(n15313), .Z(n15315) );
  XOR U14953 ( .A(n15321), .B(n15322), .Z(n15313) );
  AND U14954 ( .A(n1088), .B(n15323), .Z(n15322) );
  XNOR U14955 ( .A(n15324), .B(n15325), .Z(n15319) );
  AND U14956 ( .A(n1080), .B(n15326), .Z(n15325) );
  XOR U14957 ( .A(p_input[1530]), .B(n15324), .Z(n15326) );
  XNOR U14958 ( .A(n15327), .B(n15328), .Z(n15324) );
  AND U14959 ( .A(n1084), .B(n15323), .Z(n15328) );
  XNOR U14960 ( .A(n15327), .B(n15321), .Z(n15323) );
  XOR U14961 ( .A(n15329), .B(n15330), .Z(n15321) );
  AND U14962 ( .A(n1099), .B(n15331), .Z(n15330) );
  XNOR U14963 ( .A(n15332), .B(n15333), .Z(n15327) );
  AND U14964 ( .A(n1091), .B(n15334), .Z(n15333) );
  XOR U14965 ( .A(p_input[1546]), .B(n15332), .Z(n15334) );
  XNOR U14966 ( .A(n15335), .B(n15336), .Z(n15332) );
  AND U14967 ( .A(n1095), .B(n15331), .Z(n15336) );
  XNOR U14968 ( .A(n15335), .B(n15329), .Z(n15331) );
  XOR U14969 ( .A(n15337), .B(n15338), .Z(n15329) );
  AND U14970 ( .A(n1110), .B(n15339), .Z(n15338) );
  XNOR U14971 ( .A(n15340), .B(n15341), .Z(n15335) );
  AND U14972 ( .A(n1102), .B(n15342), .Z(n15341) );
  XOR U14973 ( .A(p_input[1562]), .B(n15340), .Z(n15342) );
  XNOR U14974 ( .A(n15343), .B(n15344), .Z(n15340) );
  AND U14975 ( .A(n1106), .B(n15339), .Z(n15344) );
  XNOR U14976 ( .A(n15343), .B(n15337), .Z(n15339) );
  XOR U14977 ( .A(n15345), .B(n15346), .Z(n15337) );
  AND U14978 ( .A(n1121), .B(n15347), .Z(n15346) );
  XNOR U14979 ( .A(n15348), .B(n15349), .Z(n15343) );
  AND U14980 ( .A(n1113), .B(n15350), .Z(n15349) );
  XOR U14981 ( .A(p_input[1578]), .B(n15348), .Z(n15350) );
  XNOR U14982 ( .A(n15351), .B(n15352), .Z(n15348) );
  AND U14983 ( .A(n1117), .B(n15347), .Z(n15352) );
  XNOR U14984 ( .A(n15351), .B(n15345), .Z(n15347) );
  XOR U14985 ( .A(n15353), .B(n15354), .Z(n15345) );
  AND U14986 ( .A(n1132), .B(n15355), .Z(n15354) );
  XNOR U14987 ( .A(n15356), .B(n15357), .Z(n15351) );
  AND U14988 ( .A(n1124), .B(n15358), .Z(n15357) );
  XOR U14989 ( .A(p_input[1594]), .B(n15356), .Z(n15358) );
  XNOR U14990 ( .A(n15359), .B(n15360), .Z(n15356) );
  AND U14991 ( .A(n1128), .B(n15355), .Z(n15360) );
  XNOR U14992 ( .A(n15359), .B(n15353), .Z(n15355) );
  XOR U14993 ( .A(n15361), .B(n15362), .Z(n15353) );
  AND U14994 ( .A(n1143), .B(n15363), .Z(n15362) );
  XNOR U14995 ( .A(n15364), .B(n15365), .Z(n15359) );
  AND U14996 ( .A(n1135), .B(n15366), .Z(n15365) );
  XOR U14997 ( .A(p_input[1610]), .B(n15364), .Z(n15366) );
  XNOR U14998 ( .A(n15367), .B(n15368), .Z(n15364) );
  AND U14999 ( .A(n1139), .B(n15363), .Z(n15368) );
  XNOR U15000 ( .A(n15367), .B(n15361), .Z(n15363) );
  XOR U15001 ( .A(n15369), .B(n15370), .Z(n15361) );
  AND U15002 ( .A(n1154), .B(n15371), .Z(n15370) );
  XNOR U15003 ( .A(n15372), .B(n15373), .Z(n15367) );
  AND U15004 ( .A(n1146), .B(n15374), .Z(n15373) );
  XOR U15005 ( .A(p_input[1626]), .B(n15372), .Z(n15374) );
  XNOR U15006 ( .A(n15375), .B(n15376), .Z(n15372) );
  AND U15007 ( .A(n1150), .B(n15371), .Z(n15376) );
  XNOR U15008 ( .A(n15375), .B(n15369), .Z(n15371) );
  XOR U15009 ( .A(n15377), .B(n15378), .Z(n15369) );
  AND U15010 ( .A(n1165), .B(n15379), .Z(n15378) );
  XNOR U15011 ( .A(n15380), .B(n15381), .Z(n15375) );
  AND U15012 ( .A(n1157), .B(n15382), .Z(n15381) );
  XOR U15013 ( .A(p_input[1642]), .B(n15380), .Z(n15382) );
  XNOR U15014 ( .A(n15383), .B(n15384), .Z(n15380) );
  AND U15015 ( .A(n1161), .B(n15379), .Z(n15384) );
  XNOR U15016 ( .A(n15383), .B(n15377), .Z(n15379) );
  XOR U15017 ( .A(n15385), .B(n15386), .Z(n15377) );
  AND U15018 ( .A(n1176), .B(n15387), .Z(n15386) );
  XNOR U15019 ( .A(n15388), .B(n15389), .Z(n15383) );
  AND U15020 ( .A(n1168), .B(n15390), .Z(n15389) );
  XOR U15021 ( .A(p_input[1658]), .B(n15388), .Z(n15390) );
  XNOR U15022 ( .A(n15391), .B(n15392), .Z(n15388) );
  AND U15023 ( .A(n1172), .B(n15387), .Z(n15392) );
  XNOR U15024 ( .A(n15391), .B(n15385), .Z(n15387) );
  XOR U15025 ( .A(n15393), .B(n15394), .Z(n15385) );
  AND U15026 ( .A(n1187), .B(n15395), .Z(n15394) );
  XNOR U15027 ( .A(n15396), .B(n15397), .Z(n15391) );
  AND U15028 ( .A(n1179), .B(n15398), .Z(n15397) );
  XOR U15029 ( .A(p_input[1674]), .B(n15396), .Z(n15398) );
  XNOR U15030 ( .A(n15399), .B(n15400), .Z(n15396) );
  AND U15031 ( .A(n1183), .B(n15395), .Z(n15400) );
  XNOR U15032 ( .A(n15399), .B(n15393), .Z(n15395) );
  XOR U15033 ( .A(n15401), .B(n15402), .Z(n15393) );
  AND U15034 ( .A(n1198), .B(n15403), .Z(n15402) );
  XNOR U15035 ( .A(n15404), .B(n15405), .Z(n15399) );
  AND U15036 ( .A(n1190), .B(n15406), .Z(n15405) );
  XOR U15037 ( .A(p_input[1690]), .B(n15404), .Z(n15406) );
  XNOR U15038 ( .A(n15407), .B(n15408), .Z(n15404) );
  AND U15039 ( .A(n1194), .B(n15403), .Z(n15408) );
  XNOR U15040 ( .A(n15407), .B(n15401), .Z(n15403) );
  XOR U15041 ( .A(n15409), .B(n15410), .Z(n15401) );
  AND U15042 ( .A(n1209), .B(n15411), .Z(n15410) );
  XNOR U15043 ( .A(n15412), .B(n15413), .Z(n15407) );
  AND U15044 ( .A(n1201), .B(n15414), .Z(n15413) );
  XOR U15045 ( .A(p_input[1706]), .B(n15412), .Z(n15414) );
  XNOR U15046 ( .A(n15415), .B(n15416), .Z(n15412) );
  AND U15047 ( .A(n1205), .B(n15411), .Z(n15416) );
  XNOR U15048 ( .A(n15415), .B(n15409), .Z(n15411) );
  XOR U15049 ( .A(n15417), .B(n15418), .Z(n15409) );
  AND U15050 ( .A(n1220), .B(n15419), .Z(n15418) );
  XNOR U15051 ( .A(n15420), .B(n15421), .Z(n15415) );
  AND U15052 ( .A(n1212), .B(n15422), .Z(n15421) );
  XOR U15053 ( .A(p_input[1722]), .B(n15420), .Z(n15422) );
  XNOR U15054 ( .A(n15423), .B(n15424), .Z(n15420) );
  AND U15055 ( .A(n1216), .B(n15419), .Z(n15424) );
  XNOR U15056 ( .A(n15423), .B(n15417), .Z(n15419) );
  XOR U15057 ( .A(n15425), .B(n15426), .Z(n15417) );
  AND U15058 ( .A(n1231), .B(n15427), .Z(n15426) );
  XNOR U15059 ( .A(n15428), .B(n15429), .Z(n15423) );
  AND U15060 ( .A(n1223), .B(n15430), .Z(n15429) );
  XOR U15061 ( .A(p_input[1738]), .B(n15428), .Z(n15430) );
  XNOR U15062 ( .A(n15431), .B(n15432), .Z(n15428) );
  AND U15063 ( .A(n1227), .B(n15427), .Z(n15432) );
  XNOR U15064 ( .A(n15431), .B(n15425), .Z(n15427) );
  XOR U15065 ( .A(n15433), .B(n15434), .Z(n15425) );
  AND U15066 ( .A(n1242), .B(n15435), .Z(n15434) );
  XNOR U15067 ( .A(n15436), .B(n15437), .Z(n15431) );
  AND U15068 ( .A(n1234), .B(n15438), .Z(n15437) );
  XOR U15069 ( .A(p_input[1754]), .B(n15436), .Z(n15438) );
  XNOR U15070 ( .A(n15439), .B(n15440), .Z(n15436) );
  AND U15071 ( .A(n1238), .B(n15435), .Z(n15440) );
  XNOR U15072 ( .A(n15439), .B(n15433), .Z(n15435) );
  XOR U15073 ( .A(n15441), .B(n15442), .Z(n15433) );
  AND U15074 ( .A(n1253), .B(n15443), .Z(n15442) );
  XNOR U15075 ( .A(n15444), .B(n15445), .Z(n15439) );
  AND U15076 ( .A(n1245), .B(n15446), .Z(n15445) );
  XOR U15077 ( .A(p_input[1770]), .B(n15444), .Z(n15446) );
  XNOR U15078 ( .A(n15447), .B(n15448), .Z(n15444) );
  AND U15079 ( .A(n1249), .B(n15443), .Z(n15448) );
  XNOR U15080 ( .A(n15447), .B(n15441), .Z(n15443) );
  XOR U15081 ( .A(n15449), .B(n15450), .Z(n15441) );
  AND U15082 ( .A(n1264), .B(n15451), .Z(n15450) );
  XNOR U15083 ( .A(n15452), .B(n15453), .Z(n15447) );
  AND U15084 ( .A(n1256), .B(n15454), .Z(n15453) );
  XOR U15085 ( .A(p_input[1786]), .B(n15452), .Z(n15454) );
  XNOR U15086 ( .A(n15455), .B(n15456), .Z(n15452) );
  AND U15087 ( .A(n1260), .B(n15451), .Z(n15456) );
  XNOR U15088 ( .A(n15455), .B(n15449), .Z(n15451) );
  XOR U15089 ( .A(n15457), .B(n15458), .Z(n15449) );
  AND U15090 ( .A(n1275), .B(n15459), .Z(n15458) );
  XNOR U15091 ( .A(n15460), .B(n15461), .Z(n15455) );
  AND U15092 ( .A(n1267), .B(n15462), .Z(n15461) );
  XOR U15093 ( .A(p_input[1802]), .B(n15460), .Z(n15462) );
  XNOR U15094 ( .A(n15463), .B(n15464), .Z(n15460) );
  AND U15095 ( .A(n1271), .B(n15459), .Z(n15464) );
  XNOR U15096 ( .A(n15463), .B(n15457), .Z(n15459) );
  XOR U15097 ( .A(n15465), .B(n15466), .Z(n15457) );
  AND U15098 ( .A(n1286), .B(n15467), .Z(n15466) );
  XNOR U15099 ( .A(n15468), .B(n15469), .Z(n15463) );
  AND U15100 ( .A(n1278), .B(n15470), .Z(n15469) );
  XOR U15101 ( .A(p_input[1818]), .B(n15468), .Z(n15470) );
  XNOR U15102 ( .A(n15471), .B(n15472), .Z(n15468) );
  AND U15103 ( .A(n1282), .B(n15467), .Z(n15472) );
  XNOR U15104 ( .A(n15471), .B(n15465), .Z(n15467) );
  XOR U15105 ( .A(n15473), .B(n15474), .Z(n15465) );
  AND U15106 ( .A(n1297), .B(n15475), .Z(n15474) );
  XNOR U15107 ( .A(n15476), .B(n15477), .Z(n15471) );
  AND U15108 ( .A(n1289), .B(n15478), .Z(n15477) );
  XOR U15109 ( .A(p_input[1834]), .B(n15476), .Z(n15478) );
  XNOR U15110 ( .A(n15479), .B(n15480), .Z(n15476) );
  AND U15111 ( .A(n1293), .B(n15475), .Z(n15480) );
  XNOR U15112 ( .A(n15479), .B(n15473), .Z(n15475) );
  XOR U15113 ( .A(n15481), .B(n15482), .Z(n15473) );
  AND U15114 ( .A(n1308), .B(n15483), .Z(n15482) );
  XNOR U15115 ( .A(n15484), .B(n15485), .Z(n15479) );
  AND U15116 ( .A(n1300), .B(n15486), .Z(n15485) );
  XOR U15117 ( .A(p_input[1850]), .B(n15484), .Z(n15486) );
  XNOR U15118 ( .A(n15487), .B(n15488), .Z(n15484) );
  AND U15119 ( .A(n1304), .B(n15483), .Z(n15488) );
  XNOR U15120 ( .A(n15487), .B(n15481), .Z(n15483) );
  XOR U15121 ( .A(n15489), .B(n15490), .Z(n15481) );
  AND U15122 ( .A(n1319), .B(n15491), .Z(n15490) );
  XNOR U15123 ( .A(n15492), .B(n15493), .Z(n15487) );
  AND U15124 ( .A(n1311), .B(n15494), .Z(n15493) );
  XOR U15125 ( .A(p_input[1866]), .B(n15492), .Z(n15494) );
  XNOR U15126 ( .A(n15495), .B(n15496), .Z(n15492) );
  AND U15127 ( .A(n1315), .B(n15491), .Z(n15496) );
  XNOR U15128 ( .A(n15495), .B(n15489), .Z(n15491) );
  XOR U15129 ( .A(n15497), .B(n15498), .Z(n15489) );
  AND U15130 ( .A(n1330), .B(n15499), .Z(n15498) );
  XNOR U15131 ( .A(n15500), .B(n15501), .Z(n15495) );
  AND U15132 ( .A(n1322), .B(n15502), .Z(n15501) );
  XOR U15133 ( .A(p_input[1882]), .B(n15500), .Z(n15502) );
  XNOR U15134 ( .A(n15503), .B(n15504), .Z(n15500) );
  AND U15135 ( .A(n1326), .B(n15499), .Z(n15504) );
  XNOR U15136 ( .A(n15503), .B(n15497), .Z(n15499) );
  XOR U15137 ( .A(n15505), .B(n15506), .Z(n15497) );
  AND U15138 ( .A(n1341), .B(n15507), .Z(n15506) );
  XNOR U15139 ( .A(n15508), .B(n15509), .Z(n15503) );
  AND U15140 ( .A(n1333), .B(n15510), .Z(n15509) );
  XOR U15141 ( .A(p_input[1898]), .B(n15508), .Z(n15510) );
  XNOR U15142 ( .A(n15511), .B(n15512), .Z(n15508) );
  AND U15143 ( .A(n1337), .B(n15507), .Z(n15512) );
  XNOR U15144 ( .A(n15511), .B(n15505), .Z(n15507) );
  XOR U15145 ( .A(n15513), .B(n15514), .Z(n15505) );
  AND U15146 ( .A(n1352), .B(n15515), .Z(n15514) );
  XNOR U15147 ( .A(n15516), .B(n15517), .Z(n15511) );
  AND U15148 ( .A(n1344), .B(n15518), .Z(n15517) );
  XOR U15149 ( .A(p_input[1914]), .B(n15516), .Z(n15518) );
  XNOR U15150 ( .A(n15519), .B(n15520), .Z(n15516) );
  AND U15151 ( .A(n1348), .B(n15515), .Z(n15520) );
  XNOR U15152 ( .A(n15519), .B(n15513), .Z(n15515) );
  XOR U15153 ( .A(n15521), .B(n15522), .Z(n15513) );
  AND U15154 ( .A(n1363), .B(n15523), .Z(n15522) );
  XNOR U15155 ( .A(n15524), .B(n15525), .Z(n15519) );
  AND U15156 ( .A(n1355), .B(n15526), .Z(n15525) );
  XOR U15157 ( .A(p_input[1930]), .B(n15524), .Z(n15526) );
  XNOR U15158 ( .A(n15527), .B(n15528), .Z(n15524) );
  AND U15159 ( .A(n1359), .B(n15523), .Z(n15528) );
  XNOR U15160 ( .A(n15527), .B(n15521), .Z(n15523) );
  XOR U15161 ( .A(n15529), .B(n15530), .Z(n15521) );
  AND U15162 ( .A(n1374), .B(n15531), .Z(n15530) );
  XNOR U15163 ( .A(n15532), .B(n15533), .Z(n15527) );
  AND U15164 ( .A(n1366), .B(n15534), .Z(n15533) );
  XOR U15165 ( .A(p_input[1946]), .B(n15532), .Z(n15534) );
  XNOR U15166 ( .A(n15535), .B(n15536), .Z(n15532) );
  AND U15167 ( .A(n1370), .B(n15531), .Z(n15536) );
  XNOR U15168 ( .A(n15535), .B(n15529), .Z(n15531) );
  XOR U15169 ( .A(n15537), .B(n15538), .Z(n15529) );
  AND U15170 ( .A(n1385), .B(n15539), .Z(n15538) );
  XNOR U15171 ( .A(n15540), .B(n15541), .Z(n15535) );
  AND U15172 ( .A(n1377), .B(n15542), .Z(n15541) );
  XOR U15173 ( .A(p_input[1962]), .B(n15540), .Z(n15542) );
  XNOR U15174 ( .A(n15543), .B(n15544), .Z(n15540) );
  AND U15175 ( .A(n1381), .B(n15539), .Z(n15544) );
  XNOR U15176 ( .A(n15543), .B(n15537), .Z(n15539) );
  XOR U15177 ( .A(n15545), .B(n15546), .Z(n15537) );
  AND U15178 ( .A(n1396), .B(n15547), .Z(n15546) );
  XNOR U15179 ( .A(n15548), .B(n15549), .Z(n15543) );
  AND U15180 ( .A(n1388), .B(n15550), .Z(n15549) );
  XOR U15181 ( .A(p_input[1978]), .B(n15548), .Z(n15550) );
  XNOR U15182 ( .A(n15551), .B(n15552), .Z(n15548) );
  AND U15183 ( .A(n1392), .B(n15547), .Z(n15552) );
  XNOR U15184 ( .A(n15551), .B(n15545), .Z(n15547) );
  XOR U15185 ( .A(n15553), .B(n15554), .Z(n15545) );
  AND U15186 ( .A(n1407), .B(n15555), .Z(n15554) );
  XNOR U15187 ( .A(n15556), .B(n15557), .Z(n15551) );
  AND U15188 ( .A(n1399), .B(n15558), .Z(n15557) );
  XOR U15189 ( .A(p_input[1994]), .B(n15556), .Z(n15558) );
  XNOR U15190 ( .A(n15559), .B(n15560), .Z(n15556) );
  AND U15191 ( .A(n1403), .B(n15555), .Z(n15560) );
  XNOR U15192 ( .A(n15559), .B(n15553), .Z(n15555) );
  XOR U15193 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n15561), .Z(n15553) );
  AND U15194 ( .A(n1417), .B(n15562), .Z(n15561) );
  XNOR U15195 ( .A(n15563), .B(n15564), .Z(n15559) );
  AND U15196 ( .A(n1410), .B(n15565), .Z(n15564) );
  XOR U15197 ( .A(p_input[2010]), .B(n15563), .Z(n15565) );
  XNOR U15198 ( .A(n15566), .B(n15567), .Z(n15563) );
  AND U15199 ( .A(n1414), .B(n15562), .Z(n15567) );
  XOR U15200 ( .A(\knn_comb_/min_val_out[0][10] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n15562) );
  XOR U15201 ( .A(n9509), .B(n15568), .Z(o[0]) );
  AND U15202 ( .A(n30), .B(n15569), .Z(n9509) );
  XOR U15203 ( .A(n9510), .B(n15568), .Z(n15569) );
  XOR U15204 ( .A(n15570), .B(n15571), .Z(n15568) );
  AND U15205 ( .A(n42), .B(n15572), .Z(n15571) );
  XOR U15206 ( .A(n15573), .B(n15574), .Z(n9510) );
  AND U15207 ( .A(n34), .B(n15575), .Z(n15574) );
  XOR U15208 ( .A(p_input[0]), .B(n15573), .Z(n15575) );
  XNOR U15209 ( .A(n15576), .B(n15577), .Z(n15573) );
  AND U15210 ( .A(n38), .B(n15572), .Z(n15577) );
  XNOR U15211 ( .A(n15576), .B(n15570), .Z(n15572) );
  XOR U15212 ( .A(n15578), .B(n15579), .Z(n15570) );
  AND U15213 ( .A(n54), .B(n15580), .Z(n15579) );
  XNOR U15214 ( .A(n15581), .B(n15582), .Z(n15576) );
  AND U15215 ( .A(n46), .B(n15583), .Z(n15582) );
  XOR U15216 ( .A(p_input[16]), .B(n15581), .Z(n15583) );
  XNOR U15217 ( .A(n15584), .B(n15585), .Z(n15581) );
  AND U15218 ( .A(n50), .B(n15580), .Z(n15585) );
  XNOR U15219 ( .A(n15584), .B(n15578), .Z(n15580) );
  XOR U15220 ( .A(n15586), .B(n15587), .Z(n15578) );
  AND U15221 ( .A(n65), .B(n15588), .Z(n15587) );
  XNOR U15222 ( .A(n15589), .B(n15590), .Z(n15584) );
  AND U15223 ( .A(n57), .B(n15591), .Z(n15590) );
  XOR U15224 ( .A(p_input[32]), .B(n15589), .Z(n15591) );
  XNOR U15225 ( .A(n15592), .B(n15593), .Z(n15589) );
  AND U15226 ( .A(n61), .B(n15588), .Z(n15593) );
  XNOR U15227 ( .A(n15592), .B(n15586), .Z(n15588) );
  XOR U15228 ( .A(n15594), .B(n15595), .Z(n15586) );
  AND U15229 ( .A(n76), .B(n15596), .Z(n15595) );
  XNOR U15230 ( .A(n15597), .B(n15598), .Z(n15592) );
  AND U15231 ( .A(n68), .B(n15599), .Z(n15598) );
  XOR U15232 ( .A(p_input[48]), .B(n15597), .Z(n15599) );
  XNOR U15233 ( .A(n15600), .B(n15601), .Z(n15597) );
  AND U15234 ( .A(n72), .B(n15596), .Z(n15601) );
  XNOR U15235 ( .A(n15600), .B(n15594), .Z(n15596) );
  XOR U15236 ( .A(n15602), .B(n15603), .Z(n15594) );
  AND U15237 ( .A(n87), .B(n15604), .Z(n15603) );
  XNOR U15238 ( .A(n15605), .B(n15606), .Z(n15600) );
  AND U15239 ( .A(n79), .B(n15607), .Z(n15606) );
  XOR U15240 ( .A(p_input[64]), .B(n15605), .Z(n15607) );
  XNOR U15241 ( .A(n15608), .B(n15609), .Z(n15605) );
  AND U15242 ( .A(n83), .B(n15604), .Z(n15609) );
  XNOR U15243 ( .A(n15608), .B(n15602), .Z(n15604) );
  XOR U15244 ( .A(n15610), .B(n15611), .Z(n15602) );
  AND U15245 ( .A(n98), .B(n15612), .Z(n15611) );
  XNOR U15246 ( .A(n15613), .B(n15614), .Z(n15608) );
  AND U15247 ( .A(n90), .B(n15615), .Z(n15614) );
  XOR U15248 ( .A(p_input[80]), .B(n15613), .Z(n15615) );
  XNOR U15249 ( .A(n15616), .B(n15617), .Z(n15613) );
  AND U15250 ( .A(n94), .B(n15612), .Z(n15617) );
  XNOR U15251 ( .A(n15616), .B(n15610), .Z(n15612) );
  XOR U15252 ( .A(n15618), .B(n15619), .Z(n15610) );
  AND U15253 ( .A(n109), .B(n15620), .Z(n15619) );
  XNOR U15254 ( .A(n15621), .B(n15622), .Z(n15616) );
  AND U15255 ( .A(n101), .B(n15623), .Z(n15622) );
  XOR U15256 ( .A(p_input[96]), .B(n15621), .Z(n15623) );
  XNOR U15257 ( .A(n15624), .B(n15625), .Z(n15621) );
  AND U15258 ( .A(n105), .B(n15620), .Z(n15625) );
  XNOR U15259 ( .A(n15624), .B(n15618), .Z(n15620) );
  XOR U15260 ( .A(n15626), .B(n15627), .Z(n15618) );
  AND U15261 ( .A(n120), .B(n15628), .Z(n15627) );
  XNOR U15262 ( .A(n15629), .B(n15630), .Z(n15624) );
  AND U15263 ( .A(n112), .B(n15631), .Z(n15630) );
  XOR U15264 ( .A(p_input[112]), .B(n15629), .Z(n15631) );
  XNOR U15265 ( .A(n15632), .B(n15633), .Z(n15629) );
  AND U15266 ( .A(n116), .B(n15628), .Z(n15633) );
  XNOR U15267 ( .A(n15632), .B(n15626), .Z(n15628) );
  XOR U15268 ( .A(n15634), .B(n15635), .Z(n15626) );
  AND U15269 ( .A(n131), .B(n15636), .Z(n15635) );
  XNOR U15270 ( .A(n15637), .B(n15638), .Z(n15632) );
  AND U15271 ( .A(n123), .B(n15639), .Z(n15638) );
  XOR U15272 ( .A(p_input[128]), .B(n15637), .Z(n15639) );
  XNOR U15273 ( .A(n15640), .B(n15641), .Z(n15637) );
  AND U15274 ( .A(n127), .B(n15636), .Z(n15641) );
  XNOR U15275 ( .A(n15640), .B(n15634), .Z(n15636) );
  XOR U15276 ( .A(n15642), .B(n15643), .Z(n15634) );
  AND U15277 ( .A(n142), .B(n15644), .Z(n15643) );
  XNOR U15278 ( .A(n15645), .B(n15646), .Z(n15640) );
  AND U15279 ( .A(n134), .B(n15647), .Z(n15646) );
  XOR U15280 ( .A(p_input[144]), .B(n15645), .Z(n15647) );
  XNOR U15281 ( .A(n15648), .B(n15649), .Z(n15645) );
  AND U15282 ( .A(n138), .B(n15644), .Z(n15649) );
  XNOR U15283 ( .A(n15648), .B(n15642), .Z(n15644) );
  XOR U15284 ( .A(n15650), .B(n15651), .Z(n15642) );
  AND U15285 ( .A(n153), .B(n15652), .Z(n15651) );
  XNOR U15286 ( .A(n15653), .B(n15654), .Z(n15648) );
  AND U15287 ( .A(n145), .B(n15655), .Z(n15654) );
  XOR U15288 ( .A(p_input[160]), .B(n15653), .Z(n15655) );
  XNOR U15289 ( .A(n15656), .B(n15657), .Z(n15653) );
  AND U15290 ( .A(n149), .B(n15652), .Z(n15657) );
  XNOR U15291 ( .A(n15656), .B(n15650), .Z(n15652) );
  XOR U15292 ( .A(n15658), .B(n15659), .Z(n15650) );
  AND U15293 ( .A(n164), .B(n15660), .Z(n15659) );
  XNOR U15294 ( .A(n15661), .B(n15662), .Z(n15656) );
  AND U15295 ( .A(n156), .B(n15663), .Z(n15662) );
  XOR U15296 ( .A(p_input[176]), .B(n15661), .Z(n15663) );
  XNOR U15297 ( .A(n15664), .B(n15665), .Z(n15661) );
  AND U15298 ( .A(n160), .B(n15660), .Z(n15665) );
  XNOR U15299 ( .A(n15664), .B(n15658), .Z(n15660) );
  XOR U15300 ( .A(n15666), .B(n15667), .Z(n15658) );
  AND U15301 ( .A(n175), .B(n15668), .Z(n15667) );
  XNOR U15302 ( .A(n15669), .B(n15670), .Z(n15664) );
  AND U15303 ( .A(n167), .B(n15671), .Z(n15670) );
  XOR U15304 ( .A(p_input[192]), .B(n15669), .Z(n15671) );
  XNOR U15305 ( .A(n15672), .B(n15673), .Z(n15669) );
  AND U15306 ( .A(n171), .B(n15668), .Z(n15673) );
  XNOR U15307 ( .A(n15672), .B(n15666), .Z(n15668) );
  XOR U15308 ( .A(n15674), .B(n15675), .Z(n15666) );
  AND U15309 ( .A(n186), .B(n15676), .Z(n15675) );
  XNOR U15310 ( .A(n15677), .B(n15678), .Z(n15672) );
  AND U15311 ( .A(n178), .B(n15679), .Z(n15678) );
  XOR U15312 ( .A(p_input[208]), .B(n15677), .Z(n15679) );
  XNOR U15313 ( .A(n15680), .B(n15681), .Z(n15677) );
  AND U15314 ( .A(n182), .B(n15676), .Z(n15681) );
  XNOR U15315 ( .A(n15680), .B(n15674), .Z(n15676) );
  XOR U15316 ( .A(n15682), .B(n15683), .Z(n15674) );
  AND U15317 ( .A(n197), .B(n15684), .Z(n15683) );
  XNOR U15318 ( .A(n15685), .B(n15686), .Z(n15680) );
  AND U15319 ( .A(n189), .B(n15687), .Z(n15686) );
  XOR U15320 ( .A(p_input[224]), .B(n15685), .Z(n15687) );
  XNOR U15321 ( .A(n15688), .B(n15689), .Z(n15685) );
  AND U15322 ( .A(n193), .B(n15684), .Z(n15689) );
  XNOR U15323 ( .A(n15688), .B(n15682), .Z(n15684) );
  XOR U15324 ( .A(n15690), .B(n15691), .Z(n15682) );
  AND U15325 ( .A(n208), .B(n15692), .Z(n15691) );
  XNOR U15326 ( .A(n15693), .B(n15694), .Z(n15688) );
  AND U15327 ( .A(n200), .B(n15695), .Z(n15694) );
  XOR U15328 ( .A(p_input[240]), .B(n15693), .Z(n15695) );
  XNOR U15329 ( .A(n15696), .B(n15697), .Z(n15693) );
  AND U15330 ( .A(n204), .B(n15692), .Z(n15697) );
  XNOR U15331 ( .A(n15696), .B(n15690), .Z(n15692) );
  XOR U15332 ( .A(n15698), .B(n15699), .Z(n15690) );
  AND U15333 ( .A(n219), .B(n15700), .Z(n15699) );
  XNOR U15334 ( .A(n15701), .B(n15702), .Z(n15696) );
  AND U15335 ( .A(n211), .B(n15703), .Z(n15702) );
  XOR U15336 ( .A(p_input[256]), .B(n15701), .Z(n15703) );
  XNOR U15337 ( .A(n15704), .B(n15705), .Z(n15701) );
  AND U15338 ( .A(n215), .B(n15700), .Z(n15705) );
  XNOR U15339 ( .A(n15704), .B(n15698), .Z(n15700) );
  XOR U15340 ( .A(n15706), .B(n15707), .Z(n15698) );
  AND U15341 ( .A(n230), .B(n15708), .Z(n15707) );
  XNOR U15342 ( .A(n15709), .B(n15710), .Z(n15704) );
  AND U15343 ( .A(n222), .B(n15711), .Z(n15710) );
  XOR U15344 ( .A(p_input[272]), .B(n15709), .Z(n15711) );
  XNOR U15345 ( .A(n15712), .B(n15713), .Z(n15709) );
  AND U15346 ( .A(n226), .B(n15708), .Z(n15713) );
  XNOR U15347 ( .A(n15712), .B(n15706), .Z(n15708) );
  XOR U15348 ( .A(n15714), .B(n15715), .Z(n15706) );
  AND U15349 ( .A(n241), .B(n15716), .Z(n15715) );
  XNOR U15350 ( .A(n15717), .B(n15718), .Z(n15712) );
  AND U15351 ( .A(n233), .B(n15719), .Z(n15718) );
  XOR U15352 ( .A(p_input[288]), .B(n15717), .Z(n15719) );
  XNOR U15353 ( .A(n15720), .B(n15721), .Z(n15717) );
  AND U15354 ( .A(n237), .B(n15716), .Z(n15721) );
  XNOR U15355 ( .A(n15720), .B(n15714), .Z(n15716) );
  XOR U15356 ( .A(n15722), .B(n15723), .Z(n15714) );
  AND U15357 ( .A(n252), .B(n15724), .Z(n15723) );
  XNOR U15358 ( .A(n15725), .B(n15726), .Z(n15720) );
  AND U15359 ( .A(n244), .B(n15727), .Z(n15726) );
  XOR U15360 ( .A(p_input[304]), .B(n15725), .Z(n15727) );
  XNOR U15361 ( .A(n15728), .B(n15729), .Z(n15725) );
  AND U15362 ( .A(n248), .B(n15724), .Z(n15729) );
  XNOR U15363 ( .A(n15728), .B(n15722), .Z(n15724) );
  XOR U15364 ( .A(n15730), .B(n15731), .Z(n15722) );
  AND U15365 ( .A(n263), .B(n15732), .Z(n15731) );
  XNOR U15366 ( .A(n15733), .B(n15734), .Z(n15728) );
  AND U15367 ( .A(n255), .B(n15735), .Z(n15734) );
  XOR U15368 ( .A(p_input[320]), .B(n15733), .Z(n15735) );
  XNOR U15369 ( .A(n15736), .B(n15737), .Z(n15733) );
  AND U15370 ( .A(n259), .B(n15732), .Z(n15737) );
  XNOR U15371 ( .A(n15736), .B(n15730), .Z(n15732) );
  XOR U15372 ( .A(n15738), .B(n15739), .Z(n15730) );
  AND U15373 ( .A(n274), .B(n15740), .Z(n15739) );
  XNOR U15374 ( .A(n15741), .B(n15742), .Z(n15736) );
  AND U15375 ( .A(n266), .B(n15743), .Z(n15742) );
  XOR U15376 ( .A(p_input[336]), .B(n15741), .Z(n15743) );
  XNOR U15377 ( .A(n15744), .B(n15745), .Z(n15741) );
  AND U15378 ( .A(n270), .B(n15740), .Z(n15745) );
  XNOR U15379 ( .A(n15744), .B(n15738), .Z(n15740) );
  XOR U15380 ( .A(n15746), .B(n15747), .Z(n15738) );
  AND U15381 ( .A(n285), .B(n15748), .Z(n15747) );
  XNOR U15382 ( .A(n15749), .B(n15750), .Z(n15744) );
  AND U15383 ( .A(n277), .B(n15751), .Z(n15750) );
  XOR U15384 ( .A(p_input[352]), .B(n15749), .Z(n15751) );
  XNOR U15385 ( .A(n15752), .B(n15753), .Z(n15749) );
  AND U15386 ( .A(n281), .B(n15748), .Z(n15753) );
  XNOR U15387 ( .A(n15752), .B(n15746), .Z(n15748) );
  XOR U15388 ( .A(n15754), .B(n15755), .Z(n15746) );
  AND U15389 ( .A(n296), .B(n15756), .Z(n15755) );
  XNOR U15390 ( .A(n15757), .B(n15758), .Z(n15752) );
  AND U15391 ( .A(n288), .B(n15759), .Z(n15758) );
  XOR U15392 ( .A(p_input[368]), .B(n15757), .Z(n15759) );
  XNOR U15393 ( .A(n15760), .B(n15761), .Z(n15757) );
  AND U15394 ( .A(n292), .B(n15756), .Z(n15761) );
  XNOR U15395 ( .A(n15760), .B(n15754), .Z(n15756) );
  XOR U15396 ( .A(n15762), .B(n15763), .Z(n15754) );
  AND U15397 ( .A(n307), .B(n15764), .Z(n15763) );
  XNOR U15398 ( .A(n15765), .B(n15766), .Z(n15760) );
  AND U15399 ( .A(n299), .B(n15767), .Z(n15766) );
  XOR U15400 ( .A(p_input[384]), .B(n15765), .Z(n15767) );
  XNOR U15401 ( .A(n15768), .B(n15769), .Z(n15765) );
  AND U15402 ( .A(n303), .B(n15764), .Z(n15769) );
  XNOR U15403 ( .A(n15768), .B(n15762), .Z(n15764) );
  XOR U15404 ( .A(n15770), .B(n15771), .Z(n15762) );
  AND U15405 ( .A(n318), .B(n15772), .Z(n15771) );
  XNOR U15406 ( .A(n15773), .B(n15774), .Z(n15768) );
  AND U15407 ( .A(n310), .B(n15775), .Z(n15774) );
  XOR U15408 ( .A(p_input[400]), .B(n15773), .Z(n15775) );
  XNOR U15409 ( .A(n15776), .B(n15777), .Z(n15773) );
  AND U15410 ( .A(n314), .B(n15772), .Z(n15777) );
  XNOR U15411 ( .A(n15776), .B(n15770), .Z(n15772) );
  XOR U15412 ( .A(n15778), .B(n15779), .Z(n15770) );
  AND U15413 ( .A(n329), .B(n15780), .Z(n15779) );
  XNOR U15414 ( .A(n15781), .B(n15782), .Z(n15776) );
  AND U15415 ( .A(n321), .B(n15783), .Z(n15782) );
  XOR U15416 ( .A(p_input[416]), .B(n15781), .Z(n15783) );
  XNOR U15417 ( .A(n15784), .B(n15785), .Z(n15781) );
  AND U15418 ( .A(n325), .B(n15780), .Z(n15785) );
  XNOR U15419 ( .A(n15784), .B(n15778), .Z(n15780) );
  XOR U15420 ( .A(n15786), .B(n15787), .Z(n15778) );
  AND U15421 ( .A(n340), .B(n15788), .Z(n15787) );
  XNOR U15422 ( .A(n15789), .B(n15790), .Z(n15784) );
  AND U15423 ( .A(n332), .B(n15791), .Z(n15790) );
  XOR U15424 ( .A(p_input[432]), .B(n15789), .Z(n15791) );
  XNOR U15425 ( .A(n15792), .B(n15793), .Z(n15789) );
  AND U15426 ( .A(n336), .B(n15788), .Z(n15793) );
  XNOR U15427 ( .A(n15792), .B(n15786), .Z(n15788) );
  XOR U15428 ( .A(n15794), .B(n15795), .Z(n15786) );
  AND U15429 ( .A(n351), .B(n15796), .Z(n15795) );
  XNOR U15430 ( .A(n15797), .B(n15798), .Z(n15792) );
  AND U15431 ( .A(n343), .B(n15799), .Z(n15798) );
  XOR U15432 ( .A(p_input[448]), .B(n15797), .Z(n15799) );
  XNOR U15433 ( .A(n15800), .B(n15801), .Z(n15797) );
  AND U15434 ( .A(n347), .B(n15796), .Z(n15801) );
  XNOR U15435 ( .A(n15800), .B(n15794), .Z(n15796) );
  XOR U15436 ( .A(n15802), .B(n15803), .Z(n15794) );
  AND U15437 ( .A(n362), .B(n15804), .Z(n15803) );
  XNOR U15438 ( .A(n15805), .B(n15806), .Z(n15800) );
  AND U15439 ( .A(n354), .B(n15807), .Z(n15806) );
  XOR U15440 ( .A(p_input[464]), .B(n15805), .Z(n15807) );
  XNOR U15441 ( .A(n15808), .B(n15809), .Z(n15805) );
  AND U15442 ( .A(n358), .B(n15804), .Z(n15809) );
  XNOR U15443 ( .A(n15808), .B(n15802), .Z(n15804) );
  XOR U15444 ( .A(n15810), .B(n15811), .Z(n15802) );
  AND U15445 ( .A(n373), .B(n15812), .Z(n15811) );
  XNOR U15446 ( .A(n15813), .B(n15814), .Z(n15808) );
  AND U15447 ( .A(n365), .B(n15815), .Z(n15814) );
  XOR U15448 ( .A(p_input[480]), .B(n15813), .Z(n15815) );
  XNOR U15449 ( .A(n15816), .B(n15817), .Z(n15813) );
  AND U15450 ( .A(n369), .B(n15812), .Z(n15817) );
  XNOR U15451 ( .A(n15816), .B(n15810), .Z(n15812) );
  XOR U15452 ( .A(n15818), .B(n15819), .Z(n15810) );
  AND U15453 ( .A(n384), .B(n15820), .Z(n15819) );
  XNOR U15454 ( .A(n15821), .B(n15822), .Z(n15816) );
  AND U15455 ( .A(n376), .B(n15823), .Z(n15822) );
  XOR U15456 ( .A(p_input[496]), .B(n15821), .Z(n15823) );
  XNOR U15457 ( .A(n15824), .B(n15825), .Z(n15821) );
  AND U15458 ( .A(n380), .B(n15820), .Z(n15825) );
  XNOR U15459 ( .A(n15824), .B(n15818), .Z(n15820) );
  XOR U15460 ( .A(n15826), .B(n15827), .Z(n15818) );
  AND U15461 ( .A(n395), .B(n15828), .Z(n15827) );
  XNOR U15462 ( .A(n15829), .B(n15830), .Z(n15824) );
  AND U15463 ( .A(n387), .B(n15831), .Z(n15830) );
  XOR U15464 ( .A(p_input[512]), .B(n15829), .Z(n15831) );
  XNOR U15465 ( .A(n15832), .B(n15833), .Z(n15829) );
  AND U15466 ( .A(n391), .B(n15828), .Z(n15833) );
  XNOR U15467 ( .A(n15832), .B(n15826), .Z(n15828) );
  XOR U15468 ( .A(n15834), .B(n15835), .Z(n15826) );
  AND U15469 ( .A(n406), .B(n15836), .Z(n15835) );
  XNOR U15470 ( .A(n15837), .B(n15838), .Z(n15832) );
  AND U15471 ( .A(n398), .B(n15839), .Z(n15838) );
  XOR U15472 ( .A(p_input[528]), .B(n15837), .Z(n15839) );
  XNOR U15473 ( .A(n15840), .B(n15841), .Z(n15837) );
  AND U15474 ( .A(n402), .B(n15836), .Z(n15841) );
  XNOR U15475 ( .A(n15840), .B(n15834), .Z(n15836) );
  XOR U15476 ( .A(n15842), .B(n15843), .Z(n15834) );
  AND U15477 ( .A(n417), .B(n15844), .Z(n15843) );
  XNOR U15478 ( .A(n15845), .B(n15846), .Z(n15840) );
  AND U15479 ( .A(n409), .B(n15847), .Z(n15846) );
  XOR U15480 ( .A(p_input[544]), .B(n15845), .Z(n15847) );
  XNOR U15481 ( .A(n15848), .B(n15849), .Z(n15845) );
  AND U15482 ( .A(n413), .B(n15844), .Z(n15849) );
  XNOR U15483 ( .A(n15848), .B(n15842), .Z(n15844) );
  XOR U15484 ( .A(n15850), .B(n15851), .Z(n15842) );
  AND U15485 ( .A(n428), .B(n15852), .Z(n15851) );
  XNOR U15486 ( .A(n15853), .B(n15854), .Z(n15848) );
  AND U15487 ( .A(n420), .B(n15855), .Z(n15854) );
  XOR U15488 ( .A(p_input[560]), .B(n15853), .Z(n15855) );
  XNOR U15489 ( .A(n15856), .B(n15857), .Z(n15853) );
  AND U15490 ( .A(n424), .B(n15852), .Z(n15857) );
  XNOR U15491 ( .A(n15856), .B(n15850), .Z(n15852) );
  XOR U15492 ( .A(n15858), .B(n15859), .Z(n15850) );
  AND U15493 ( .A(n439), .B(n15860), .Z(n15859) );
  XNOR U15494 ( .A(n15861), .B(n15862), .Z(n15856) );
  AND U15495 ( .A(n431), .B(n15863), .Z(n15862) );
  XOR U15496 ( .A(p_input[576]), .B(n15861), .Z(n15863) );
  XNOR U15497 ( .A(n15864), .B(n15865), .Z(n15861) );
  AND U15498 ( .A(n435), .B(n15860), .Z(n15865) );
  XNOR U15499 ( .A(n15864), .B(n15858), .Z(n15860) );
  XOR U15500 ( .A(n15866), .B(n15867), .Z(n15858) );
  AND U15501 ( .A(n450), .B(n15868), .Z(n15867) );
  XNOR U15502 ( .A(n15869), .B(n15870), .Z(n15864) );
  AND U15503 ( .A(n442), .B(n15871), .Z(n15870) );
  XOR U15504 ( .A(p_input[592]), .B(n15869), .Z(n15871) );
  XNOR U15505 ( .A(n15872), .B(n15873), .Z(n15869) );
  AND U15506 ( .A(n446), .B(n15868), .Z(n15873) );
  XNOR U15507 ( .A(n15872), .B(n15866), .Z(n15868) );
  XOR U15508 ( .A(n15874), .B(n15875), .Z(n15866) );
  AND U15509 ( .A(n461), .B(n15876), .Z(n15875) );
  XNOR U15510 ( .A(n15877), .B(n15878), .Z(n15872) );
  AND U15511 ( .A(n453), .B(n15879), .Z(n15878) );
  XOR U15512 ( .A(p_input[608]), .B(n15877), .Z(n15879) );
  XNOR U15513 ( .A(n15880), .B(n15881), .Z(n15877) );
  AND U15514 ( .A(n457), .B(n15876), .Z(n15881) );
  XNOR U15515 ( .A(n15880), .B(n15874), .Z(n15876) );
  XOR U15516 ( .A(n15882), .B(n15883), .Z(n15874) );
  AND U15517 ( .A(n472), .B(n15884), .Z(n15883) );
  XNOR U15518 ( .A(n15885), .B(n15886), .Z(n15880) );
  AND U15519 ( .A(n464), .B(n15887), .Z(n15886) );
  XOR U15520 ( .A(p_input[624]), .B(n15885), .Z(n15887) );
  XNOR U15521 ( .A(n15888), .B(n15889), .Z(n15885) );
  AND U15522 ( .A(n468), .B(n15884), .Z(n15889) );
  XNOR U15523 ( .A(n15888), .B(n15882), .Z(n15884) );
  XOR U15524 ( .A(n15890), .B(n15891), .Z(n15882) );
  AND U15525 ( .A(n483), .B(n15892), .Z(n15891) );
  XNOR U15526 ( .A(n15893), .B(n15894), .Z(n15888) );
  AND U15527 ( .A(n475), .B(n15895), .Z(n15894) );
  XOR U15528 ( .A(p_input[640]), .B(n15893), .Z(n15895) );
  XNOR U15529 ( .A(n15896), .B(n15897), .Z(n15893) );
  AND U15530 ( .A(n479), .B(n15892), .Z(n15897) );
  XNOR U15531 ( .A(n15896), .B(n15890), .Z(n15892) );
  XOR U15532 ( .A(n15898), .B(n15899), .Z(n15890) );
  AND U15533 ( .A(n494), .B(n15900), .Z(n15899) );
  XNOR U15534 ( .A(n15901), .B(n15902), .Z(n15896) );
  AND U15535 ( .A(n486), .B(n15903), .Z(n15902) );
  XOR U15536 ( .A(p_input[656]), .B(n15901), .Z(n15903) );
  XNOR U15537 ( .A(n15904), .B(n15905), .Z(n15901) );
  AND U15538 ( .A(n490), .B(n15900), .Z(n15905) );
  XNOR U15539 ( .A(n15904), .B(n15898), .Z(n15900) );
  XOR U15540 ( .A(n15906), .B(n15907), .Z(n15898) );
  AND U15541 ( .A(n505), .B(n15908), .Z(n15907) );
  XNOR U15542 ( .A(n15909), .B(n15910), .Z(n15904) );
  AND U15543 ( .A(n497), .B(n15911), .Z(n15910) );
  XOR U15544 ( .A(p_input[672]), .B(n15909), .Z(n15911) );
  XNOR U15545 ( .A(n15912), .B(n15913), .Z(n15909) );
  AND U15546 ( .A(n501), .B(n15908), .Z(n15913) );
  XNOR U15547 ( .A(n15912), .B(n15906), .Z(n15908) );
  XOR U15548 ( .A(n15914), .B(n15915), .Z(n15906) );
  AND U15549 ( .A(n516), .B(n15916), .Z(n15915) );
  XNOR U15550 ( .A(n15917), .B(n15918), .Z(n15912) );
  AND U15551 ( .A(n508), .B(n15919), .Z(n15918) );
  XOR U15552 ( .A(p_input[688]), .B(n15917), .Z(n15919) );
  XNOR U15553 ( .A(n15920), .B(n15921), .Z(n15917) );
  AND U15554 ( .A(n512), .B(n15916), .Z(n15921) );
  XNOR U15555 ( .A(n15920), .B(n15914), .Z(n15916) );
  XOR U15556 ( .A(n15922), .B(n15923), .Z(n15914) );
  AND U15557 ( .A(n527), .B(n15924), .Z(n15923) );
  XNOR U15558 ( .A(n15925), .B(n15926), .Z(n15920) );
  AND U15559 ( .A(n519), .B(n15927), .Z(n15926) );
  XOR U15560 ( .A(p_input[704]), .B(n15925), .Z(n15927) );
  XNOR U15561 ( .A(n15928), .B(n15929), .Z(n15925) );
  AND U15562 ( .A(n523), .B(n15924), .Z(n15929) );
  XNOR U15563 ( .A(n15928), .B(n15922), .Z(n15924) );
  XOR U15564 ( .A(n15930), .B(n15931), .Z(n15922) );
  AND U15565 ( .A(n538), .B(n15932), .Z(n15931) );
  XNOR U15566 ( .A(n15933), .B(n15934), .Z(n15928) );
  AND U15567 ( .A(n530), .B(n15935), .Z(n15934) );
  XOR U15568 ( .A(p_input[720]), .B(n15933), .Z(n15935) );
  XNOR U15569 ( .A(n15936), .B(n15937), .Z(n15933) );
  AND U15570 ( .A(n534), .B(n15932), .Z(n15937) );
  XNOR U15571 ( .A(n15936), .B(n15930), .Z(n15932) );
  XOR U15572 ( .A(n15938), .B(n15939), .Z(n15930) );
  AND U15573 ( .A(n549), .B(n15940), .Z(n15939) );
  XNOR U15574 ( .A(n15941), .B(n15942), .Z(n15936) );
  AND U15575 ( .A(n541), .B(n15943), .Z(n15942) );
  XOR U15576 ( .A(p_input[736]), .B(n15941), .Z(n15943) );
  XNOR U15577 ( .A(n15944), .B(n15945), .Z(n15941) );
  AND U15578 ( .A(n545), .B(n15940), .Z(n15945) );
  XNOR U15579 ( .A(n15944), .B(n15938), .Z(n15940) );
  XOR U15580 ( .A(n15946), .B(n15947), .Z(n15938) );
  AND U15581 ( .A(n560), .B(n15948), .Z(n15947) );
  XNOR U15582 ( .A(n15949), .B(n15950), .Z(n15944) );
  AND U15583 ( .A(n552), .B(n15951), .Z(n15950) );
  XOR U15584 ( .A(p_input[752]), .B(n15949), .Z(n15951) );
  XNOR U15585 ( .A(n15952), .B(n15953), .Z(n15949) );
  AND U15586 ( .A(n556), .B(n15948), .Z(n15953) );
  XNOR U15587 ( .A(n15952), .B(n15946), .Z(n15948) );
  XOR U15588 ( .A(n15954), .B(n15955), .Z(n15946) );
  AND U15589 ( .A(n571), .B(n15956), .Z(n15955) );
  XNOR U15590 ( .A(n15957), .B(n15958), .Z(n15952) );
  AND U15591 ( .A(n563), .B(n15959), .Z(n15958) );
  XOR U15592 ( .A(p_input[768]), .B(n15957), .Z(n15959) );
  XNOR U15593 ( .A(n15960), .B(n15961), .Z(n15957) );
  AND U15594 ( .A(n567), .B(n15956), .Z(n15961) );
  XNOR U15595 ( .A(n15960), .B(n15954), .Z(n15956) );
  XOR U15596 ( .A(n15962), .B(n15963), .Z(n15954) );
  AND U15597 ( .A(n582), .B(n15964), .Z(n15963) );
  XNOR U15598 ( .A(n15965), .B(n15966), .Z(n15960) );
  AND U15599 ( .A(n574), .B(n15967), .Z(n15966) );
  XOR U15600 ( .A(p_input[784]), .B(n15965), .Z(n15967) );
  XNOR U15601 ( .A(n15968), .B(n15969), .Z(n15965) );
  AND U15602 ( .A(n578), .B(n15964), .Z(n15969) );
  XNOR U15603 ( .A(n15968), .B(n15962), .Z(n15964) );
  XOR U15604 ( .A(n15970), .B(n15971), .Z(n15962) );
  AND U15605 ( .A(n593), .B(n15972), .Z(n15971) );
  XNOR U15606 ( .A(n15973), .B(n15974), .Z(n15968) );
  AND U15607 ( .A(n585), .B(n15975), .Z(n15974) );
  XOR U15608 ( .A(p_input[800]), .B(n15973), .Z(n15975) );
  XNOR U15609 ( .A(n15976), .B(n15977), .Z(n15973) );
  AND U15610 ( .A(n589), .B(n15972), .Z(n15977) );
  XNOR U15611 ( .A(n15976), .B(n15970), .Z(n15972) );
  XOR U15612 ( .A(n15978), .B(n15979), .Z(n15970) );
  AND U15613 ( .A(n604), .B(n15980), .Z(n15979) );
  XNOR U15614 ( .A(n15981), .B(n15982), .Z(n15976) );
  AND U15615 ( .A(n596), .B(n15983), .Z(n15982) );
  XOR U15616 ( .A(p_input[816]), .B(n15981), .Z(n15983) );
  XNOR U15617 ( .A(n15984), .B(n15985), .Z(n15981) );
  AND U15618 ( .A(n600), .B(n15980), .Z(n15985) );
  XNOR U15619 ( .A(n15984), .B(n15978), .Z(n15980) );
  XOR U15620 ( .A(n15986), .B(n15987), .Z(n15978) );
  AND U15621 ( .A(n615), .B(n15988), .Z(n15987) );
  XNOR U15622 ( .A(n15989), .B(n15990), .Z(n15984) );
  AND U15623 ( .A(n607), .B(n15991), .Z(n15990) );
  XOR U15624 ( .A(p_input[832]), .B(n15989), .Z(n15991) );
  XNOR U15625 ( .A(n15992), .B(n15993), .Z(n15989) );
  AND U15626 ( .A(n611), .B(n15988), .Z(n15993) );
  XNOR U15627 ( .A(n15992), .B(n15986), .Z(n15988) );
  XOR U15628 ( .A(n15994), .B(n15995), .Z(n15986) );
  AND U15629 ( .A(n626), .B(n15996), .Z(n15995) );
  XNOR U15630 ( .A(n15997), .B(n15998), .Z(n15992) );
  AND U15631 ( .A(n618), .B(n15999), .Z(n15998) );
  XOR U15632 ( .A(p_input[848]), .B(n15997), .Z(n15999) );
  XNOR U15633 ( .A(n16000), .B(n16001), .Z(n15997) );
  AND U15634 ( .A(n622), .B(n15996), .Z(n16001) );
  XNOR U15635 ( .A(n16000), .B(n15994), .Z(n15996) );
  XOR U15636 ( .A(n16002), .B(n16003), .Z(n15994) );
  AND U15637 ( .A(n637), .B(n16004), .Z(n16003) );
  XNOR U15638 ( .A(n16005), .B(n16006), .Z(n16000) );
  AND U15639 ( .A(n629), .B(n16007), .Z(n16006) );
  XOR U15640 ( .A(p_input[864]), .B(n16005), .Z(n16007) );
  XNOR U15641 ( .A(n16008), .B(n16009), .Z(n16005) );
  AND U15642 ( .A(n633), .B(n16004), .Z(n16009) );
  XNOR U15643 ( .A(n16008), .B(n16002), .Z(n16004) );
  XOR U15644 ( .A(n16010), .B(n16011), .Z(n16002) );
  AND U15645 ( .A(n648), .B(n16012), .Z(n16011) );
  XNOR U15646 ( .A(n16013), .B(n16014), .Z(n16008) );
  AND U15647 ( .A(n640), .B(n16015), .Z(n16014) );
  XOR U15648 ( .A(p_input[880]), .B(n16013), .Z(n16015) );
  XNOR U15649 ( .A(n16016), .B(n16017), .Z(n16013) );
  AND U15650 ( .A(n644), .B(n16012), .Z(n16017) );
  XNOR U15651 ( .A(n16016), .B(n16010), .Z(n16012) );
  XOR U15652 ( .A(n16018), .B(n16019), .Z(n16010) );
  AND U15653 ( .A(n659), .B(n16020), .Z(n16019) );
  XNOR U15654 ( .A(n16021), .B(n16022), .Z(n16016) );
  AND U15655 ( .A(n651), .B(n16023), .Z(n16022) );
  XOR U15656 ( .A(p_input[896]), .B(n16021), .Z(n16023) );
  XNOR U15657 ( .A(n16024), .B(n16025), .Z(n16021) );
  AND U15658 ( .A(n655), .B(n16020), .Z(n16025) );
  XNOR U15659 ( .A(n16024), .B(n16018), .Z(n16020) );
  XOR U15660 ( .A(n16026), .B(n16027), .Z(n16018) );
  AND U15661 ( .A(n670), .B(n16028), .Z(n16027) );
  XNOR U15662 ( .A(n16029), .B(n16030), .Z(n16024) );
  AND U15663 ( .A(n662), .B(n16031), .Z(n16030) );
  XOR U15664 ( .A(p_input[912]), .B(n16029), .Z(n16031) );
  XNOR U15665 ( .A(n16032), .B(n16033), .Z(n16029) );
  AND U15666 ( .A(n666), .B(n16028), .Z(n16033) );
  XNOR U15667 ( .A(n16032), .B(n16026), .Z(n16028) );
  XOR U15668 ( .A(n16034), .B(n16035), .Z(n16026) );
  AND U15669 ( .A(n681), .B(n16036), .Z(n16035) );
  XNOR U15670 ( .A(n16037), .B(n16038), .Z(n16032) );
  AND U15671 ( .A(n673), .B(n16039), .Z(n16038) );
  XOR U15672 ( .A(p_input[928]), .B(n16037), .Z(n16039) );
  XNOR U15673 ( .A(n16040), .B(n16041), .Z(n16037) );
  AND U15674 ( .A(n677), .B(n16036), .Z(n16041) );
  XNOR U15675 ( .A(n16040), .B(n16034), .Z(n16036) );
  XOR U15676 ( .A(n16042), .B(n16043), .Z(n16034) );
  AND U15677 ( .A(n692), .B(n16044), .Z(n16043) );
  XNOR U15678 ( .A(n16045), .B(n16046), .Z(n16040) );
  AND U15679 ( .A(n684), .B(n16047), .Z(n16046) );
  XOR U15680 ( .A(p_input[944]), .B(n16045), .Z(n16047) );
  XNOR U15681 ( .A(n16048), .B(n16049), .Z(n16045) );
  AND U15682 ( .A(n688), .B(n16044), .Z(n16049) );
  XNOR U15683 ( .A(n16048), .B(n16042), .Z(n16044) );
  XOR U15684 ( .A(n16050), .B(n16051), .Z(n16042) );
  AND U15685 ( .A(n703), .B(n16052), .Z(n16051) );
  XNOR U15686 ( .A(n16053), .B(n16054), .Z(n16048) );
  AND U15687 ( .A(n695), .B(n16055), .Z(n16054) );
  XOR U15688 ( .A(p_input[960]), .B(n16053), .Z(n16055) );
  XNOR U15689 ( .A(n16056), .B(n16057), .Z(n16053) );
  AND U15690 ( .A(n699), .B(n16052), .Z(n16057) );
  XNOR U15691 ( .A(n16056), .B(n16050), .Z(n16052) );
  XOR U15692 ( .A(n16058), .B(n16059), .Z(n16050) );
  AND U15693 ( .A(n714), .B(n16060), .Z(n16059) );
  XNOR U15694 ( .A(n16061), .B(n16062), .Z(n16056) );
  AND U15695 ( .A(n706), .B(n16063), .Z(n16062) );
  XOR U15696 ( .A(p_input[976]), .B(n16061), .Z(n16063) );
  XNOR U15697 ( .A(n16064), .B(n16065), .Z(n16061) );
  AND U15698 ( .A(n710), .B(n16060), .Z(n16065) );
  XNOR U15699 ( .A(n16064), .B(n16058), .Z(n16060) );
  XOR U15700 ( .A(n16066), .B(n16067), .Z(n16058) );
  AND U15701 ( .A(n725), .B(n16068), .Z(n16067) );
  XNOR U15702 ( .A(n16069), .B(n16070), .Z(n16064) );
  AND U15703 ( .A(n717), .B(n16071), .Z(n16070) );
  XOR U15704 ( .A(p_input[992]), .B(n16069), .Z(n16071) );
  XNOR U15705 ( .A(n16072), .B(n16073), .Z(n16069) );
  AND U15706 ( .A(n721), .B(n16068), .Z(n16073) );
  XNOR U15707 ( .A(n16072), .B(n16066), .Z(n16068) );
  XOR U15708 ( .A(n16074), .B(n16075), .Z(n16066) );
  AND U15709 ( .A(n736), .B(n16076), .Z(n16075) );
  XNOR U15710 ( .A(n16077), .B(n16078), .Z(n16072) );
  AND U15711 ( .A(n728), .B(n16079), .Z(n16078) );
  XOR U15712 ( .A(p_input[1008]), .B(n16077), .Z(n16079) );
  XNOR U15713 ( .A(n16080), .B(n16081), .Z(n16077) );
  AND U15714 ( .A(n732), .B(n16076), .Z(n16081) );
  XNOR U15715 ( .A(n16080), .B(n16074), .Z(n16076) );
  XOR U15716 ( .A(n16082), .B(n16083), .Z(n16074) );
  AND U15717 ( .A(n747), .B(n16084), .Z(n16083) );
  XNOR U15718 ( .A(n16085), .B(n16086), .Z(n16080) );
  AND U15719 ( .A(n739), .B(n16087), .Z(n16086) );
  XOR U15720 ( .A(p_input[1024]), .B(n16085), .Z(n16087) );
  XNOR U15721 ( .A(n16088), .B(n16089), .Z(n16085) );
  AND U15722 ( .A(n743), .B(n16084), .Z(n16089) );
  XNOR U15723 ( .A(n16088), .B(n16082), .Z(n16084) );
  XOR U15724 ( .A(n16090), .B(n16091), .Z(n16082) );
  AND U15725 ( .A(n758), .B(n16092), .Z(n16091) );
  XNOR U15726 ( .A(n16093), .B(n16094), .Z(n16088) );
  AND U15727 ( .A(n750), .B(n16095), .Z(n16094) );
  XOR U15728 ( .A(p_input[1040]), .B(n16093), .Z(n16095) );
  XNOR U15729 ( .A(n16096), .B(n16097), .Z(n16093) );
  AND U15730 ( .A(n754), .B(n16092), .Z(n16097) );
  XNOR U15731 ( .A(n16096), .B(n16090), .Z(n16092) );
  XOR U15732 ( .A(n16098), .B(n16099), .Z(n16090) );
  AND U15733 ( .A(n769), .B(n16100), .Z(n16099) );
  XNOR U15734 ( .A(n16101), .B(n16102), .Z(n16096) );
  AND U15735 ( .A(n761), .B(n16103), .Z(n16102) );
  XOR U15736 ( .A(p_input[1056]), .B(n16101), .Z(n16103) );
  XNOR U15737 ( .A(n16104), .B(n16105), .Z(n16101) );
  AND U15738 ( .A(n765), .B(n16100), .Z(n16105) );
  XNOR U15739 ( .A(n16104), .B(n16098), .Z(n16100) );
  XOR U15740 ( .A(n16106), .B(n16107), .Z(n16098) );
  AND U15741 ( .A(n780), .B(n16108), .Z(n16107) );
  XNOR U15742 ( .A(n16109), .B(n16110), .Z(n16104) );
  AND U15743 ( .A(n772), .B(n16111), .Z(n16110) );
  XOR U15744 ( .A(p_input[1072]), .B(n16109), .Z(n16111) );
  XNOR U15745 ( .A(n16112), .B(n16113), .Z(n16109) );
  AND U15746 ( .A(n776), .B(n16108), .Z(n16113) );
  XNOR U15747 ( .A(n16112), .B(n16106), .Z(n16108) );
  XOR U15748 ( .A(n16114), .B(n16115), .Z(n16106) );
  AND U15749 ( .A(n791), .B(n16116), .Z(n16115) );
  XNOR U15750 ( .A(n16117), .B(n16118), .Z(n16112) );
  AND U15751 ( .A(n783), .B(n16119), .Z(n16118) );
  XOR U15752 ( .A(p_input[1088]), .B(n16117), .Z(n16119) );
  XNOR U15753 ( .A(n16120), .B(n16121), .Z(n16117) );
  AND U15754 ( .A(n787), .B(n16116), .Z(n16121) );
  XNOR U15755 ( .A(n16120), .B(n16114), .Z(n16116) );
  XOR U15756 ( .A(n16122), .B(n16123), .Z(n16114) );
  AND U15757 ( .A(n802), .B(n16124), .Z(n16123) );
  XNOR U15758 ( .A(n16125), .B(n16126), .Z(n16120) );
  AND U15759 ( .A(n794), .B(n16127), .Z(n16126) );
  XOR U15760 ( .A(p_input[1104]), .B(n16125), .Z(n16127) );
  XNOR U15761 ( .A(n16128), .B(n16129), .Z(n16125) );
  AND U15762 ( .A(n798), .B(n16124), .Z(n16129) );
  XNOR U15763 ( .A(n16128), .B(n16122), .Z(n16124) );
  XOR U15764 ( .A(n16130), .B(n16131), .Z(n16122) );
  AND U15765 ( .A(n813), .B(n16132), .Z(n16131) );
  XNOR U15766 ( .A(n16133), .B(n16134), .Z(n16128) );
  AND U15767 ( .A(n805), .B(n16135), .Z(n16134) );
  XOR U15768 ( .A(p_input[1120]), .B(n16133), .Z(n16135) );
  XNOR U15769 ( .A(n16136), .B(n16137), .Z(n16133) );
  AND U15770 ( .A(n809), .B(n16132), .Z(n16137) );
  XNOR U15771 ( .A(n16136), .B(n16130), .Z(n16132) );
  XOR U15772 ( .A(n16138), .B(n16139), .Z(n16130) );
  AND U15773 ( .A(n824), .B(n16140), .Z(n16139) );
  XNOR U15774 ( .A(n16141), .B(n16142), .Z(n16136) );
  AND U15775 ( .A(n816), .B(n16143), .Z(n16142) );
  XOR U15776 ( .A(p_input[1136]), .B(n16141), .Z(n16143) );
  XNOR U15777 ( .A(n16144), .B(n16145), .Z(n16141) );
  AND U15778 ( .A(n820), .B(n16140), .Z(n16145) );
  XNOR U15779 ( .A(n16144), .B(n16138), .Z(n16140) );
  XOR U15780 ( .A(n16146), .B(n16147), .Z(n16138) );
  AND U15781 ( .A(n835), .B(n16148), .Z(n16147) );
  XNOR U15782 ( .A(n16149), .B(n16150), .Z(n16144) );
  AND U15783 ( .A(n827), .B(n16151), .Z(n16150) );
  XOR U15784 ( .A(p_input[1152]), .B(n16149), .Z(n16151) );
  XNOR U15785 ( .A(n16152), .B(n16153), .Z(n16149) );
  AND U15786 ( .A(n831), .B(n16148), .Z(n16153) );
  XNOR U15787 ( .A(n16152), .B(n16146), .Z(n16148) );
  XOR U15788 ( .A(n16154), .B(n16155), .Z(n16146) );
  AND U15789 ( .A(n846), .B(n16156), .Z(n16155) );
  XNOR U15790 ( .A(n16157), .B(n16158), .Z(n16152) );
  AND U15791 ( .A(n838), .B(n16159), .Z(n16158) );
  XOR U15792 ( .A(p_input[1168]), .B(n16157), .Z(n16159) );
  XNOR U15793 ( .A(n16160), .B(n16161), .Z(n16157) );
  AND U15794 ( .A(n842), .B(n16156), .Z(n16161) );
  XNOR U15795 ( .A(n16160), .B(n16154), .Z(n16156) );
  XOR U15796 ( .A(n16162), .B(n16163), .Z(n16154) );
  AND U15797 ( .A(n857), .B(n16164), .Z(n16163) );
  XNOR U15798 ( .A(n16165), .B(n16166), .Z(n16160) );
  AND U15799 ( .A(n849), .B(n16167), .Z(n16166) );
  XOR U15800 ( .A(p_input[1184]), .B(n16165), .Z(n16167) );
  XNOR U15801 ( .A(n16168), .B(n16169), .Z(n16165) );
  AND U15802 ( .A(n853), .B(n16164), .Z(n16169) );
  XNOR U15803 ( .A(n16168), .B(n16162), .Z(n16164) );
  XOR U15804 ( .A(n16170), .B(n16171), .Z(n16162) );
  AND U15805 ( .A(n868), .B(n16172), .Z(n16171) );
  XNOR U15806 ( .A(n16173), .B(n16174), .Z(n16168) );
  AND U15807 ( .A(n860), .B(n16175), .Z(n16174) );
  XOR U15808 ( .A(p_input[1200]), .B(n16173), .Z(n16175) );
  XNOR U15809 ( .A(n16176), .B(n16177), .Z(n16173) );
  AND U15810 ( .A(n864), .B(n16172), .Z(n16177) );
  XNOR U15811 ( .A(n16176), .B(n16170), .Z(n16172) );
  XOR U15812 ( .A(n16178), .B(n16179), .Z(n16170) );
  AND U15813 ( .A(n879), .B(n16180), .Z(n16179) );
  XNOR U15814 ( .A(n16181), .B(n16182), .Z(n16176) );
  AND U15815 ( .A(n871), .B(n16183), .Z(n16182) );
  XOR U15816 ( .A(p_input[1216]), .B(n16181), .Z(n16183) );
  XNOR U15817 ( .A(n16184), .B(n16185), .Z(n16181) );
  AND U15818 ( .A(n875), .B(n16180), .Z(n16185) );
  XNOR U15819 ( .A(n16184), .B(n16178), .Z(n16180) );
  XOR U15820 ( .A(n16186), .B(n16187), .Z(n16178) );
  AND U15821 ( .A(n890), .B(n16188), .Z(n16187) );
  XNOR U15822 ( .A(n16189), .B(n16190), .Z(n16184) );
  AND U15823 ( .A(n882), .B(n16191), .Z(n16190) );
  XOR U15824 ( .A(p_input[1232]), .B(n16189), .Z(n16191) );
  XNOR U15825 ( .A(n16192), .B(n16193), .Z(n16189) );
  AND U15826 ( .A(n886), .B(n16188), .Z(n16193) );
  XNOR U15827 ( .A(n16192), .B(n16186), .Z(n16188) );
  XOR U15828 ( .A(n16194), .B(n16195), .Z(n16186) );
  AND U15829 ( .A(n901), .B(n16196), .Z(n16195) );
  XNOR U15830 ( .A(n16197), .B(n16198), .Z(n16192) );
  AND U15831 ( .A(n893), .B(n16199), .Z(n16198) );
  XOR U15832 ( .A(p_input[1248]), .B(n16197), .Z(n16199) );
  XNOR U15833 ( .A(n16200), .B(n16201), .Z(n16197) );
  AND U15834 ( .A(n897), .B(n16196), .Z(n16201) );
  XNOR U15835 ( .A(n16200), .B(n16194), .Z(n16196) );
  XOR U15836 ( .A(n16202), .B(n16203), .Z(n16194) );
  AND U15837 ( .A(n912), .B(n16204), .Z(n16203) );
  XNOR U15838 ( .A(n16205), .B(n16206), .Z(n16200) );
  AND U15839 ( .A(n904), .B(n16207), .Z(n16206) );
  XOR U15840 ( .A(p_input[1264]), .B(n16205), .Z(n16207) );
  XNOR U15841 ( .A(n16208), .B(n16209), .Z(n16205) );
  AND U15842 ( .A(n908), .B(n16204), .Z(n16209) );
  XNOR U15843 ( .A(n16208), .B(n16202), .Z(n16204) );
  XOR U15844 ( .A(n16210), .B(n16211), .Z(n16202) );
  AND U15845 ( .A(n923), .B(n16212), .Z(n16211) );
  XNOR U15846 ( .A(n16213), .B(n16214), .Z(n16208) );
  AND U15847 ( .A(n915), .B(n16215), .Z(n16214) );
  XOR U15848 ( .A(p_input[1280]), .B(n16213), .Z(n16215) );
  XNOR U15849 ( .A(n16216), .B(n16217), .Z(n16213) );
  AND U15850 ( .A(n919), .B(n16212), .Z(n16217) );
  XNOR U15851 ( .A(n16216), .B(n16210), .Z(n16212) );
  XOR U15852 ( .A(n16218), .B(n16219), .Z(n16210) );
  AND U15853 ( .A(n934), .B(n16220), .Z(n16219) );
  XNOR U15854 ( .A(n16221), .B(n16222), .Z(n16216) );
  AND U15855 ( .A(n926), .B(n16223), .Z(n16222) );
  XOR U15856 ( .A(p_input[1296]), .B(n16221), .Z(n16223) );
  XNOR U15857 ( .A(n16224), .B(n16225), .Z(n16221) );
  AND U15858 ( .A(n930), .B(n16220), .Z(n16225) );
  XNOR U15859 ( .A(n16224), .B(n16218), .Z(n16220) );
  XOR U15860 ( .A(n16226), .B(n16227), .Z(n16218) );
  AND U15861 ( .A(n945), .B(n16228), .Z(n16227) );
  XNOR U15862 ( .A(n16229), .B(n16230), .Z(n16224) );
  AND U15863 ( .A(n937), .B(n16231), .Z(n16230) );
  XOR U15864 ( .A(p_input[1312]), .B(n16229), .Z(n16231) );
  XNOR U15865 ( .A(n16232), .B(n16233), .Z(n16229) );
  AND U15866 ( .A(n941), .B(n16228), .Z(n16233) );
  XNOR U15867 ( .A(n16232), .B(n16226), .Z(n16228) );
  XOR U15868 ( .A(n16234), .B(n16235), .Z(n16226) );
  AND U15869 ( .A(n956), .B(n16236), .Z(n16235) );
  XNOR U15870 ( .A(n16237), .B(n16238), .Z(n16232) );
  AND U15871 ( .A(n948), .B(n16239), .Z(n16238) );
  XOR U15872 ( .A(p_input[1328]), .B(n16237), .Z(n16239) );
  XNOR U15873 ( .A(n16240), .B(n16241), .Z(n16237) );
  AND U15874 ( .A(n952), .B(n16236), .Z(n16241) );
  XNOR U15875 ( .A(n16240), .B(n16234), .Z(n16236) );
  XOR U15876 ( .A(n16242), .B(n16243), .Z(n16234) );
  AND U15877 ( .A(n967), .B(n16244), .Z(n16243) );
  XNOR U15878 ( .A(n16245), .B(n16246), .Z(n16240) );
  AND U15879 ( .A(n959), .B(n16247), .Z(n16246) );
  XOR U15880 ( .A(p_input[1344]), .B(n16245), .Z(n16247) );
  XNOR U15881 ( .A(n16248), .B(n16249), .Z(n16245) );
  AND U15882 ( .A(n963), .B(n16244), .Z(n16249) );
  XNOR U15883 ( .A(n16248), .B(n16242), .Z(n16244) );
  XOR U15884 ( .A(n16250), .B(n16251), .Z(n16242) );
  AND U15885 ( .A(n978), .B(n16252), .Z(n16251) );
  XNOR U15886 ( .A(n16253), .B(n16254), .Z(n16248) );
  AND U15887 ( .A(n970), .B(n16255), .Z(n16254) );
  XOR U15888 ( .A(p_input[1360]), .B(n16253), .Z(n16255) );
  XNOR U15889 ( .A(n16256), .B(n16257), .Z(n16253) );
  AND U15890 ( .A(n974), .B(n16252), .Z(n16257) );
  XNOR U15891 ( .A(n16256), .B(n16250), .Z(n16252) );
  XOR U15892 ( .A(n16258), .B(n16259), .Z(n16250) );
  AND U15893 ( .A(n989), .B(n16260), .Z(n16259) );
  XNOR U15894 ( .A(n16261), .B(n16262), .Z(n16256) );
  AND U15895 ( .A(n981), .B(n16263), .Z(n16262) );
  XOR U15896 ( .A(p_input[1376]), .B(n16261), .Z(n16263) );
  XNOR U15897 ( .A(n16264), .B(n16265), .Z(n16261) );
  AND U15898 ( .A(n985), .B(n16260), .Z(n16265) );
  XNOR U15899 ( .A(n16264), .B(n16258), .Z(n16260) );
  XOR U15900 ( .A(n16266), .B(n16267), .Z(n16258) );
  AND U15901 ( .A(n1000), .B(n16268), .Z(n16267) );
  XNOR U15902 ( .A(n16269), .B(n16270), .Z(n16264) );
  AND U15903 ( .A(n992), .B(n16271), .Z(n16270) );
  XOR U15904 ( .A(p_input[1392]), .B(n16269), .Z(n16271) );
  XNOR U15905 ( .A(n16272), .B(n16273), .Z(n16269) );
  AND U15906 ( .A(n996), .B(n16268), .Z(n16273) );
  XNOR U15907 ( .A(n16272), .B(n16266), .Z(n16268) );
  XOR U15908 ( .A(n16274), .B(n16275), .Z(n16266) );
  AND U15909 ( .A(n1011), .B(n16276), .Z(n16275) );
  XNOR U15910 ( .A(n16277), .B(n16278), .Z(n16272) );
  AND U15911 ( .A(n1003), .B(n16279), .Z(n16278) );
  XOR U15912 ( .A(p_input[1408]), .B(n16277), .Z(n16279) );
  XNOR U15913 ( .A(n16280), .B(n16281), .Z(n16277) );
  AND U15914 ( .A(n1007), .B(n16276), .Z(n16281) );
  XNOR U15915 ( .A(n16280), .B(n16274), .Z(n16276) );
  XOR U15916 ( .A(n16282), .B(n16283), .Z(n16274) );
  AND U15917 ( .A(n1022), .B(n16284), .Z(n16283) );
  XNOR U15918 ( .A(n16285), .B(n16286), .Z(n16280) );
  AND U15919 ( .A(n1014), .B(n16287), .Z(n16286) );
  XOR U15920 ( .A(p_input[1424]), .B(n16285), .Z(n16287) );
  XNOR U15921 ( .A(n16288), .B(n16289), .Z(n16285) );
  AND U15922 ( .A(n1018), .B(n16284), .Z(n16289) );
  XNOR U15923 ( .A(n16288), .B(n16282), .Z(n16284) );
  XOR U15924 ( .A(n16290), .B(n16291), .Z(n16282) );
  AND U15925 ( .A(n1033), .B(n16292), .Z(n16291) );
  XNOR U15926 ( .A(n16293), .B(n16294), .Z(n16288) );
  AND U15927 ( .A(n1025), .B(n16295), .Z(n16294) );
  XOR U15928 ( .A(p_input[1440]), .B(n16293), .Z(n16295) );
  XNOR U15929 ( .A(n16296), .B(n16297), .Z(n16293) );
  AND U15930 ( .A(n1029), .B(n16292), .Z(n16297) );
  XNOR U15931 ( .A(n16296), .B(n16290), .Z(n16292) );
  XOR U15932 ( .A(n16298), .B(n16299), .Z(n16290) );
  AND U15933 ( .A(n1044), .B(n16300), .Z(n16299) );
  XNOR U15934 ( .A(n16301), .B(n16302), .Z(n16296) );
  AND U15935 ( .A(n1036), .B(n16303), .Z(n16302) );
  XOR U15936 ( .A(p_input[1456]), .B(n16301), .Z(n16303) );
  XNOR U15937 ( .A(n16304), .B(n16305), .Z(n16301) );
  AND U15938 ( .A(n1040), .B(n16300), .Z(n16305) );
  XNOR U15939 ( .A(n16304), .B(n16298), .Z(n16300) );
  XOR U15940 ( .A(n16306), .B(n16307), .Z(n16298) );
  AND U15941 ( .A(n1055), .B(n16308), .Z(n16307) );
  XNOR U15942 ( .A(n16309), .B(n16310), .Z(n16304) );
  AND U15943 ( .A(n1047), .B(n16311), .Z(n16310) );
  XOR U15944 ( .A(p_input[1472]), .B(n16309), .Z(n16311) );
  XNOR U15945 ( .A(n16312), .B(n16313), .Z(n16309) );
  AND U15946 ( .A(n1051), .B(n16308), .Z(n16313) );
  XNOR U15947 ( .A(n16312), .B(n16306), .Z(n16308) );
  XOR U15948 ( .A(n16314), .B(n16315), .Z(n16306) );
  AND U15949 ( .A(n1066), .B(n16316), .Z(n16315) );
  XNOR U15950 ( .A(n16317), .B(n16318), .Z(n16312) );
  AND U15951 ( .A(n1058), .B(n16319), .Z(n16318) );
  XOR U15952 ( .A(p_input[1488]), .B(n16317), .Z(n16319) );
  XNOR U15953 ( .A(n16320), .B(n16321), .Z(n16317) );
  AND U15954 ( .A(n1062), .B(n16316), .Z(n16321) );
  XNOR U15955 ( .A(n16320), .B(n16314), .Z(n16316) );
  XOR U15956 ( .A(n16322), .B(n16323), .Z(n16314) );
  AND U15957 ( .A(n1077), .B(n16324), .Z(n16323) );
  XNOR U15958 ( .A(n16325), .B(n16326), .Z(n16320) );
  AND U15959 ( .A(n1069), .B(n16327), .Z(n16326) );
  XOR U15960 ( .A(p_input[1504]), .B(n16325), .Z(n16327) );
  XNOR U15961 ( .A(n16328), .B(n16329), .Z(n16325) );
  AND U15962 ( .A(n1073), .B(n16324), .Z(n16329) );
  XNOR U15963 ( .A(n16328), .B(n16322), .Z(n16324) );
  XOR U15964 ( .A(n16330), .B(n16331), .Z(n16322) );
  AND U15965 ( .A(n1088), .B(n16332), .Z(n16331) );
  XNOR U15966 ( .A(n16333), .B(n16334), .Z(n16328) );
  AND U15967 ( .A(n1080), .B(n16335), .Z(n16334) );
  XOR U15968 ( .A(p_input[1520]), .B(n16333), .Z(n16335) );
  XNOR U15969 ( .A(n16336), .B(n16337), .Z(n16333) );
  AND U15970 ( .A(n1084), .B(n16332), .Z(n16337) );
  XNOR U15971 ( .A(n16336), .B(n16330), .Z(n16332) );
  XOR U15972 ( .A(n16338), .B(n16339), .Z(n16330) );
  AND U15973 ( .A(n1099), .B(n16340), .Z(n16339) );
  XNOR U15974 ( .A(n16341), .B(n16342), .Z(n16336) );
  AND U15975 ( .A(n1091), .B(n16343), .Z(n16342) );
  XOR U15976 ( .A(p_input[1536]), .B(n16341), .Z(n16343) );
  XNOR U15977 ( .A(n16344), .B(n16345), .Z(n16341) );
  AND U15978 ( .A(n1095), .B(n16340), .Z(n16345) );
  XNOR U15979 ( .A(n16344), .B(n16338), .Z(n16340) );
  XOR U15980 ( .A(n16346), .B(n16347), .Z(n16338) );
  AND U15981 ( .A(n1110), .B(n16348), .Z(n16347) );
  XNOR U15982 ( .A(n16349), .B(n16350), .Z(n16344) );
  AND U15983 ( .A(n1102), .B(n16351), .Z(n16350) );
  XOR U15984 ( .A(p_input[1552]), .B(n16349), .Z(n16351) );
  XNOR U15985 ( .A(n16352), .B(n16353), .Z(n16349) );
  AND U15986 ( .A(n1106), .B(n16348), .Z(n16353) );
  XNOR U15987 ( .A(n16352), .B(n16346), .Z(n16348) );
  XOR U15988 ( .A(n16354), .B(n16355), .Z(n16346) );
  AND U15989 ( .A(n1121), .B(n16356), .Z(n16355) );
  XNOR U15990 ( .A(n16357), .B(n16358), .Z(n16352) );
  AND U15991 ( .A(n1113), .B(n16359), .Z(n16358) );
  XOR U15992 ( .A(p_input[1568]), .B(n16357), .Z(n16359) );
  XNOR U15993 ( .A(n16360), .B(n16361), .Z(n16357) );
  AND U15994 ( .A(n1117), .B(n16356), .Z(n16361) );
  XNOR U15995 ( .A(n16360), .B(n16354), .Z(n16356) );
  XOR U15996 ( .A(n16362), .B(n16363), .Z(n16354) );
  AND U15997 ( .A(n1132), .B(n16364), .Z(n16363) );
  XNOR U15998 ( .A(n16365), .B(n16366), .Z(n16360) );
  AND U15999 ( .A(n1124), .B(n16367), .Z(n16366) );
  XOR U16000 ( .A(p_input[1584]), .B(n16365), .Z(n16367) );
  XNOR U16001 ( .A(n16368), .B(n16369), .Z(n16365) );
  AND U16002 ( .A(n1128), .B(n16364), .Z(n16369) );
  XNOR U16003 ( .A(n16368), .B(n16362), .Z(n16364) );
  XOR U16004 ( .A(n16370), .B(n16371), .Z(n16362) );
  AND U16005 ( .A(n1143), .B(n16372), .Z(n16371) );
  XNOR U16006 ( .A(n16373), .B(n16374), .Z(n16368) );
  AND U16007 ( .A(n1135), .B(n16375), .Z(n16374) );
  XOR U16008 ( .A(p_input[1600]), .B(n16373), .Z(n16375) );
  XNOR U16009 ( .A(n16376), .B(n16377), .Z(n16373) );
  AND U16010 ( .A(n1139), .B(n16372), .Z(n16377) );
  XNOR U16011 ( .A(n16376), .B(n16370), .Z(n16372) );
  XOR U16012 ( .A(n16378), .B(n16379), .Z(n16370) );
  AND U16013 ( .A(n1154), .B(n16380), .Z(n16379) );
  XNOR U16014 ( .A(n16381), .B(n16382), .Z(n16376) );
  AND U16015 ( .A(n1146), .B(n16383), .Z(n16382) );
  XOR U16016 ( .A(p_input[1616]), .B(n16381), .Z(n16383) );
  XNOR U16017 ( .A(n16384), .B(n16385), .Z(n16381) );
  AND U16018 ( .A(n1150), .B(n16380), .Z(n16385) );
  XNOR U16019 ( .A(n16384), .B(n16378), .Z(n16380) );
  XOR U16020 ( .A(n16386), .B(n16387), .Z(n16378) );
  AND U16021 ( .A(n1165), .B(n16388), .Z(n16387) );
  XNOR U16022 ( .A(n16389), .B(n16390), .Z(n16384) );
  AND U16023 ( .A(n1157), .B(n16391), .Z(n16390) );
  XOR U16024 ( .A(p_input[1632]), .B(n16389), .Z(n16391) );
  XNOR U16025 ( .A(n16392), .B(n16393), .Z(n16389) );
  AND U16026 ( .A(n1161), .B(n16388), .Z(n16393) );
  XNOR U16027 ( .A(n16392), .B(n16386), .Z(n16388) );
  XOR U16028 ( .A(n16394), .B(n16395), .Z(n16386) );
  AND U16029 ( .A(n1176), .B(n16396), .Z(n16395) );
  XNOR U16030 ( .A(n16397), .B(n16398), .Z(n16392) );
  AND U16031 ( .A(n1168), .B(n16399), .Z(n16398) );
  XOR U16032 ( .A(p_input[1648]), .B(n16397), .Z(n16399) );
  XNOR U16033 ( .A(n16400), .B(n16401), .Z(n16397) );
  AND U16034 ( .A(n1172), .B(n16396), .Z(n16401) );
  XNOR U16035 ( .A(n16400), .B(n16394), .Z(n16396) );
  XOR U16036 ( .A(n16402), .B(n16403), .Z(n16394) );
  AND U16037 ( .A(n1187), .B(n16404), .Z(n16403) );
  XNOR U16038 ( .A(n16405), .B(n16406), .Z(n16400) );
  AND U16039 ( .A(n1179), .B(n16407), .Z(n16406) );
  XOR U16040 ( .A(p_input[1664]), .B(n16405), .Z(n16407) );
  XNOR U16041 ( .A(n16408), .B(n16409), .Z(n16405) );
  AND U16042 ( .A(n1183), .B(n16404), .Z(n16409) );
  XNOR U16043 ( .A(n16408), .B(n16402), .Z(n16404) );
  XOR U16044 ( .A(n16410), .B(n16411), .Z(n16402) );
  AND U16045 ( .A(n1198), .B(n16412), .Z(n16411) );
  XNOR U16046 ( .A(n16413), .B(n16414), .Z(n16408) );
  AND U16047 ( .A(n1190), .B(n16415), .Z(n16414) );
  XOR U16048 ( .A(p_input[1680]), .B(n16413), .Z(n16415) );
  XNOR U16049 ( .A(n16416), .B(n16417), .Z(n16413) );
  AND U16050 ( .A(n1194), .B(n16412), .Z(n16417) );
  XNOR U16051 ( .A(n16416), .B(n16410), .Z(n16412) );
  XOR U16052 ( .A(n16418), .B(n16419), .Z(n16410) );
  AND U16053 ( .A(n1209), .B(n16420), .Z(n16419) );
  XNOR U16054 ( .A(n16421), .B(n16422), .Z(n16416) );
  AND U16055 ( .A(n1201), .B(n16423), .Z(n16422) );
  XOR U16056 ( .A(p_input[1696]), .B(n16421), .Z(n16423) );
  XNOR U16057 ( .A(n16424), .B(n16425), .Z(n16421) );
  AND U16058 ( .A(n1205), .B(n16420), .Z(n16425) );
  XNOR U16059 ( .A(n16424), .B(n16418), .Z(n16420) );
  XOR U16060 ( .A(n16426), .B(n16427), .Z(n16418) );
  AND U16061 ( .A(n1220), .B(n16428), .Z(n16427) );
  XNOR U16062 ( .A(n16429), .B(n16430), .Z(n16424) );
  AND U16063 ( .A(n1212), .B(n16431), .Z(n16430) );
  XOR U16064 ( .A(p_input[1712]), .B(n16429), .Z(n16431) );
  XNOR U16065 ( .A(n16432), .B(n16433), .Z(n16429) );
  AND U16066 ( .A(n1216), .B(n16428), .Z(n16433) );
  XNOR U16067 ( .A(n16432), .B(n16426), .Z(n16428) );
  XOR U16068 ( .A(n16434), .B(n16435), .Z(n16426) );
  AND U16069 ( .A(n1231), .B(n16436), .Z(n16435) );
  XNOR U16070 ( .A(n16437), .B(n16438), .Z(n16432) );
  AND U16071 ( .A(n1223), .B(n16439), .Z(n16438) );
  XOR U16072 ( .A(p_input[1728]), .B(n16437), .Z(n16439) );
  XNOR U16073 ( .A(n16440), .B(n16441), .Z(n16437) );
  AND U16074 ( .A(n1227), .B(n16436), .Z(n16441) );
  XNOR U16075 ( .A(n16440), .B(n16434), .Z(n16436) );
  XOR U16076 ( .A(n16442), .B(n16443), .Z(n16434) );
  AND U16077 ( .A(n1242), .B(n16444), .Z(n16443) );
  XNOR U16078 ( .A(n16445), .B(n16446), .Z(n16440) );
  AND U16079 ( .A(n1234), .B(n16447), .Z(n16446) );
  XOR U16080 ( .A(p_input[1744]), .B(n16445), .Z(n16447) );
  XNOR U16081 ( .A(n16448), .B(n16449), .Z(n16445) );
  AND U16082 ( .A(n1238), .B(n16444), .Z(n16449) );
  XNOR U16083 ( .A(n16448), .B(n16442), .Z(n16444) );
  XOR U16084 ( .A(n16450), .B(n16451), .Z(n16442) );
  AND U16085 ( .A(n1253), .B(n16452), .Z(n16451) );
  XNOR U16086 ( .A(n16453), .B(n16454), .Z(n16448) );
  AND U16087 ( .A(n1245), .B(n16455), .Z(n16454) );
  XOR U16088 ( .A(p_input[1760]), .B(n16453), .Z(n16455) );
  XNOR U16089 ( .A(n16456), .B(n16457), .Z(n16453) );
  AND U16090 ( .A(n1249), .B(n16452), .Z(n16457) );
  XNOR U16091 ( .A(n16456), .B(n16450), .Z(n16452) );
  XOR U16092 ( .A(n16458), .B(n16459), .Z(n16450) );
  AND U16093 ( .A(n1264), .B(n16460), .Z(n16459) );
  XNOR U16094 ( .A(n16461), .B(n16462), .Z(n16456) );
  AND U16095 ( .A(n1256), .B(n16463), .Z(n16462) );
  XOR U16096 ( .A(p_input[1776]), .B(n16461), .Z(n16463) );
  XNOR U16097 ( .A(n16464), .B(n16465), .Z(n16461) );
  AND U16098 ( .A(n1260), .B(n16460), .Z(n16465) );
  XNOR U16099 ( .A(n16464), .B(n16458), .Z(n16460) );
  XOR U16100 ( .A(n16466), .B(n16467), .Z(n16458) );
  AND U16101 ( .A(n1275), .B(n16468), .Z(n16467) );
  XNOR U16102 ( .A(n16469), .B(n16470), .Z(n16464) );
  AND U16103 ( .A(n1267), .B(n16471), .Z(n16470) );
  XOR U16104 ( .A(p_input[1792]), .B(n16469), .Z(n16471) );
  XNOR U16105 ( .A(n16472), .B(n16473), .Z(n16469) );
  AND U16106 ( .A(n1271), .B(n16468), .Z(n16473) );
  XNOR U16107 ( .A(n16472), .B(n16466), .Z(n16468) );
  XOR U16108 ( .A(n16474), .B(n16475), .Z(n16466) );
  AND U16109 ( .A(n1286), .B(n16476), .Z(n16475) );
  XNOR U16110 ( .A(n16477), .B(n16478), .Z(n16472) );
  AND U16111 ( .A(n1278), .B(n16479), .Z(n16478) );
  XOR U16112 ( .A(p_input[1808]), .B(n16477), .Z(n16479) );
  XNOR U16113 ( .A(n16480), .B(n16481), .Z(n16477) );
  AND U16114 ( .A(n1282), .B(n16476), .Z(n16481) );
  XNOR U16115 ( .A(n16480), .B(n16474), .Z(n16476) );
  XOR U16116 ( .A(n16482), .B(n16483), .Z(n16474) );
  AND U16117 ( .A(n1297), .B(n16484), .Z(n16483) );
  XNOR U16118 ( .A(n16485), .B(n16486), .Z(n16480) );
  AND U16119 ( .A(n1289), .B(n16487), .Z(n16486) );
  XOR U16120 ( .A(p_input[1824]), .B(n16485), .Z(n16487) );
  XNOR U16121 ( .A(n16488), .B(n16489), .Z(n16485) );
  AND U16122 ( .A(n1293), .B(n16484), .Z(n16489) );
  XNOR U16123 ( .A(n16488), .B(n16482), .Z(n16484) );
  XOR U16124 ( .A(n16490), .B(n16491), .Z(n16482) );
  AND U16125 ( .A(n1308), .B(n16492), .Z(n16491) );
  XNOR U16126 ( .A(n16493), .B(n16494), .Z(n16488) );
  AND U16127 ( .A(n1300), .B(n16495), .Z(n16494) );
  XOR U16128 ( .A(p_input[1840]), .B(n16493), .Z(n16495) );
  XNOR U16129 ( .A(n16496), .B(n16497), .Z(n16493) );
  AND U16130 ( .A(n1304), .B(n16492), .Z(n16497) );
  XNOR U16131 ( .A(n16496), .B(n16490), .Z(n16492) );
  XOR U16132 ( .A(n16498), .B(n16499), .Z(n16490) );
  AND U16133 ( .A(n1319), .B(n16500), .Z(n16499) );
  XNOR U16134 ( .A(n16501), .B(n16502), .Z(n16496) );
  AND U16135 ( .A(n1311), .B(n16503), .Z(n16502) );
  XOR U16136 ( .A(p_input[1856]), .B(n16501), .Z(n16503) );
  XNOR U16137 ( .A(n16504), .B(n16505), .Z(n16501) );
  AND U16138 ( .A(n1315), .B(n16500), .Z(n16505) );
  XNOR U16139 ( .A(n16504), .B(n16498), .Z(n16500) );
  XOR U16140 ( .A(n16506), .B(n16507), .Z(n16498) );
  AND U16141 ( .A(n1330), .B(n16508), .Z(n16507) );
  XNOR U16142 ( .A(n16509), .B(n16510), .Z(n16504) );
  AND U16143 ( .A(n1322), .B(n16511), .Z(n16510) );
  XOR U16144 ( .A(p_input[1872]), .B(n16509), .Z(n16511) );
  XNOR U16145 ( .A(n16512), .B(n16513), .Z(n16509) );
  AND U16146 ( .A(n1326), .B(n16508), .Z(n16513) );
  XNOR U16147 ( .A(n16512), .B(n16506), .Z(n16508) );
  XOR U16148 ( .A(n16514), .B(n16515), .Z(n16506) );
  AND U16149 ( .A(n1341), .B(n16516), .Z(n16515) );
  XNOR U16150 ( .A(n16517), .B(n16518), .Z(n16512) );
  AND U16151 ( .A(n1333), .B(n16519), .Z(n16518) );
  XOR U16152 ( .A(p_input[1888]), .B(n16517), .Z(n16519) );
  XNOR U16153 ( .A(n16520), .B(n16521), .Z(n16517) );
  AND U16154 ( .A(n1337), .B(n16516), .Z(n16521) );
  XNOR U16155 ( .A(n16520), .B(n16514), .Z(n16516) );
  XOR U16156 ( .A(n16522), .B(n16523), .Z(n16514) );
  AND U16157 ( .A(n1352), .B(n16524), .Z(n16523) );
  XNOR U16158 ( .A(n16525), .B(n16526), .Z(n16520) );
  AND U16159 ( .A(n1344), .B(n16527), .Z(n16526) );
  XOR U16160 ( .A(p_input[1904]), .B(n16525), .Z(n16527) );
  XNOR U16161 ( .A(n16528), .B(n16529), .Z(n16525) );
  AND U16162 ( .A(n1348), .B(n16524), .Z(n16529) );
  XNOR U16163 ( .A(n16528), .B(n16522), .Z(n16524) );
  XOR U16164 ( .A(n16530), .B(n16531), .Z(n16522) );
  AND U16165 ( .A(n1363), .B(n16532), .Z(n16531) );
  XNOR U16166 ( .A(n16533), .B(n16534), .Z(n16528) );
  AND U16167 ( .A(n1355), .B(n16535), .Z(n16534) );
  XOR U16168 ( .A(p_input[1920]), .B(n16533), .Z(n16535) );
  XNOR U16169 ( .A(n16536), .B(n16537), .Z(n16533) );
  AND U16170 ( .A(n1359), .B(n16532), .Z(n16537) );
  XNOR U16171 ( .A(n16536), .B(n16530), .Z(n16532) );
  XOR U16172 ( .A(n16538), .B(n16539), .Z(n16530) );
  AND U16173 ( .A(n1374), .B(n16540), .Z(n16539) );
  XNOR U16174 ( .A(n16541), .B(n16542), .Z(n16536) );
  AND U16175 ( .A(n1366), .B(n16543), .Z(n16542) );
  XOR U16176 ( .A(p_input[1936]), .B(n16541), .Z(n16543) );
  XNOR U16177 ( .A(n16544), .B(n16545), .Z(n16541) );
  AND U16178 ( .A(n1370), .B(n16540), .Z(n16545) );
  XNOR U16179 ( .A(n16544), .B(n16538), .Z(n16540) );
  XOR U16180 ( .A(n16546), .B(n16547), .Z(n16538) );
  AND U16181 ( .A(n1385), .B(n16548), .Z(n16547) );
  XNOR U16182 ( .A(n16549), .B(n16550), .Z(n16544) );
  AND U16183 ( .A(n1377), .B(n16551), .Z(n16550) );
  XOR U16184 ( .A(p_input[1952]), .B(n16549), .Z(n16551) );
  XNOR U16185 ( .A(n16552), .B(n16553), .Z(n16549) );
  AND U16186 ( .A(n1381), .B(n16548), .Z(n16553) );
  XNOR U16187 ( .A(n16552), .B(n16546), .Z(n16548) );
  XOR U16188 ( .A(n16554), .B(n16555), .Z(n16546) );
  AND U16189 ( .A(n1396), .B(n16556), .Z(n16555) );
  XNOR U16190 ( .A(n16557), .B(n16558), .Z(n16552) );
  AND U16191 ( .A(n1388), .B(n16559), .Z(n16558) );
  XOR U16192 ( .A(p_input[1968]), .B(n16557), .Z(n16559) );
  XNOR U16193 ( .A(n16560), .B(n16561), .Z(n16557) );
  AND U16194 ( .A(n1392), .B(n16556), .Z(n16561) );
  XNOR U16195 ( .A(n16560), .B(n16554), .Z(n16556) );
  XOR U16196 ( .A(n16562), .B(n16563), .Z(n16554) );
  AND U16197 ( .A(n1407), .B(n16564), .Z(n16563) );
  XNOR U16198 ( .A(n16565), .B(n16566), .Z(n16560) );
  AND U16199 ( .A(n1399), .B(n16567), .Z(n16566) );
  XOR U16200 ( .A(p_input[1984]), .B(n16565), .Z(n16567) );
  XNOR U16201 ( .A(n16568), .B(n16569), .Z(n16565) );
  AND U16202 ( .A(n1403), .B(n16564), .Z(n16569) );
  XNOR U16203 ( .A(n16568), .B(n16562), .Z(n16564) );
  XOR U16204 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n16570), .Z(n16562) );
  AND U16205 ( .A(n1417), .B(n16571), .Z(n16570) );
  XNOR U16206 ( .A(n16572), .B(n16573), .Z(n16568) );
  AND U16207 ( .A(n1410), .B(n16574), .Z(n16573) );
  XOR U16208 ( .A(p_input[2000]), .B(n16572), .Z(n16574) );
  XNOR U16209 ( .A(n16575), .B(n16576), .Z(n16572) );
  AND U16210 ( .A(n1414), .B(n16571), .Z(n16576) );
  XOR U16211 ( .A(\knn_comb_/min_val_out[0][0] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n16571) );
  IV U16212 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n16575) );
  XNOR U16213 ( .A(n16577), .B(n16578), .Z(n30) );
  AND U16214 ( .A(n16579), .B(n16580), .Z(n16578) );
  XNOR U16215 ( .A(n16577), .B(n16581), .Z(n16580) );
  XOR U16216 ( .A(n16582), .B(n16583), .Z(n16581) );
  AND U16217 ( .A(n34), .B(n16584), .Z(n16583) );
  XNOR U16218 ( .A(n16582), .B(n16585), .Z(n16584) );
  XNOR U16219 ( .A(n16577), .B(n16586), .Z(n16579) );
  XOR U16220 ( .A(n16587), .B(n16588), .Z(n16586) );
  AND U16221 ( .A(n42), .B(n16589), .Z(n16588) );
  XOR U16222 ( .A(n16590), .B(n16591), .Z(n16577) );
  AND U16223 ( .A(n16592), .B(n16593), .Z(n16591) );
  XOR U16224 ( .A(n16594), .B(n16590), .Z(n16593) );
  XOR U16225 ( .A(n16595), .B(n16596), .Z(n16594) );
  AND U16226 ( .A(n34), .B(n16597), .Z(n16596) );
  XOR U16227 ( .A(n16598), .B(n16595), .Z(n16597) );
  XNOR U16228 ( .A(n16590), .B(n16599), .Z(n16592) );
  XOR U16229 ( .A(n16600), .B(n16601), .Z(n16599) );
  AND U16230 ( .A(n42), .B(n16602), .Z(n16601) );
  XOR U16231 ( .A(n16603), .B(n16604), .Z(n16590) );
  AND U16232 ( .A(n16605), .B(n16606), .Z(n16604) );
  XOR U16233 ( .A(n16607), .B(n16603), .Z(n16606) );
  XOR U16234 ( .A(n16608), .B(n16609), .Z(n16607) );
  AND U16235 ( .A(n34), .B(n16610), .Z(n16609) );
  XNOR U16236 ( .A(n16611), .B(n16608), .Z(n16610) );
  XNOR U16237 ( .A(n16603), .B(n16612), .Z(n16605) );
  XOR U16238 ( .A(n16613), .B(n16614), .Z(n16612) );
  AND U16239 ( .A(n42), .B(n16615), .Z(n16614) );
  XOR U16240 ( .A(n16616), .B(n16617), .Z(n16603) );
  AND U16241 ( .A(n16618), .B(n16619), .Z(n16617) );
  XOR U16242 ( .A(n16616), .B(n16620), .Z(n16619) );
  XOR U16243 ( .A(n16621), .B(n16622), .Z(n16620) );
  AND U16244 ( .A(n34), .B(n16623), .Z(n16622) );
  XOR U16245 ( .A(n16624), .B(n16621), .Z(n16623) );
  XNOR U16246 ( .A(n16625), .B(n16616), .Z(n16618) );
  XNOR U16247 ( .A(n16626), .B(n16627), .Z(n16625) );
  AND U16248 ( .A(n42), .B(n16628), .Z(n16627) );
  AND U16249 ( .A(n16629), .B(n16630), .Z(n16616) );
  XNOR U16250 ( .A(n16631), .B(n16632), .Z(n16630) );
  AND U16251 ( .A(n34), .B(n16633), .Z(n16632) );
  XNOR U16252 ( .A(n16634), .B(n16631), .Z(n16633) );
  XNOR U16253 ( .A(n16635), .B(n16636), .Z(n34) );
  AND U16254 ( .A(n16637), .B(n16638), .Z(n16636) );
  XOR U16255 ( .A(n16585), .B(n16635), .Z(n16638) );
  AND U16256 ( .A(n16639), .B(n16640), .Z(n16585) );
  XOR U16257 ( .A(n16635), .B(n16582), .Z(n16637) );
  XNOR U16258 ( .A(n16641), .B(n16642), .Z(n16582) );
  AND U16259 ( .A(n38), .B(n16589), .Z(n16642) );
  XOR U16260 ( .A(n16587), .B(n16641), .Z(n16589) );
  XOR U16261 ( .A(n16643), .B(n16644), .Z(n16635) );
  AND U16262 ( .A(n16645), .B(n16646), .Z(n16644) );
  XNOR U16263 ( .A(n16643), .B(n16639), .Z(n16646) );
  IV U16264 ( .A(n16598), .Z(n16639) );
  XOR U16265 ( .A(n16647), .B(n16648), .Z(n16598) );
  XOR U16266 ( .A(n16649), .B(n16640), .Z(n16648) );
  AND U16267 ( .A(n16611), .B(n16650), .Z(n16640) );
  AND U16268 ( .A(n16651), .B(n16652), .Z(n16649) );
  XOR U16269 ( .A(n16653), .B(n16647), .Z(n16651) );
  XNOR U16270 ( .A(n16595), .B(n16643), .Z(n16645) );
  XNOR U16271 ( .A(n16654), .B(n16655), .Z(n16595) );
  AND U16272 ( .A(n38), .B(n16602), .Z(n16655) );
  XOR U16273 ( .A(n16654), .B(n16656), .Z(n16602) );
  XOR U16274 ( .A(n16657), .B(n16658), .Z(n16643) );
  AND U16275 ( .A(n16659), .B(n16660), .Z(n16658) );
  XNOR U16276 ( .A(n16657), .B(n16611), .Z(n16660) );
  XOR U16277 ( .A(n16661), .B(n16652), .Z(n16611) );
  XNOR U16278 ( .A(n16662), .B(n16647), .Z(n16652) );
  XOR U16279 ( .A(n16663), .B(n16664), .Z(n16647) );
  AND U16280 ( .A(n16665), .B(n16666), .Z(n16664) );
  XOR U16281 ( .A(n16667), .B(n16663), .Z(n16665) );
  XNOR U16282 ( .A(n16668), .B(n16669), .Z(n16662) );
  AND U16283 ( .A(n16670), .B(n16671), .Z(n16669) );
  XOR U16284 ( .A(n16668), .B(n16672), .Z(n16670) );
  XNOR U16285 ( .A(n16653), .B(n16650), .Z(n16661) );
  AND U16286 ( .A(n16673), .B(n16674), .Z(n16650) );
  XOR U16287 ( .A(n16675), .B(n16676), .Z(n16653) );
  AND U16288 ( .A(n16677), .B(n16678), .Z(n16676) );
  XOR U16289 ( .A(n16675), .B(n16679), .Z(n16677) );
  XNOR U16290 ( .A(n16608), .B(n16657), .Z(n16659) );
  XNOR U16291 ( .A(n16680), .B(n16681), .Z(n16608) );
  AND U16292 ( .A(n38), .B(n16615), .Z(n16681) );
  XOR U16293 ( .A(n16680), .B(n16682), .Z(n16615) );
  XOR U16294 ( .A(n16683), .B(n16684), .Z(n16657) );
  AND U16295 ( .A(n16685), .B(n16686), .Z(n16684) );
  XNOR U16296 ( .A(n16683), .B(n16673), .Z(n16686) );
  IV U16297 ( .A(n16624), .Z(n16673) );
  XNOR U16298 ( .A(n16687), .B(n16666), .Z(n16624) );
  XNOR U16299 ( .A(n16688), .B(n16672), .Z(n16666) );
  XNOR U16300 ( .A(n16689), .B(n16690), .Z(n16672) );
  NOR U16301 ( .A(n16691), .B(n16692), .Z(n16690) );
  XOR U16302 ( .A(n16689), .B(n16693), .Z(n16691) );
  XNOR U16303 ( .A(n16671), .B(n16663), .Z(n16688) );
  XOR U16304 ( .A(n16694), .B(n16695), .Z(n16663) );
  AND U16305 ( .A(n16696), .B(n16697), .Z(n16695) );
  XNOR U16306 ( .A(n16694), .B(n16698), .Z(n16696) );
  XNOR U16307 ( .A(n16699), .B(n16668), .Z(n16671) );
  XOR U16308 ( .A(n16700), .B(n16701), .Z(n16668) );
  AND U16309 ( .A(n16702), .B(n16703), .Z(n16701) );
  XOR U16310 ( .A(n16700), .B(n16704), .Z(n16702) );
  XNOR U16311 ( .A(n16705), .B(n16706), .Z(n16699) );
  NOR U16312 ( .A(n16707), .B(n16708), .Z(n16706) );
  XNOR U16313 ( .A(n16705), .B(n16709), .Z(n16707) );
  XNOR U16314 ( .A(n16667), .B(n16674), .Z(n16687) );
  NOR U16315 ( .A(n16634), .B(n16710), .Z(n16674) );
  XOR U16316 ( .A(n16679), .B(n16678), .Z(n16667) );
  XNOR U16317 ( .A(n16711), .B(n16675), .Z(n16678) );
  XOR U16318 ( .A(n16712), .B(n16713), .Z(n16675) );
  AND U16319 ( .A(n16714), .B(n16715), .Z(n16713) );
  XOR U16320 ( .A(n16712), .B(n16716), .Z(n16714) );
  XNOR U16321 ( .A(n16717), .B(n16718), .Z(n16711) );
  NOR U16322 ( .A(n16719), .B(n16720), .Z(n16718) );
  XNOR U16323 ( .A(n16717), .B(n16721), .Z(n16719) );
  XOR U16324 ( .A(n16722), .B(n16723), .Z(n16679) );
  NOR U16325 ( .A(n16724), .B(n16725), .Z(n16723) );
  XNOR U16326 ( .A(n16722), .B(n16726), .Z(n16724) );
  XNOR U16327 ( .A(n16621), .B(n16683), .Z(n16685) );
  XNOR U16328 ( .A(n16727), .B(n16728), .Z(n16621) );
  AND U16329 ( .A(n38), .B(n16628), .Z(n16728) );
  XOR U16330 ( .A(n16727), .B(n16626), .Z(n16628) );
  AND U16331 ( .A(n16631), .B(n16634), .Z(n16683) );
  XOR U16332 ( .A(n16729), .B(n16710), .Z(n16634) );
  XNOR U16333 ( .A(p_input[0]), .B(p_input[2048]), .Z(n16710) );
  XOR U16334 ( .A(n16698), .B(n16697), .Z(n16729) );
  XNOR U16335 ( .A(n16730), .B(n16704), .Z(n16697) );
  XNOR U16336 ( .A(n16693), .B(n16692), .Z(n16704) );
  XNOR U16337 ( .A(n16731), .B(n16689), .Z(n16692) );
  XNOR U16338 ( .A(p_input[10]), .B(p_input[2058]), .Z(n16689) );
  XOR U16339 ( .A(p_input[11]), .B(n16732), .Z(n16731) );
  XOR U16340 ( .A(p_input[12]), .B(p_input[2060]), .Z(n16693) );
  XOR U16341 ( .A(n16703), .B(n16733), .Z(n16730) );
  IV U16342 ( .A(n16694), .Z(n16733) );
  XOR U16343 ( .A(p_input[1]), .B(p_input[2049]), .Z(n16694) );
  XNOR U16344 ( .A(n16734), .B(n16709), .Z(n16703) );
  XNOR U16345 ( .A(p_input[15]), .B(n16735), .Z(n16709) );
  XOR U16346 ( .A(n16700), .B(n16708), .Z(n16734) );
  XOR U16347 ( .A(n16736), .B(n16705), .Z(n16708) );
  XOR U16348 ( .A(p_input[13]), .B(p_input[2061]), .Z(n16705) );
  XOR U16349 ( .A(p_input[14]), .B(n16737), .Z(n16736) );
  XNOR U16350 ( .A(n16738), .B(p_input[9]), .Z(n16700) );
  XNOR U16351 ( .A(n16716), .B(n16715), .Z(n16698) );
  XNOR U16352 ( .A(n16739), .B(n16721), .Z(n16715) );
  XOR U16353 ( .A(p_input[2056]), .B(p_input[8]), .Z(n16721) );
  XOR U16354 ( .A(n16712), .B(n16720), .Z(n16739) );
  XOR U16355 ( .A(n16740), .B(n16717), .Z(n16720) );
  XOR U16356 ( .A(p_input[2054]), .B(p_input[6]), .Z(n16717) );
  XNOR U16357 ( .A(p_input[2055]), .B(p_input[7]), .Z(n16740) );
  XNOR U16358 ( .A(n16741), .B(p_input[2]), .Z(n16712) );
  XNOR U16359 ( .A(n16726), .B(n16725), .Z(n16716) );
  XOR U16360 ( .A(n16742), .B(n16722), .Z(n16725) );
  XOR U16361 ( .A(p_input[2051]), .B(p_input[3]), .Z(n16722) );
  XNOR U16362 ( .A(p_input[2052]), .B(p_input[4]), .Z(n16742) );
  XOR U16363 ( .A(p_input[2053]), .B(p_input[5]), .Z(n16726) );
  XNOR U16364 ( .A(n16743), .B(n16744), .Z(n16631) );
  AND U16365 ( .A(n38), .B(n16745), .Z(n16744) );
  XNOR U16366 ( .A(n16746), .B(n16747), .Z(n38) );
  AND U16367 ( .A(n16748), .B(n16749), .Z(n16747) );
  XOR U16368 ( .A(n16746), .B(n16641), .Z(n16749) );
  XNOR U16369 ( .A(n16746), .B(n16587), .Z(n16748) );
  XOR U16370 ( .A(n16750), .B(n16751), .Z(n16746) );
  AND U16371 ( .A(n16752), .B(n16753), .Z(n16751) );
  XNOR U16372 ( .A(n16654), .B(n16750), .Z(n16753) );
  XOR U16373 ( .A(n16750), .B(n16656), .Z(n16752) );
  XOR U16374 ( .A(n16754), .B(n16755), .Z(n16750) );
  AND U16375 ( .A(n16756), .B(n16757), .Z(n16755) );
  XOR U16376 ( .A(n16754), .B(n16682), .Z(n16756) );
  IV U16377 ( .A(n16613), .Z(n16682) );
  XOR U16378 ( .A(n16758), .B(n16759), .Z(n16629) );
  AND U16379 ( .A(n42), .B(n16745), .Z(n16759) );
  XNOR U16380 ( .A(n16743), .B(n16758), .Z(n16745) );
  XNOR U16381 ( .A(n16760), .B(n16761), .Z(n42) );
  AND U16382 ( .A(n16762), .B(n16763), .Z(n16761) );
  XNOR U16383 ( .A(n16764), .B(n16760), .Z(n16763) );
  IV U16384 ( .A(n16641), .Z(n16764) );
  XNOR U16385 ( .A(n16765), .B(n16766), .Z(n16641) );
  AND U16386 ( .A(n46), .B(n16767), .Z(n16766) );
  XNOR U16387 ( .A(n16765), .B(n16768), .Z(n16767) );
  XNOR U16388 ( .A(n16587), .B(n16760), .Z(n16762) );
  XOR U16389 ( .A(n16769), .B(n16770), .Z(n16587) );
  AND U16390 ( .A(n54), .B(n16771), .Z(n16770) );
  XOR U16391 ( .A(n16772), .B(n16773), .Z(n16760) );
  AND U16392 ( .A(n16774), .B(n16775), .Z(n16773) );
  XNOR U16393 ( .A(n16772), .B(n16654), .Z(n16775) );
  XNOR U16394 ( .A(n16776), .B(n16777), .Z(n16654) );
  AND U16395 ( .A(n46), .B(n16778), .Z(n16777) );
  XOR U16396 ( .A(n16779), .B(n16776), .Z(n16778) );
  XNOR U16397 ( .A(n16600), .B(n16772), .Z(n16774) );
  IV U16398 ( .A(n16656), .Z(n16600) );
  XOR U16399 ( .A(n16780), .B(n16781), .Z(n16656) );
  AND U16400 ( .A(n54), .B(n16782), .Z(n16781) );
  XOR U16401 ( .A(n16754), .B(n16783), .Z(n16772) );
  AND U16402 ( .A(n16784), .B(n16757), .Z(n16783) );
  XNOR U16403 ( .A(n16680), .B(n16754), .Z(n16757) );
  XNOR U16404 ( .A(n16785), .B(n16786), .Z(n16680) );
  AND U16405 ( .A(n46), .B(n16787), .Z(n16786) );
  XNOR U16406 ( .A(n16788), .B(n16785), .Z(n16787) );
  XNOR U16407 ( .A(n16613), .B(n16754), .Z(n16784) );
  XNOR U16408 ( .A(n16789), .B(n16790), .Z(n16613) );
  AND U16409 ( .A(n54), .B(n16791), .Z(n16790) );
  XOR U16410 ( .A(n16792), .B(n16793), .Z(n16754) );
  AND U16411 ( .A(n16794), .B(n16795), .Z(n16793) );
  XNOR U16412 ( .A(n16792), .B(n16727), .Z(n16795) );
  XNOR U16413 ( .A(n16796), .B(n16797), .Z(n16727) );
  AND U16414 ( .A(n46), .B(n16798), .Z(n16797) );
  XOR U16415 ( .A(n16799), .B(n16796), .Z(n16798) );
  XNOR U16416 ( .A(n16800), .B(n16792), .Z(n16794) );
  IV U16417 ( .A(n16626), .Z(n16800) );
  XOR U16418 ( .A(n16801), .B(n16802), .Z(n16626) );
  AND U16419 ( .A(n54), .B(n16803), .Z(n16802) );
  AND U16420 ( .A(n16758), .B(n16743), .Z(n16792) );
  XNOR U16421 ( .A(n16804), .B(n16805), .Z(n16743) );
  AND U16422 ( .A(n46), .B(n16806), .Z(n16805) );
  XNOR U16423 ( .A(n16807), .B(n16804), .Z(n16806) );
  XNOR U16424 ( .A(n16808), .B(n16809), .Z(n46) );
  AND U16425 ( .A(n16810), .B(n16811), .Z(n16809) );
  XOR U16426 ( .A(n16768), .B(n16808), .Z(n16811) );
  AND U16427 ( .A(n16812), .B(n16813), .Z(n16768) );
  XOR U16428 ( .A(n16808), .B(n16765), .Z(n16810) );
  XNOR U16429 ( .A(n16814), .B(n16815), .Z(n16765) );
  AND U16430 ( .A(n50), .B(n16771), .Z(n16815) );
  XOR U16431 ( .A(n16769), .B(n16814), .Z(n16771) );
  XOR U16432 ( .A(n16816), .B(n16817), .Z(n16808) );
  AND U16433 ( .A(n16818), .B(n16819), .Z(n16817) );
  XNOR U16434 ( .A(n16816), .B(n16812), .Z(n16819) );
  IV U16435 ( .A(n16779), .Z(n16812) );
  XOR U16436 ( .A(n16820), .B(n16821), .Z(n16779) );
  XOR U16437 ( .A(n16822), .B(n16813), .Z(n16821) );
  AND U16438 ( .A(n16788), .B(n16823), .Z(n16813) );
  AND U16439 ( .A(n16824), .B(n16825), .Z(n16822) );
  XOR U16440 ( .A(n16826), .B(n16820), .Z(n16824) );
  XNOR U16441 ( .A(n16776), .B(n16816), .Z(n16818) );
  XNOR U16442 ( .A(n16827), .B(n16828), .Z(n16776) );
  AND U16443 ( .A(n50), .B(n16782), .Z(n16828) );
  XOR U16444 ( .A(n16827), .B(n16780), .Z(n16782) );
  XOR U16445 ( .A(n16829), .B(n16830), .Z(n16816) );
  AND U16446 ( .A(n16831), .B(n16832), .Z(n16830) );
  XNOR U16447 ( .A(n16829), .B(n16788), .Z(n16832) );
  XOR U16448 ( .A(n16833), .B(n16825), .Z(n16788) );
  XNOR U16449 ( .A(n16834), .B(n16820), .Z(n16825) );
  XOR U16450 ( .A(n16835), .B(n16836), .Z(n16820) );
  AND U16451 ( .A(n16837), .B(n16838), .Z(n16836) );
  XOR U16452 ( .A(n16839), .B(n16835), .Z(n16837) );
  XNOR U16453 ( .A(n16840), .B(n16841), .Z(n16834) );
  AND U16454 ( .A(n16842), .B(n16843), .Z(n16841) );
  XOR U16455 ( .A(n16840), .B(n16844), .Z(n16842) );
  XNOR U16456 ( .A(n16826), .B(n16823), .Z(n16833) );
  AND U16457 ( .A(n16845), .B(n16846), .Z(n16823) );
  XOR U16458 ( .A(n16847), .B(n16848), .Z(n16826) );
  AND U16459 ( .A(n16849), .B(n16850), .Z(n16848) );
  XOR U16460 ( .A(n16847), .B(n16851), .Z(n16849) );
  XNOR U16461 ( .A(n16785), .B(n16829), .Z(n16831) );
  XNOR U16462 ( .A(n16852), .B(n16853), .Z(n16785) );
  AND U16463 ( .A(n50), .B(n16791), .Z(n16853) );
  XOR U16464 ( .A(n16852), .B(n16789), .Z(n16791) );
  XOR U16465 ( .A(n16854), .B(n16855), .Z(n16829) );
  AND U16466 ( .A(n16856), .B(n16857), .Z(n16855) );
  XNOR U16467 ( .A(n16854), .B(n16845), .Z(n16857) );
  IV U16468 ( .A(n16799), .Z(n16845) );
  XNOR U16469 ( .A(n16858), .B(n16838), .Z(n16799) );
  XNOR U16470 ( .A(n16859), .B(n16844), .Z(n16838) );
  XOR U16471 ( .A(n16860), .B(n16861), .Z(n16844) );
  NOR U16472 ( .A(n16862), .B(n16863), .Z(n16861) );
  XNOR U16473 ( .A(n16860), .B(n16864), .Z(n16862) );
  XNOR U16474 ( .A(n16843), .B(n16835), .Z(n16859) );
  XOR U16475 ( .A(n16865), .B(n16866), .Z(n16835) );
  AND U16476 ( .A(n16867), .B(n16868), .Z(n16866) );
  XNOR U16477 ( .A(n16865), .B(n16869), .Z(n16867) );
  XNOR U16478 ( .A(n16870), .B(n16840), .Z(n16843) );
  XOR U16479 ( .A(n16871), .B(n16872), .Z(n16840) );
  AND U16480 ( .A(n16873), .B(n16874), .Z(n16872) );
  XOR U16481 ( .A(n16871), .B(n16875), .Z(n16873) );
  XNOR U16482 ( .A(n16876), .B(n16877), .Z(n16870) );
  NOR U16483 ( .A(n16878), .B(n16879), .Z(n16877) );
  XOR U16484 ( .A(n16876), .B(n16880), .Z(n16878) );
  XNOR U16485 ( .A(n16839), .B(n16846), .Z(n16858) );
  NOR U16486 ( .A(n16807), .B(n16881), .Z(n16846) );
  XOR U16487 ( .A(n16851), .B(n16850), .Z(n16839) );
  XNOR U16488 ( .A(n16882), .B(n16847), .Z(n16850) );
  XOR U16489 ( .A(n16883), .B(n16884), .Z(n16847) );
  AND U16490 ( .A(n16885), .B(n16886), .Z(n16884) );
  XNOR U16491 ( .A(n16887), .B(n16888), .Z(n16885) );
  IV U16492 ( .A(n16883), .Z(n16887) );
  XNOR U16493 ( .A(n16889), .B(n16890), .Z(n16882) );
  NOR U16494 ( .A(n16891), .B(n16892), .Z(n16890) );
  XNOR U16495 ( .A(n16889), .B(n16893), .Z(n16891) );
  XOR U16496 ( .A(n16894), .B(n16895), .Z(n16851) );
  NOR U16497 ( .A(n16896), .B(n16897), .Z(n16895) );
  XNOR U16498 ( .A(n16894), .B(n16898), .Z(n16896) );
  XNOR U16499 ( .A(n16796), .B(n16854), .Z(n16856) );
  XNOR U16500 ( .A(n16899), .B(n16900), .Z(n16796) );
  AND U16501 ( .A(n50), .B(n16803), .Z(n16900) );
  XOR U16502 ( .A(n16899), .B(n16801), .Z(n16803) );
  AND U16503 ( .A(n16804), .B(n16807), .Z(n16854) );
  XOR U16504 ( .A(n16901), .B(n16881), .Z(n16807) );
  XNOR U16505 ( .A(p_input[16]), .B(p_input[2048]), .Z(n16881) );
  XOR U16506 ( .A(n16869), .B(n16868), .Z(n16901) );
  XNOR U16507 ( .A(n16902), .B(n16875), .Z(n16868) );
  XNOR U16508 ( .A(n16864), .B(n16863), .Z(n16875) );
  XOR U16509 ( .A(n16903), .B(n16860), .Z(n16863) );
  XNOR U16510 ( .A(n16904), .B(p_input[26]), .Z(n16860) );
  XNOR U16511 ( .A(p_input[2059]), .B(p_input[27]), .Z(n16903) );
  XOR U16512 ( .A(p_input[2060]), .B(p_input[28]), .Z(n16864) );
  XOR U16513 ( .A(n16874), .B(n16905), .Z(n16902) );
  IV U16514 ( .A(n16865), .Z(n16905) );
  XOR U16515 ( .A(p_input[17]), .B(p_input[2049]), .Z(n16865) );
  XOR U16516 ( .A(n16906), .B(n16880), .Z(n16874) );
  XNOR U16517 ( .A(p_input[2063]), .B(p_input[31]), .Z(n16880) );
  XOR U16518 ( .A(n16871), .B(n16879), .Z(n16906) );
  XOR U16519 ( .A(n16907), .B(n16876), .Z(n16879) );
  XOR U16520 ( .A(p_input[2061]), .B(p_input[29]), .Z(n16876) );
  XNOR U16521 ( .A(p_input[2062]), .B(p_input[30]), .Z(n16907) );
  XNOR U16522 ( .A(n16738), .B(p_input[25]), .Z(n16871) );
  XNOR U16523 ( .A(n16888), .B(n16886), .Z(n16869) );
  XNOR U16524 ( .A(n16908), .B(n16893), .Z(n16886) );
  XOR U16525 ( .A(p_input[2056]), .B(p_input[24]), .Z(n16893) );
  XOR U16526 ( .A(n16883), .B(n16892), .Z(n16908) );
  XOR U16527 ( .A(n16909), .B(n16889), .Z(n16892) );
  XOR U16528 ( .A(p_input[2054]), .B(p_input[22]), .Z(n16889) );
  XNOR U16529 ( .A(p_input[2055]), .B(p_input[23]), .Z(n16909) );
  XOR U16530 ( .A(p_input[18]), .B(p_input[2050]), .Z(n16883) );
  XNOR U16531 ( .A(n16898), .B(n16897), .Z(n16888) );
  XOR U16532 ( .A(n16910), .B(n16894), .Z(n16897) );
  XOR U16533 ( .A(p_input[19]), .B(p_input[2051]), .Z(n16894) );
  XNOR U16534 ( .A(p_input[2052]), .B(p_input[20]), .Z(n16910) );
  XOR U16535 ( .A(p_input[2053]), .B(p_input[21]), .Z(n16898) );
  XNOR U16536 ( .A(n16911), .B(n16912), .Z(n16804) );
  AND U16537 ( .A(n50), .B(n16913), .Z(n16912) );
  XNOR U16538 ( .A(n16914), .B(n16915), .Z(n50) );
  AND U16539 ( .A(n16916), .B(n16917), .Z(n16915) );
  XOR U16540 ( .A(n16914), .B(n16814), .Z(n16917) );
  XNOR U16541 ( .A(n16914), .B(n16769), .Z(n16916) );
  XOR U16542 ( .A(n16918), .B(n16919), .Z(n16914) );
  AND U16543 ( .A(n16920), .B(n16921), .Z(n16919) );
  XOR U16544 ( .A(n16918), .B(n16780), .Z(n16920) );
  XOR U16545 ( .A(n16922), .B(n16923), .Z(n16758) );
  AND U16546 ( .A(n54), .B(n16913), .Z(n16923) );
  XNOR U16547 ( .A(n16911), .B(n16922), .Z(n16913) );
  XNOR U16548 ( .A(n16924), .B(n16925), .Z(n54) );
  AND U16549 ( .A(n16926), .B(n16927), .Z(n16925) );
  XNOR U16550 ( .A(n16928), .B(n16924), .Z(n16927) );
  IV U16551 ( .A(n16814), .Z(n16928) );
  XNOR U16552 ( .A(n16929), .B(n16930), .Z(n16814) );
  AND U16553 ( .A(n57), .B(n16931), .Z(n16930) );
  XNOR U16554 ( .A(n16929), .B(n16932), .Z(n16931) );
  XNOR U16555 ( .A(n16769), .B(n16924), .Z(n16926) );
  XOR U16556 ( .A(n16933), .B(n16934), .Z(n16769) );
  AND U16557 ( .A(n65), .B(n16935), .Z(n16934) );
  XOR U16558 ( .A(n16918), .B(n16936), .Z(n16924) );
  AND U16559 ( .A(n16937), .B(n16921), .Z(n16936) );
  XNOR U16560 ( .A(n16827), .B(n16918), .Z(n16921) );
  XNOR U16561 ( .A(n16938), .B(n16939), .Z(n16827) );
  AND U16562 ( .A(n57), .B(n16940), .Z(n16939) );
  XOR U16563 ( .A(n16941), .B(n16938), .Z(n16940) );
  XNOR U16564 ( .A(n16942), .B(n16918), .Z(n16937) );
  IV U16565 ( .A(n16780), .Z(n16942) );
  XOR U16566 ( .A(n16943), .B(n16944), .Z(n16780) );
  AND U16567 ( .A(n65), .B(n16945), .Z(n16944) );
  XOR U16568 ( .A(n16946), .B(n16947), .Z(n16918) );
  AND U16569 ( .A(n16948), .B(n16949), .Z(n16947) );
  XNOR U16570 ( .A(n16852), .B(n16946), .Z(n16949) );
  XNOR U16571 ( .A(n16950), .B(n16951), .Z(n16852) );
  AND U16572 ( .A(n57), .B(n16952), .Z(n16951) );
  XNOR U16573 ( .A(n16953), .B(n16950), .Z(n16952) );
  XOR U16574 ( .A(n16946), .B(n16789), .Z(n16948) );
  XOR U16575 ( .A(n16954), .B(n16955), .Z(n16789) );
  AND U16576 ( .A(n65), .B(n16956), .Z(n16955) );
  XOR U16577 ( .A(n16957), .B(n16958), .Z(n16946) );
  AND U16578 ( .A(n16959), .B(n16960), .Z(n16958) );
  XNOR U16579 ( .A(n16957), .B(n16899), .Z(n16960) );
  XNOR U16580 ( .A(n16961), .B(n16962), .Z(n16899) );
  AND U16581 ( .A(n57), .B(n16963), .Z(n16962) );
  XOR U16582 ( .A(n16964), .B(n16961), .Z(n16963) );
  XNOR U16583 ( .A(n16965), .B(n16957), .Z(n16959) );
  IV U16584 ( .A(n16801), .Z(n16965) );
  XOR U16585 ( .A(n16966), .B(n16967), .Z(n16801) );
  AND U16586 ( .A(n65), .B(n16968), .Z(n16967) );
  AND U16587 ( .A(n16922), .B(n16911), .Z(n16957) );
  XNOR U16588 ( .A(n16969), .B(n16970), .Z(n16911) );
  AND U16589 ( .A(n57), .B(n16971), .Z(n16970) );
  XNOR U16590 ( .A(n16972), .B(n16969), .Z(n16971) );
  XNOR U16591 ( .A(n16973), .B(n16974), .Z(n57) );
  AND U16592 ( .A(n16975), .B(n16976), .Z(n16974) );
  XOR U16593 ( .A(n16932), .B(n16973), .Z(n16976) );
  AND U16594 ( .A(n16977), .B(n16978), .Z(n16932) );
  XOR U16595 ( .A(n16973), .B(n16929), .Z(n16975) );
  XNOR U16596 ( .A(n16979), .B(n16980), .Z(n16929) );
  AND U16597 ( .A(n61), .B(n16935), .Z(n16980) );
  XOR U16598 ( .A(n16933), .B(n16979), .Z(n16935) );
  XOR U16599 ( .A(n16981), .B(n16982), .Z(n16973) );
  AND U16600 ( .A(n16983), .B(n16984), .Z(n16982) );
  XNOR U16601 ( .A(n16981), .B(n16977), .Z(n16984) );
  IV U16602 ( .A(n16941), .Z(n16977) );
  XOR U16603 ( .A(n16985), .B(n16986), .Z(n16941) );
  XOR U16604 ( .A(n16987), .B(n16978), .Z(n16986) );
  AND U16605 ( .A(n16953), .B(n16988), .Z(n16978) );
  AND U16606 ( .A(n16989), .B(n16990), .Z(n16987) );
  XOR U16607 ( .A(n16991), .B(n16985), .Z(n16989) );
  XNOR U16608 ( .A(n16938), .B(n16981), .Z(n16983) );
  XNOR U16609 ( .A(n16992), .B(n16993), .Z(n16938) );
  AND U16610 ( .A(n61), .B(n16945), .Z(n16993) );
  XOR U16611 ( .A(n16992), .B(n16943), .Z(n16945) );
  XOR U16612 ( .A(n16994), .B(n16995), .Z(n16981) );
  AND U16613 ( .A(n16996), .B(n16997), .Z(n16995) );
  XNOR U16614 ( .A(n16994), .B(n16953), .Z(n16997) );
  XOR U16615 ( .A(n16998), .B(n16990), .Z(n16953) );
  XNOR U16616 ( .A(n16999), .B(n16985), .Z(n16990) );
  XOR U16617 ( .A(n17000), .B(n17001), .Z(n16985) );
  AND U16618 ( .A(n17002), .B(n17003), .Z(n17001) );
  XOR U16619 ( .A(n17004), .B(n17000), .Z(n17002) );
  XNOR U16620 ( .A(n17005), .B(n17006), .Z(n16999) );
  AND U16621 ( .A(n17007), .B(n17008), .Z(n17006) );
  XOR U16622 ( .A(n17005), .B(n17009), .Z(n17007) );
  XNOR U16623 ( .A(n16991), .B(n16988), .Z(n16998) );
  AND U16624 ( .A(n17010), .B(n17011), .Z(n16988) );
  XOR U16625 ( .A(n17012), .B(n17013), .Z(n16991) );
  AND U16626 ( .A(n17014), .B(n17015), .Z(n17013) );
  XOR U16627 ( .A(n17012), .B(n17016), .Z(n17014) );
  XNOR U16628 ( .A(n16950), .B(n16994), .Z(n16996) );
  XNOR U16629 ( .A(n17017), .B(n17018), .Z(n16950) );
  AND U16630 ( .A(n61), .B(n16956), .Z(n17018) );
  XOR U16631 ( .A(n17017), .B(n16954), .Z(n16956) );
  XOR U16632 ( .A(n17019), .B(n17020), .Z(n16994) );
  AND U16633 ( .A(n17021), .B(n17022), .Z(n17020) );
  XNOR U16634 ( .A(n17019), .B(n17010), .Z(n17022) );
  IV U16635 ( .A(n16964), .Z(n17010) );
  XNOR U16636 ( .A(n17023), .B(n17003), .Z(n16964) );
  XNOR U16637 ( .A(n17024), .B(n17009), .Z(n17003) );
  XOR U16638 ( .A(n17025), .B(n17026), .Z(n17009) );
  NOR U16639 ( .A(n17027), .B(n17028), .Z(n17026) );
  XNOR U16640 ( .A(n17025), .B(n17029), .Z(n17027) );
  XNOR U16641 ( .A(n17008), .B(n17000), .Z(n17024) );
  XOR U16642 ( .A(n17030), .B(n17031), .Z(n17000) );
  AND U16643 ( .A(n17032), .B(n17033), .Z(n17031) );
  XNOR U16644 ( .A(n17030), .B(n17034), .Z(n17032) );
  XNOR U16645 ( .A(n17035), .B(n17005), .Z(n17008) );
  XOR U16646 ( .A(n17036), .B(n17037), .Z(n17005) );
  AND U16647 ( .A(n17038), .B(n17039), .Z(n17037) );
  XOR U16648 ( .A(n17036), .B(n17040), .Z(n17038) );
  XNOR U16649 ( .A(n17041), .B(n17042), .Z(n17035) );
  NOR U16650 ( .A(n17043), .B(n17044), .Z(n17042) );
  XOR U16651 ( .A(n17041), .B(n17045), .Z(n17043) );
  XNOR U16652 ( .A(n17004), .B(n17011), .Z(n17023) );
  NOR U16653 ( .A(n16972), .B(n17046), .Z(n17011) );
  XOR U16654 ( .A(n17016), .B(n17015), .Z(n17004) );
  XNOR U16655 ( .A(n17047), .B(n17012), .Z(n17015) );
  XOR U16656 ( .A(n17048), .B(n17049), .Z(n17012) );
  AND U16657 ( .A(n17050), .B(n17051), .Z(n17049) );
  XOR U16658 ( .A(n17048), .B(n17052), .Z(n17050) );
  XNOR U16659 ( .A(n17053), .B(n17054), .Z(n17047) );
  NOR U16660 ( .A(n17055), .B(n17056), .Z(n17054) );
  XNOR U16661 ( .A(n17053), .B(n17057), .Z(n17055) );
  XOR U16662 ( .A(n17058), .B(n17059), .Z(n17016) );
  NOR U16663 ( .A(n17060), .B(n17061), .Z(n17059) );
  XNOR U16664 ( .A(n17058), .B(n17062), .Z(n17060) );
  XNOR U16665 ( .A(n16961), .B(n17019), .Z(n17021) );
  XNOR U16666 ( .A(n17063), .B(n17064), .Z(n16961) );
  AND U16667 ( .A(n61), .B(n16968), .Z(n17064) );
  XOR U16668 ( .A(n17063), .B(n16966), .Z(n16968) );
  AND U16669 ( .A(n16969), .B(n16972), .Z(n17019) );
  XOR U16670 ( .A(n17065), .B(n17046), .Z(n16972) );
  XNOR U16671 ( .A(p_input[2048]), .B(p_input[32]), .Z(n17046) );
  XOR U16672 ( .A(n17034), .B(n17033), .Z(n17065) );
  XNOR U16673 ( .A(n17066), .B(n17040), .Z(n17033) );
  XNOR U16674 ( .A(n17029), .B(n17028), .Z(n17040) );
  XOR U16675 ( .A(n17067), .B(n17025), .Z(n17028) );
  XNOR U16676 ( .A(n16904), .B(p_input[42]), .Z(n17025) );
  XNOR U16677 ( .A(p_input[2059]), .B(p_input[43]), .Z(n17067) );
  XOR U16678 ( .A(p_input[2060]), .B(p_input[44]), .Z(n17029) );
  XNOR U16679 ( .A(n17039), .B(n17030), .Z(n17066) );
  XNOR U16680 ( .A(n17068), .B(p_input[33]), .Z(n17030) );
  XOR U16681 ( .A(n17069), .B(n17045), .Z(n17039) );
  XNOR U16682 ( .A(p_input[2063]), .B(p_input[47]), .Z(n17045) );
  XOR U16683 ( .A(n17036), .B(n17044), .Z(n17069) );
  XOR U16684 ( .A(n17070), .B(n17041), .Z(n17044) );
  XOR U16685 ( .A(p_input[2061]), .B(p_input[45]), .Z(n17041) );
  XNOR U16686 ( .A(p_input[2062]), .B(p_input[46]), .Z(n17070) );
  XNOR U16687 ( .A(n16738), .B(p_input[41]), .Z(n17036) );
  XNOR U16688 ( .A(n17052), .B(n17051), .Z(n17034) );
  XNOR U16689 ( .A(n17071), .B(n17057), .Z(n17051) );
  XOR U16690 ( .A(p_input[2056]), .B(p_input[40]), .Z(n17057) );
  XOR U16691 ( .A(n17048), .B(n17056), .Z(n17071) );
  XOR U16692 ( .A(n17072), .B(n17053), .Z(n17056) );
  XOR U16693 ( .A(p_input[2054]), .B(p_input[38]), .Z(n17053) );
  XNOR U16694 ( .A(p_input[2055]), .B(p_input[39]), .Z(n17072) );
  XNOR U16695 ( .A(n16741), .B(p_input[34]), .Z(n17048) );
  XNOR U16696 ( .A(n17062), .B(n17061), .Z(n17052) );
  XOR U16697 ( .A(n17073), .B(n17058), .Z(n17061) );
  XOR U16698 ( .A(p_input[2051]), .B(p_input[35]), .Z(n17058) );
  XNOR U16699 ( .A(p_input[2052]), .B(p_input[36]), .Z(n17073) );
  XOR U16700 ( .A(p_input[2053]), .B(p_input[37]), .Z(n17062) );
  XNOR U16701 ( .A(n17074), .B(n17075), .Z(n16969) );
  AND U16702 ( .A(n61), .B(n17076), .Z(n17075) );
  XNOR U16703 ( .A(n17077), .B(n17078), .Z(n61) );
  AND U16704 ( .A(n17079), .B(n17080), .Z(n17078) );
  XOR U16705 ( .A(n17077), .B(n16979), .Z(n17080) );
  XNOR U16706 ( .A(n17077), .B(n16933), .Z(n17079) );
  XOR U16707 ( .A(n17081), .B(n17082), .Z(n17077) );
  AND U16708 ( .A(n17083), .B(n17084), .Z(n17082) );
  XOR U16709 ( .A(n17081), .B(n16943), .Z(n17083) );
  XOR U16710 ( .A(n17085), .B(n17086), .Z(n16922) );
  AND U16711 ( .A(n65), .B(n17076), .Z(n17086) );
  XNOR U16712 ( .A(n17074), .B(n17085), .Z(n17076) );
  XNOR U16713 ( .A(n17087), .B(n17088), .Z(n65) );
  AND U16714 ( .A(n17089), .B(n17090), .Z(n17088) );
  XNOR U16715 ( .A(n17091), .B(n17087), .Z(n17090) );
  IV U16716 ( .A(n16979), .Z(n17091) );
  XNOR U16717 ( .A(n17092), .B(n17093), .Z(n16979) );
  AND U16718 ( .A(n68), .B(n17094), .Z(n17093) );
  XNOR U16719 ( .A(n17092), .B(n17095), .Z(n17094) );
  XNOR U16720 ( .A(n16933), .B(n17087), .Z(n17089) );
  XOR U16721 ( .A(n17096), .B(n17097), .Z(n16933) );
  AND U16722 ( .A(n76), .B(n17098), .Z(n17097) );
  XOR U16723 ( .A(n17081), .B(n17099), .Z(n17087) );
  AND U16724 ( .A(n17100), .B(n17084), .Z(n17099) );
  XNOR U16725 ( .A(n16992), .B(n17081), .Z(n17084) );
  XNOR U16726 ( .A(n17101), .B(n17102), .Z(n16992) );
  AND U16727 ( .A(n68), .B(n17103), .Z(n17102) );
  XOR U16728 ( .A(n17104), .B(n17101), .Z(n17103) );
  XNOR U16729 ( .A(n17105), .B(n17081), .Z(n17100) );
  IV U16730 ( .A(n16943), .Z(n17105) );
  XOR U16731 ( .A(n17106), .B(n17107), .Z(n16943) );
  AND U16732 ( .A(n76), .B(n17108), .Z(n17107) );
  XOR U16733 ( .A(n17109), .B(n17110), .Z(n17081) );
  AND U16734 ( .A(n17111), .B(n17112), .Z(n17110) );
  XNOR U16735 ( .A(n17017), .B(n17109), .Z(n17112) );
  XNOR U16736 ( .A(n17113), .B(n17114), .Z(n17017) );
  AND U16737 ( .A(n68), .B(n17115), .Z(n17114) );
  XNOR U16738 ( .A(n17116), .B(n17113), .Z(n17115) );
  XOR U16739 ( .A(n17109), .B(n16954), .Z(n17111) );
  XOR U16740 ( .A(n17117), .B(n17118), .Z(n16954) );
  AND U16741 ( .A(n76), .B(n17119), .Z(n17118) );
  XOR U16742 ( .A(n17120), .B(n17121), .Z(n17109) );
  AND U16743 ( .A(n17122), .B(n17123), .Z(n17121) );
  XNOR U16744 ( .A(n17120), .B(n17063), .Z(n17123) );
  XNOR U16745 ( .A(n17124), .B(n17125), .Z(n17063) );
  AND U16746 ( .A(n68), .B(n17126), .Z(n17125) );
  XOR U16747 ( .A(n17127), .B(n17124), .Z(n17126) );
  XNOR U16748 ( .A(n17128), .B(n17120), .Z(n17122) );
  IV U16749 ( .A(n16966), .Z(n17128) );
  XOR U16750 ( .A(n17129), .B(n17130), .Z(n16966) );
  AND U16751 ( .A(n76), .B(n17131), .Z(n17130) );
  AND U16752 ( .A(n17085), .B(n17074), .Z(n17120) );
  XNOR U16753 ( .A(n17132), .B(n17133), .Z(n17074) );
  AND U16754 ( .A(n68), .B(n17134), .Z(n17133) );
  XNOR U16755 ( .A(n17135), .B(n17132), .Z(n17134) );
  XNOR U16756 ( .A(n17136), .B(n17137), .Z(n68) );
  AND U16757 ( .A(n17138), .B(n17139), .Z(n17137) );
  XOR U16758 ( .A(n17095), .B(n17136), .Z(n17139) );
  AND U16759 ( .A(n17140), .B(n17141), .Z(n17095) );
  XOR U16760 ( .A(n17136), .B(n17092), .Z(n17138) );
  XNOR U16761 ( .A(n17142), .B(n17143), .Z(n17092) );
  AND U16762 ( .A(n72), .B(n17098), .Z(n17143) );
  XOR U16763 ( .A(n17096), .B(n17142), .Z(n17098) );
  XOR U16764 ( .A(n17144), .B(n17145), .Z(n17136) );
  AND U16765 ( .A(n17146), .B(n17147), .Z(n17145) );
  XNOR U16766 ( .A(n17144), .B(n17140), .Z(n17147) );
  IV U16767 ( .A(n17104), .Z(n17140) );
  XOR U16768 ( .A(n17148), .B(n17149), .Z(n17104) );
  XOR U16769 ( .A(n17150), .B(n17141), .Z(n17149) );
  AND U16770 ( .A(n17116), .B(n17151), .Z(n17141) );
  AND U16771 ( .A(n17152), .B(n17153), .Z(n17150) );
  XOR U16772 ( .A(n17154), .B(n17148), .Z(n17152) );
  XNOR U16773 ( .A(n17101), .B(n17144), .Z(n17146) );
  XNOR U16774 ( .A(n17155), .B(n17156), .Z(n17101) );
  AND U16775 ( .A(n72), .B(n17108), .Z(n17156) );
  XOR U16776 ( .A(n17155), .B(n17106), .Z(n17108) );
  XOR U16777 ( .A(n17157), .B(n17158), .Z(n17144) );
  AND U16778 ( .A(n17159), .B(n17160), .Z(n17158) );
  XNOR U16779 ( .A(n17157), .B(n17116), .Z(n17160) );
  XOR U16780 ( .A(n17161), .B(n17153), .Z(n17116) );
  XNOR U16781 ( .A(n17162), .B(n17148), .Z(n17153) );
  XOR U16782 ( .A(n17163), .B(n17164), .Z(n17148) );
  AND U16783 ( .A(n17165), .B(n17166), .Z(n17164) );
  XOR U16784 ( .A(n17167), .B(n17163), .Z(n17165) );
  XNOR U16785 ( .A(n17168), .B(n17169), .Z(n17162) );
  AND U16786 ( .A(n17170), .B(n17171), .Z(n17169) );
  XOR U16787 ( .A(n17168), .B(n17172), .Z(n17170) );
  XNOR U16788 ( .A(n17154), .B(n17151), .Z(n17161) );
  AND U16789 ( .A(n17173), .B(n17174), .Z(n17151) );
  XOR U16790 ( .A(n17175), .B(n17176), .Z(n17154) );
  AND U16791 ( .A(n17177), .B(n17178), .Z(n17176) );
  XOR U16792 ( .A(n17175), .B(n17179), .Z(n17177) );
  XNOR U16793 ( .A(n17113), .B(n17157), .Z(n17159) );
  XNOR U16794 ( .A(n17180), .B(n17181), .Z(n17113) );
  AND U16795 ( .A(n72), .B(n17119), .Z(n17181) );
  XOR U16796 ( .A(n17180), .B(n17117), .Z(n17119) );
  XOR U16797 ( .A(n17182), .B(n17183), .Z(n17157) );
  AND U16798 ( .A(n17184), .B(n17185), .Z(n17183) );
  XNOR U16799 ( .A(n17182), .B(n17173), .Z(n17185) );
  IV U16800 ( .A(n17127), .Z(n17173) );
  XNOR U16801 ( .A(n17186), .B(n17166), .Z(n17127) );
  XNOR U16802 ( .A(n17187), .B(n17172), .Z(n17166) );
  XOR U16803 ( .A(n17188), .B(n17189), .Z(n17172) );
  NOR U16804 ( .A(n17190), .B(n17191), .Z(n17189) );
  XNOR U16805 ( .A(n17188), .B(n17192), .Z(n17190) );
  XNOR U16806 ( .A(n17171), .B(n17163), .Z(n17187) );
  XOR U16807 ( .A(n17193), .B(n17194), .Z(n17163) );
  AND U16808 ( .A(n17195), .B(n17196), .Z(n17194) );
  XNOR U16809 ( .A(n17193), .B(n17197), .Z(n17195) );
  XNOR U16810 ( .A(n17198), .B(n17168), .Z(n17171) );
  XOR U16811 ( .A(n17199), .B(n17200), .Z(n17168) );
  AND U16812 ( .A(n17201), .B(n17202), .Z(n17200) );
  XOR U16813 ( .A(n17199), .B(n17203), .Z(n17201) );
  XNOR U16814 ( .A(n17204), .B(n17205), .Z(n17198) );
  NOR U16815 ( .A(n17206), .B(n17207), .Z(n17205) );
  XOR U16816 ( .A(n17204), .B(n17208), .Z(n17206) );
  XNOR U16817 ( .A(n17167), .B(n17174), .Z(n17186) );
  NOR U16818 ( .A(n17135), .B(n17209), .Z(n17174) );
  XOR U16819 ( .A(n17179), .B(n17178), .Z(n17167) );
  XNOR U16820 ( .A(n17210), .B(n17175), .Z(n17178) );
  XOR U16821 ( .A(n17211), .B(n17212), .Z(n17175) );
  AND U16822 ( .A(n17213), .B(n17214), .Z(n17212) );
  XOR U16823 ( .A(n17211), .B(n17215), .Z(n17213) );
  XNOR U16824 ( .A(n17216), .B(n17217), .Z(n17210) );
  NOR U16825 ( .A(n17218), .B(n17219), .Z(n17217) );
  XNOR U16826 ( .A(n17216), .B(n17220), .Z(n17218) );
  XOR U16827 ( .A(n17221), .B(n17222), .Z(n17179) );
  NOR U16828 ( .A(n17223), .B(n17224), .Z(n17222) );
  XNOR U16829 ( .A(n17221), .B(n17225), .Z(n17223) );
  XNOR U16830 ( .A(n17124), .B(n17182), .Z(n17184) );
  XNOR U16831 ( .A(n17226), .B(n17227), .Z(n17124) );
  AND U16832 ( .A(n72), .B(n17131), .Z(n17227) );
  XOR U16833 ( .A(n17226), .B(n17129), .Z(n17131) );
  AND U16834 ( .A(n17132), .B(n17135), .Z(n17182) );
  XOR U16835 ( .A(n17228), .B(n17209), .Z(n17135) );
  XNOR U16836 ( .A(p_input[2048]), .B(p_input[48]), .Z(n17209) );
  XOR U16837 ( .A(n17197), .B(n17196), .Z(n17228) );
  XNOR U16838 ( .A(n17229), .B(n17203), .Z(n17196) );
  XNOR U16839 ( .A(n17192), .B(n17191), .Z(n17203) );
  XOR U16840 ( .A(n17230), .B(n17188), .Z(n17191) );
  XNOR U16841 ( .A(n16904), .B(p_input[58]), .Z(n17188) );
  XNOR U16842 ( .A(p_input[2059]), .B(p_input[59]), .Z(n17230) );
  XOR U16843 ( .A(p_input[2060]), .B(p_input[60]), .Z(n17192) );
  XNOR U16844 ( .A(n17202), .B(n17193), .Z(n17229) );
  XNOR U16845 ( .A(n17068), .B(p_input[49]), .Z(n17193) );
  XOR U16846 ( .A(n17231), .B(n17208), .Z(n17202) );
  XNOR U16847 ( .A(p_input[2063]), .B(p_input[63]), .Z(n17208) );
  XOR U16848 ( .A(n17199), .B(n17207), .Z(n17231) );
  XOR U16849 ( .A(n17232), .B(n17204), .Z(n17207) );
  XOR U16850 ( .A(p_input[2061]), .B(p_input[61]), .Z(n17204) );
  XNOR U16851 ( .A(p_input[2062]), .B(p_input[62]), .Z(n17232) );
  XNOR U16852 ( .A(n16738), .B(p_input[57]), .Z(n17199) );
  XNOR U16853 ( .A(n17215), .B(n17214), .Z(n17197) );
  XNOR U16854 ( .A(n17233), .B(n17220), .Z(n17214) );
  XOR U16855 ( .A(p_input[2056]), .B(p_input[56]), .Z(n17220) );
  XOR U16856 ( .A(n17211), .B(n17219), .Z(n17233) );
  XOR U16857 ( .A(n17234), .B(n17216), .Z(n17219) );
  XOR U16858 ( .A(p_input[2054]), .B(p_input[54]), .Z(n17216) );
  XNOR U16859 ( .A(p_input[2055]), .B(p_input[55]), .Z(n17234) );
  XNOR U16860 ( .A(n16741), .B(p_input[50]), .Z(n17211) );
  XNOR U16861 ( .A(n17225), .B(n17224), .Z(n17215) );
  XOR U16862 ( .A(n17235), .B(n17221), .Z(n17224) );
  XOR U16863 ( .A(p_input[2051]), .B(p_input[51]), .Z(n17221) );
  XNOR U16864 ( .A(p_input[2052]), .B(p_input[52]), .Z(n17235) );
  XOR U16865 ( .A(p_input[2053]), .B(p_input[53]), .Z(n17225) );
  XNOR U16866 ( .A(n17236), .B(n17237), .Z(n17132) );
  AND U16867 ( .A(n72), .B(n17238), .Z(n17237) );
  XNOR U16868 ( .A(n17239), .B(n17240), .Z(n72) );
  AND U16869 ( .A(n17241), .B(n17242), .Z(n17240) );
  XOR U16870 ( .A(n17239), .B(n17142), .Z(n17242) );
  XNOR U16871 ( .A(n17239), .B(n17096), .Z(n17241) );
  XOR U16872 ( .A(n17243), .B(n17244), .Z(n17239) );
  AND U16873 ( .A(n17245), .B(n17246), .Z(n17244) );
  XOR U16874 ( .A(n17243), .B(n17106), .Z(n17245) );
  XOR U16875 ( .A(n17247), .B(n17248), .Z(n17085) );
  AND U16876 ( .A(n76), .B(n17238), .Z(n17248) );
  XNOR U16877 ( .A(n17236), .B(n17247), .Z(n17238) );
  XNOR U16878 ( .A(n17249), .B(n17250), .Z(n76) );
  AND U16879 ( .A(n17251), .B(n17252), .Z(n17250) );
  XNOR U16880 ( .A(n17253), .B(n17249), .Z(n17252) );
  IV U16881 ( .A(n17142), .Z(n17253) );
  XNOR U16882 ( .A(n17254), .B(n17255), .Z(n17142) );
  AND U16883 ( .A(n79), .B(n17256), .Z(n17255) );
  XNOR U16884 ( .A(n17254), .B(n17257), .Z(n17256) );
  XNOR U16885 ( .A(n17096), .B(n17249), .Z(n17251) );
  XOR U16886 ( .A(n17258), .B(n17259), .Z(n17096) );
  AND U16887 ( .A(n87), .B(n17260), .Z(n17259) );
  XOR U16888 ( .A(n17243), .B(n17261), .Z(n17249) );
  AND U16889 ( .A(n17262), .B(n17246), .Z(n17261) );
  XNOR U16890 ( .A(n17155), .B(n17243), .Z(n17246) );
  XNOR U16891 ( .A(n17263), .B(n17264), .Z(n17155) );
  AND U16892 ( .A(n79), .B(n17265), .Z(n17264) );
  XOR U16893 ( .A(n17266), .B(n17263), .Z(n17265) );
  XNOR U16894 ( .A(n17267), .B(n17243), .Z(n17262) );
  IV U16895 ( .A(n17106), .Z(n17267) );
  XOR U16896 ( .A(n17268), .B(n17269), .Z(n17106) );
  AND U16897 ( .A(n87), .B(n17270), .Z(n17269) );
  XOR U16898 ( .A(n17271), .B(n17272), .Z(n17243) );
  AND U16899 ( .A(n17273), .B(n17274), .Z(n17272) );
  XNOR U16900 ( .A(n17180), .B(n17271), .Z(n17274) );
  XNOR U16901 ( .A(n17275), .B(n17276), .Z(n17180) );
  AND U16902 ( .A(n79), .B(n17277), .Z(n17276) );
  XNOR U16903 ( .A(n17278), .B(n17275), .Z(n17277) );
  XOR U16904 ( .A(n17271), .B(n17117), .Z(n17273) );
  XOR U16905 ( .A(n17279), .B(n17280), .Z(n17117) );
  AND U16906 ( .A(n87), .B(n17281), .Z(n17280) );
  XOR U16907 ( .A(n17282), .B(n17283), .Z(n17271) );
  AND U16908 ( .A(n17284), .B(n17285), .Z(n17283) );
  XNOR U16909 ( .A(n17282), .B(n17226), .Z(n17285) );
  XNOR U16910 ( .A(n17286), .B(n17287), .Z(n17226) );
  AND U16911 ( .A(n79), .B(n17288), .Z(n17287) );
  XOR U16912 ( .A(n17289), .B(n17286), .Z(n17288) );
  XNOR U16913 ( .A(n17290), .B(n17282), .Z(n17284) );
  IV U16914 ( .A(n17129), .Z(n17290) );
  XOR U16915 ( .A(n17291), .B(n17292), .Z(n17129) );
  AND U16916 ( .A(n87), .B(n17293), .Z(n17292) );
  AND U16917 ( .A(n17247), .B(n17236), .Z(n17282) );
  XNOR U16918 ( .A(n17294), .B(n17295), .Z(n17236) );
  AND U16919 ( .A(n79), .B(n17296), .Z(n17295) );
  XNOR U16920 ( .A(n17297), .B(n17294), .Z(n17296) );
  XNOR U16921 ( .A(n17298), .B(n17299), .Z(n79) );
  AND U16922 ( .A(n17300), .B(n17301), .Z(n17299) );
  XOR U16923 ( .A(n17257), .B(n17298), .Z(n17301) );
  AND U16924 ( .A(n17302), .B(n17303), .Z(n17257) );
  XOR U16925 ( .A(n17298), .B(n17254), .Z(n17300) );
  XNOR U16926 ( .A(n17304), .B(n17305), .Z(n17254) );
  AND U16927 ( .A(n83), .B(n17260), .Z(n17305) );
  XOR U16928 ( .A(n17258), .B(n17304), .Z(n17260) );
  XOR U16929 ( .A(n17306), .B(n17307), .Z(n17298) );
  AND U16930 ( .A(n17308), .B(n17309), .Z(n17307) );
  XNOR U16931 ( .A(n17306), .B(n17302), .Z(n17309) );
  IV U16932 ( .A(n17266), .Z(n17302) );
  XOR U16933 ( .A(n17310), .B(n17311), .Z(n17266) );
  XOR U16934 ( .A(n17312), .B(n17303), .Z(n17311) );
  AND U16935 ( .A(n17278), .B(n17313), .Z(n17303) );
  AND U16936 ( .A(n17314), .B(n17315), .Z(n17312) );
  XOR U16937 ( .A(n17316), .B(n17310), .Z(n17314) );
  XNOR U16938 ( .A(n17263), .B(n17306), .Z(n17308) );
  XNOR U16939 ( .A(n17317), .B(n17318), .Z(n17263) );
  AND U16940 ( .A(n83), .B(n17270), .Z(n17318) );
  XOR U16941 ( .A(n17317), .B(n17268), .Z(n17270) );
  XOR U16942 ( .A(n17319), .B(n17320), .Z(n17306) );
  AND U16943 ( .A(n17321), .B(n17322), .Z(n17320) );
  XNOR U16944 ( .A(n17319), .B(n17278), .Z(n17322) );
  XOR U16945 ( .A(n17323), .B(n17315), .Z(n17278) );
  XNOR U16946 ( .A(n17324), .B(n17310), .Z(n17315) );
  XOR U16947 ( .A(n17325), .B(n17326), .Z(n17310) );
  AND U16948 ( .A(n17327), .B(n17328), .Z(n17326) );
  XOR U16949 ( .A(n17329), .B(n17325), .Z(n17327) );
  XNOR U16950 ( .A(n17330), .B(n17331), .Z(n17324) );
  AND U16951 ( .A(n17332), .B(n17333), .Z(n17331) );
  XOR U16952 ( .A(n17330), .B(n17334), .Z(n17332) );
  XNOR U16953 ( .A(n17316), .B(n17313), .Z(n17323) );
  AND U16954 ( .A(n17335), .B(n17336), .Z(n17313) );
  XOR U16955 ( .A(n17337), .B(n17338), .Z(n17316) );
  AND U16956 ( .A(n17339), .B(n17340), .Z(n17338) );
  XOR U16957 ( .A(n17337), .B(n17341), .Z(n17339) );
  XNOR U16958 ( .A(n17275), .B(n17319), .Z(n17321) );
  XNOR U16959 ( .A(n17342), .B(n17343), .Z(n17275) );
  AND U16960 ( .A(n83), .B(n17281), .Z(n17343) );
  XOR U16961 ( .A(n17342), .B(n17279), .Z(n17281) );
  XOR U16962 ( .A(n17344), .B(n17345), .Z(n17319) );
  AND U16963 ( .A(n17346), .B(n17347), .Z(n17345) );
  XNOR U16964 ( .A(n17344), .B(n17335), .Z(n17347) );
  IV U16965 ( .A(n17289), .Z(n17335) );
  XNOR U16966 ( .A(n17348), .B(n17328), .Z(n17289) );
  XNOR U16967 ( .A(n17349), .B(n17334), .Z(n17328) );
  XOR U16968 ( .A(n17350), .B(n17351), .Z(n17334) );
  NOR U16969 ( .A(n17352), .B(n17353), .Z(n17351) );
  XNOR U16970 ( .A(n17350), .B(n17354), .Z(n17352) );
  XNOR U16971 ( .A(n17333), .B(n17325), .Z(n17349) );
  XOR U16972 ( .A(n17355), .B(n17356), .Z(n17325) );
  AND U16973 ( .A(n17357), .B(n17358), .Z(n17356) );
  XNOR U16974 ( .A(n17355), .B(n17359), .Z(n17357) );
  XNOR U16975 ( .A(n17360), .B(n17330), .Z(n17333) );
  XOR U16976 ( .A(n17361), .B(n17362), .Z(n17330) );
  AND U16977 ( .A(n17363), .B(n17364), .Z(n17362) );
  XOR U16978 ( .A(n17361), .B(n17365), .Z(n17363) );
  XNOR U16979 ( .A(n17366), .B(n17367), .Z(n17360) );
  NOR U16980 ( .A(n17368), .B(n17369), .Z(n17367) );
  XOR U16981 ( .A(n17366), .B(n17370), .Z(n17368) );
  XNOR U16982 ( .A(n17329), .B(n17336), .Z(n17348) );
  NOR U16983 ( .A(n17297), .B(n17371), .Z(n17336) );
  XOR U16984 ( .A(n17341), .B(n17340), .Z(n17329) );
  XNOR U16985 ( .A(n17372), .B(n17337), .Z(n17340) );
  XOR U16986 ( .A(n17373), .B(n17374), .Z(n17337) );
  AND U16987 ( .A(n17375), .B(n17376), .Z(n17374) );
  XOR U16988 ( .A(n17373), .B(n17377), .Z(n17375) );
  XNOR U16989 ( .A(n17378), .B(n17379), .Z(n17372) );
  NOR U16990 ( .A(n17380), .B(n17381), .Z(n17379) );
  XNOR U16991 ( .A(n17378), .B(n17382), .Z(n17380) );
  XOR U16992 ( .A(n17383), .B(n17384), .Z(n17341) );
  NOR U16993 ( .A(n17385), .B(n17386), .Z(n17384) );
  XNOR U16994 ( .A(n17383), .B(n17387), .Z(n17385) );
  XNOR U16995 ( .A(n17286), .B(n17344), .Z(n17346) );
  XNOR U16996 ( .A(n17388), .B(n17389), .Z(n17286) );
  AND U16997 ( .A(n83), .B(n17293), .Z(n17389) );
  XOR U16998 ( .A(n17388), .B(n17291), .Z(n17293) );
  AND U16999 ( .A(n17294), .B(n17297), .Z(n17344) );
  XOR U17000 ( .A(n17390), .B(n17371), .Z(n17297) );
  XNOR U17001 ( .A(p_input[2048]), .B(p_input[64]), .Z(n17371) );
  XOR U17002 ( .A(n17359), .B(n17358), .Z(n17390) );
  XNOR U17003 ( .A(n17391), .B(n17365), .Z(n17358) );
  XNOR U17004 ( .A(n17354), .B(n17353), .Z(n17365) );
  XOR U17005 ( .A(n17392), .B(n17350), .Z(n17353) );
  XNOR U17006 ( .A(n16904), .B(p_input[74]), .Z(n17350) );
  XNOR U17007 ( .A(p_input[2059]), .B(p_input[75]), .Z(n17392) );
  XOR U17008 ( .A(p_input[2060]), .B(p_input[76]), .Z(n17354) );
  XNOR U17009 ( .A(n17364), .B(n17355), .Z(n17391) );
  XNOR U17010 ( .A(n17068), .B(p_input[65]), .Z(n17355) );
  XOR U17011 ( .A(n17393), .B(n17370), .Z(n17364) );
  XNOR U17012 ( .A(p_input[2063]), .B(p_input[79]), .Z(n17370) );
  XOR U17013 ( .A(n17361), .B(n17369), .Z(n17393) );
  XOR U17014 ( .A(n17394), .B(n17366), .Z(n17369) );
  XOR U17015 ( .A(p_input[2061]), .B(p_input[77]), .Z(n17366) );
  XNOR U17016 ( .A(p_input[2062]), .B(p_input[78]), .Z(n17394) );
  XNOR U17017 ( .A(n16738), .B(p_input[73]), .Z(n17361) );
  XNOR U17018 ( .A(n17377), .B(n17376), .Z(n17359) );
  XNOR U17019 ( .A(n17395), .B(n17382), .Z(n17376) );
  XOR U17020 ( .A(p_input[2056]), .B(p_input[72]), .Z(n17382) );
  XOR U17021 ( .A(n17373), .B(n17381), .Z(n17395) );
  XOR U17022 ( .A(n17396), .B(n17378), .Z(n17381) );
  XOR U17023 ( .A(p_input[2054]), .B(p_input[70]), .Z(n17378) );
  XNOR U17024 ( .A(p_input[2055]), .B(p_input[71]), .Z(n17396) );
  XNOR U17025 ( .A(n16741), .B(p_input[66]), .Z(n17373) );
  XNOR U17026 ( .A(n17387), .B(n17386), .Z(n17377) );
  XOR U17027 ( .A(n17397), .B(n17383), .Z(n17386) );
  XOR U17028 ( .A(p_input[2051]), .B(p_input[67]), .Z(n17383) );
  XNOR U17029 ( .A(p_input[2052]), .B(p_input[68]), .Z(n17397) );
  XOR U17030 ( .A(p_input[2053]), .B(p_input[69]), .Z(n17387) );
  XNOR U17031 ( .A(n17398), .B(n17399), .Z(n17294) );
  AND U17032 ( .A(n83), .B(n17400), .Z(n17399) );
  XNOR U17033 ( .A(n17401), .B(n17402), .Z(n83) );
  AND U17034 ( .A(n17403), .B(n17404), .Z(n17402) );
  XOR U17035 ( .A(n17401), .B(n17304), .Z(n17404) );
  XNOR U17036 ( .A(n17401), .B(n17258), .Z(n17403) );
  XOR U17037 ( .A(n17405), .B(n17406), .Z(n17401) );
  AND U17038 ( .A(n17407), .B(n17408), .Z(n17406) );
  XOR U17039 ( .A(n17405), .B(n17268), .Z(n17407) );
  XOR U17040 ( .A(n17409), .B(n17410), .Z(n17247) );
  AND U17041 ( .A(n87), .B(n17400), .Z(n17410) );
  XNOR U17042 ( .A(n17398), .B(n17409), .Z(n17400) );
  XNOR U17043 ( .A(n17411), .B(n17412), .Z(n87) );
  AND U17044 ( .A(n17413), .B(n17414), .Z(n17412) );
  XNOR U17045 ( .A(n17415), .B(n17411), .Z(n17414) );
  IV U17046 ( .A(n17304), .Z(n17415) );
  XNOR U17047 ( .A(n17416), .B(n17417), .Z(n17304) );
  AND U17048 ( .A(n90), .B(n17418), .Z(n17417) );
  XNOR U17049 ( .A(n17416), .B(n17419), .Z(n17418) );
  XNOR U17050 ( .A(n17258), .B(n17411), .Z(n17413) );
  XOR U17051 ( .A(n17420), .B(n17421), .Z(n17258) );
  AND U17052 ( .A(n98), .B(n17422), .Z(n17421) );
  XOR U17053 ( .A(n17405), .B(n17423), .Z(n17411) );
  AND U17054 ( .A(n17424), .B(n17408), .Z(n17423) );
  XNOR U17055 ( .A(n17317), .B(n17405), .Z(n17408) );
  XNOR U17056 ( .A(n17425), .B(n17426), .Z(n17317) );
  AND U17057 ( .A(n90), .B(n17427), .Z(n17426) );
  XOR U17058 ( .A(n17428), .B(n17425), .Z(n17427) );
  XNOR U17059 ( .A(n17429), .B(n17405), .Z(n17424) );
  IV U17060 ( .A(n17268), .Z(n17429) );
  XOR U17061 ( .A(n17430), .B(n17431), .Z(n17268) );
  AND U17062 ( .A(n98), .B(n17432), .Z(n17431) );
  XOR U17063 ( .A(n17433), .B(n17434), .Z(n17405) );
  AND U17064 ( .A(n17435), .B(n17436), .Z(n17434) );
  XNOR U17065 ( .A(n17342), .B(n17433), .Z(n17436) );
  XNOR U17066 ( .A(n17437), .B(n17438), .Z(n17342) );
  AND U17067 ( .A(n90), .B(n17439), .Z(n17438) );
  XNOR U17068 ( .A(n17440), .B(n17437), .Z(n17439) );
  XOR U17069 ( .A(n17433), .B(n17279), .Z(n17435) );
  XOR U17070 ( .A(n17441), .B(n17442), .Z(n17279) );
  AND U17071 ( .A(n98), .B(n17443), .Z(n17442) );
  XOR U17072 ( .A(n17444), .B(n17445), .Z(n17433) );
  AND U17073 ( .A(n17446), .B(n17447), .Z(n17445) );
  XNOR U17074 ( .A(n17444), .B(n17388), .Z(n17447) );
  XNOR U17075 ( .A(n17448), .B(n17449), .Z(n17388) );
  AND U17076 ( .A(n90), .B(n17450), .Z(n17449) );
  XOR U17077 ( .A(n17451), .B(n17448), .Z(n17450) );
  XNOR U17078 ( .A(n17452), .B(n17444), .Z(n17446) );
  IV U17079 ( .A(n17291), .Z(n17452) );
  XOR U17080 ( .A(n17453), .B(n17454), .Z(n17291) );
  AND U17081 ( .A(n98), .B(n17455), .Z(n17454) );
  AND U17082 ( .A(n17409), .B(n17398), .Z(n17444) );
  XNOR U17083 ( .A(n17456), .B(n17457), .Z(n17398) );
  AND U17084 ( .A(n90), .B(n17458), .Z(n17457) );
  XNOR U17085 ( .A(n17459), .B(n17456), .Z(n17458) );
  XNOR U17086 ( .A(n17460), .B(n17461), .Z(n90) );
  AND U17087 ( .A(n17462), .B(n17463), .Z(n17461) );
  XOR U17088 ( .A(n17419), .B(n17460), .Z(n17463) );
  AND U17089 ( .A(n17464), .B(n17465), .Z(n17419) );
  XOR U17090 ( .A(n17460), .B(n17416), .Z(n17462) );
  XNOR U17091 ( .A(n17466), .B(n17467), .Z(n17416) );
  AND U17092 ( .A(n94), .B(n17422), .Z(n17467) );
  XOR U17093 ( .A(n17420), .B(n17466), .Z(n17422) );
  XOR U17094 ( .A(n17468), .B(n17469), .Z(n17460) );
  AND U17095 ( .A(n17470), .B(n17471), .Z(n17469) );
  XNOR U17096 ( .A(n17468), .B(n17464), .Z(n17471) );
  IV U17097 ( .A(n17428), .Z(n17464) );
  XOR U17098 ( .A(n17472), .B(n17473), .Z(n17428) );
  XOR U17099 ( .A(n17474), .B(n17465), .Z(n17473) );
  AND U17100 ( .A(n17440), .B(n17475), .Z(n17465) );
  AND U17101 ( .A(n17476), .B(n17477), .Z(n17474) );
  XOR U17102 ( .A(n17478), .B(n17472), .Z(n17476) );
  XNOR U17103 ( .A(n17425), .B(n17468), .Z(n17470) );
  XNOR U17104 ( .A(n17479), .B(n17480), .Z(n17425) );
  AND U17105 ( .A(n94), .B(n17432), .Z(n17480) );
  XOR U17106 ( .A(n17479), .B(n17430), .Z(n17432) );
  XOR U17107 ( .A(n17481), .B(n17482), .Z(n17468) );
  AND U17108 ( .A(n17483), .B(n17484), .Z(n17482) );
  XNOR U17109 ( .A(n17481), .B(n17440), .Z(n17484) );
  XOR U17110 ( .A(n17485), .B(n17477), .Z(n17440) );
  XNOR U17111 ( .A(n17486), .B(n17472), .Z(n17477) );
  XOR U17112 ( .A(n17487), .B(n17488), .Z(n17472) );
  AND U17113 ( .A(n17489), .B(n17490), .Z(n17488) );
  XOR U17114 ( .A(n17491), .B(n17487), .Z(n17489) );
  XNOR U17115 ( .A(n17492), .B(n17493), .Z(n17486) );
  AND U17116 ( .A(n17494), .B(n17495), .Z(n17493) );
  XOR U17117 ( .A(n17492), .B(n17496), .Z(n17494) );
  XNOR U17118 ( .A(n17478), .B(n17475), .Z(n17485) );
  AND U17119 ( .A(n17497), .B(n17498), .Z(n17475) );
  XOR U17120 ( .A(n17499), .B(n17500), .Z(n17478) );
  AND U17121 ( .A(n17501), .B(n17502), .Z(n17500) );
  XOR U17122 ( .A(n17499), .B(n17503), .Z(n17501) );
  XNOR U17123 ( .A(n17437), .B(n17481), .Z(n17483) );
  XNOR U17124 ( .A(n17504), .B(n17505), .Z(n17437) );
  AND U17125 ( .A(n94), .B(n17443), .Z(n17505) );
  XOR U17126 ( .A(n17504), .B(n17441), .Z(n17443) );
  XOR U17127 ( .A(n17506), .B(n17507), .Z(n17481) );
  AND U17128 ( .A(n17508), .B(n17509), .Z(n17507) );
  XNOR U17129 ( .A(n17506), .B(n17497), .Z(n17509) );
  IV U17130 ( .A(n17451), .Z(n17497) );
  XNOR U17131 ( .A(n17510), .B(n17490), .Z(n17451) );
  XNOR U17132 ( .A(n17511), .B(n17496), .Z(n17490) );
  XOR U17133 ( .A(n17512), .B(n17513), .Z(n17496) );
  NOR U17134 ( .A(n17514), .B(n17515), .Z(n17513) );
  XNOR U17135 ( .A(n17512), .B(n17516), .Z(n17514) );
  XNOR U17136 ( .A(n17495), .B(n17487), .Z(n17511) );
  XOR U17137 ( .A(n17517), .B(n17518), .Z(n17487) );
  AND U17138 ( .A(n17519), .B(n17520), .Z(n17518) );
  XNOR U17139 ( .A(n17517), .B(n17521), .Z(n17519) );
  XNOR U17140 ( .A(n17522), .B(n17492), .Z(n17495) );
  XOR U17141 ( .A(n17523), .B(n17524), .Z(n17492) );
  AND U17142 ( .A(n17525), .B(n17526), .Z(n17524) );
  XOR U17143 ( .A(n17523), .B(n17527), .Z(n17525) );
  XNOR U17144 ( .A(n17528), .B(n17529), .Z(n17522) );
  NOR U17145 ( .A(n17530), .B(n17531), .Z(n17529) );
  XOR U17146 ( .A(n17528), .B(n17532), .Z(n17530) );
  XNOR U17147 ( .A(n17491), .B(n17498), .Z(n17510) );
  NOR U17148 ( .A(n17459), .B(n17533), .Z(n17498) );
  XOR U17149 ( .A(n17503), .B(n17502), .Z(n17491) );
  XNOR U17150 ( .A(n17534), .B(n17499), .Z(n17502) );
  XOR U17151 ( .A(n17535), .B(n17536), .Z(n17499) );
  AND U17152 ( .A(n17537), .B(n17538), .Z(n17536) );
  XOR U17153 ( .A(n17535), .B(n17539), .Z(n17537) );
  XNOR U17154 ( .A(n17540), .B(n17541), .Z(n17534) );
  NOR U17155 ( .A(n17542), .B(n17543), .Z(n17541) );
  XNOR U17156 ( .A(n17540), .B(n17544), .Z(n17542) );
  XOR U17157 ( .A(n17545), .B(n17546), .Z(n17503) );
  NOR U17158 ( .A(n17547), .B(n17548), .Z(n17546) );
  XNOR U17159 ( .A(n17545), .B(n17549), .Z(n17547) );
  XNOR U17160 ( .A(n17448), .B(n17506), .Z(n17508) );
  XNOR U17161 ( .A(n17550), .B(n17551), .Z(n17448) );
  AND U17162 ( .A(n94), .B(n17455), .Z(n17551) );
  XOR U17163 ( .A(n17550), .B(n17453), .Z(n17455) );
  AND U17164 ( .A(n17456), .B(n17459), .Z(n17506) );
  XOR U17165 ( .A(n17552), .B(n17533), .Z(n17459) );
  XNOR U17166 ( .A(p_input[2048]), .B(p_input[80]), .Z(n17533) );
  XOR U17167 ( .A(n17521), .B(n17520), .Z(n17552) );
  XNOR U17168 ( .A(n17553), .B(n17527), .Z(n17520) );
  XNOR U17169 ( .A(n17516), .B(n17515), .Z(n17527) );
  XOR U17170 ( .A(n17554), .B(n17512), .Z(n17515) );
  XNOR U17171 ( .A(n16904), .B(p_input[90]), .Z(n17512) );
  XNOR U17172 ( .A(p_input[2059]), .B(p_input[91]), .Z(n17554) );
  XOR U17173 ( .A(p_input[2060]), .B(p_input[92]), .Z(n17516) );
  XNOR U17174 ( .A(n17526), .B(n17517), .Z(n17553) );
  XNOR U17175 ( .A(n17068), .B(p_input[81]), .Z(n17517) );
  XOR U17176 ( .A(n17555), .B(n17532), .Z(n17526) );
  XNOR U17177 ( .A(p_input[2063]), .B(p_input[95]), .Z(n17532) );
  XOR U17178 ( .A(n17523), .B(n17531), .Z(n17555) );
  XOR U17179 ( .A(n17556), .B(n17528), .Z(n17531) );
  XOR U17180 ( .A(p_input[2061]), .B(p_input[93]), .Z(n17528) );
  XNOR U17181 ( .A(p_input[2062]), .B(p_input[94]), .Z(n17556) );
  XNOR U17182 ( .A(n16738), .B(p_input[89]), .Z(n17523) );
  XNOR U17183 ( .A(n17539), .B(n17538), .Z(n17521) );
  XNOR U17184 ( .A(n17557), .B(n17544), .Z(n17538) );
  XOR U17185 ( .A(p_input[2056]), .B(p_input[88]), .Z(n17544) );
  XOR U17186 ( .A(n17535), .B(n17543), .Z(n17557) );
  XOR U17187 ( .A(n17558), .B(n17540), .Z(n17543) );
  XOR U17188 ( .A(p_input[2054]), .B(p_input[86]), .Z(n17540) );
  XNOR U17189 ( .A(p_input[2055]), .B(p_input[87]), .Z(n17558) );
  XNOR U17190 ( .A(n16741), .B(p_input[82]), .Z(n17535) );
  XNOR U17191 ( .A(n17549), .B(n17548), .Z(n17539) );
  XOR U17192 ( .A(n17559), .B(n17545), .Z(n17548) );
  XOR U17193 ( .A(p_input[2051]), .B(p_input[83]), .Z(n17545) );
  XNOR U17194 ( .A(p_input[2052]), .B(p_input[84]), .Z(n17559) );
  XOR U17195 ( .A(p_input[2053]), .B(p_input[85]), .Z(n17549) );
  XNOR U17196 ( .A(n17560), .B(n17561), .Z(n17456) );
  AND U17197 ( .A(n94), .B(n17562), .Z(n17561) );
  XNOR U17198 ( .A(n17563), .B(n17564), .Z(n94) );
  AND U17199 ( .A(n17565), .B(n17566), .Z(n17564) );
  XOR U17200 ( .A(n17563), .B(n17466), .Z(n17566) );
  XNOR U17201 ( .A(n17563), .B(n17420), .Z(n17565) );
  XOR U17202 ( .A(n17567), .B(n17568), .Z(n17563) );
  AND U17203 ( .A(n17569), .B(n17570), .Z(n17568) );
  XOR U17204 ( .A(n17567), .B(n17430), .Z(n17569) );
  XOR U17205 ( .A(n17571), .B(n17572), .Z(n17409) );
  AND U17206 ( .A(n98), .B(n17562), .Z(n17572) );
  XNOR U17207 ( .A(n17560), .B(n17571), .Z(n17562) );
  XNOR U17208 ( .A(n17573), .B(n17574), .Z(n98) );
  AND U17209 ( .A(n17575), .B(n17576), .Z(n17574) );
  XNOR U17210 ( .A(n17577), .B(n17573), .Z(n17576) );
  IV U17211 ( .A(n17466), .Z(n17577) );
  XNOR U17212 ( .A(n17578), .B(n17579), .Z(n17466) );
  AND U17213 ( .A(n101), .B(n17580), .Z(n17579) );
  XNOR U17214 ( .A(n17578), .B(n17581), .Z(n17580) );
  XNOR U17215 ( .A(n17420), .B(n17573), .Z(n17575) );
  XOR U17216 ( .A(n17582), .B(n17583), .Z(n17420) );
  AND U17217 ( .A(n109), .B(n17584), .Z(n17583) );
  XOR U17218 ( .A(n17567), .B(n17585), .Z(n17573) );
  AND U17219 ( .A(n17586), .B(n17570), .Z(n17585) );
  XNOR U17220 ( .A(n17479), .B(n17567), .Z(n17570) );
  XNOR U17221 ( .A(n17587), .B(n17588), .Z(n17479) );
  AND U17222 ( .A(n101), .B(n17589), .Z(n17588) );
  XOR U17223 ( .A(n17590), .B(n17587), .Z(n17589) );
  XNOR U17224 ( .A(n17591), .B(n17567), .Z(n17586) );
  IV U17225 ( .A(n17430), .Z(n17591) );
  XOR U17226 ( .A(n17592), .B(n17593), .Z(n17430) );
  AND U17227 ( .A(n109), .B(n17594), .Z(n17593) );
  XOR U17228 ( .A(n17595), .B(n17596), .Z(n17567) );
  AND U17229 ( .A(n17597), .B(n17598), .Z(n17596) );
  XNOR U17230 ( .A(n17504), .B(n17595), .Z(n17598) );
  XNOR U17231 ( .A(n17599), .B(n17600), .Z(n17504) );
  AND U17232 ( .A(n101), .B(n17601), .Z(n17600) );
  XNOR U17233 ( .A(n17602), .B(n17599), .Z(n17601) );
  XOR U17234 ( .A(n17595), .B(n17441), .Z(n17597) );
  XOR U17235 ( .A(n17603), .B(n17604), .Z(n17441) );
  AND U17236 ( .A(n109), .B(n17605), .Z(n17604) );
  XOR U17237 ( .A(n17606), .B(n17607), .Z(n17595) );
  AND U17238 ( .A(n17608), .B(n17609), .Z(n17607) );
  XNOR U17239 ( .A(n17606), .B(n17550), .Z(n17609) );
  XNOR U17240 ( .A(n17610), .B(n17611), .Z(n17550) );
  AND U17241 ( .A(n101), .B(n17612), .Z(n17611) );
  XOR U17242 ( .A(n17613), .B(n17610), .Z(n17612) );
  XNOR U17243 ( .A(n17614), .B(n17606), .Z(n17608) );
  IV U17244 ( .A(n17453), .Z(n17614) );
  XOR U17245 ( .A(n17615), .B(n17616), .Z(n17453) );
  AND U17246 ( .A(n109), .B(n17617), .Z(n17616) );
  AND U17247 ( .A(n17571), .B(n17560), .Z(n17606) );
  XNOR U17248 ( .A(n17618), .B(n17619), .Z(n17560) );
  AND U17249 ( .A(n101), .B(n17620), .Z(n17619) );
  XNOR U17250 ( .A(n17621), .B(n17618), .Z(n17620) );
  XNOR U17251 ( .A(n17622), .B(n17623), .Z(n101) );
  AND U17252 ( .A(n17624), .B(n17625), .Z(n17623) );
  XOR U17253 ( .A(n17581), .B(n17622), .Z(n17625) );
  AND U17254 ( .A(n17626), .B(n17627), .Z(n17581) );
  XOR U17255 ( .A(n17622), .B(n17578), .Z(n17624) );
  XNOR U17256 ( .A(n17628), .B(n17629), .Z(n17578) );
  AND U17257 ( .A(n105), .B(n17584), .Z(n17629) );
  XOR U17258 ( .A(n17582), .B(n17628), .Z(n17584) );
  XOR U17259 ( .A(n17630), .B(n17631), .Z(n17622) );
  AND U17260 ( .A(n17632), .B(n17633), .Z(n17631) );
  XNOR U17261 ( .A(n17630), .B(n17626), .Z(n17633) );
  IV U17262 ( .A(n17590), .Z(n17626) );
  XOR U17263 ( .A(n17634), .B(n17635), .Z(n17590) );
  XOR U17264 ( .A(n17636), .B(n17627), .Z(n17635) );
  AND U17265 ( .A(n17602), .B(n17637), .Z(n17627) );
  AND U17266 ( .A(n17638), .B(n17639), .Z(n17636) );
  XOR U17267 ( .A(n17640), .B(n17634), .Z(n17638) );
  XNOR U17268 ( .A(n17587), .B(n17630), .Z(n17632) );
  XNOR U17269 ( .A(n17641), .B(n17642), .Z(n17587) );
  AND U17270 ( .A(n105), .B(n17594), .Z(n17642) );
  XOR U17271 ( .A(n17641), .B(n17592), .Z(n17594) );
  XOR U17272 ( .A(n17643), .B(n17644), .Z(n17630) );
  AND U17273 ( .A(n17645), .B(n17646), .Z(n17644) );
  XNOR U17274 ( .A(n17643), .B(n17602), .Z(n17646) );
  XOR U17275 ( .A(n17647), .B(n17639), .Z(n17602) );
  XNOR U17276 ( .A(n17648), .B(n17634), .Z(n17639) );
  XOR U17277 ( .A(n17649), .B(n17650), .Z(n17634) );
  AND U17278 ( .A(n17651), .B(n17652), .Z(n17650) );
  XOR U17279 ( .A(n17653), .B(n17649), .Z(n17651) );
  XNOR U17280 ( .A(n17654), .B(n17655), .Z(n17648) );
  AND U17281 ( .A(n17656), .B(n17657), .Z(n17655) );
  XOR U17282 ( .A(n17654), .B(n17658), .Z(n17656) );
  XNOR U17283 ( .A(n17640), .B(n17637), .Z(n17647) );
  AND U17284 ( .A(n17659), .B(n17660), .Z(n17637) );
  XOR U17285 ( .A(n17661), .B(n17662), .Z(n17640) );
  AND U17286 ( .A(n17663), .B(n17664), .Z(n17662) );
  XOR U17287 ( .A(n17661), .B(n17665), .Z(n17663) );
  XNOR U17288 ( .A(n17599), .B(n17643), .Z(n17645) );
  XNOR U17289 ( .A(n17666), .B(n17667), .Z(n17599) );
  AND U17290 ( .A(n105), .B(n17605), .Z(n17667) );
  XOR U17291 ( .A(n17666), .B(n17603), .Z(n17605) );
  XOR U17292 ( .A(n17668), .B(n17669), .Z(n17643) );
  AND U17293 ( .A(n17670), .B(n17671), .Z(n17669) );
  XNOR U17294 ( .A(n17668), .B(n17659), .Z(n17671) );
  IV U17295 ( .A(n17613), .Z(n17659) );
  XNOR U17296 ( .A(n17672), .B(n17652), .Z(n17613) );
  XNOR U17297 ( .A(n17673), .B(n17658), .Z(n17652) );
  XNOR U17298 ( .A(n17674), .B(n17675), .Z(n17658) );
  NOR U17299 ( .A(n17676), .B(n17677), .Z(n17675) );
  XOR U17300 ( .A(n17674), .B(n17678), .Z(n17676) );
  XNOR U17301 ( .A(n17657), .B(n17649), .Z(n17673) );
  XOR U17302 ( .A(n17679), .B(n17680), .Z(n17649) );
  AND U17303 ( .A(n17681), .B(n17682), .Z(n17680) );
  XOR U17304 ( .A(n17679), .B(n17683), .Z(n17681) );
  XNOR U17305 ( .A(n17684), .B(n17654), .Z(n17657) );
  XOR U17306 ( .A(n17685), .B(n17686), .Z(n17654) );
  AND U17307 ( .A(n17687), .B(n17688), .Z(n17686) );
  XNOR U17308 ( .A(n17689), .B(n17690), .Z(n17687) );
  IV U17309 ( .A(n17685), .Z(n17689) );
  XNOR U17310 ( .A(n17691), .B(n17692), .Z(n17684) );
  NOR U17311 ( .A(n17693), .B(n17694), .Z(n17692) );
  XNOR U17312 ( .A(n17691), .B(n17695), .Z(n17693) );
  XNOR U17313 ( .A(n17653), .B(n17660), .Z(n17672) );
  NOR U17314 ( .A(n17621), .B(n17696), .Z(n17660) );
  XOR U17315 ( .A(n17665), .B(n17664), .Z(n17653) );
  XNOR U17316 ( .A(n17697), .B(n17661), .Z(n17664) );
  XOR U17317 ( .A(n17698), .B(n17699), .Z(n17661) );
  AND U17318 ( .A(n17700), .B(n17701), .Z(n17699) );
  XOR U17319 ( .A(n17698), .B(n17702), .Z(n17700) );
  XNOR U17320 ( .A(n17703), .B(n17704), .Z(n17697) );
  NOR U17321 ( .A(n17705), .B(n17706), .Z(n17704) );
  XNOR U17322 ( .A(n17703), .B(n17707), .Z(n17705) );
  XOR U17323 ( .A(n17708), .B(n17709), .Z(n17665) );
  NOR U17324 ( .A(n17710), .B(n17711), .Z(n17709) );
  XNOR U17325 ( .A(n17708), .B(n17712), .Z(n17710) );
  XNOR U17326 ( .A(n17610), .B(n17668), .Z(n17670) );
  XNOR U17327 ( .A(n17713), .B(n17714), .Z(n17610) );
  AND U17328 ( .A(n105), .B(n17617), .Z(n17714) );
  XOR U17329 ( .A(n17713), .B(n17615), .Z(n17617) );
  AND U17330 ( .A(n17618), .B(n17621), .Z(n17668) );
  XOR U17331 ( .A(n17715), .B(n17696), .Z(n17621) );
  XNOR U17332 ( .A(p_input[2048]), .B(p_input[96]), .Z(n17696) );
  XNOR U17333 ( .A(n17683), .B(n17682), .Z(n17715) );
  XNOR U17334 ( .A(n17716), .B(n17690), .Z(n17682) );
  XNOR U17335 ( .A(n17678), .B(n17677), .Z(n17690) );
  XNOR U17336 ( .A(n17717), .B(n17674), .Z(n17677) );
  XNOR U17337 ( .A(p_input[106]), .B(p_input[2058]), .Z(n17674) );
  XOR U17338 ( .A(p_input[107]), .B(n16732), .Z(n17717) );
  XOR U17339 ( .A(p_input[108]), .B(p_input[2060]), .Z(n17678) );
  XNOR U17340 ( .A(n17688), .B(n17679), .Z(n17716) );
  XNOR U17341 ( .A(n17068), .B(p_input[97]), .Z(n17679) );
  XNOR U17342 ( .A(n17718), .B(n17695), .Z(n17688) );
  XNOR U17343 ( .A(p_input[111]), .B(n16735), .Z(n17695) );
  XOR U17344 ( .A(n17685), .B(n17694), .Z(n17718) );
  XOR U17345 ( .A(n17719), .B(n17691), .Z(n17694) );
  XOR U17346 ( .A(p_input[109]), .B(p_input[2061]), .Z(n17691) );
  XOR U17347 ( .A(p_input[110]), .B(n16737), .Z(n17719) );
  XOR U17348 ( .A(p_input[105]), .B(p_input[2057]), .Z(n17685) );
  XOR U17349 ( .A(n17702), .B(n17701), .Z(n17683) );
  XNOR U17350 ( .A(n17720), .B(n17707), .Z(n17701) );
  XOR U17351 ( .A(p_input[104]), .B(p_input[2056]), .Z(n17707) );
  XOR U17352 ( .A(n17698), .B(n17706), .Z(n17720) );
  XOR U17353 ( .A(n17721), .B(n17703), .Z(n17706) );
  XOR U17354 ( .A(p_input[102]), .B(p_input[2054]), .Z(n17703) );
  XOR U17355 ( .A(p_input[103]), .B(n17722), .Z(n17721) );
  XNOR U17356 ( .A(n16741), .B(p_input[98]), .Z(n17698) );
  XNOR U17357 ( .A(n17712), .B(n17711), .Z(n17702) );
  XOR U17358 ( .A(n17723), .B(n17708), .Z(n17711) );
  XOR U17359 ( .A(p_input[2051]), .B(p_input[99]), .Z(n17708) );
  XOR U17360 ( .A(p_input[100]), .B(n17724), .Z(n17723) );
  XOR U17361 ( .A(p_input[101]), .B(p_input[2053]), .Z(n17712) );
  XNOR U17362 ( .A(n17725), .B(n17726), .Z(n17618) );
  AND U17363 ( .A(n105), .B(n17727), .Z(n17726) );
  XNOR U17364 ( .A(n17728), .B(n17729), .Z(n105) );
  AND U17365 ( .A(n17730), .B(n17731), .Z(n17729) );
  XOR U17366 ( .A(n17728), .B(n17628), .Z(n17731) );
  XNOR U17367 ( .A(n17728), .B(n17582), .Z(n17730) );
  XOR U17368 ( .A(n17732), .B(n17733), .Z(n17728) );
  AND U17369 ( .A(n17734), .B(n17735), .Z(n17733) );
  XOR U17370 ( .A(n17732), .B(n17592), .Z(n17734) );
  XOR U17371 ( .A(n17736), .B(n17737), .Z(n17571) );
  AND U17372 ( .A(n109), .B(n17727), .Z(n17737) );
  XNOR U17373 ( .A(n17725), .B(n17736), .Z(n17727) );
  XNOR U17374 ( .A(n17738), .B(n17739), .Z(n109) );
  AND U17375 ( .A(n17740), .B(n17741), .Z(n17739) );
  XNOR U17376 ( .A(n17742), .B(n17738), .Z(n17741) );
  IV U17377 ( .A(n17628), .Z(n17742) );
  XNOR U17378 ( .A(n17743), .B(n17744), .Z(n17628) );
  AND U17379 ( .A(n112), .B(n17745), .Z(n17744) );
  XNOR U17380 ( .A(n17743), .B(n17746), .Z(n17745) );
  XNOR U17381 ( .A(n17582), .B(n17738), .Z(n17740) );
  XOR U17382 ( .A(n17747), .B(n17748), .Z(n17582) );
  AND U17383 ( .A(n120), .B(n17749), .Z(n17748) );
  XOR U17384 ( .A(n17732), .B(n17750), .Z(n17738) );
  AND U17385 ( .A(n17751), .B(n17735), .Z(n17750) );
  XNOR U17386 ( .A(n17641), .B(n17732), .Z(n17735) );
  XNOR U17387 ( .A(n17752), .B(n17753), .Z(n17641) );
  AND U17388 ( .A(n112), .B(n17754), .Z(n17753) );
  XOR U17389 ( .A(n17755), .B(n17752), .Z(n17754) );
  XNOR U17390 ( .A(n17756), .B(n17732), .Z(n17751) );
  IV U17391 ( .A(n17592), .Z(n17756) );
  XOR U17392 ( .A(n17757), .B(n17758), .Z(n17592) );
  AND U17393 ( .A(n120), .B(n17759), .Z(n17758) );
  XOR U17394 ( .A(n17760), .B(n17761), .Z(n17732) );
  AND U17395 ( .A(n17762), .B(n17763), .Z(n17761) );
  XNOR U17396 ( .A(n17666), .B(n17760), .Z(n17763) );
  XNOR U17397 ( .A(n17764), .B(n17765), .Z(n17666) );
  AND U17398 ( .A(n112), .B(n17766), .Z(n17765) );
  XNOR U17399 ( .A(n17767), .B(n17764), .Z(n17766) );
  XOR U17400 ( .A(n17760), .B(n17603), .Z(n17762) );
  XOR U17401 ( .A(n17768), .B(n17769), .Z(n17603) );
  AND U17402 ( .A(n120), .B(n17770), .Z(n17769) );
  XOR U17403 ( .A(n17771), .B(n17772), .Z(n17760) );
  AND U17404 ( .A(n17773), .B(n17774), .Z(n17772) );
  XNOR U17405 ( .A(n17771), .B(n17713), .Z(n17774) );
  XNOR U17406 ( .A(n17775), .B(n17776), .Z(n17713) );
  AND U17407 ( .A(n112), .B(n17777), .Z(n17776) );
  XOR U17408 ( .A(n17778), .B(n17775), .Z(n17777) );
  XNOR U17409 ( .A(n17779), .B(n17771), .Z(n17773) );
  IV U17410 ( .A(n17615), .Z(n17779) );
  XOR U17411 ( .A(n17780), .B(n17781), .Z(n17615) );
  AND U17412 ( .A(n120), .B(n17782), .Z(n17781) );
  AND U17413 ( .A(n17736), .B(n17725), .Z(n17771) );
  XNOR U17414 ( .A(n17783), .B(n17784), .Z(n17725) );
  AND U17415 ( .A(n112), .B(n17785), .Z(n17784) );
  XNOR U17416 ( .A(n17786), .B(n17783), .Z(n17785) );
  XNOR U17417 ( .A(n17787), .B(n17788), .Z(n112) );
  AND U17418 ( .A(n17789), .B(n17790), .Z(n17788) );
  XOR U17419 ( .A(n17746), .B(n17787), .Z(n17790) );
  AND U17420 ( .A(n17791), .B(n17792), .Z(n17746) );
  XOR U17421 ( .A(n17787), .B(n17743), .Z(n17789) );
  XNOR U17422 ( .A(n17793), .B(n17794), .Z(n17743) );
  AND U17423 ( .A(n116), .B(n17749), .Z(n17794) );
  XOR U17424 ( .A(n17747), .B(n17793), .Z(n17749) );
  XOR U17425 ( .A(n17795), .B(n17796), .Z(n17787) );
  AND U17426 ( .A(n17797), .B(n17798), .Z(n17796) );
  XNOR U17427 ( .A(n17795), .B(n17791), .Z(n17798) );
  IV U17428 ( .A(n17755), .Z(n17791) );
  XOR U17429 ( .A(n17799), .B(n17800), .Z(n17755) );
  XOR U17430 ( .A(n17801), .B(n17792), .Z(n17800) );
  AND U17431 ( .A(n17767), .B(n17802), .Z(n17792) );
  AND U17432 ( .A(n17803), .B(n17804), .Z(n17801) );
  XOR U17433 ( .A(n17805), .B(n17799), .Z(n17803) );
  XNOR U17434 ( .A(n17752), .B(n17795), .Z(n17797) );
  XNOR U17435 ( .A(n17806), .B(n17807), .Z(n17752) );
  AND U17436 ( .A(n116), .B(n17759), .Z(n17807) );
  XOR U17437 ( .A(n17806), .B(n17757), .Z(n17759) );
  XOR U17438 ( .A(n17808), .B(n17809), .Z(n17795) );
  AND U17439 ( .A(n17810), .B(n17811), .Z(n17809) );
  XNOR U17440 ( .A(n17808), .B(n17767), .Z(n17811) );
  XOR U17441 ( .A(n17812), .B(n17804), .Z(n17767) );
  XNOR U17442 ( .A(n17813), .B(n17799), .Z(n17804) );
  XOR U17443 ( .A(n17814), .B(n17815), .Z(n17799) );
  AND U17444 ( .A(n17816), .B(n17817), .Z(n17815) );
  XOR U17445 ( .A(n17818), .B(n17814), .Z(n17816) );
  XNOR U17446 ( .A(n17819), .B(n17820), .Z(n17813) );
  AND U17447 ( .A(n17821), .B(n17822), .Z(n17820) );
  XOR U17448 ( .A(n17819), .B(n17823), .Z(n17821) );
  XNOR U17449 ( .A(n17805), .B(n17802), .Z(n17812) );
  AND U17450 ( .A(n17824), .B(n17825), .Z(n17802) );
  XOR U17451 ( .A(n17826), .B(n17827), .Z(n17805) );
  AND U17452 ( .A(n17828), .B(n17829), .Z(n17827) );
  XOR U17453 ( .A(n17826), .B(n17830), .Z(n17828) );
  XNOR U17454 ( .A(n17764), .B(n17808), .Z(n17810) );
  XNOR U17455 ( .A(n17831), .B(n17832), .Z(n17764) );
  AND U17456 ( .A(n116), .B(n17770), .Z(n17832) );
  XOR U17457 ( .A(n17831), .B(n17768), .Z(n17770) );
  XOR U17458 ( .A(n17833), .B(n17834), .Z(n17808) );
  AND U17459 ( .A(n17835), .B(n17836), .Z(n17834) );
  XNOR U17460 ( .A(n17833), .B(n17824), .Z(n17836) );
  IV U17461 ( .A(n17778), .Z(n17824) );
  XNOR U17462 ( .A(n17837), .B(n17817), .Z(n17778) );
  XNOR U17463 ( .A(n17838), .B(n17823), .Z(n17817) );
  XNOR U17464 ( .A(n17839), .B(n17840), .Z(n17823) );
  NOR U17465 ( .A(n17841), .B(n17842), .Z(n17840) );
  XOR U17466 ( .A(n17839), .B(n17843), .Z(n17841) );
  XNOR U17467 ( .A(n17822), .B(n17814), .Z(n17838) );
  XOR U17468 ( .A(n17844), .B(n17845), .Z(n17814) );
  AND U17469 ( .A(n17846), .B(n17847), .Z(n17845) );
  XOR U17470 ( .A(n17844), .B(n17848), .Z(n17846) );
  XNOR U17471 ( .A(n17849), .B(n17819), .Z(n17822) );
  XOR U17472 ( .A(n17850), .B(n17851), .Z(n17819) );
  AND U17473 ( .A(n17852), .B(n17853), .Z(n17851) );
  XNOR U17474 ( .A(n17854), .B(n17855), .Z(n17852) );
  IV U17475 ( .A(n17850), .Z(n17854) );
  XNOR U17476 ( .A(n17856), .B(n17857), .Z(n17849) );
  NOR U17477 ( .A(n17858), .B(n17859), .Z(n17857) );
  XNOR U17478 ( .A(n17856), .B(n17860), .Z(n17858) );
  XNOR U17479 ( .A(n17818), .B(n17825), .Z(n17837) );
  NOR U17480 ( .A(n17786), .B(n17861), .Z(n17825) );
  XOR U17481 ( .A(n17830), .B(n17829), .Z(n17818) );
  XNOR U17482 ( .A(n17862), .B(n17826), .Z(n17829) );
  XOR U17483 ( .A(n17863), .B(n17864), .Z(n17826) );
  AND U17484 ( .A(n17865), .B(n17866), .Z(n17864) );
  XNOR U17485 ( .A(n17867), .B(n17868), .Z(n17865) );
  IV U17486 ( .A(n17863), .Z(n17867) );
  XNOR U17487 ( .A(n17869), .B(n17870), .Z(n17862) );
  NOR U17488 ( .A(n17871), .B(n17872), .Z(n17870) );
  XNOR U17489 ( .A(n17869), .B(n17873), .Z(n17871) );
  XOR U17490 ( .A(n17874), .B(n17875), .Z(n17830) );
  NOR U17491 ( .A(n17876), .B(n17877), .Z(n17875) );
  XNOR U17492 ( .A(n17874), .B(n17878), .Z(n17876) );
  XNOR U17493 ( .A(n17775), .B(n17833), .Z(n17835) );
  XNOR U17494 ( .A(n17879), .B(n17880), .Z(n17775) );
  AND U17495 ( .A(n116), .B(n17782), .Z(n17880) );
  XOR U17496 ( .A(n17879), .B(n17780), .Z(n17782) );
  AND U17497 ( .A(n17783), .B(n17786), .Z(n17833) );
  XOR U17498 ( .A(n17881), .B(n17861), .Z(n17786) );
  XNOR U17499 ( .A(p_input[112]), .B(p_input[2048]), .Z(n17861) );
  XNOR U17500 ( .A(n17848), .B(n17847), .Z(n17881) );
  XNOR U17501 ( .A(n17882), .B(n17855), .Z(n17847) );
  XNOR U17502 ( .A(n17843), .B(n17842), .Z(n17855) );
  XNOR U17503 ( .A(n17883), .B(n17839), .Z(n17842) );
  XNOR U17504 ( .A(p_input[122]), .B(p_input[2058]), .Z(n17839) );
  XOR U17505 ( .A(p_input[123]), .B(n16732), .Z(n17883) );
  XOR U17506 ( .A(p_input[124]), .B(p_input[2060]), .Z(n17843) );
  XOR U17507 ( .A(n17853), .B(n17884), .Z(n17882) );
  IV U17508 ( .A(n17844), .Z(n17884) );
  XOR U17509 ( .A(p_input[113]), .B(p_input[2049]), .Z(n17844) );
  XNOR U17510 ( .A(n17885), .B(n17860), .Z(n17853) );
  XNOR U17511 ( .A(p_input[127]), .B(n16735), .Z(n17860) );
  XOR U17512 ( .A(n17850), .B(n17859), .Z(n17885) );
  XOR U17513 ( .A(n17886), .B(n17856), .Z(n17859) );
  XOR U17514 ( .A(p_input[125]), .B(p_input[2061]), .Z(n17856) );
  XOR U17515 ( .A(p_input[126]), .B(n16737), .Z(n17886) );
  XOR U17516 ( .A(p_input[121]), .B(p_input[2057]), .Z(n17850) );
  XOR U17517 ( .A(n17868), .B(n17866), .Z(n17848) );
  XNOR U17518 ( .A(n17887), .B(n17873), .Z(n17866) );
  XOR U17519 ( .A(p_input[120]), .B(p_input[2056]), .Z(n17873) );
  XOR U17520 ( .A(n17863), .B(n17872), .Z(n17887) );
  XOR U17521 ( .A(n17888), .B(n17869), .Z(n17872) );
  XOR U17522 ( .A(p_input[118]), .B(p_input[2054]), .Z(n17869) );
  XOR U17523 ( .A(p_input[119]), .B(n17722), .Z(n17888) );
  XOR U17524 ( .A(p_input[114]), .B(p_input[2050]), .Z(n17863) );
  XNOR U17525 ( .A(n17878), .B(n17877), .Z(n17868) );
  XOR U17526 ( .A(n17889), .B(n17874), .Z(n17877) );
  XOR U17527 ( .A(p_input[115]), .B(p_input[2051]), .Z(n17874) );
  XOR U17528 ( .A(p_input[116]), .B(n17724), .Z(n17889) );
  XOR U17529 ( .A(p_input[117]), .B(p_input[2053]), .Z(n17878) );
  XNOR U17530 ( .A(n17890), .B(n17891), .Z(n17783) );
  AND U17531 ( .A(n116), .B(n17892), .Z(n17891) );
  XNOR U17532 ( .A(n17893), .B(n17894), .Z(n116) );
  AND U17533 ( .A(n17895), .B(n17896), .Z(n17894) );
  XOR U17534 ( .A(n17893), .B(n17793), .Z(n17896) );
  XNOR U17535 ( .A(n17893), .B(n17747), .Z(n17895) );
  XOR U17536 ( .A(n17897), .B(n17898), .Z(n17893) );
  AND U17537 ( .A(n17899), .B(n17900), .Z(n17898) );
  XOR U17538 ( .A(n17897), .B(n17757), .Z(n17899) );
  XOR U17539 ( .A(n17901), .B(n17902), .Z(n17736) );
  AND U17540 ( .A(n120), .B(n17892), .Z(n17902) );
  XNOR U17541 ( .A(n17890), .B(n17901), .Z(n17892) );
  XNOR U17542 ( .A(n17903), .B(n17904), .Z(n120) );
  AND U17543 ( .A(n17905), .B(n17906), .Z(n17904) );
  XNOR U17544 ( .A(n17907), .B(n17903), .Z(n17906) );
  IV U17545 ( .A(n17793), .Z(n17907) );
  XNOR U17546 ( .A(n17908), .B(n17909), .Z(n17793) );
  AND U17547 ( .A(n123), .B(n17910), .Z(n17909) );
  XNOR U17548 ( .A(n17908), .B(n17911), .Z(n17910) );
  XNOR U17549 ( .A(n17747), .B(n17903), .Z(n17905) );
  XOR U17550 ( .A(n17912), .B(n17913), .Z(n17747) );
  AND U17551 ( .A(n131), .B(n17914), .Z(n17913) );
  XOR U17552 ( .A(n17897), .B(n17915), .Z(n17903) );
  AND U17553 ( .A(n17916), .B(n17900), .Z(n17915) );
  XNOR U17554 ( .A(n17806), .B(n17897), .Z(n17900) );
  XNOR U17555 ( .A(n17917), .B(n17918), .Z(n17806) );
  AND U17556 ( .A(n123), .B(n17919), .Z(n17918) );
  XOR U17557 ( .A(n17920), .B(n17917), .Z(n17919) );
  XNOR U17558 ( .A(n17921), .B(n17897), .Z(n17916) );
  IV U17559 ( .A(n17757), .Z(n17921) );
  XOR U17560 ( .A(n17922), .B(n17923), .Z(n17757) );
  AND U17561 ( .A(n131), .B(n17924), .Z(n17923) );
  XOR U17562 ( .A(n17925), .B(n17926), .Z(n17897) );
  AND U17563 ( .A(n17927), .B(n17928), .Z(n17926) );
  XNOR U17564 ( .A(n17831), .B(n17925), .Z(n17928) );
  XNOR U17565 ( .A(n17929), .B(n17930), .Z(n17831) );
  AND U17566 ( .A(n123), .B(n17931), .Z(n17930) );
  XNOR U17567 ( .A(n17932), .B(n17929), .Z(n17931) );
  XOR U17568 ( .A(n17925), .B(n17768), .Z(n17927) );
  XOR U17569 ( .A(n17933), .B(n17934), .Z(n17768) );
  AND U17570 ( .A(n131), .B(n17935), .Z(n17934) );
  XOR U17571 ( .A(n17936), .B(n17937), .Z(n17925) );
  AND U17572 ( .A(n17938), .B(n17939), .Z(n17937) );
  XNOR U17573 ( .A(n17936), .B(n17879), .Z(n17939) );
  XNOR U17574 ( .A(n17940), .B(n17941), .Z(n17879) );
  AND U17575 ( .A(n123), .B(n17942), .Z(n17941) );
  XOR U17576 ( .A(n17943), .B(n17940), .Z(n17942) );
  XNOR U17577 ( .A(n17944), .B(n17936), .Z(n17938) );
  IV U17578 ( .A(n17780), .Z(n17944) );
  XOR U17579 ( .A(n17945), .B(n17946), .Z(n17780) );
  AND U17580 ( .A(n131), .B(n17947), .Z(n17946) );
  AND U17581 ( .A(n17901), .B(n17890), .Z(n17936) );
  XNOR U17582 ( .A(n17948), .B(n17949), .Z(n17890) );
  AND U17583 ( .A(n123), .B(n17950), .Z(n17949) );
  XNOR U17584 ( .A(n17951), .B(n17948), .Z(n17950) );
  XNOR U17585 ( .A(n17952), .B(n17953), .Z(n123) );
  AND U17586 ( .A(n17954), .B(n17955), .Z(n17953) );
  XOR U17587 ( .A(n17911), .B(n17952), .Z(n17955) );
  AND U17588 ( .A(n17956), .B(n17957), .Z(n17911) );
  XOR U17589 ( .A(n17952), .B(n17908), .Z(n17954) );
  XNOR U17590 ( .A(n17958), .B(n17959), .Z(n17908) );
  AND U17591 ( .A(n127), .B(n17914), .Z(n17959) );
  XOR U17592 ( .A(n17912), .B(n17958), .Z(n17914) );
  XOR U17593 ( .A(n17960), .B(n17961), .Z(n17952) );
  AND U17594 ( .A(n17962), .B(n17963), .Z(n17961) );
  XNOR U17595 ( .A(n17960), .B(n17956), .Z(n17963) );
  IV U17596 ( .A(n17920), .Z(n17956) );
  XOR U17597 ( .A(n17964), .B(n17965), .Z(n17920) );
  XOR U17598 ( .A(n17966), .B(n17957), .Z(n17965) );
  AND U17599 ( .A(n17932), .B(n17967), .Z(n17957) );
  AND U17600 ( .A(n17968), .B(n17969), .Z(n17966) );
  XOR U17601 ( .A(n17970), .B(n17964), .Z(n17968) );
  XNOR U17602 ( .A(n17917), .B(n17960), .Z(n17962) );
  XNOR U17603 ( .A(n17971), .B(n17972), .Z(n17917) );
  AND U17604 ( .A(n127), .B(n17924), .Z(n17972) );
  XOR U17605 ( .A(n17971), .B(n17922), .Z(n17924) );
  XOR U17606 ( .A(n17973), .B(n17974), .Z(n17960) );
  AND U17607 ( .A(n17975), .B(n17976), .Z(n17974) );
  XNOR U17608 ( .A(n17973), .B(n17932), .Z(n17976) );
  XOR U17609 ( .A(n17977), .B(n17969), .Z(n17932) );
  XNOR U17610 ( .A(n17978), .B(n17964), .Z(n17969) );
  XOR U17611 ( .A(n17979), .B(n17980), .Z(n17964) );
  AND U17612 ( .A(n17981), .B(n17982), .Z(n17980) );
  XOR U17613 ( .A(n17983), .B(n17979), .Z(n17981) );
  XNOR U17614 ( .A(n17984), .B(n17985), .Z(n17978) );
  AND U17615 ( .A(n17986), .B(n17987), .Z(n17985) );
  XOR U17616 ( .A(n17984), .B(n17988), .Z(n17986) );
  XNOR U17617 ( .A(n17970), .B(n17967), .Z(n17977) );
  AND U17618 ( .A(n17989), .B(n17990), .Z(n17967) );
  XOR U17619 ( .A(n17991), .B(n17992), .Z(n17970) );
  AND U17620 ( .A(n17993), .B(n17994), .Z(n17992) );
  XOR U17621 ( .A(n17991), .B(n17995), .Z(n17993) );
  XNOR U17622 ( .A(n17929), .B(n17973), .Z(n17975) );
  XNOR U17623 ( .A(n17996), .B(n17997), .Z(n17929) );
  AND U17624 ( .A(n127), .B(n17935), .Z(n17997) );
  XOR U17625 ( .A(n17996), .B(n17933), .Z(n17935) );
  XOR U17626 ( .A(n17998), .B(n17999), .Z(n17973) );
  AND U17627 ( .A(n18000), .B(n18001), .Z(n17999) );
  XNOR U17628 ( .A(n17998), .B(n17989), .Z(n18001) );
  IV U17629 ( .A(n17943), .Z(n17989) );
  XNOR U17630 ( .A(n18002), .B(n17982), .Z(n17943) );
  XNOR U17631 ( .A(n18003), .B(n17988), .Z(n17982) );
  XNOR U17632 ( .A(n18004), .B(n18005), .Z(n17988) );
  NOR U17633 ( .A(n18006), .B(n18007), .Z(n18005) );
  XOR U17634 ( .A(n18004), .B(n18008), .Z(n18006) );
  XNOR U17635 ( .A(n17987), .B(n17979), .Z(n18003) );
  XOR U17636 ( .A(n18009), .B(n18010), .Z(n17979) );
  AND U17637 ( .A(n18011), .B(n18012), .Z(n18010) );
  XOR U17638 ( .A(n18009), .B(n18013), .Z(n18011) );
  XNOR U17639 ( .A(n18014), .B(n17984), .Z(n17987) );
  XOR U17640 ( .A(n18015), .B(n18016), .Z(n17984) );
  AND U17641 ( .A(n18017), .B(n18018), .Z(n18016) );
  XNOR U17642 ( .A(n18019), .B(n18020), .Z(n18017) );
  IV U17643 ( .A(n18015), .Z(n18019) );
  XNOR U17644 ( .A(n18021), .B(n18022), .Z(n18014) );
  NOR U17645 ( .A(n18023), .B(n18024), .Z(n18022) );
  XNOR U17646 ( .A(n18021), .B(n18025), .Z(n18023) );
  XNOR U17647 ( .A(n17983), .B(n17990), .Z(n18002) );
  NOR U17648 ( .A(n17951), .B(n18026), .Z(n17990) );
  XOR U17649 ( .A(n17995), .B(n17994), .Z(n17983) );
  XNOR U17650 ( .A(n18027), .B(n17991), .Z(n17994) );
  XOR U17651 ( .A(n18028), .B(n18029), .Z(n17991) );
  AND U17652 ( .A(n18030), .B(n18031), .Z(n18029) );
  XNOR U17653 ( .A(n18032), .B(n18033), .Z(n18030) );
  IV U17654 ( .A(n18028), .Z(n18032) );
  XNOR U17655 ( .A(n18034), .B(n18035), .Z(n18027) );
  NOR U17656 ( .A(n18036), .B(n18037), .Z(n18035) );
  XNOR U17657 ( .A(n18034), .B(n18038), .Z(n18036) );
  XOR U17658 ( .A(n18039), .B(n18040), .Z(n17995) );
  NOR U17659 ( .A(n18041), .B(n18042), .Z(n18040) );
  XNOR U17660 ( .A(n18039), .B(n18043), .Z(n18041) );
  XNOR U17661 ( .A(n17940), .B(n17998), .Z(n18000) );
  XNOR U17662 ( .A(n18044), .B(n18045), .Z(n17940) );
  AND U17663 ( .A(n127), .B(n17947), .Z(n18045) );
  XOR U17664 ( .A(n18044), .B(n17945), .Z(n17947) );
  AND U17665 ( .A(n17948), .B(n17951), .Z(n17998) );
  XOR U17666 ( .A(n18046), .B(n18026), .Z(n17951) );
  XNOR U17667 ( .A(p_input[128]), .B(p_input[2048]), .Z(n18026) );
  XNOR U17668 ( .A(n18013), .B(n18012), .Z(n18046) );
  XNOR U17669 ( .A(n18047), .B(n18020), .Z(n18012) );
  XNOR U17670 ( .A(n18008), .B(n18007), .Z(n18020) );
  XNOR U17671 ( .A(n18048), .B(n18004), .Z(n18007) );
  XNOR U17672 ( .A(p_input[138]), .B(p_input[2058]), .Z(n18004) );
  XOR U17673 ( .A(p_input[139]), .B(n16732), .Z(n18048) );
  XOR U17674 ( .A(p_input[140]), .B(p_input[2060]), .Z(n18008) );
  XOR U17675 ( .A(n18018), .B(n18049), .Z(n18047) );
  IV U17676 ( .A(n18009), .Z(n18049) );
  XOR U17677 ( .A(p_input[129]), .B(p_input[2049]), .Z(n18009) );
  XNOR U17678 ( .A(n18050), .B(n18025), .Z(n18018) );
  XNOR U17679 ( .A(p_input[143]), .B(n16735), .Z(n18025) );
  XOR U17680 ( .A(n18015), .B(n18024), .Z(n18050) );
  XOR U17681 ( .A(n18051), .B(n18021), .Z(n18024) );
  XOR U17682 ( .A(p_input[141]), .B(p_input[2061]), .Z(n18021) );
  XOR U17683 ( .A(p_input[142]), .B(n16737), .Z(n18051) );
  XOR U17684 ( .A(p_input[137]), .B(p_input[2057]), .Z(n18015) );
  XOR U17685 ( .A(n18033), .B(n18031), .Z(n18013) );
  XNOR U17686 ( .A(n18052), .B(n18038), .Z(n18031) );
  XOR U17687 ( .A(p_input[136]), .B(p_input[2056]), .Z(n18038) );
  XOR U17688 ( .A(n18028), .B(n18037), .Z(n18052) );
  XOR U17689 ( .A(n18053), .B(n18034), .Z(n18037) );
  XOR U17690 ( .A(p_input[134]), .B(p_input[2054]), .Z(n18034) );
  XOR U17691 ( .A(p_input[135]), .B(n17722), .Z(n18053) );
  XOR U17692 ( .A(p_input[130]), .B(p_input[2050]), .Z(n18028) );
  XNOR U17693 ( .A(n18043), .B(n18042), .Z(n18033) );
  XOR U17694 ( .A(n18054), .B(n18039), .Z(n18042) );
  XOR U17695 ( .A(p_input[131]), .B(p_input[2051]), .Z(n18039) );
  XOR U17696 ( .A(p_input[132]), .B(n17724), .Z(n18054) );
  XOR U17697 ( .A(p_input[133]), .B(p_input[2053]), .Z(n18043) );
  XNOR U17698 ( .A(n18055), .B(n18056), .Z(n17948) );
  AND U17699 ( .A(n127), .B(n18057), .Z(n18056) );
  XNOR U17700 ( .A(n18058), .B(n18059), .Z(n127) );
  AND U17701 ( .A(n18060), .B(n18061), .Z(n18059) );
  XOR U17702 ( .A(n18058), .B(n17958), .Z(n18061) );
  XNOR U17703 ( .A(n18058), .B(n17912), .Z(n18060) );
  XOR U17704 ( .A(n18062), .B(n18063), .Z(n18058) );
  AND U17705 ( .A(n18064), .B(n18065), .Z(n18063) );
  XOR U17706 ( .A(n18062), .B(n17922), .Z(n18064) );
  XOR U17707 ( .A(n18066), .B(n18067), .Z(n17901) );
  AND U17708 ( .A(n131), .B(n18057), .Z(n18067) );
  XNOR U17709 ( .A(n18055), .B(n18066), .Z(n18057) );
  XNOR U17710 ( .A(n18068), .B(n18069), .Z(n131) );
  AND U17711 ( .A(n18070), .B(n18071), .Z(n18069) );
  XNOR U17712 ( .A(n18072), .B(n18068), .Z(n18071) );
  IV U17713 ( .A(n17958), .Z(n18072) );
  XNOR U17714 ( .A(n18073), .B(n18074), .Z(n17958) );
  AND U17715 ( .A(n134), .B(n18075), .Z(n18074) );
  XNOR U17716 ( .A(n18073), .B(n18076), .Z(n18075) );
  XNOR U17717 ( .A(n17912), .B(n18068), .Z(n18070) );
  XOR U17718 ( .A(n18077), .B(n18078), .Z(n17912) );
  AND U17719 ( .A(n142), .B(n18079), .Z(n18078) );
  XOR U17720 ( .A(n18062), .B(n18080), .Z(n18068) );
  AND U17721 ( .A(n18081), .B(n18065), .Z(n18080) );
  XNOR U17722 ( .A(n17971), .B(n18062), .Z(n18065) );
  XNOR U17723 ( .A(n18082), .B(n18083), .Z(n17971) );
  AND U17724 ( .A(n134), .B(n18084), .Z(n18083) );
  XOR U17725 ( .A(n18085), .B(n18082), .Z(n18084) );
  XNOR U17726 ( .A(n18086), .B(n18062), .Z(n18081) );
  IV U17727 ( .A(n17922), .Z(n18086) );
  XOR U17728 ( .A(n18087), .B(n18088), .Z(n17922) );
  AND U17729 ( .A(n142), .B(n18089), .Z(n18088) );
  XOR U17730 ( .A(n18090), .B(n18091), .Z(n18062) );
  AND U17731 ( .A(n18092), .B(n18093), .Z(n18091) );
  XNOR U17732 ( .A(n17996), .B(n18090), .Z(n18093) );
  XNOR U17733 ( .A(n18094), .B(n18095), .Z(n17996) );
  AND U17734 ( .A(n134), .B(n18096), .Z(n18095) );
  XNOR U17735 ( .A(n18097), .B(n18094), .Z(n18096) );
  XOR U17736 ( .A(n18090), .B(n17933), .Z(n18092) );
  XOR U17737 ( .A(n18098), .B(n18099), .Z(n17933) );
  AND U17738 ( .A(n142), .B(n18100), .Z(n18099) );
  XOR U17739 ( .A(n18101), .B(n18102), .Z(n18090) );
  AND U17740 ( .A(n18103), .B(n18104), .Z(n18102) );
  XNOR U17741 ( .A(n18101), .B(n18044), .Z(n18104) );
  XNOR U17742 ( .A(n18105), .B(n18106), .Z(n18044) );
  AND U17743 ( .A(n134), .B(n18107), .Z(n18106) );
  XOR U17744 ( .A(n18108), .B(n18105), .Z(n18107) );
  XNOR U17745 ( .A(n18109), .B(n18101), .Z(n18103) );
  IV U17746 ( .A(n17945), .Z(n18109) );
  XOR U17747 ( .A(n18110), .B(n18111), .Z(n17945) );
  AND U17748 ( .A(n142), .B(n18112), .Z(n18111) );
  AND U17749 ( .A(n18066), .B(n18055), .Z(n18101) );
  XNOR U17750 ( .A(n18113), .B(n18114), .Z(n18055) );
  AND U17751 ( .A(n134), .B(n18115), .Z(n18114) );
  XNOR U17752 ( .A(n18116), .B(n18113), .Z(n18115) );
  XNOR U17753 ( .A(n18117), .B(n18118), .Z(n134) );
  AND U17754 ( .A(n18119), .B(n18120), .Z(n18118) );
  XOR U17755 ( .A(n18076), .B(n18117), .Z(n18120) );
  AND U17756 ( .A(n18121), .B(n18122), .Z(n18076) );
  XOR U17757 ( .A(n18117), .B(n18073), .Z(n18119) );
  XNOR U17758 ( .A(n18123), .B(n18124), .Z(n18073) );
  AND U17759 ( .A(n138), .B(n18079), .Z(n18124) );
  XOR U17760 ( .A(n18077), .B(n18123), .Z(n18079) );
  XOR U17761 ( .A(n18125), .B(n18126), .Z(n18117) );
  AND U17762 ( .A(n18127), .B(n18128), .Z(n18126) );
  XNOR U17763 ( .A(n18125), .B(n18121), .Z(n18128) );
  IV U17764 ( .A(n18085), .Z(n18121) );
  XOR U17765 ( .A(n18129), .B(n18130), .Z(n18085) );
  XOR U17766 ( .A(n18131), .B(n18122), .Z(n18130) );
  AND U17767 ( .A(n18097), .B(n18132), .Z(n18122) );
  AND U17768 ( .A(n18133), .B(n18134), .Z(n18131) );
  XOR U17769 ( .A(n18135), .B(n18129), .Z(n18133) );
  XNOR U17770 ( .A(n18082), .B(n18125), .Z(n18127) );
  XNOR U17771 ( .A(n18136), .B(n18137), .Z(n18082) );
  AND U17772 ( .A(n138), .B(n18089), .Z(n18137) );
  XOR U17773 ( .A(n18136), .B(n18087), .Z(n18089) );
  XOR U17774 ( .A(n18138), .B(n18139), .Z(n18125) );
  AND U17775 ( .A(n18140), .B(n18141), .Z(n18139) );
  XNOR U17776 ( .A(n18138), .B(n18097), .Z(n18141) );
  XOR U17777 ( .A(n18142), .B(n18134), .Z(n18097) );
  XNOR U17778 ( .A(n18143), .B(n18129), .Z(n18134) );
  XOR U17779 ( .A(n18144), .B(n18145), .Z(n18129) );
  AND U17780 ( .A(n18146), .B(n18147), .Z(n18145) );
  XOR U17781 ( .A(n18148), .B(n18144), .Z(n18146) );
  XNOR U17782 ( .A(n18149), .B(n18150), .Z(n18143) );
  AND U17783 ( .A(n18151), .B(n18152), .Z(n18150) );
  XOR U17784 ( .A(n18149), .B(n18153), .Z(n18151) );
  XNOR U17785 ( .A(n18135), .B(n18132), .Z(n18142) );
  AND U17786 ( .A(n18154), .B(n18155), .Z(n18132) );
  XOR U17787 ( .A(n18156), .B(n18157), .Z(n18135) );
  AND U17788 ( .A(n18158), .B(n18159), .Z(n18157) );
  XOR U17789 ( .A(n18156), .B(n18160), .Z(n18158) );
  XNOR U17790 ( .A(n18094), .B(n18138), .Z(n18140) );
  XNOR U17791 ( .A(n18161), .B(n18162), .Z(n18094) );
  AND U17792 ( .A(n138), .B(n18100), .Z(n18162) );
  XOR U17793 ( .A(n18161), .B(n18098), .Z(n18100) );
  XOR U17794 ( .A(n18163), .B(n18164), .Z(n18138) );
  AND U17795 ( .A(n18165), .B(n18166), .Z(n18164) );
  XNOR U17796 ( .A(n18163), .B(n18154), .Z(n18166) );
  IV U17797 ( .A(n18108), .Z(n18154) );
  XNOR U17798 ( .A(n18167), .B(n18147), .Z(n18108) );
  XNOR U17799 ( .A(n18168), .B(n18153), .Z(n18147) );
  XNOR U17800 ( .A(n18169), .B(n18170), .Z(n18153) );
  NOR U17801 ( .A(n18171), .B(n18172), .Z(n18170) );
  XOR U17802 ( .A(n18169), .B(n18173), .Z(n18171) );
  XNOR U17803 ( .A(n18152), .B(n18144), .Z(n18168) );
  XOR U17804 ( .A(n18174), .B(n18175), .Z(n18144) );
  AND U17805 ( .A(n18176), .B(n18177), .Z(n18175) );
  XOR U17806 ( .A(n18174), .B(n18178), .Z(n18176) );
  XNOR U17807 ( .A(n18179), .B(n18149), .Z(n18152) );
  XOR U17808 ( .A(n18180), .B(n18181), .Z(n18149) );
  AND U17809 ( .A(n18182), .B(n18183), .Z(n18181) );
  XNOR U17810 ( .A(n18184), .B(n18185), .Z(n18182) );
  IV U17811 ( .A(n18180), .Z(n18184) );
  XNOR U17812 ( .A(n18186), .B(n18187), .Z(n18179) );
  NOR U17813 ( .A(n18188), .B(n18189), .Z(n18187) );
  XNOR U17814 ( .A(n18186), .B(n18190), .Z(n18188) );
  XNOR U17815 ( .A(n18148), .B(n18155), .Z(n18167) );
  NOR U17816 ( .A(n18116), .B(n18191), .Z(n18155) );
  XOR U17817 ( .A(n18160), .B(n18159), .Z(n18148) );
  XNOR U17818 ( .A(n18192), .B(n18156), .Z(n18159) );
  XOR U17819 ( .A(n18193), .B(n18194), .Z(n18156) );
  AND U17820 ( .A(n18195), .B(n18196), .Z(n18194) );
  XNOR U17821 ( .A(n18197), .B(n18198), .Z(n18195) );
  IV U17822 ( .A(n18193), .Z(n18197) );
  XNOR U17823 ( .A(n18199), .B(n18200), .Z(n18192) );
  NOR U17824 ( .A(n18201), .B(n18202), .Z(n18200) );
  XNOR U17825 ( .A(n18199), .B(n18203), .Z(n18201) );
  XOR U17826 ( .A(n18204), .B(n18205), .Z(n18160) );
  NOR U17827 ( .A(n18206), .B(n18207), .Z(n18205) );
  XNOR U17828 ( .A(n18204), .B(n18208), .Z(n18206) );
  XNOR U17829 ( .A(n18105), .B(n18163), .Z(n18165) );
  XNOR U17830 ( .A(n18209), .B(n18210), .Z(n18105) );
  AND U17831 ( .A(n138), .B(n18112), .Z(n18210) );
  XOR U17832 ( .A(n18209), .B(n18110), .Z(n18112) );
  AND U17833 ( .A(n18113), .B(n18116), .Z(n18163) );
  XOR U17834 ( .A(n18211), .B(n18191), .Z(n18116) );
  XNOR U17835 ( .A(p_input[144]), .B(p_input[2048]), .Z(n18191) );
  XNOR U17836 ( .A(n18178), .B(n18177), .Z(n18211) );
  XNOR U17837 ( .A(n18212), .B(n18185), .Z(n18177) );
  XNOR U17838 ( .A(n18173), .B(n18172), .Z(n18185) );
  XNOR U17839 ( .A(n18213), .B(n18169), .Z(n18172) );
  XNOR U17840 ( .A(p_input[154]), .B(p_input[2058]), .Z(n18169) );
  XOR U17841 ( .A(p_input[155]), .B(n16732), .Z(n18213) );
  XOR U17842 ( .A(p_input[156]), .B(p_input[2060]), .Z(n18173) );
  XOR U17843 ( .A(n18183), .B(n18214), .Z(n18212) );
  IV U17844 ( .A(n18174), .Z(n18214) );
  XOR U17845 ( .A(p_input[145]), .B(p_input[2049]), .Z(n18174) );
  XNOR U17846 ( .A(n18215), .B(n18190), .Z(n18183) );
  XNOR U17847 ( .A(p_input[159]), .B(n16735), .Z(n18190) );
  XOR U17848 ( .A(n18180), .B(n18189), .Z(n18215) );
  XOR U17849 ( .A(n18216), .B(n18186), .Z(n18189) );
  XOR U17850 ( .A(p_input[157]), .B(p_input[2061]), .Z(n18186) );
  XOR U17851 ( .A(p_input[158]), .B(n16737), .Z(n18216) );
  XOR U17852 ( .A(p_input[153]), .B(p_input[2057]), .Z(n18180) );
  XOR U17853 ( .A(n18198), .B(n18196), .Z(n18178) );
  XNOR U17854 ( .A(n18217), .B(n18203), .Z(n18196) );
  XOR U17855 ( .A(p_input[152]), .B(p_input[2056]), .Z(n18203) );
  XOR U17856 ( .A(n18193), .B(n18202), .Z(n18217) );
  XOR U17857 ( .A(n18218), .B(n18199), .Z(n18202) );
  XOR U17858 ( .A(p_input[150]), .B(p_input[2054]), .Z(n18199) );
  XOR U17859 ( .A(p_input[151]), .B(n17722), .Z(n18218) );
  XOR U17860 ( .A(p_input[146]), .B(p_input[2050]), .Z(n18193) );
  XNOR U17861 ( .A(n18208), .B(n18207), .Z(n18198) );
  XOR U17862 ( .A(n18219), .B(n18204), .Z(n18207) );
  XOR U17863 ( .A(p_input[147]), .B(p_input[2051]), .Z(n18204) );
  XOR U17864 ( .A(p_input[148]), .B(n17724), .Z(n18219) );
  XOR U17865 ( .A(p_input[149]), .B(p_input[2053]), .Z(n18208) );
  XNOR U17866 ( .A(n18220), .B(n18221), .Z(n18113) );
  AND U17867 ( .A(n138), .B(n18222), .Z(n18221) );
  XNOR U17868 ( .A(n18223), .B(n18224), .Z(n138) );
  AND U17869 ( .A(n18225), .B(n18226), .Z(n18224) );
  XOR U17870 ( .A(n18223), .B(n18123), .Z(n18226) );
  XNOR U17871 ( .A(n18223), .B(n18077), .Z(n18225) );
  XOR U17872 ( .A(n18227), .B(n18228), .Z(n18223) );
  AND U17873 ( .A(n18229), .B(n18230), .Z(n18228) );
  XOR U17874 ( .A(n18227), .B(n18087), .Z(n18229) );
  XOR U17875 ( .A(n18231), .B(n18232), .Z(n18066) );
  AND U17876 ( .A(n142), .B(n18222), .Z(n18232) );
  XNOR U17877 ( .A(n18220), .B(n18231), .Z(n18222) );
  XNOR U17878 ( .A(n18233), .B(n18234), .Z(n142) );
  AND U17879 ( .A(n18235), .B(n18236), .Z(n18234) );
  XNOR U17880 ( .A(n18237), .B(n18233), .Z(n18236) );
  IV U17881 ( .A(n18123), .Z(n18237) );
  XNOR U17882 ( .A(n18238), .B(n18239), .Z(n18123) );
  AND U17883 ( .A(n145), .B(n18240), .Z(n18239) );
  XNOR U17884 ( .A(n18238), .B(n18241), .Z(n18240) );
  XNOR U17885 ( .A(n18077), .B(n18233), .Z(n18235) );
  XOR U17886 ( .A(n18242), .B(n18243), .Z(n18077) );
  AND U17887 ( .A(n153), .B(n18244), .Z(n18243) );
  XOR U17888 ( .A(n18227), .B(n18245), .Z(n18233) );
  AND U17889 ( .A(n18246), .B(n18230), .Z(n18245) );
  XNOR U17890 ( .A(n18136), .B(n18227), .Z(n18230) );
  XNOR U17891 ( .A(n18247), .B(n18248), .Z(n18136) );
  AND U17892 ( .A(n145), .B(n18249), .Z(n18248) );
  XOR U17893 ( .A(n18250), .B(n18247), .Z(n18249) );
  XNOR U17894 ( .A(n18251), .B(n18227), .Z(n18246) );
  IV U17895 ( .A(n18087), .Z(n18251) );
  XOR U17896 ( .A(n18252), .B(n18253), .Z(n18087) );
  AND U17897 ( .A(n153), .B(n18254), .Z(n18253) );
  XOR U17898 ( .A(n18255), .B(n18256), .Z(n18227) );
  AND U17899 ( .A(n18257), .B(n18258), .Z(n18256) );
  XNOR U17900 ( .A(n18161), .B(n18255), .Z(n18258) );
  XNOR U17901 ( .A(n18259), .B(n18260), .Z(n18161) );
  AND U17902 ( .A(n145), .B(n18261), .Z(n18260) );
  XNOR U17903 ( .A(n18262), .B(n18259), .Z(n18261) );
  XOR U17904 ( .A(n18255), .B(n18098), .Z(n18257) );
  XOR U17905 ( .A(n18263), .B(n18264), .Z(n18098) );
  AND U17906 ( .A(n153), .B(n18265), .Z(n18264) );
  XOR U17907 ( .A(n18266), .B(n18267), .Z(n18255) );
  AND U17908 ( .A(n18268), .B(n18269), .Z(n18267) );
  XNOR U17909 ( .A(n18266), .B(n18209), .Z(n18269) );
  XNOR U17910 ( .A(n18270), .B(n18271), .Z(n18209) );
  AND U17911 ( .A(n145), .B(n18272), .Z(n18271) );
  XOR U17912 ( .A(n18273), .B(n18270), .Z(n18272) );
  XNOR U17913 ( .A(n18274), .B(n18266), .Z(n18268) );
  IV U17914 ( .A(n18110), .Z(n18274) );
  XOR U17915 ( .A(n18275), .B(n18276), .Z(n18110) );
  AND U17916 ( .A(n153), .B(n18277), .Z(n18276) );
  AND U17917 ( .A(n18231), .B(n18220), .Z(n18266) );
  XNOR U17918 ( .A(n18278), .B(n18279), .Z(n18220) );
  AND U17919 ( .A(n145), .B(n18280), .Z(n18279) );
  XNOR U17920 ( .A(n18281), .B(n18278), .Z(n18280) );
  XNOR U17921 ( .A(n18282), .B(n18283), .Z(n145) );
  AND U17922 ( .A(n18284), .B(n18285), .Z(n18283) );
  XOR U17923 ( .A(n18241), .B(n18282), .Z(n18285) );
  AND U17924 ( .A(n18286), .B(n18287), .Z(n18241) );
  XOR U17925 ( .A(n18282), .B(n18238), .Z(n18284) );
  XNOR U17926 ( .A(n18288), .B(n18289), .Z(n18238) );
  AND U17927 ( .A(n149), .B(n18244), .Z(n18289) );
  XOR U17928 ( .A(n18242), .B(n18288), .Z(n18244) );
  XOR U17929 ( .A(n18290), .B(n18291), .Z(n18282) );
  AND U17930 ( .A(n18292), .B(n18293), .Z(n18291) );
  XNOR U17931 ( .A(n18290), .B(n18286), .Z(n18293) );
  IV U17932 ( .A(n18250), .Z(n18286) );
  XOR U17933 ( .A(n18294), .B(n18295), .Z(n18250) );
  XOR U17934 ( .A(n18296), .B(n18287), .Z(n18295) );
  AND U17935 ( .A(n18262), .B(n18297), .Z(n18287) );
  AND U17936 ( .A(n18298), .B(n18299), .Z(n18296) );
  XOR U17937 ( .A(n18300), .B(n18294), .Z(n18298) );
  XNOR U17938 ( .A(n18247), .B(n18290), .Z(n18292) );
  XNOR U17939 ( .A(n18301), .B(n18302), .Z(n18247) );
  AND U17940 ( .A(n149), .B(n18254), .Z(n18302) );
  XOR U17941 ( .A(n18301), .B(n18252), .Z(n18254) );
  XOR U17942 ( .A(n18303), .B(n18304), .Z(n18290) );
  AND U17943 ( .A(n18305), .B(n18306), .Z(n18304) );
  XNOR U17944 ( .A(n18303), .B(n18262), .Z(n18306) );
  XOR U17945 ( .A(n18307), .B(n18299), .Z(n18262) );
  XNOR U17946 ( .A(n18308), .B(n18294), .Z(n18299) );
  XOR U17947 ( .A(n18309), .B(n18310), .Z(n18294) );
  AND U17948 ( .A(n18311), .B(n18312), .Z(n18310) );
  XOR U17949 ( .A(n18313), .B(n18309), .Z(n18311) );
  XNOR U17950 ( .A(n18314), .B(n18315), .Z(n18308) );
  AND U17951 ( .A(n18316), .B(n18317), .Z(n18315) );
  XOR U17952 ( .A(n18314), .B(n18318), .Z(n18316) );
  XNOR U17953 ( .A(n18300), .B(n18297), .Z(n18307) );
  AND U17954 ( .A(n18319), .B(n18320), .Z(n18297) );
  XOR U17955 ( .A(n18321), .B(n18322), .Z(n18300) );
  AND U17956 ( .A(n18323), .B(n18324), .Z(n18322) );
  XOR U17957 ( .A(n18321), .B(n18325), .Z(n18323) );
  XNOR U17958 ( .A(n18259), .B(n18303), .Z(n18305) );
  XNOR U17959 ( .A(n18326), .B(n18327), .Z(n18259) );
  AND U17960 ( .A(n149), .B(n18265), .Z(n18327) );
  XOR U17961 ( .A(n18326), .B(n18263), .Z(n18265) );
  XOR U17962 ( .A(n18328), .B(n18329), .Z(n18303) );
  AND U17963 ( .A(n18330), .B(n18331), .Z(n18329) );
  XNOR U17964 ( .A(n18328), .B(n18319), .Z(n18331) );
  IV U17965 ( .A(n18273), .Z(n18319) );
  XNOR U17966 ( .A(n18332), .B(n18312), .Z(n18273) );
  XNOR U17967 ( .A(n18333), .B(n18318), .Z(n18312) );
  XNOR U17968 ( .A(n18334), .B(n18335), .Z(n18318) );
  NOR U17969 ( .A(n18336), .B(n18337), .Z(n18335) );
  XOR U17970 ( .A(n18334), .B(n18338), .Z(n18336) );
  XNOR U17971 ( .A(n18317), .B(n18309), .Z(n18333) );
  XOR U17972 ( .A(n18339), .B(n18340), .Z(n18309) );
  AND U17973 ( .A(n18341), .B(n18342), .Z(n18340) );
  XOR U17974 ( .A(n18339), .B(n18343), .Z(n18341) );
  XNOR U17975 ( .A(n18344), .B(n18314), .Z(n18317) );
  XOR U17976 ( .A(n18345), .B(n18346), .Z(n18314) );
  AND U17977 ( .A(n18347), .B(n18348), .Z(n18346) );
  XNOR U17978 ( .A(n18349), .B(n18350), .Z(n18347) );
  IV U17979 ( .A(n18345), .Z(n18349) );
  XNOR U17980 ( .A(n18351), .B(n18352), .Z(n18344) );
  NOR U17981 ( .A(n18353), .B(n18354), .Z(n18352) );
  XNOR U17982 ( .A(n18351), .B(n18355), .Z(n18353) );
  XNOR U17983 ( .A(n18313), .B(n18320), .Z(n18332) );
  NOR U17984 ( .A(n18281), .B(n18356), .Z(n18320) );
  XOR U17985 ( .A(n18325), .B(n18324), .Z(n18313) );
  XNOR U17986 ( .A(n18357), .B(n18321), .Z(n18324) );
  XOR U17987 ( .A(n18358), .B(n18359), .Z(n18321) );
  AND U17988 ( .A(n18360), .B(n18361), .Z(n18359) );
  XNOR U17989 ( .A(n18362), .B(n18363), .Z(n18360) );
  IV U17990 ( .A(n18358), .Z(n18362) );
  XNOR U17991 ( .A(n18364), .B(n18365), .Z(n18357) );
  NOR U17992 ( .A(n18366), .B(n18367), .Z(n18365) );
  XNOR U17993 ( .A(n18364), .B(n18368), .Z(n18366) );
  XOR U17994 ( .A(n18369), .B(n18370), .Z(n18325) );
  NOR U17995 ( .A(n18371), .B(n18372), .Z(n18370) );
  XNOR U17996 ( .A(n18369), .B(n18373), .Z(n18371) );
  XNOR U17997 ( .A(n18270), .B(n18328), .Z(n18330) );
  XNOR U17998 ( .A(n18374), .B(n18375), .Z(n18270) );
  AND U17999 ( .A(n149), .B(n18277), .Z(n18375) );
  XOR U18000 ( .A(n18374), .B(n18275), .Z(n18277) );
  AND U18001 ( .A(n18278), .B(n18281), .Z(n18328) );
  XOR U18002 ( .A(n18376), .B(n18356), .Z(n18281) );
  XNOR U18003 ( .A(p_input[160]), .B(p_input[2048]), .Z(n18356) );
  XNOR U18004 ( .A(n18343), .B(n18342), .Z(n18376) );
  XNOR U18005 ( .A(n18377), .B(n18350), .Z(n18342) );
  XNOR U18006 ( .A(n18338), .B(n18337), .Z(n18350) );
  XNOR U18007 ( .A(n18378), .B(n18334), .Z(n18337) );
  XNOR U18008 ( .A(p_input[170]), .B(p_input[2058]), .Z(n18334) );
  XOR U18009 ( .A(p_input[171]), .B(n16732), .Z(n18378) );
  XOR U18010 ( .A(p_input[172]), .B(p_input[2060]), .Z(n18338) );
  XOR U18011 ( .A(n18348), .B(n18379), .Z(n18377) );
  IV U18012 ( .A(n18339), .Z(n18379) );
  XOR U18013 ( .A(p_input[161]), .B(p_input[2049]), .Z(n18339) );
  XNOR U18014 ( .A(n18380), .B(n18355), .Z(n18348) );
  XNOR U18015 ( .A(p_input[175]), .B(n16735), .Z(n18355) );
  XOR U18016 ( .A(n18345), .B(n18354), .Z(n18380) );
  XOR U18017 ( .A(n18381), .B(n18351), .Z(n18354) );
  XOR U18018 ( .A(p_input[173]), .B(p_input[2061]), .Z(n18351) );
  XOR U18019 ( .A(p_input[174]), .B(n16737), .Z(n18381) );
  XOR U18020 ( .A(p_input[169]), .B(p_input[2057]), .Z(n18345) );
  XOR U18021 ( .A(n18363), .B(n18361), .Z(n18343) );
  XNOR U18022 ( .A(n18382), .B(n18368), .Z(n18361) );
  XOR U18023 ( .A(p_input[168]), .B(p_input[2056]), .Z(n18368) );
  XOR U18024 ( .A(n18358), .B(n18367), .Z(n18382) );
  XOR U18025 ( .A(n18383), .B(n18364), .Z(n18367) );
  XOR U18026 ( .A(p_input[166]), .B(p_input[2054]), .Z(n18364) );
  XOR U18027 ( .A(p_input[167]), .B(n17722), .Z(n18383) );
  XOR U18028 ( .A(p_input[162]), .B(p_input[2050]), .Z(n18358) );
  XNOR U18029 ( .A(n18373), .B(n18372), .Z(n18363) );
  XOR U18030 ( .A(n18384), .B(n18369), .Z(n18372) );
  XOR U18031 ( .A(p_input[163]), .B(p_input[2051]), .Z(n18369) );
  XOR U18032 ( .A(p_input[164]), .B(n17724), .Z(n18384) );
  XOR U18033 ( .A(p_input[165]), .B(p_input[2053]), .Z(n18373) );
  XNOR U18034 ( .A(n18385), .B(n18386), .Z(n18278) );
  AND U18035 ( .A(n149), .B(n18387), .Z(n18386) );
  XNOR U18036 ( .A(n18388), .B(n18389), .Z(n149) );
  AND U18037 ( .A(n18390), .B(n18391), .Z(n18389) );
  XOR U18038 ( .A(n18388), .B(n18288), .Z(n18391) );
  XNOR U18039 ( .A(n18388), .B(n18242), .Z(n18390) );
  XOR U18040 ( .A(n18392), .B(n18393), .Z(n18388) );
  AND U18041 ( .A(n18394), .B(n18395), .Z(n18393) );
  XOR U18042 ( .A(n18392), .B(n18252), .Z(n18394) );
  XOR U18043 ( .A(n18396), .B(n18397), .Z(n18231) );
  AND U18044 ( .A(n153), .B(n18387), .Z(n18397) );
  XNOR U18045 ( .A(n18385), .B(n18396), .Z(n18387) );
  XNOR U18046 ( .A(n18398), .B(n18399), .Z(n153) );
  AND U18047 ( .A(n18400), .B(n18401), .Z(n18399) );
  XNOR U18048 ( .A(n18402), .B(n18398), .Z(n18401) );
  IV U18049 ( .A(n18288), .Z(n18402) );
  XNOR U18050 ( .A(n18403), .B(n18404), .Z(n18288) );
  AND U18051 ( .A(n156), .B(n18405), .Z(n18404) );
  XNOR U18052 ( .A(n18403), .B(n18406), .Z(n18405) );
  XNOR U18053 ( .A(n18242), .B(n18398), .Z(n18400) );
  XOR U18054 ( .A(n18407), .B(n18408), .Z(n18242) );
  AND U18055 ( .A(n164), .B(n18409), .Z(n18408) );
  XOR U18056 ( .A(n18392), .B(n18410), .Z(n18398) );
  AND U18057 ( .A(n18411), .B(n18395), .Z(n18410) );
  XNOR U18058 ( .A(n18301), .B(n18392), .Z(n18395) );
  XNOR U18059 ( .A(n18412), .B(n18413), .Z(n18301) );
  AND U18060 ( .A(n156), .B(n18414), .Z(n18413) );
  XOR U18061 ( .A(n18415), .B(n18412), .Z(n18414) );
  XNOR U18062 ( .A(n18416), .B(n18392), .Z(n18411) );
  IV U18063 ( .A(n18252), .Z(n18416) );
  XOR U18064 ( .A(n18417), .B(n18418), .Z(n18252) );
  AND U18065 ( .A(n164), .B(n18419), .Z(n18418) );
  XOR U18066 ( .A(n18420), .B(n18421), .Z(n18392) );
  AND U18067 ( .A(n18422), .B(n18423), .Z(n18421) );
  XNOR U18068 ( .A(n18326), .B(n18420), .Z(n18423) );
  XNOR U18069 ( .A(n18424), .B(n18425), .Z(n18326) );
  AND U18070 ( .A(n156), .B(n18426), .Z(n18425) );
  XNOR U18071 ( .A(n18427), .B(n18424), .Z(n18426) );
  XOR U18072 ( .A(n18420), .B(n18263), .Z(n18422) );
  XOR U18073 ( .A(n18428), .B(n18429), .Z(n18263) );
  AND U18074 ( .A(n164), .B(n18430), .Z(n18429) );
  XOR U18075 ( .A(n18431), .B(n18432), .Z(n18420) );
  AND U18076 ( .A(n18433), .B(n18434), .Z(n18432) );
  XNOR U18077 ( .A(n18431), .B(n18374), .Z(n18434) );
  XNOR U18078 ( .A(n18435), .B(n18436), .Z(n18374) );
  AND U18079 ( .A(n156), .B(n18437), .Z(n18436) );
  XOR U18080 ( .A(n18438), .B(n18435), .Z(n18437) );
  XNOR U18081 ( .A(n18439), .B(n18431), .Z(n18433) );
  IV U18082 ( .A(n18275), .Z(n18439) );
  XOR U18083 ( .A(n18440), .B(n18441), .Z(n18275) );
  AND U18084 ( .A(n164), .B(n18442), .Z(n18441) );
  AND U18085 ( .A(n18396), .B(n18385), .Z(n18431) );
  XNOR U18086 ( .A(n18443), .B(n18444), .Z(n18385) );
  AND U18087 ( .A(n156), .B(n18445), .Z(n18444) );
  XNOR U18088 ( .A(n18446), .B(n18443), .Z(n18445) );
  XNOR U18089 ( .A(n18447), .B(n18448), .Z(n156) );
  AND U18090 ( .A(n18449), .B(n18450), .Z(n18448) );
  XOR U18091 ( .A(n18406), .B(n18447), .Z(n18450) );
  AND U18092 ( .A(n18451), .B(n18452), .Z(n18406) );
  XOR U18093 ( .A(n18447), .B(n18403), .Z(n18449) );
  XNOR U18094 ( .A(n18453), .B(n18454), .Z(n18403) );
  AND U18095 ( .A(n160), .B(n18409), .Z(n18454) );
  XOR U18096 ( .A(n18407), .B(n18453), .Z(n18409) );
  XOR U18097 ( .A(n18455), .B(n18456), .Z(n18447) );
  AND U18098 ( .A(n18457), .B(n18458), .Z(n18456) );
  XNOR U18099 ( .A(n18455), .B(n18451), .Z(n18458) );
  IV U18100 ( .A(n18415), .Z(n18451) );
  XOR U18101 ( .A(n18459), .B(n18460), .Z(n18415) );
  XOR U18102 ( .A(n18461), .B(n18452), .Z(n18460) );
  AND U18103 ( .A(n18427), .B(n18462), .Z(n18452) );
  AND U18104 ( .A(n18463), .B(n18464), .Z(n18461) );
  XOR U18105 ( .A(n18465), .B(n18459), .Z(n18463) );
  XNOR U18106 ( .A(n18412), .B(n18455), .Z(n18457) );
  XNOR U18107 ( .A(n18466), .B(n18467), .Z(n18412) );
  AND U18108 ( .A(n160), .B(n18419), .Z(n18467) );
  XOR U18109 ( .A(n18466), .B(n18417), .Z(n18419) );
  XOR U18110 ( .A(n18468), .B(n18469), .Z(n18455) );
  AND U18111 ( .A(n18470), .B(n18471), .Z(n18469) );
  XNOR U18112 ( .A(n18468), .B(n18427), .Z(n18471) );
  XOR U18113 ( .A(n18472), .B(n18464), .Z(n18427) );
  XNOR U18114 ( .A(n18473), .B(n18459), .Z(n18464) );
  XOR U18115 ( .A(n18474), .B(n18475), .Z(n18459) );
  AND U18116 ( .A(n18476), .B(n18477), .Z(n18475) );
  XOR U18117 ( .A(n18478), .B(n18474), .Z(n18476) );
  XNOR U18118 ( .A(n18479), .B(n18480), .Z(n18473) );
  AND U18119 ( .A(n18481), .B(n18482), .Z(n18480) );
  XOR U18120 ( .A(n18479), .B(n18483), .Z(n18481) );
  XNOR U18121 ( .A(n18465), .B(n18462), .Z(n18472) );
  AND U18122 ( .A(n18484), .B(n18485), .Z(n18462) );
  XOR U18123 ( .A(n18486), .B(n18487), .Z(n18465) );
  AND U18124 ( .A(n18488), .B(n18489), .Z(n18487) );
  XOR U18125 ( .A(n18486), .B(n18490), .Z(n18488) );
  XNOR U18126 ( .A(n18424), .B(n18468), .Z(n18470) );
  XNOR U18127 ( .A(n18491), .B(n18492), .Z(n18424) );
  AND U18128 ( .A(n160), .B(n18430), .Z(n18492) );
  XOR U18129 ( .A(n18491), .B(n18428), .Z(n18430) );
  XOR U18130 ( .A(n18493), .B(n18494), .Z(n18468) );
  AND U18131 ( .A(n18495), .B(n18496), .Z(n18494) );
  XNOR U18132 ( .A(n18493), .B(n18484), .Z(n18496) );
  IV U18133 ( .A(n18438), .Z(n18484) );
  XNOR U18134 ( .A(n18497), .B(n18477), .Z(n18438) );
  XNOR U18135 ( .A(n18498), .B(n18483), .Z(n18477) );
  XNOR U18136 ( .A(n18499), .B(n18500), .Z(n18483) );
  NOR U18137 ( .A(n18501), .B(n18502), .Z(n18500) );
  XOR U18138 ( .A(n18499), .B(n18503), .Z(n18501) );
  XNOR U18139 ( .A(n18482), .B(n18474), .Z(n18498) );
  XOR U18140 ( .A(n18504), .B(n18505), .Z(n18474) );
  AND U18141 ( .A(n18506), .B(n18507), .Z(n18505) );
  XOR U18142 ( .A(n18504), .B(n18508), .Z(n18506) );
  XNOR U18143 ( .A(n18509), .B(n18479), .Z(n18482) );
  XOR U18144 ( .A(n18510), .B(n18511), .Z(n18479) );
  AND U18145 ( .A(n18512), .B(n18513), .Z(n18511) );
  XNOR U18146 ( .A(n18514), .B(n18515), .Z(n18512) );
  IV U18147 ( .A(n18510), .Z(n18514) );
  XNOR U18148 ( .A(n18516), .B(n18517), .Z(n18509) );
  NOR U18149 ( .A(n18518), .B(n18519), .Z(n18517) );
  XNOR U18150 ( .A(n18516), .B(n18520), .Z(n18518) );
  XNOR U18151 ( .A(n18478), .B(n18485), .Z(n18497) );
  NOR U18152 ( .A(n18446), .B(n18521), .Z(n18485) );
  XOR U18153 ( .A(n18490), .B(n18489), .Z(n18478) );
  XNOR U18154 ( .A(n18522), .B(n18486), .Z(n18489) );
  XOR U18155 ( .A(n18523), .B(n18524), .Z(n18486) );
  AND U18156 ( .A(n18525), .B(n18526), .Z(n18524) );
  XNOR U18157 ( .A(n18527), .B(n18528), .Z(n18525) );
  IV U18158 ( .A(n18523), .Z(n18527) );
  XNOR U18159 ( .A(n18529), .B(n18530), .Z(n18522) );
  NOR U18160 ( .A(n18531), .B(n18532), .Z(n18530) );
  XNOR U18161 ( .A(n18529), .B(n18533), .Z(n18531) );
  XOR U18162 ( .A(n18534), .B(n18535), .Z(n18490) );
  NOR U18163 ( .A(n18536), .B(n18537), .Z(n18535) );
  XNOR U18164 ( .A(n18534), .B(n18538), .Z(n18536) );
  XNOR U18165 ( .A(n18435), .B(n18493), .Z(n18495) );
  XNOR U18166 ( .A(n18539), .B(n18540), .Z(n18435) );
  AND U18167 ( .A(n160), .B(n18442), .Z(n18540) );
  XOR U18168 ( .A(n18539), .B(n18440), .Z(n18442) );
  AND U18169 ( .A(n18443), .B(n18446), .Z(n18493) );
  XOR U18170 ( .A(n18541), .B(n18521), .Z(n18446) );
  XNOR U18171 ( .A(p_input[176]), .B(p_input[2048]), .Z(n18521) );
  XNOR U18172 ( .A(n18508), .B(n18507), .Z(n18541) );
  XNOR U18173 ( .A(n18542), .B(n18515), .Z(n18507) );
  XNOR U18174 ( .A(n18503), .B(n18502), .Z(n18515) );
  XNOR U18175 ( .A(n18543), .B(n18499), .Z(n18502) );
  XNOR U18176 ( .A(p_input[186]), .B(p_input[2058]), .Z(n18499) );
  XOR U18177 ( .A(p_input[187]), .B(n16732), .Z(n18543) );
  XOR U18178 ( .A(p_input[188]), .B(p_input[2060]), .Z(n18503) );
  XOR U18179 ( .A(n18513), .B(n18544), .Z(n18542) );
  IV U18180 ( .A(n18504), .Z(n18544) );
  XOR U18181 ( .A(p_input[177]), .B(p_input[2049]), .Z(n18504) );
  XNOR U18182 ( .A(n18545), .B(n18520), .Z(n18513) );
  XNOR U18183 ( .A(p_input[191]), .B(n16735), .Z(n18520) );
  XOR U18184 ( .A(n18510), .B(n18519), .Z(n18545) );
  XOR U18185 ( .A(n18546), .B(n18516), .Z(n18519) );
  XOR U18186 ( .A(p_input[189]), .B(p_input[2061]), .Z(n18516) );
  XOR U18187 ( .A(p_input[190]), .B(n16737), .Z(n18546) );
  XOR U18188 ( .A(p_input[185]), .B(p_input[2057]), .Z(n18510) );
  XOR U18189 ( .A(n18528), .B(n18526), .Z(n18508) );
  XNOR U18190 ( .A(n18547), .B(n18533), .Z(n18526) );
  XOR U18191 ( .A(p_input[184]), .B(p_input[2056]), .Z(n18533) );
  XOR U18192 ( .A(n18523), .B(n18532), .Z(n18547) );
  XOR U18193 ( .A(n18548), .B(n18529), .Z(n18532) );
  XOR U18194 ( .A(p_input[182]), .B(p_input[2054]), .Z(n18529) );
  XOR U18195 ( .A(p_input[183]), .B(n17722), .Z(n18548) );
  XOR U18196 ( .A(p_input[178]), .B(p_input[2050]), .Z(n18523) );
  XNOR U18197 ( .A(n18538), .B(n18537), .Z(n18528) );
  XOR U18198 ( .A(n18549), .B(n18534), .Z(n18537) );
  XOR U18199 ( .A(p_input[179]), .B(p_input[2051]), .Z(n18534) );
  XOR U18200 ( .A(p_input[180]), .B(n17724), .Z(n18549) );
  XOR U18201 ( .A(p_input[181]), .B(p_input[2053]), .Z(n18538) );
  XNOR U18202 ( .A(n18550), .B(n18551), .Z(n18443) );
  AND U18203 ( .A(n160), .B(n18552), .Z(n18551) );
  XNOR U18204 ( .A(n18553), .B(n18554), .Z(n160) );
  AND U18205 ( .A(n18555), .B(n18556), .Z(n18554) );
  XOR U18206 ( .A(n18553), .B(n18453), .Z(n18556) );
  XNOR U18207 ( .A(n18553), .B(n18407), .Z(n18555) );
  XOR U18208 ( .A(n18557), .B(n18558), .Z(n18553) );
  AND U18209 ( .A(n18559), .B(n18560), .Z(n18558) );
  XOR U18210 ( .A(n18557), .B(n18417), .Z(n18559) );
  XOR U18211 ( .A(n18561), .B(n18562), .Z(n18396) );
  AND U18212 ( .A(n164), .B(n18552), .Z(n18562) );
  XNOR U18213 ( .A(n18550), .B(n18561), .Z(n18552) );
  XNOR U18214 ( .A(n18563), .B(n18564), .Z(n164) );
  AND U18215 ( .A(n18565), .B(n18566), .Z(n18564) );
  XNOR U18216 ( .A(n18567), .B(n18563), .Z(n18566) );
  IV U18217 ( .A(n18453), .Z(n18567) );
  XNOR U18218 ( .A(n18568), .B(n18569), .Z(n18453) );
  AND U18219 ( .A(n167), .B(n18570), .Z(n18569) );
  XNOR U18220 ( .A(n18568), .B(n18571), .Z(n18570) );
  XNOR U18221 ( .A(n18407), .B(n18563), .Z(n18565) );
  XOR U18222 ( .A(n18572), .B(n18573), .Z(n18407) );
  AND U18223 ( .A(n175), .B(n18574), .Z(n18573) );
  XOR U18224 ( .A(n18557), .B(n18575), .Z(n18563) );
  AND U18225 ( .A(n18576), .B(n18560), .Z(n18575) );
  XNOR U18226 ( .A(n18466), .B(n18557), .Z(n18560) );
  XNOR U18227 ( .A(n18577), .B(n18578), .Z(n18466) );
  AND U18228 ( .A(n167), .B(n18579), .Z(n18578) );
  XOR U18229 ( .A(n18580), .B(n18577), .Z(n18579) );
  XNOR U18230 ( .A(n18581), .B(n18557), .Z(n18576) );
  IV U18231 ( .A(n18417), .Z(n18581) );
  XOR U18232 ( .A(n18582), .B(n18583), .Z(n18417) );
  AND U18233 ( .A(n175), .B(n18584), .Z(n18583) );
  XOR U18234 ( .A(n18585), .B(n18586), .Z(n18557) );
  AND U18235 ( .A(n18587), .B(n18588), .Z(n18586) );
  XNOR U18236 ( .A(n18491), .B(n18585), .Z(n18588) );
  XNOR U18237 ( .A(n18589), .B(n18590), .Z(n18491) );
  AND U18238 ( .A(n167), .B(n18591), .Z(n18590) );
  XNOR U18239 ( .A(n18592), .B(n18589), .Z(n18591) );
  XOR U18240 ( .A(n18585), .B(n18428), .Z(n18587) );
  XOR U18241 ( .A(n18593), .B(n18594), .Z(n18428) );
  AND U18242 ( .A(n175), .B(n18595), .Z(n18594) );
  XOR U18243 ( .A(n18596), .B(n18597), .Z(n18585) );
  AND U18244 ( .A(n18598), .B(n18599), .Z(n18597) );
  XNOR U18245 ( .A(n18596), .B(n18539), .Z(n18599) );
  XNOR U18246 ( .A(n18600), .B(n18601), .Z(n18539) );
  AND U18247 ( .A(n167), .B(n18602), .Z(n18601) );
  XOR U18248 ( .A(n18603), .B(n18600), .Z(n18602) );
  XNOR U18249 ( .A(n18604), .B(n18596), .Z(n18598) );
  IV U18250 ( .A(n18440), .Z(n18604) );
  XOR U18251 ( .A(n18605), .B(n18606), .Z(n18440) );
  AND U18252 ( .A(n175), .B(n18607), .Z(n18606) );
  AND U18253 ( .A(n18561), .B(n18550), .Z(n18596) );
  XNOR U18254 ( .A(n18608), .B(n18609), .Z(n18550) );
  AND U18255 ( .A(n167), .B(n18610), .Z(n18609) );
  XNOR U18256 ( .A(n18611), .B(n18608), .Z(n18610) );
  XNOR U18257 ( .A(n18612), .B(n18613), .Z(n167) );
  AND U18258 ( .A(n18614), .B(n18615), .Z(n18613) );
  XOR U18259 ( .A(n18571), .B(n18612), .Z(n18615) );
  AND U18260 ( .A(n18616), .B(n18617), .Z(n18571) );
  XOR U18261 ( .A(n18612), .B(n18568), .Z(n18614) );
  XNOR U18262 ( .A(n18618), .B(n18619), .Z(n18568) );
  AND U18263 ( .A(n171), .B(n18574), .Z(n18619) );
  XOR U18264 ( .A(n18572), .B(n18618), .Z(n18574) );
  XOR U18265 ( .A(n18620), .B(n18621), .Z(n18612) );
  AND U18266 ( .A(n18622), .B(n18623), .Z(n18621) );
  XNOR U18267 ( .A(n18620), .B(n18616), .Z(n18623) );
  IV U18268 ( .A(n18580), .Z(n18616) );
  XOR U18269 ( .A(n18624), .B(n18625), .Z(n18580) );
  XOR U18270 ( .A(n18626), .B(n18617), .Z(n18625) );
  AND U18271 ( .A(n18592), .B(n18627), .Z(n18617) );
  AND U18272 ( .A(n18628), .B(n18629), .Z(n18626) );
  XOR U18273 ( .A(n18630), .B(n18624), .Z(n18628) );
  XNOR U18274 ( .A(n18577), .B(n18620), .Z(n18622) );
  XNOR U18275 ( .A(n18631), .B(n18632), .Z(n18577) );
  AND U18276 ( .A(n171), .B(n18584), .Z(n18632) );
  XOR U18277 ( .A(n18631), .B(n18582), .Z(n18584) );
  XOR U18278 ( .A(n18633), .B(n18634), .Z(n18620) );
  AND U18279 ( .A(n18635), .B(n18636), .Z(n18634) );
  XNOR U18280 ( .A(n18633), .B(n18592), .Z(n18636) );
  XOR U18281 ( .A(n18637), .B(n18629), .Z(n18592) );
  XNOR U18282 ( .A(n18638), .B(n18624), .Z(n18629) );
  XOR U18283 ( .A(n18639), .B(n18640), .Z(n18624) );
  AND U18284 ( .A(n18641), .B(n18642), .Z(n18640) );
  XOR U18285 ( .A(n18643), .B(n18639), .Z(n18641) );
  XNOR U18286 ( .A(n18644), .B(n18645), .Z(n18638) );
  AND U18287 ( .A(n18646), .B(n18647), .Z(n18645) );
  XOR U18288 ( .A(n18644), .B(n18648), .Z(n18646) );
  XNOR U18289 ( .A(n18630), .B(n18627), .Z(n18637) );
  AND U18290 ( .A(n18649), .B(n18650), .Z(n18627) );
  XOR U18291 ( .A(n18651), .B(n18652), .Z(n18630) );
  AND U18292 ( .A(n18653), .B(n18654), .Z(n18652) );
  XOR U18293 ( .A(n18651), .B(n18655), .Z(n18653) );
  XNOR U18294 ( .A(n18589), .B(n18633), .Z(n18635) );
  XNOR U18295 ( .A(n18656), .B(n18657), .Z(n18589) );
  AND U18296 ( .A(n171), .B(n18595), .Z(n18657) );
  XOR U18297 ( .A(n18656), .B(n18593), .Z(n18595) );
  XOR U18298 ( .A(n18658), .B(n18659), .Z(n18633) );
  AND U18299 ( .A(n18660), .B(n18661), .Z(n18659) );
  XNOR U18300 ( .A(n18658), .B(n18649), .Z(n18661) );
  IV U18301 ( .A(n18603), .Z(n18649) );
  XNOR U18302 ( .A(n18662), .B(n18642), .Z(n18603) );
  XNOR U18303 ( .A(n18663), .B(n18648), .Z(n18642) );
  XNOR U18304 ( .A(n18664), .B(n18665), .Z(n18648) );
  NOR U18305 ( .A(n18666), .B(n18667), .Z(n18665) );
  XOR U18306 ( .A(n18664), .B(n18668), .Z(n18666) );
  XNOR U18307 ( .A(n18647), .B(n18639), .Z(n18663) );
  XOR U18308 ( .A(n18669), .B(n18670), .Z(n18639) );
  AND U18309 ( .A(n18671), .B(n18672), .Z(n18670) );
  XOR U18310 ( .A(n18669), .B(n18673), .Z(n18671) );
  XNOR U18311 ( .A(n18674), .B(n18644), .Z(n18647) );
  XOR U18312 ( .A(n18675), .B(n18676), .Z(n18644) );
  AND U18313 ( .A(n18677), .B(n18678), .Z(n18676) );
  XNOR U18314 ( .A(n18679), .B(n18680), .Z(n18677) );
  IV U18315 ( .A(n18675), .Z(n18679) );
  XNOR U18316 ( .A(n18681), .B(n18682), .Z(n18674) );
  NOR U18317 ( .A(n18683), .B(n18684), .Z(n18682) );
  XOR U18318 ( .A(n18681), .B(n18685), .Z(n18683) );
  XNOR U18319 ( .A(n18643), .B(n18650), .Z(n18662) );
  NOR U18320 ( .A(n18611), .B(n18686), .Z(n18650) );
  XOR U18321 ( .A(n18655), .B(n18654), .Z(n18643) );
  XNOR U18322 ( .A(n18687), .B(n18651), .Z(n18654) );
  XOR U18323 ( .A(n18688), .B(n18689), .Z(n18651) );
  AND U18324 ( .A(n18690), .B(n18691), .Z(n18689) );
  XNOR U18325 ( .A(n18692), .B(n18693), .Z(n18690) );
  IV U18326 ( .A(n18688), .Z(n18692) );
  XNOR U18327 ( .A(n18694), .B(n18695), .Z(n18687) );
  NOR U18328 ( .A(n18696), .B(n18697), .Z(n18695) );
  XNOR U18329 ( .A(n18694), .B(n18698), .Z(n18696) );
  XOR U18330 ( .A(n18699), .B(n18700), .Z(n18655) );
  NOR U18331 ( .A(n18701), .B(n18702), .Z(n18700) );
  XNOR U18332 ( .A(n18699), .B(n18703), .Z(n18701) );
  XNOR U18333 ( .A(n18600), .B(n18658), .Z(n18660) );
  XNOR U18334 ( .A(n18704), .B(n18705), .Z(n18600) );
  AND U18335 ( .A(n171), .B(n18607), .Z(n18705) );
  XOR U18336 ( .A(n18704), .B(n18605), .Z(n18607) );
  AND U18337 ( .A(n18608), .B(n18611), .Z(n18658) );
  XOR U18338 ( .A(n18706), .B(n18686), .Z(n18611) );
  XNOR U18339 ( .A(p_input[192]), .B(p_input[2048]), .Z(n18686) );
  XNOR U18340 ( .A(n18673), .B(n18672), .Z(n18706) );
  XNOR U18341 ( .A(n18707), .B(n18680), .Z(n18672) );
  XNOR U18342 ( .A(n18668), .B(n18667), .Z(n18680) );
  XNOR U18343 ( .A(n18708), .B(n18664), .Z(n18667) );
  XNOR U18344 ( .A(p_input[202]), .B(p_input[2058]), .Z(n18664) );
  XOR U18345 ( .A(p_input[203]), .B(n16732), .Z(n18708) );
  XOR U18346 ( .A(p_input[204]), .B(p_input[2060]), .Z(n18668) );
  XOR U18347 ( .A(n18678), .B(n18709), .Z(n18707) );
  IV U18348 ( .A(n18669), .Z(n18709) );
  XOR U18349 ( .A(p_input[193]), .B(p_input[2049]), .Z(n18669) );
  XOR U18350 ( .A(n18710), .B(n18685), .Z(n18678) );
  XNOR U18351 ( .A(p_input[2063]), .B(p_input[207]), .Z(n18685) );
  XOR U18352 ( .A(n18675), .B(n18684), .Z(n18710) );
  XOR U18353 ( .A(n18711), .B(n18681), .Z(n18684) );
  XOR U18354 ( .A(p_input[205]), .B(p_input[2061]), .Z(n18681) );
  XNOR U18355 ( .A(p_input[2062]), .B(p_input[206]), .Z(n18711) );
  XOR U18356 ( .A(p_input[201]), .B(p_input[2057]), .Z(n18675) );
  XOR U18357 ( .A(n18693), .B(n18691), .Z(n18673) );
  XNOR U18358 ( .A(n18712), .B(n18698), .Z(n18691) );
  XOR U18359 ( .A(p_input[200]), .B(p_input[2056]), .Z(n18698) );
  XOR U18360 ( .A(n18688), .B(n18697), .Z(n18712) );
  XOR U18361 ( .A(n18713), .B(n18694), .Z(n18697) );
  XOR U18362 ( .A(p_input[198]), .B(p_input[2054]), .Z(n18694) );
  XOR U18363 ( .A(p_input[199]), .B(n17722), .Z(n18713) );
  XOR U18364 ( .A(p_input[194]), .B(p_input[2050]), .Z(n18688) );
  XNOR U18365 ( .A(n18703), .B(n18702), .Z(n18693) );
  XOR U18366 ( .A(n18714), .B(n18699), .Z(n18702) );
  XOR U18367 ( .A(p_input[195]), .B(p_input[2051]), .Z(n18699) );
  XOR U18368 ( .A(p_input[196]), .B(n17724), .Z(n18714) );
  XOR U18369 ( .A(p_input[197]), .B(p_input[2053]), .Z(n18703) );
  XNOR U18370 ( .A(n18715), .B(n18716), .Z(n18608) );
  AND U18371 ( .A(n171), .B(n18717), .Z(n18716) );
  XNOR U18372 ( .A(n18718), .B(n18719), .Z(n171) );
  AND U18373 ( .A(n18720), .B(n18721), .Z(n18719) );
  XOR U18374 ( .A(n18718), .B(n18618), .Z(n18721) );
  XNOR U18375 ( .A(n18718), .B(n18572), .Z(n18720) );
  XOR U18376 ( .A(n18722), .B(n18723), .Z(n18718) );
  AND U18377 ( .A(n18724), .B(n18725), .Z(n18723) );
  XOR U18378 ( .A(n18722), .B(n18582), .Z(n18724) );
  XOR U18379 ( .A(n18726), .B(n18727), .Z(n18561) );
  AND U18380 ( .A(n175), .B(n18717), .Z(n18727) );
  XNOR U18381 ( .A(n18715), .B(n18726), .Z(n18717) );
  XNOR U18382 ( .A(n18728), .B(n18729), .Z(n175) );
  AND U18383 ( .A(n18730), .B(n18731), .Z(n18729) );
  XNOR U18384 ( .A(n18732), .B(n18728), .Z(n18731) );
  IV U18385 ( .A(n18618), .Z(n18732) );
  XNOR U18386 ( .A(n18733), .B(n18734), .Z(n18618) );
  AND U18387 ( .A(n178), .B(n18735), .Z(n18734) );
  XNOR U18388 ( .A(n18733), .B(n18736), .Z(n18735) );
  XNOR U18389 ( .A(n18572), .B(n18728), .Z(n18730) );
  XOR U18390 ( .A(n18737), .B(n18738), .Z(n18572) );
  AND U18391 ( .A(n186), .B(n18739), .Z(n18738) );
  XOR U18392 ( .A(n18722), .B(n18740), .Z(n18728) );
  AND U18393 ( .A(n18741), .B(n18725), .Z(n18740) );
  XNOR U18394 ( .A(n18631), .B(n18722), .Z(n18725) );
  XNOR U18395 ( .A(n18742), .B(n18743), .Z(n18631) );
  AND U18396 ( .A(n178), .B(n18744), .Z(n18743) );
  XOR U18397 ( .A(n18745), .B(n18742), .Z(n18744) );
  XNOR U18398 ( .A(n18746), .B(n18722), .Z(n18741) );
  IV U18399 ( .A(n18582), .Z(n18746) );
  XOR U18400 ( .A(n18747), .B(n18748), .Z(n18582) );
  AND U18401 ( .A(n186), .B(n18749), .Z(n18748) );
  XOR U18402 ( .A(n18750), .B(n18751), .Z(n18722) );
  AND U18403 ( .A(n18752), .B(n18753), .Z(n18751) );
  XNOR U18404 ( .A(n18656), .B(n18750), .Z(n18753) );
  XNOR U18405 ( .A(n18754), .B(n18755), .Z(n18656) );
  AND U18406 ( .A(n178), .B(n18756), .Z(n18755) );
  XNOR U18407 ( .A(n18757), .B(n18754), .Z(n18756) );
  XOR U18408 ( .A(n18750), .B(n18593), .Z(n18752) );
  XOR U18409 ( .A(n18758), .B(n18759), .Z(n18593) );
  AND U18410 ( .A(n186), .B(n18760), .Z(n18759) );
  XOR U18411 ( .A(n18761), .B(n18762), .Z(n18750) );
  AND U18412 ( .A(n18763), .B(n18764), .Z(n18762) );
  XNOR U18413 ( .A(n18761), .B(n18704), .Z(n18764) );
  XNOR U18414 ( .A(n18765), .B(n18766), .Z(n18704) );
  AND U18415 ( .A(n178), .B(n18767), .Z(n18766) );
  XOR U18416 ( .A(n18768), .B(n18765), .Z(n18767) );
  XNOR U18417 ( .A(n18769), .B(n18761), .Z(n18763) );
  IV U18418 ( .A(n18605), .Z(n18769) );
  XOR U18419 ( .A(n18770), .B(n18771), .Z(n18605) );
  AND U18420 ( .A(n186), .B(n18772), .Z(n18771) );
  AND U18421 ( .A(n18726), .B(n18715), .Z(n18761) );
  XNOR U18422 ( .A(n18773), .B(n18774), .Z(n18715) );
  AND U18423 ( .A(n178), .B(n18775), .Z(n18774) );
  XNOR U18424 ( .A(n18776), .B(n18773), .Z(n18775) );
  XNOR U18425 ( .A(n18777), .B(n18778), .Z(n178) );
  AND U18426 ( .A(n18779), .B(n18780), .Z(n18778) );
  XOR U18427 ( .A(n18736), .B(n18777), .Z(n18780) );
  AND U18428 ( .A(n18781), .B(n18782), .Z(n18736) );
  XOR U18429 ( .A(n18777), .B(n18733), .Z(n18779) );
  XNOR U18430 ( .A(n18783), .B(n18784), .Z(n18733) );
  AND U18431 ( .A(n182), .B(n18739), .Z(n18784) );
  XOR U18432 ( .A(n18737), .B(n18783), .Z(n18739) );
  XOR U18433 ( .A(n18785), .B(n18786), .Z(n18777) );
  AND U18434 ( .A(n18787), .B(n18788), .Z(n18786) );
  XNOR U18435 ( .A(n18785), .B(n18781), .Z(n18788) );
  IV U18436 ( .A(n18745), .Z(n18781) );
  XOR U18437 ( .A(n18789), .B(n18790), .Z(n18745) );
  XOR U18438 ( .A(n18791), .B(n18782), .Z(n18790) );
  AND U18439 ( .A(n18757), .B(n18792), .Z(n18782) );
  AND U18440 ( .A(n18793), .B(n18794), .Z(n18791) );
  XOR U18441 ( .A(n18795), .B(n18789), .Z(n18793) );
  XNOR U18442 ( .A(n18742), .B(n18785), .Z(n18787) );
  XNOR U18443 ( .A(n18796), .B(n18797), .Z(n18742) );
  AND U18444 ( .A(n182), .B(n18749), .Z(n18797) );
  XOR U18445 ( .A(n18796), .B(n18747), .Z(n18749) );
  XOR U18446 ( .A(n18798), .B(n18799), .Z(n18785) );
  AND U18447 ( .A(n18800), .B(n18801), .Z(n18799) );
  XNOR U18448 ( .A(n18798), .B(n18757), .Z(n18801) );
  XOR U18449 ( .A(n18802), .B(n18794), .Z(n18757) );
  XNOR U18450 ( .A(n18803), .B(n18789), .Z(n18794) );
  XOR U18451 ( .A(n18804), .B(n18805), .Z(n18789) );
  AND U18452 ( .A(n18806), .B(n18807), .Z(n18805) );
  XOR U18453 ( .A(n18808), .B(n18804), .Z(n18806) );
  XNOR U18454 ( .A(n18809), .B(n18810), .Z(n18803) );
  AND U18455 ( .A(n18811), .B(n18812), .Z(n18810) );
  XOR U18456 ( .A(n18809), .B(n18813), .Z(n18811) );
  XNOR U18457 ( .A(n18795), .B(n18792), .Z(n18802) );
  AND U18458 ( .A(n18814), .B(n18815), .Z(n18792) );
  XOR U18459 ( .A(n18816), .B(n18817), .Z(n18795) );
  AND U18460 ( .A(n18818), .B(n18819), .Z(n18817) );
  XOR U18461 ( .A(n18816), .B(n18820), .Z(n18818) );
  XNOR U18462 ( .A(n18754), .B(n18798), .Z(n18800) );
  XNOR U18463 ( .A(n18821), .B(n18822), .Z(n18754) );
  AND U18464 ( .A(n182), .B(n18760), .Z(n18822) );
  XOR U18465 ( .A(n18821), .B(n18758), .Z(n18760) );
  XOR U18466 ( .A(n18823), .B(n18824), .Z(n18798) );
  AND U18467 ( .A(n18825), .B(n18826), .Z(n18824) );
  XNOR U18468 ( .A(n18823), .B(n18814), .Z(n18826) );
  IV U18469 ( .A(n18768), .Z(n18814) );
  XNOR U18470 ( .A(n18827), .B(n18807), .Z(n18768) );
  XNOR U18471 ( .A(n18828), .B(n18813), .Z(n18807) );
  XOR U18472 ( .A(n18829), .B(n18830), .Z(n18813) );
  NOR U18473 ( .A(n18831), .B(n18832), .Z(n18830) );
  XNOR U18474 ( .A(n18829), .B(n18833), .Z(n18831) );
  XNOR U18475 ( .A(n18812), .B(n18804), .Z(n18828) );
  XOR U18476 ( .A(n18834), .B(n18835), .Z(n18804) );
  AND U18477 ( .A(n18836), .B(n18837), .Z(n18835) );
  XNOR U18478 ( .A(n18834), .B(n18838), .Z(n18836) );
  XNOR U18479 ( .A(n18839), .B(n18809), .Z(n18812) );
  XOR U18480 ( .A(n18840), .B(n18841), .Z(n18809) );
  AND U18481 ( .A(n18842), .B(n18843), .Z(n18841) );
  XOR U18482 ( .A(n18840), .B(n18844), .Z(n18842) );
  XNOR U18483 ( .A(n18845), .B(n18846), .Z(n18839) );
  NOR U18484 ( .A(n18847), .B(n18848), .Z(n18846) );
  XOR U18485 ( .A(n18845), .B(n18849), .Z(n18847) );
  XNOR U18486 ( .A(n18808), .B(n18815), .Z(n18827) );
  NOR U18487 ( .A(n18776), .B(n18850), .Z(n18815) );
  XOR U18488 ( .A(n18820), .B(n18819), .Z(n18808) );
  XNOR U18489 ( .A(n18851), .B(n18816), .Z(n18819) );
  XOR U18490 ( .A(n18852), .B(n18853), .Z(n18816) );
  AND U18491 ( .A(n18854), .B(n18855), .Z(n18853) );
  XOR U18492 ( .A(n18852), .B(n18856), .Z(n18854) );
  XNOR U18493 ( .A(n18857), .B(n18858), .Z(n18851) );
  NOR U18494 ( .A(n18859), .B(n18860), .Z(n18858) );
  XNOR U18495 ( .A(n18857), .B(n18861), .Z(n18859) );
  XOR U18496 ( .A(n18862), .B(n18863), .Z(n18820) );
  NOR U18497 ( .A(n18864), .B(n18865), .Z(n18863) );
  XNOR U18498 ( .A(n18862), .B(n18866), .Z(n18864) );
  XNOR U18499 ( .A(n18765), .B(n18823), .Z(n18825) );
  XNOR U18500 ( .A(n18867), .B(n18868), .Z(n18765) );
  AND U18501 ( .A(n182), .B(n18772), .Z(n18868) );
  XOR U18502 ( .A(n18867), .B(n18770), .Z(n18772) );
  AND U18503 ( .A(n18773), .B(n18776), .Z(n18823) );
  XOR U18504 ( .A(n18869), .B(n18850), .Z(n18776) );
  XNOR U18505 ( .A(p_input[2048]), .B(p_input[208]), .Z(n18850) );
  XOR U18506 ( .A(n18838), .B(n18837), .Z(n18869) );
  XNOR U18507 ( .A(n18870), .B(n18844), .Z(n18837) );
  XNOR U18508 ( .A(n18833), .B(n18832), .Z(n18844) );
  XOR U18509 ( .A(n18871), .B(n18829), .Z(n18832) );
  XNOR U18510 ( .A(n16904), .B(p_input[218]), .Z(n18829) );
  XNOR U18511 ( .A(p_input[2059]), .B(p_input[219]), .Z(n18871) );
  XOR U18512 ( .A(p_input[2060]), .B(p_input[220]), .Z(n18833) );
  XNOR U18513 ( .A(n18843), .B(n18834), .Z(n18870) );
  XNOR U18514 ( .A(n17068), .B(p_input[209]), .Z(n18834) );
  XOR U18515 ( .A(n18872), .B(n18849), .Z(n18843) );
  XNOR U18516 ( .A(p_input[2063]), .B(p_input[223]), .Z(n18849) );
  XOR U18517 ( .A(n18840), .B(n18848), .Z(n18872) );
  XOR U18518 ( .A(n18873), .B(n18845), .Z(n18848) );
  XOR U18519 ( .A(p_input[2061]), .B(p_input[221]), .Z(n18845) );
  XNOR U18520 ( .A(p_input[2062]), .B(p_input[222]), .Z(n18873) );
  XNOR U18521 ( .A(n16738), .B(p_input[217]), .Z(n18840) );
  XNOR U18522 ( .A(n18856), .B(n18855), .Z(n18838) );
  XNOR U18523 ( .A(n18874), .B(n18861), .Z(n18855) );
  XOR U18524 ( .A(p_input[2056]), .B(p_input[216]), .Z(n18861) );
  XOR U18525 ( .A(n18852), .B(n18860), .Z(n18874) );
  XOR U18526 ( .A(n18875), .B(n18857), .Z(n18860) );
  XOR U18527 ( .A(p_input[2054]), .B(p_input[214]), .Z(n18857) );
  XNOR U18528 ( .A(p_input[2055]), .B(p_input[215]), .Z(n18875) );
  XNOR U18529 ( .A(n16741), .B(p_input[210]), .Z(n18852) );
  XNOR U18530 ( .A(n18866), .B(n18865), .Z(n18856) );
  XOR U18531 ( .A(n18876), .B(n18862), .Z(n18865) );
  XOR U18532 ( .A(p_input[2051]), .B(p_input[211]), .Z(n18862) );
  XNOR U18533 ( .A(p_input[2052]), .B(p_input[212]), .Z(n18876) );
  XOR U18534 ( .A(p_input[2053]), .B(p_input[213]), .Z(n18866) );
  XNOR U18535 ( .A(n18877), .B(n18878), .Z(n18773) );
  AND U18536 ( .A(n182), .B(n18879), .Z(n18878) );
  XNOR U18537 ( .A(n18880), .B(n18881), .Z(n182) );
  AND U18538 ( .A(n18882), .B(n18883), .Z(n18881) );
  XOR U18539 ( .A(n18880), .B(n18783), .Z(n18883) );
  XNOR U18540 ( .A(n18880), .B(n18737), .Z(n18882) );
  XOR U18541 ( .A(n18884), .B(n18885), .Z(n18880) );
  AND U18542 ( .A(n18886), .B(n18887), .Z(n18885) );
  XOR U18543 ( .A(n18884), .B(n18747), .Z(n18886) );
  XOR U18544 ( .A(n18888), .B(n18889), .Z(n18726) );
  AND U18545 ( .A(n186), .B(n18879), .Z(n18889) );
  XNOR U18546 ( .A(n18877), .B(n18888), .Z(n18879) );
  XNOR U18547 ( .A(n18890), .B(n18891), .Z(n186) );
  AND U18548 ( .A(n18892), .B(n18893), .Z(n18891) );
  XNOR U18549 ( .A(n18894), .B(n18890), .Z(n18893) );
  IV U18550 ( .A(n18783), .Z(n18894) );
  XNOR U18551 ( .A(n18895), .B(n18896), .Z(n18783) );
  AND U18552 ( .A(n189), .B(n18897), .Z(n18896) );
  XNOR U18553 ( .A(n18895), .B(n18898), .Z(n18897) );
  XNOR U18554 ( .A(n18737), .B(n18890), .Z(n18892) );
  XOR U18555 ( .A(n18899), .B(n18900), .Z(n18737) );
  AND U18556 ( .A(n197), .B(n18901), .Z(n18900) );
  XOR U18557 ( .A(n18884), .B(n18902), .Z(n18890) );
  AND U18558 ( .A(n18903), .B(n18887), .Z(n18902) );
  XNOR U18559 ( .A(n18796), .B(n18884), .Z(n18887) );
  XNOR U18560 ( .A(n18904), .B(n18905), .Z(n18796) );
  AND U18561 ( .A(n189), .B(n18906), .Z(n18905) );
  XOR U18562 ( .A(n18907), .B(n18904), .Z(n18906) );
  XNOR U18563 ( .A(n18908), .B(n18884), .Z(n18903) );
  IV U18564 ( .A(n18747), .Z(n18908) );
  XOR U18565 ( .A(n18909), .B(n18910), .Z(n18747) );
  AND U18566 ( .A(n197), .B(n18911), .Z(n18910) );
  XOR U18567 ( .A(n18912), .B(n18913), .Z(n18884) );
  AND U18568 ( .A(n18914), .B(n18915), .Z(n18913) );
  XNOR U18569 ( .A(n18821), .B(n18912), .Z(n18915) );
  XNOR U18570 ( .A(n18916), .B(n18917), .Z(n18821) );
  AND U18571 ( .A(n189), .B(n18918), .Z(n18917) );
  XNOR U18572 ( .A(n18919), .B(n18916), .Z(n18918) );
  XOR U18573 ( .A(n18912), .B(n18758), .Z(n18914) );
  XOR U18574 ( .A(n18920), .B(n18921), .Z(n18758) );
  AND U18575 ( .A(n197), .B(n18922), .Z(n18921) );
  XOR U18576 ( .A(n18923), .B(n18924), .Z(n18912) );
  AND U18577 ( .A(n18925), .B(n18926), .Z(n18924) );
  XNOR U18578 ( .A(n18923), .B(n18867), .Z(n18926) );
  XNOR U18579 ( .A(n18927), .B(n18928), .Z(n18867) );
  AND U18580 ( .A(n189), .B(n18929), .Z(n18928) );
  XOR U18581 ( .A(n18930), .B(n18927), .Z(n18929) );
  XNOR U18582 ( .A(n18931), .B(n18923), .Z(n18925) );
  IV U18583 ( .A(n18770), .Z(n18931) );
  XOR U18584 ( .A(n18932), .B(n18933), .Z(n18770) );
  AND U18585 ( .A(n197), .B(n18934), .Z(n18933) );
  AND U18586 ( .A(n18888), .B(n18877), .Z(n18923) );
  XNOR U18587 ( .A(n18935), .B(n18936), .Z(n18877) );
  AND U18588 ( .A(n189), .B(n18937), .Z(n18936) );
  XNOR U18589 ( .A(n18938), .B(n18935), .Z(n18937) );
  XNOR U18590 ( .A(n18939), .B(n18940), .Z(n189) );
  AND U18591 ( .A(n18941), .B(n18942), .Z(n18940) );
  XOR U18592 ( .A(n18898), .B(n18939), .Z(n18942) );
  AND U18593 ( .A(n18943), .B(n18944), .Z(n18898) );
  XOR U18594 ( .A(n18939), .B(n18895), .Z(n18941) );
  XNOR U18595 ( .A(n18945), .B(n18946), .Z(n18895) );
  AND U18596 ( .A(n193), .B(n18901), .Z(n18946) );
  XOR U18597 ( .A(n18899), .B(n18945), .Z(n18901) );
  XOR U18598 ( .A(n18947), .B(n18948), .Z(n18939) );
  AND U18599 ( .A(n18949), .B(n18950), .Z(n18948) );
  XNOR U18600 ( .A(n18947), .B(n18943), .Z(n18950) );
  IV U18601 ( .A(n18907), .Z(n18943) );
  XOR U18602 ( .A(n18951), .B(n18952), .Z(n18907) );
  XOR U18603 ( .A(n18953), .B(n18944), .Z(n18952) );
  AND U18604 ( .A(n18919), .B(n18954), .Z(n18944) );
  AND U18605 ( .A(n18955), .B(n18956), .Z(n18953) );
  XOR U18606 ( .A(n18957), .B(n18951), .Z(n18955) );
  XNOR U18607 ( .A(n18904), .B(n18947), .Z(n18949) );
  XNOR U18608 ( .A(n18958), .B(n18959), .Z(n18904) );
  AND U18609 ( .A(n193), .B(n18911), .Z(n18959) );
  XOR U18610 ( .A(n18958), .B(n18909), .Z(n18911) );
  XOR U18611 ( .A(n18960), .B(n18961), .Z(n18947) );
  AND U18612 ( .A(n18962), .B(n18963), .Z(n18961) );
  XNOR U18613 ( .A(n18960), .B(n18919), .Z(n18963) );
  XOR U18614 ( .A(n18964), .B(n18956), .Z(n18919) );
  XNOR U18615 ( .A(n18965), .B(n18951), .Z(n18956) );
  XOR U18616 ( .A(n18966), .B(n18967), .Z(n18951) );
  AND U18617 ( .A(n18968), .B(n18969), .Z(n18967) );
  XOR U18618 ( .A(n18970), .B(n18966), .Z(n18968) );
  XNOR U18619 ( .A(n18971), .B(n18972), .Z(n18965) );
  AND U18620 ( .A(n18973), .B(n18974), .Z(n18972) );
  XOR U18621 ( .A(n18971), .B(n18975), .Z(n18973) );
  XNOR U18622 ( .A(n18957), .B(n18954), .Z(n18964) );
  AND U18623 ( .A(n18976), .B(n18977), .Z(n18954) );
  XOR U18624 ( .A(n18978), .B(n18979), .Z(n18957) );
  AND U18625 ( .A(n18980), .B(n18981), .Z(n18979) );
  XOR U18626 ( .A(n18978), .B(n18982), .Z(n18980) );
  XNOR U18627 ( .A(n18916), .B(n18960), .Z(n18962) );
  XNOR U18628 ( .A(n18983), .B(n18984), .Z(n18916) );
  AND U18629 ( .A(n193), .B(n18922), .Z(n18984) );
  XOR U18630 ( .A(n18983), .B(n18920), .Z(n18922) );
  XOR U18631 ( .A(n18985), .B(n18986), .Z(n18960) );
  AND U18632 ( .A(n18987), .B(n18988), .Z(n18986) );
  XNOR U18633 ( .A(n18985), .B(n18976), .Z(n18988) );
  IV U18634 ( .A(n18930), .Z(n18976) );
  XNOR U18635 ( .A(n18989), .B(n18969), .Z(n18930) );
  XNOR U18636 ( .A(n18990), .B(n18975), .Z(n18969) );
  XOR U18637 ( .A(n18991), .B(n18992), .Z(n18975) );
  NOR U18638 ( .A(n18993), .B(n18994), .Z(n18992) );
  XNOR U18639 ( .A(n18991), .B(n18995), .Z(n18993) );
  XNOR U18640 ( .A(n18974), .B(n18966), .Z(n18990) );
  XOR U18641 ( .A(n18996), .B(n18997), .Z(n18966) );
  AND U18642 ( .A(n18998), .B(n18999), .Z(n18997) );
  XNOR U18643 ( .A(n18996), .B(n19000), .Z(n18998) );
  XNOR U18644 ( .A(n19001), .B(n18971), .Z(n18974) );
  XOR U18645 ( .A(n19002), .B(n19003), .Z(n18971) );
  AND U18646 ( .A(n19004), .B(n19005), .Z(n19003) );
  XOR U18647 ( .A(n19002), .B(n19006), .Z(n19004) );
  XNOR U18648 ( .A(n19007), .B(n19008), .Z(n19001) );
  NOR U18649 ( .A(n19009), .B(n19010), .Z(n19008) );
  XOR U18650 ( .A(n19007), .B(n19011), .Z(n19009) );
  XNOR U18651 ( .A(n18970), .B(n18977), .Z(n18989) );
  NOR U18652 ( .A(n18938), .B(n19012), .Z(n18977) );
  XOR U18653 ( .A(n18982), .B(n18981), .Z(n18970) );
  XNOR U18654 ( .A(n19013), .B(n18978), .Z(n18981) );
  XOR U18655 ( .A(n19014), .B(n19015), .Z(n18978) );
  AND U18656 ( .A(n19016), .B(n19017), .Z(n19015) );
  XOR U18657 ( .A(n19014), .B(n19018), .Z(n19016) );
  XNOR U18658 ( .A(n19019), .B(n19020), .Z(n19013) );
  NOR U18659 ( .A(n19021), .B(n19022), .Z(n19020) );
  XNOR U18660 ( .A(n19019), .B(n19023), .Z(n19021) );
  XOR U18661 ( .A(n19024), .B(n19025), .Z(n18982) );
  NOR U18662 ( .A(n19026), .B(n19027), .Z(n19025) );
  XNOR U18663 ( .A(n19024), .B(n19028), .Z(n19026) );
  XNOR U18664 ( .A(n18927), .B(n18985), .Z(n18987) );
  XNOR U18665 ( .A(n19029), .B(n19030), .Z(n18927) );
  AND U18666 ( .A(n193), .B(n18934), .Z(n19030) );
  XOR U18667 ( .A(n19029), .B(n18932), .Z(n18934) );
  AND U18668 ( .A(n18935), .B(n18938), .Z(n18985) );
  XOR U18669 ( .A(n19031), .B(n19012), .Z(n18938) );
  XNOR U18670 ( .A(p_input[2048]), .B(p_input[224]), .Z(n19012) );
  XOR U18671 ( .A(n19000), .B(n18999), .Z(n19031) );
  XNOR U18672 ( .A(n19032), .B(n19006), .Z(n18999) );
  XNOR U18673 ( .A(n18995), .B(n18994), .Z(n19006) );
  XOR U18674 ( .A(n19033), .B(n18991), .Z(n18994) );
  XNOR U18675 ( .A(n16904), .B(p_input[234]), .Z(n18991) );
  XNOR U18676 ( .A(p_input[2059]), .B(p_input[235]), .Z(n19033) );
  XOR U18677 ( .A(p_input[2060]), .B(p_input[236]), .Z(n18995) );
  XNOR U18678 ( .A(n19005), .B(n18996), .Z(n19032) );
  XNOR U18679 ( .A(n17068), .B(p_input[225]), .Z(n18996) );
  XOR U18680 ( .A(n19034), .B(n19011), .Z(n19005) );
  XNOR U18681 ( .A(p_input[2063]), .B(p_input[239]), .Z(n19011) );
  XOR U18682 ( .A(n19002), .B(n19010), .Z(n19034) );
  XOR U18683 ( .A(n19035), .B(n19007), .Z(n19010) );
  XOR U18684 ( .A(p_input[2061]), .B(p_input[237]), .Z(n19007) );
  XNOR U18685 ( .A(p_input[2062]), .B(p_input[238]), .Z(n19035) );
  XNOR U18686 ( .A(n16738), .B(p_input[233]), .Z(n19002) );
  XNOR U18687 ( .A(n19018), .B(n19017), .Z(n19000) );
  XNOR U18688 ( .A(n19036), .B(n19023), .Z(n19017) );
  XOR U18689 ( .A(p_input[2056]), .B(p_input[232]), .Z(n19023) );
  XOR U18690 ( .A(n19014), .B(n19022), .Z(n19036) );
  XOR U18691 ( .A(n19037), .B(n19019), .Z(n19022) );
  XOR U18692 ( .A(p_input[2054]), .B(p_input[230]), .Z(n19019) );
  XNOR U18693 ( .A(p_input[2055]), .B(p_input[231]), .Z(n19037) );
  XNOR U18694 ( .A(n16741), .B(p_input[226]), .Z(n19014) );
  XNOR U18695 ( .A(n19028), .B(n19027), .Z(n19018) );
  XOR U18696 ( .A(n19038), .B(n19024), .Z(n19027) );
  XOR U18697 ( .A(p_input[2051]), .B(p_input[227]), .Z(n19024) );
  XNOR U18698 ( .A(p_input[2052]), .B(p_input[228]), .Z(n19038) );
  XOR U18699 ( .A(p_input[2053]), .B(p_input[229]), .Z(n19028) );
  XNOR U18700 ( .A(n19039), .B(n19040), .Z(n18935) );
  AND U18701 ( .A(n193), .B(n19041), .Z(n19040) );
  XNOR U18702 ( .A(n19042), .B(n19043), .Z(n193) );
  AND U18703 ( .A(n19044), .B(n19045), .Z(n19043) );
  XOR U18704 ( .A(n19042), .B(n18945), .Z(n19045) );
  XNOR U18705 ( .A(n19042), .B(n18899), .Z(n19044) );
  XOR U18706 ( .A(n19046), .B(n19047), .Z(n19042) );
  AND U18707 ( .A(n19048), .B(n19049), .Z(n19047) );
  XOR U18708 ( .A(n19046), .B(n18909), .Z(n19048) );
  XOR U18709 ( .A(n19050), .B(n19051), .Z(n18888) );
  AND U18710 ( .A(n197), .B(n19041), .Z(n19051) );
  XNOR U18711 ( .A(n19039), .B(n19050), .Z(n19041) );
  XNOR U18712 ( .A(n19052), .B(n19053), .Z(n197) );
  AND U18713 ( .A(n19054), .B(n19055), .Z(n19053) );
  XNOR U18714 ( .A(n19056), .B(n19052), .Z(n19055) );
  IV U18715 ( .A(n18945), .Z(n19056) );
  XNOR U18716 ( .A(n19057), .B(n19058), .Z(n18945) );
  AND U18717 ( .A(n200), .B(n19059), .Z(n19058) );
  XNOR U18718 ( .A(n19057), .B(n19060), .Z(n19059) );
  XNOR U18719 ( .A(n18899), .B(n19052), .Z(n19054) );
  XOR U18720 ( .A(n19061), .B(n19062), .Z(n18899) );
  AND U18721 ( .A(n208), .B(n19063), .Z(n19062) );
  XOR U18722 ( .A(n19046), .B(n19064), .Z(n19052) );
  AND U18723 ( .A(n19065), .B(n19049), .Z(n19064) );
  XNOR U18724 ( .A(n18958), .B(n19046), .Z(n19049) );
  XNOR U18725 ( .A(n19066), .B(n19067), .Z(n18958) );
  AND U18726 ( .A(n200), .B(n19068), .Z(n19067) );
  XOR U18727 ( .A(n19069), .B(n19066), .Z(n19068) );
  XNOR U18728 ( .A(n19070), .B(n19046), .Z(n19065) );
  IV U18729 ( .A(n18909), .Z(n19070) );
  XOR U18730 ( .A(n19071), .B(n19072), .Z(n18909) );
  AND U18731 ( .A(n208), .B(n19073), .Z(n19072) );
  XOR U18732 ( .A(n19074), .B(n19075), .Z(n19046) );
  AND U18733 ( .A(n19076), .B(n19077), .Z(n19075) );
  XNOR U18734 ( .A(n18983), .B(n19074), .Z(n19077) );
  XNOR U18735 ( .A(n19078), .B(n19079), .Z(n18983) );
  AND U18736 ( .A(n200), .B(n19080), .Z(n19079) );
  XNOR U18737 ( .A(n19081), .B(n19078), .Z(n19080) );
  XOR U18738 ( .A(n19074), .B(n18920), .Z(n19076) );
  XOR U18739 ( .A(n19082), .B(n19083), .Z(n18920) );
  AND U18740 ( .A(n208), .B(n19084), .Z(n19083) );
  XOR U18741 ( .A(n19085), .B(n19086), .Z(n19074) );
  AND U18742 ( .A(n19087), .B(n19088), .Z(n19086) );
  XNOR U18743 ( .A(n19085), .B(n19029), .Z(n19088) );
  XNOR U18744 ( .A(n19089), .B(n19090), .Z(n19029) );
  AND U18745 ( .A(n200), .B(n19091), .Z(n19090) );
  XOR U18746 ( .A(n19092), .B(n19089), .Z(n19091) );
  XNOR U18747 ( .A(n19093), .B(n19085), .Z(n19087) );
  IV U18748 ( .A(n18932), .Z(n19093) );
  XOR U18749 ( .A(n19094), .B(n19095), .Z(n18932) );
  AND U18750 ( .A(n208), .B(n19096), .Z(n19095) );
  AND U18751 ( .A(n19050), .B(n19039), .Z(n19085) );
  XNOR U18752 ( .A(n19097), .B(n19098), .Z(n19039) );
  AND U18753 ( .A(n200), .B(n19099), .Z(n19098) );
  XNOR U18754 ( .A(n19100), .B(n19097), .Z(n19099) );
  XNOR U18755 ( .A(n19101), .B(n19102), .Z(n200) );
  AND U18756 ( .A(n19103), .B(n19104), .Z(n19102) );
  XOR U18757 ( .A(n19060), .B(n19101), .Z(n19104) );
  AND U18758 ( .A(n19105), .B(n19106), .Z(n19060) );
  XOR U18759 ( .A(n19101), .B(n19057), .Z(n19103) );
  XNOR U18760 ( .A(n19107), .B(n19108), .Z(n19057) );
  AND U18761 ( .A(n204), .B(n19063), .Z(n19108) );
  XOR U18762 ( .A(n19061), .B(n19107), .Z(n19063) );
  XOR U18763 ( .A(n19109), .B(n19110), .Z(n19101) );
  AND U18764 ( .A(n19111), .B(n19112), .Z(n19110) );
  XNOR U18765 ( .A(n19109), .B(n19105), .Z(n19112) );
  IV U18766 ( .A(n19069), .Z(n19105) );
  XOR U18767 ( .A(n19113), .B(n19114), .Z(n19069) );
  XOR U18768 ( .A(n19115), .B(n19106), .Z(n19114) );
  AND U18769 ( .A(n19081), .B(n19116), .Z(n19106) );
  AND U18770 ( .A(n19117), .B(n19118), .Z(n19115) );
  XOR U18771 ( .A(n19119), .B(n19113), .Z(n19117) );
  XNOR U18772 ( .A(n19066), .B(n19109), .Z(n19111) );
  XNOR U18773 ( .A(n19120), .B(n19121), .Z(n19066) );
  AND U18774 ( .A(n204), .B(n19073), .Z(n19121) );
  XOR U18775 ( .A(n19120), .B(n19071), .Z(n19073) );
  XOR U18776 ( .A(n19122), .B(n19123), .Z(n19109) );
  AND U18777 ( .A(n19124), .B(n19125), .Z(n19123) );
  XNOR U18778 ( .A(n19122), .B(n19081), .Z(n19125) );
  XOR U18779 ( .A(n19126), .B(n19118), .Z(n19081) );
  XNOR U18780 ( .A(n19127), .B(n19113), .Z(n19118) );
  XOR U18781 ( .A(n19128), .B(n19129), .Z(n19113) );
  AND U18782 ( .A(n19130), .B(n19131), .Z(n19129) );
  XOR U18783 ( .A(n19132), .B(n19128), .Z(n19130) );
  XNOR U18784 ( .A(n19133), .B(n19134), .Z(n19127) );
  AND U18785 ( .A(n19135), .B(n19136), .Z(n19134) );
  XOR U18786 ( .A(n19133), .B(n19137), .Z(n19135) );
  XNOR U18787 ( .A(n19119), .B(n19116), .Z(n19126) );
  AND U18788 ( .A(n19138), .B(n19139), .Z(n19116) );
  XOR U18789 ( .A(n19140), .B(n19141), .Z(n19119) );
  AND U18790 ( .A(n19142), .B(n19143), .Z(n19141) );
  XOR U18791 ( .A(n19140), .B(n19144), .Z(n19142) );
  XNOR U18792 ( .A(n19078), .B(n19122), .Z(n19124) );
  XNOR U18793 ( .A(n19145), .B(n19146), .Z(n19078) );
  AND U18794 ( .A(n204), .B(n19084), .Z(n19146) );
  XOR U18795 ( .A(n19145), .B(n19082), .Z(n19084) );
  XOR U18796 ( .A(n19147), .B(n19148), .Z(n19122) );
  AND U18797 ( .A(n19149), .B(n19150), .Z(n19148) );
  XNOR U18798 ( .A(n19147), .B(n19138), .Z(n19150) );
  IV U18799 ( .A(n19092), .Z(n19138) );
  XNOR U18800 ( .A(n19151), .B(n19131), .Z(n19092) );
  XNOR U18801 ( .A(n19152), .B(n19137), .Z(n19131) );
  XOR U18802 ( .A(n19153), .B(n19154), .Z(n19137) );
  NOR U18803 ( .A(n19155), .B(n19156), .Z(n19154) );
  XNOR U18804 ( .A(n19153), .B(n19157), .Z(n19155) );
  XNOR U18805 ( .A(n19136), .B(n19128), .Z(n19152) );
  XOR U18806 ( .A(n19158), .B(n19159), .Z(n19128) );
  AND U18807 ( .A(n19160), .B(n19161), .Z(n19159) );
  XNOR U18808 ( .A(n19158), .B(n19162), .Z(n19160) );
  XNOR U18809 ( .A(n19163), .B(n19133), .Z(n19136) );
  XOR U18810 ( .A(n19164), .B(n19165), .Z(n19133) );
  AND U18811 ( .A(n19166), .B(n19167), .Z(n19165) );
  XOR U18812 ( .A(n19164), .B(n19168), .Z(n19166) );
  XNOR U18813 ( .A(n19169), .B(n19170), .Z(n19163) );
  NOR U18814 ( .A(n19171), .B(n19172), .Z(n19170) );
  XOR U18815 ( .A(n19169), .B(n19173), .Z(n19171) );
  XNOR U18816 ( .A(n19132), .B(n19139), .Z(n19151) );
  NOR U18817 ( .A(n19100), .B(n19174), .Z(n19139) );
  XOR U18818 ( .A(n19144), .B(n19143), .Z(n19132) );
  XNOR U18819 ( .A(n19175), .B(n19140), .Z(n19143) );
  XOR U18820 ( .A(n19176), .B(n19177), .Z(n19140) );
  AND U18821 ( .A(n19178), .B(n19179), .Z(n19177) );
  XOR U18822 ( .A(n19176), .B(n19180), .Z(n19178) );
  XNOR U18823 ( .A(n19181), .B(n19182), .Z(n19175) );
  NOR U18824 ( .A(n19183), .B(n19184), .Z(n19182) );
  XNOR U18825 ( .A(n19181), .B(n19185), .Z(n19183) );
  XOR U18826 ( .A(n19186), .B(n19187), .Z(n19144) );
  NOR U18827 ( .A(n19188), .B(n19189), .Z(n19187) );
  XNOR U18828 ( .A(n19186), .B(n19190), .Z(n19188) );
  XNOR U18829 ( .A(n19089), .B(n19147), .Z(n19149) );
  XNOR U18830 ( .A(n19191), .B(n19192), .Z(n19089) );
  AND U18831 ( .A(n204), .B(n19096), .Z(n19192) );
  XOR U18832 ( .A(n19191), .B(n19094), .Z(n19096) );
  AND U18833 ( .A(n19097), .B(n19100), .Z(n19147) );
  XOR U18834 ( .A(n19193), .B(n19174), .Z(n19100) );
  XNOR U18835 ( .A(p_input[2048]), .B(p_input[240]), .Z(n19174) );
  XOR U18836 ( .A(n19162), .B(n19161), .Z(n19193) );
  XNOR U18837 ( .A(n19194), .B(n19168), .Z(n19161) );
  XNOR U18838 ( .A(n19157), .B(n19156), .Z(n19168) );
  XOR U18839 ( .A(n19195), .B(n19153), .Z(n19156) );
  XNOR U18840 ( .A(n16904), .B(p_input[250]), .Z(n19153) );
  XNOR U18841 ( .A(p_input[2059]), .B(p_input[251]), .Z(n19195) );
  XOR U18842 ( .A(p_input[2060]), .B(p_input[252]), .Z(n19157) );
  XNOR U18843 ( .A(n19167), .B(n19158), .Z(n19194) );
  XNOR U18844 ( .A(n17068), .B(p_input[241]), .Z(n19158) );
  XOR U18845 ( .A(n19196), .B(n19173), .Z(n19167) );
  XNOR U18846 ( .A(p_input[2063]), .B(p_input[255]), .Z(n19173) );
  XOR U18847 ( .A(n19164), .B(n19172), .Z(n19196) );
  XOR U18848 ( .A(n19197), .B(n19169), .Z(n19172) );
  XOR U18849 ( .A(p_input[2061]), .B(p_input[253]), .Z(n19169) );
  XNOR U18850 ( .A(p_input[2062]), .B(p_input[254]), .Z(n19197) );
  XNOR U18851 ( .A(n16738), .B(p_input[249]), .Z(n19164) );
  XNOR U18852 ( .A(n19180), .B(n19179), .Z(n19162) );
  XNOR U18853 ( .A(n19198), .B(n19185), .Z(n19179) );
  XOR U18854 ( .A(p_input[2056]), .B(p_input[248]), .Z(n19185) );
  XOR U18855 ( .A(n19176), .B(n19184), .Z(n19198) );
  XOR U18856 ( .A(n19199), .B(n19181), .Z(n19184) );
  XOR U18857 ( .A(p_input[2054]), .B(p_input[246]), .Z(n19181) );
  XNOR U18858 ( .A(p_input[2055]), .B(p_input[247]), .Z(n19199) );
  XNOR U18859 ( .A(n16741), .B(p_input[242]), .Z(n19176) );
  XNOR U18860 ( .A(n19190), .B(n19189), .Z(n19180) );
  XOR U18861 ( .A(n19200), .B(n19186), .Z(n19189) );
  XOR U18862 ( .A(p_input[2051]), .B(p_input[243]), .Z(n19186) );
  XNOR U18863 ( .A(p_input[2052]), .B(p_input[244]), .Z(n19200) );
  XOR U18864 ( .A(p_input[2053]), .B(p_input[245]), .Z(n19190) );
  XNOR U18865 ( .A(n19201), .B(n19202), .Z(n19097) );
  AND U18866 ( .A(n204), .B(n19203), .Z(n19202) );
  XNOR U18867 ( .A(n19204), .B(n19205), .Z(n204) );
  AND U18868 ( .A(n19206), .B(n19207), .Z(n19205) );
  XOR U18869 ( .A(n19204), .B(n19107), .Z(n19207) );
  XNOR U18870 ( .A(n19204), .B(n19061), .Z(n19206) );
  XOR U18871 ( .A(n19208), .B(n19209), .Z(n19204) );
  AND U18872 ( .A(n19210), .B(n19211), .Z(n19209) );
  XOR U18873 ( .A(n19208), .B(n19071), .Z(n19210) );
  XOR U18874 ( .A(n19212), .B(n19213), .Z(n19050) );
  AND U18875 ( .A(n208), .B(n19203), .Z(n19213) );
  XNOR U18876 ( .A(n19201), .B(n19212), .Z(n19203) );
  XNOR U18877 ( .A(n19214), .B(n19215), .Z(n208) );
  AND U18878 ( .A(n19216), .B(n19217), .Z(n19215) );
  XNOR U18879 ( .A(n19218), .B(n19214), .Z(n19217) );
  IV U18880 ( .A(n19107), .Z(n19218) );
  XNOR U18881 ( .A(n19219), .B(n19220), .Z(n19107) );
  AND U18882 ( .A(n211), .B(n19221), .Z(n19220) );
  XNOR U18883 ( .A(n19219), .B(n19222), .Z(n19221) );
  XNOR U18884 ( .A(n19061), .B(n19214), .Z(n19216) );
  XOR U18885 ( .A(n19223), .B(n19224), .Z(n19061) );
  AND U18886 ( .A(n219), .B(n19225), .Z(n19224) );
  XOR U18887 ( .A(n19208), .B(n19226), .Z(n19214) );
  AND U18888 ( .A(n19227), .B(n19211), .Z(n19226) );
  XNOR U18889 ( .A(n19120), .B(n19208), .Z(n19211) );
  XNOR U18890 ( .A(n19228), .B(n19229), .Z(n19120) );
  AND U18891 ( .A(n211), .B(n19230), .Z(n19229) );
  XOR U18892 ( .A(n19231), .B(n19228), .Z(n19230) );
  XNOR U18893 ( .A(n19232), .B(n19208), .Z(n19227) );
  IV U18894 ( .A(n19071), .Z(n19232) );
  XOR U18895 ( .A(n19233), .B(n19234), .Z(n19071) );
  AND U18896 ( .A(n219), .B(n19235), .Z(n19234) );
  XOR U18897 ( .A(n19236), .B(n19237), .Z(n19208) );
  AND U18898 ( .A(n19238), .B(n19239), .Z(n19237) );
  XNOR U18899 ( .A(n19145), .B(n19236), .Z(n19239) );
  XNOR U18900 ( .A(n19240), .B(n19241), .Z(n19145) );
  AND U18901 ( .A(n211), .B(n19242), .Z(n19241) );
  XNOR U18902 ( .A(n19243), .B(n19240), .Z(n19242) );
  XOR U18903 ( .A(n19236), .B(n19082), .Z(n19238) );
  XOR U18904 ( .A(n19244), .B(n19245), .Z(n19082) );
  AND U18905 ( .A(n219), .B(n19246), .Z(n19245) );
  XOR U18906 ( .A(n19247), .B(n19248), .Z(n19236) );
  AND U18907 ( .A(n19249), .B(n19250), .Z(n19248) );
  XNOR U18908 ( .A(n19247), .B(n19191), .Z(n19250) );
  XNOR U18909 ( .A(n19251), .B(n19252), .Z(n19191) );
  AND U18910 ( .A(n211), .B(n19253), .Z(n19252) );
  XOR U18911 ( .A(n19254), .B(n19251), .Z(n19253) );
  XNOR U18912 ( .A(n19255), .B(n19247), .Z(n19249) );
  IV U18913 ( .A(n19094), .Z(n19255) );
  XOR U18914 ( .A(n19256), .B(n19257), .Z(n19094) );
  AND U18915 ( .A(n219), .B(n19258), .Z(n19257) );
  AND U18916 ( .A(n19212), .B(n19201), .Z(n19247) );
  XNOR U18917 ( .A(n19259), .B(n19260), .Z(n19201) );
  AND U18918 ( .A(n211), .B(n19261), .Z(n19260) );
  XNOR U18919 ( .A(n19262), .B(n19259), .Z(n19261) );
  XNOR U18920 ( .A(n19263), .B(n19264), .Z(n211) );
  AND U18921 ( .A(n19265), .B(n19266), .Z(n19264) );
  XOR U18922 ( .A(n19222), .B(n19263), .Z(n19266) );
  AND U18923 ( .A(n19267), .B(n19268), .Z(n19222) );
  XOR U18924 ( .A(n19263), .B(n19219), .Z(n19265) );
  XNOR U18925 ( .A(n19269), .B(n19270), .Z(n19219) );
  AND U18926 ( .A(n215), .B(n19225), .Z(n19270) );
  XOR U18927 ( .A(n19223), .B(n19269), .Z(n19225) );
  XOR U18928 ( .A(n19271), .B(n19272), .Z(n19263) );
  AND U18929 ( .A(n19273), .B(n19274), .Z(n19272) );
  XNOR U18930 ( .A(n19271), .B(n19267), .Z(n19274) );
  IV U18931 ( .A(n19231), .Z(n19267) );
  XOR U18932 ( .A(n19275), .B(n19276), .Z(n19231) );
  XOR U18933 ( .A(n19277), .B(n19268), .Z(n19276) );
  AND U18934 ( .A(n19243), .B(n19278), .Z(n19268) );
  AND U18935 ( .A(n19279), .B(n19280), .Z(n19277) );
  XOR U18936 ( .A(n19281), .B(n19275), .Z(n19279) );
  XNOR U18937 ( .A(n19228), .B(n19271), .Z(n19273) );
  XNOR U18938 ( .A(n19282), .B(n19283), .Z(n19228) );
  AND U18939 ( .A(n215), .B(n19235), .Z(n19283) );
  XOR U18940 ( .A(n19282), .B(n19233), .Z(n19235) );
  XOR U18941 ( .A(n19284), .B(n19285), .Z(n19271) );
  AND U18942 ( .A(n19286), .B(n19287), .Z(n19285) );
  XNOR U18943 ( .A(n19284), .B(n19243), .Z(n19287) );
  XOR U18944 ( .A(n19288), .B(n19280), .Z(n19243) );
  XNOR U18945 ( .A(n19289), .B(n19275), .Z(n19280) );
  XOR U18946 ( .A(n19290), .B(n19291), .Z(n19275) );
  AND U18947 ( .A(n19292), .B(n19293), .Z(n19291) );
  XOR U18948 ( .A(n19294), .B(n19290), .Z(n19292) );
  XNOR U18949 ( .A(n19295), .B(n19296), .Z(n19289) );
  AND U18950 ( .A(n19297), .B(n19298), .Z(n19296) );
  XOR U18951 ( .A(n19295), .B(n19299), .Z(n19297) );
  XNOR U18952 ( .A(n19281), .B(n19278), .Z(n19288) );
  AND U18953 ( .A(n19300), .B(n19301), .Z(n19278) );
  XOR U18954 ( .A(n19302), .B(n19303), .Z(n19281) );
  AND U18955 ( .A(n19304), .B(n19305), .Z(n19303) );
  XOR U18956 ( .A(n19302), .B(n19306), .Z(n19304) );
  XNOR U18957 ( .A(n19240), .B(n19284), .Z(n19286) );
  XNOR U18958 ( .A(n19307), .B(n19308), .Z(n19240) );
  AND U18959 ( .A(n215), .B(n19246), .Z(n19308) );
  XOR U18960 ( .A(n19307), .B(n19244), .Z(n19246) );
  XOR U18961 ( .A(n19309), .B(n19310), .Z(n19284) );
  AND U18962 ( .A(n19311), .B(n19312), .Z(n19310) );
  XNOR U18963 ( .A(n19309), .B(n19300), .Z(n19312) );
  IV U18964 ( .A(n19254), .Z(n19300) );
  XNOR U18965 ( .A(n19313), .B(n19293), .Z(n19254) );
  XNOR U18966 ( .A(n19314), .B(n19299), .Z(n19293) );
  XOR U18967 ( .A(n19315), .B(n19316), .Z(n19299) );
  NOR U18968 ( .A(n19317), .B(n19318), .Z(n19316) );
  XNOR U18969 ( .A(n19315), .B(n19319), .Z(n19317) );
  XNOR U18970 ( .A(n19298), .B(n19290), .Z(n19314) );
  XOR U18971 ( .A(n19320), .B(n19321), .Z(n19290) );
  AND U18972 ( .A(n19322), .B(n19323), .Z(n19321) );
  XNOR U18973 ( .A(n19320), .B(n19324), .Z(n19322) );
  XNOR U18974 ( .A(n19325), .B(n19295), .Z(n19298) );
  XOR U18975 ( .A(n19326), .B(n19327), .Z(n19295) );
  AND U18976 ( .A(n19328), .B(n19329), .Z(n19327) );
  XOR U18977 ( .A(n19326), .B(n19330), .Z(n19328) );
  XNOR U18978 ( .A(n19331), .B(n19332), .Z(n19325) );
  NOR U18979 ( .A(n19333), .B(n19334), .Z(n19332) );
  XOR U18980 ( .A(n19331), .B(n19335), .Z(n19333) );
  XNOR U18981 ( .A(n19294), .B(n19301), .Z(n19313) );
  NOR U18982 ( .A(n19262), .B(n19336), .Z(n19301) );
  XOR U18983 ( .A(n19306), .B(n19305), .Z(n19294) );
  XNOR U18984 ( .A(n19337), .B(n19302), .Z(n19305) );
  XOR U18985 ( .A(n19338), .B(n19339), .Z(n19302) );
  AND U18986 ( .A(n19340), .B(n19341), .Z(n19339) );
  XOR U18987 ( .A(n19338), .B(n19342), .Z(n19340) );
  XNOR U18988 ( .A(n19343), .B(n19344), .Z(n19337) );
  NOR U18989 ( .A(n19345), .B(n19346), .Z(n19344) );
  XNOR U18990 ( .A(n19343), .B(n19347), .Z(n19345) );
  XOR U18991 ( .A(n19348), .B(n19349), .Z(n19306) );
  NOR U18992 ( .A(n19350), .B(n19351), .Z(n19349) );
  XNOR U18993 ( .A(n19348), .B(n19352), .Z(n19350) );
  XNOR U18994 ( .A(n19251), .B(n19309), .Z(n19311) );
  XNOR U18995 ( .A(n19353), .B(n19354), .Z(n19251) );
  AND U18996 ( .A(n215), .B(n19258), .Z(n19354) );
  XOR U18997 ( .A(n19353), .B(n19256), .Z(n19258) );
  AND U18998 ( .A(n19259), .B(n19262), .Z(n19309) );
  XOR U18999 ( .A(n19355), .B(n19336), .Z(n19262) );
  XNOR U19000 ( .A(p_input[2048]), .B(p_input[256]), .Z(n19336) );
  XOR U19001 ( .A(n19324), .B(n19323), .Z(n19355) );
  XNOR U19002 ( .A(n19356), .B(n19330), .Z(n19323) );
  XNOR U19003 ( .A(n19319), .B(n19318), .Z(n19330) );
  XOR U19004 ( .A(n19357), .B(n19315), .Z(n19318) );
  XNOR U19005 ( .A(n16904), .B(p_input[266]), .Z(n19315) );
  XNOR U19006 ( .A(p_input[2059]), .B(p_input[267]), .Z(n19357) );
  XOR U19007 ( .A(p_input[2060]), .B(p_input[268]), .Z(n19319) );
  XNOR U19008 ( .A(n19329), .B(n19320), .Z(n19356) );
  XNOR U19009 ( .A(n17068), .B(p_input[257]), .Z(n19320) );
  XOR U19010 ( .A(n19358), .B(n19335), .Z(n19329) );
  XNOR U19011 ( .A(p_input[2063]), .B(p_input[271]), .Z(n19335) );
  XOR U19012 ( .A(n19326), .B(n19334), .Z(n19358) );
  XOR U19013 ( .A(n19359), .B(n19331), .Z(n19334) );
  XOR U19014 ( .A(p_input[2061]), .B(p_input[269]), .Z(n19331) );
  XNOR U19015 ( .A(p_input[2062]), .B(p_input[270]), .Z(n19359) );
  XNOR U19016 ( .A(n16738), .B(p_input[265]), .Z(n19326) );
  XNOR U19017 ( .A(n19342), .B(n19341), .Z(n19324) );
  XNOR U19018 ( .A(n19360), .B(n19347), .Z(n19341) );
  XOR U19019 ( .A(p_input[2056]), .B(p_input[264]), .Z(n19347) );
  XOR U19020 ( .A(n19338), .B(n19346), .Z(n19360) );
  XOR U19021 ( .A(n19361), .B(n19343), .Z(n19346) );
  XOR U19022 ( .A(p_input[2054]), .B(p_input[262]), .Z(n19343) );
  XNOR U19023 ( .A(p_input[2055]), .B(p_input[263]), .Z(n19361) );
  XNOR U19024 ( .A(n16741), .B(p_input[258]), .Z(n19338) );
  XNOR U19025 ( .A(n19352), .B(n19351), .Z(n19342) );
  XOR U19026 ( .A(n19362), .B(n19348), .Z(n19351) );
  XOR U19027 ( .A(p_input[2051]), .B(p_input[259]), .Z(n19348) );
  XNOR U19028 ( .A(p_input[2052]), .B(p_input[260]), .Z(n19362) );
  XOR U19029 ( .A(p_input[2053]), .B(p_input[261]), .Z(n19352) );
  XNOR U19030 ( .A(n19363), .B(n19364), .Z(n19259) );
  AND U19031 ( .A(n215), .B(n19365), .Z(n19364) );
  XNOR U19032 ( .A(n19366), .B(n19367), .Z(n215) );
  AND U19033 ( .A(n19368), .B(n19369), .Z(n19367) );
  XOR U19034 ( .A(n19366), .B(n19269), .Z(n19369) );
  XNOR U19035 ( .A(n19366), .B(n19223), .Z(n19368) );
  XOR U19036 ( .A(n19370), .B(n19371), .Z(n19366) );
  AND U19037 ( .A(n19372), .B(n19373), .Z(n19371) );
  XOR U19038 ( .A(n19370), .B(n19233), .Z(n19372) );
  XOR U19039 ( .A(n19374), .B(n19375), .Z(n19212) );
  AND U19040 ( .A(n219), .B(n19365), .Z(n19375) );
  XNOR U19041 ( .A(n19363), .B(n19374), .Z(n19365) );
  XNOR U19042 ( .A(n19376), .B(n19377), .Z(n219) );
  AND U19043 ( .A(n19378), .B(n19379), .Z(n19377) );
  XNOR U19044 ( .A(n19380), .B(n19376), .Z(n19379) );
  IV U19045 ( .A(n19269), .Z(n19380) );
  XNOR U19046 ( .A(n19381), .B(n19382), .Z(n19269) );
  AND U19047 ( .A(n222), .B(n19383), .Z(n19382) );
  XNOR U19048 ( .A(n19381), .B(n19384), .Z(n19383) );
  XNOR U19049 ( .A(n19223), .B(n19376), .Z(n19378) );
  XOR U19050 ( .A(n19385), .B(n19386), .Z(n19223) );
  AND U19051 ( .A(n230), .B(n19387), .Z(n19386) );
  XOR U19052 ( .A(n19370), .B(n19388), .Z(n19376) );
  AND U19053 ( .A(n19389), .B(n19373), .Z(n19388) );
  XNOR U19054 ( .A(n19282), .B(n19370), .Z(n19373) );
  XNOR U19055 ( .A(n19390), .B(n19391), .Z(n19282) );
  AND U19056 ( .A(n222), .B(n19392), .Z(n19391) );
  XOR U19057 ( .A(n19393), .B(n19390), .Z(n19392) );
  XNOR U19058 ( .A(n19394), .B(n19370), .Z(n19389) );
  IV U19059 ( .A(n19233), .Z(n19394) );
  XOR U19060 ( .A(n19395), .B(n19396), .Z(n19233) );
  AND U19061 ( .A(n230), .B(n19397), .Z(n19396) );
  XOR U19062 ( .A(n19398), .B(n19399), .Z(n19370) );
  AND U19063 ( .A(n19400), .B(n19401), .Z(n19399) );
  XNOR U19064 ( .A(n19307), .B(n19398), .Z(n19401) );
  XNOR U19065 ( .A(n19402), .B(n19403), .Z(n19307) );
  AND U19066 ( .A(n222), .B(n19404), .Z(n19403) );
  XNOR U19067 ( .A(n19405), .B(n19402), .Z(n19404) );
  XOR U19068 ( .A(n19398), .B(n19244), .Z(n19400) );
  XOR U19069 ( .A(n19406), .B(n19407), .Z(n19244) );
  AND U19070 ( .A(n230), .B(n19408), .Z(n19407) );
  XOR U19071 ( .A(n19409), .B(n19410), .Z(n19398) );
  AND U19072 ( .A(n19411), .B(n19412), .Z(n19410) );
  XNOR U19073 ( .A(n19409), .B(n19353), .Z(n19412) );
  XNOR U19074 ( .A(n19413), .B(n19414), .Z(n19353) );
  AND U19075 ( .A(n222), .B(n19415), .Z(n19414) );
  XOR U19076 ( .A(n19416), .B(n19413), .Z(n19415) );
  XNOR U19077 ( .A(n19417), .B(n19409), .Z(n19411) );
  IV U19078 ( .A(n19256), .Z(n19417) );
  XOR U19079 ( .A(n19418), .B(n19419), .Z(n19256) );
  AND U19080 ( .A(n230), .B(n19420), .Z(n19419) );
  AND U19081 ( .A(n19374), .B(n19363), .Z(n19409) );
  XNOR U19082 ( .A(n19421), .B(n19422), .Z(n19363) );
  AND U19083 ( .A(n222), .B(n19423), .Z(n19422) );
  XNOR U19084 ( .A(n19424), .B(n19421), .Z(n19423) );
  XNOR U19085 ( .A(n19425), .B(n19426), .Z(n222) );
  AND U19086 ( .A(n19427), .B(n19428), .Z(n19426) );
  XOR U19087 ( .A(n19384), .B(n19425), .Z(n19428) );
  AND U19088 ( .A(n19429), .B(n19430), .Z(n19384) );
  XOR U19089 ( .A(n19425), .B(n19381), .Z(n19427) );
  XNOR U19090 ( .A(n19431), .B(n19432), .Z(n19381) );
  AND U19091 ( .A(n226), .B(n19387), .Z(n19432) );
  XOR U19092 ( .A(n19385), .B(n19431), .Z(n19387) );
  XOR U19093 ( .A(n19433), .B(n19434), .Z(n19425) );
  AND U19094 ( .A(n19435), .B(n19436), .Z(n19434) );
  XNOR U19095 ( .A(n19433), .B(n19429), .Z(n19436) );
  IV U19096 ( .A(n19393), .Z(n19429) );
  XOR U19097 ( .A(n19437), .B(n19438), .Z(n19393) );
  XOR U19098 ( .A(n19439), .B(n19430), .Z(n19438) );
  AND U19099 ( .A(n19405), .B(n19440), .Z(n19430) );
  AND U19100 ( .A(n19441), .B(n19442), .Z(n19439) );
  XOR U19101 ( .A(n19443), .B(n19437), .Z(n19441) );
  XNOR U19102 ( .A(n19390), .B(n19433), .Z(n19435) );
  XNOR U19103 ( .A(n19444), .B(n19445), .Z(n19390) );
  AND U19104 ( .A(n226), .B(n19397), .Z(n19445) );
  XOR U19105 ( .A(n19444), .B(n19395), .Z(n19397) );
  XOR U19106 ( .A(n19446), .B(n19447), .Z(n19433) );
  AND U19107 ( .A(n19448), .B(n19449), .Z(n19447) );
  XNOR U19108 ( .A(n19446), .B(n19405), .Z(n19449) );
  XOR U19109 ( .A(n19450), .B(n19442), .Z(n19405) );
  XNOR U19110 ( .A(n19451), .B(n19437), .Z(n19442) );
  XOR U19111 ( .A(n19452), .B(n19453), .Z(n19437) );
  AND U19112 ( .A(n19454), .B(n19455), .Z(n19453) );
  XOR U19113 ( .A(n19456), .B(n19452), .Z(n19454) );
  XNOR U19114 ( .A(n19457), .B(n19458), .Z(n19451) );
  AND U19115 ( .A(n19459), .B(n19460), .Z(n19458) );
  XOR U19116 ( .A(n19457), .B(n19461), .Z(n19459) );
  XNOR U19117 ( .A(n19443), .B(n19440), .Z(n19450) );
  AND U19118 ( .A(n19462), .B(n19463), .Z(n19440) );
  XOR U19119 ( .A(n19464), .B(n19465), .Z(n19443) );
  AND U19120 ( .A(n19466), .B(n19467), .Z(n19465) );
  XOR U19121 ( .A(n19464), .B(n19468), .Z(n19466) );
  XNOR U19122 ( .A(n19402), .B(n19446), .Z(n19448) );
  XNOR U19123 ( .A(n19469), .B(n19470), .Z(n19402) );
  AND U19124 ( .A(n226), .B(n19408), .Z(n19470) );
  XOR U19125 ( .A(n19469), .B(n19406), .Z(n19408) );
  XOR U19126 ( .A(n19471), .B(n19472), .Z(n19446) );
  AND U19127 ( .A(n19473), .B(n19474), .Z(n19472) );
  XNOR U19128 ( .A(n19471), .B(n19462), .Z(n19474) );
  IV U19129 ( .A(n19416), .Z(n19462) );
  XNOR U19130 ( .A(n19475), .B(n19455), .Z(n19416) );
  XNOR U19131 ( .A(n19476), .B(n19461), .Z(n19455) );
  XOR U19132 ( .A(n19477), .B(n19478), .Z(n19461) );
  NOR U19133 ( .A(n19479), .B(n19480), .Z(n19478) );
  XNOR U19134 ( .A(n19477), .B(n19481), .Z(n19479) );
  XNOR U19135 ( .A(n19460), .B(n19452), .Z(n19476) );
  XOR U19136 ( .A(n19482), .B(n19483), .Z(n19452) );
  AND U19137 ( .A(n19484), .B(n19485), .Z(n19483) );
  XNOR U19138 ( .A(n19482), .B(n19486), .Z(n19484) );
  XNOR U19139 ( .A(n19487), .B(n19457), .Z(n19460) );
  XOR U19140 ( .A(n19488), .B(n19489), .Z(n19457) );
  AND U19141 ( .A(n19490), .B(n19491), .Z(n19489) );
  XOR U19142 ( .A(n19488), .B(n19492), .Z(n19490) );
  XNOR U19143 ( .A(n19493), .B(n19494), .Z(n19487) );
  NOR U19144 ( .A(n19495), .B(n19496), .Z(n19494) );
  XOR U19145 ( .A(n19493), .B(n19497), .Z(n19495) );
  XNOR U19146 ( .A(n19456), .B(n19463), .Z(n19475) );
  NOR U19147 ( .A(n19424), .B(n19498), .Z(n19463) );
  XOR U19148 ( .A(n19468), .B(n19467), .Z(n19456) );
  XNOR U19149 ( .A(n19499), .B(n19464), .Z(n19467) );
  XOR U19150 ( .A(n19500), .B(n19501), .Z(n19464) );
  AND U19151 ( .A(n19502), .B(n19503), .Z(n19501) );
  XOR U19152 ( .A(n19500), .B(n19504), .Z(n19502) );
  XNOR U19153 ( .A(n19505), .B(n19506), .Z(n19499) );
  NOR U19154 ( .A(n19507), .B(n19508), .Z(n19506) );
  XNOR U19155 ( .A(n19505), .B(n19509), .Z(n19507) );
  XOR U19156 ( .A(n19510), .B(n19511), .Z(n19468) );
  NOR U19157 ( .A(n19512), .B(n19513), .Z(n19511) );
  XNOR U19158 ( .A(n19510), .B(n19514), .Z(n19512) );
  XNOR U19159 ( .A(n19413), .B(n19471), .Z(n19473) );
  XNOR U19160 ( .A(n19515), .B(n19516), .Z(n19413) );
  AND U19161 ( .A(n226), .B(n19420), .Z(n19516) );
  XOR U19162 ( .A(n19515), .B(n19418), .Z(n19420) );
  AND U19163 ( .A(n19421), .B(n19424), .Z(n19471) );
  XOR U19164 ( .A(n19517), .B(n19498), .Z(n19424) );
  XNOR U19165 ( .A(p_input[2048]), .B(p_input[272]), .Z(n19498) );
  XOR U19166 ( .A(n19486), .B(n19485), .Z(n19517) );
  XNOR U19167 ( .A(n19518), .B(n19492), .Z(n19485) );
  XNOR U19168 ( .A(n19481), .B(n19480), .Z(n19492) );
  XOR U19169 ( .A(n19519), .B(n19477), .Z(n19480) );
  XNOR U19170 ( .A(n16904), .B(p_input[282]), .Z(n19477) );
  XNOR U19171 ( .A(p_input[2059]), .B(p_input[283]), .Z(n19519) );
  XOR U19172 ( .A(p_input[2060]), .B(p_input[284]), .Z(n19481) );
  XNOR U19173 ( .A(n19491), .B(n19482), .Z(n19518) );
  XNOR U19174 ( .A(n17068), .B(p_input[273]), .Z(n19482) );
  XOR U19175 ( .A(n19520), .B(n19497), .Z(n19491) );
  XNOR U19176 ( .A(p_input[2063]), .B(p_input[287]), .Z(n19497) );
  XOR U19177 ( .A(n19488), .B(n19496), .Z(n19520) );
  XOR U19178 ( .A(n19521), .B(n19493), .Z(n19496) );
  XOR U19179 ( .A(p_input[2061]), .B(p_input[285]), .Z(n19493) );
  XNOR U19180 ( .A(p_input[2062]), .B(p_input[286]), .Z(n19521) );
  XNOR U19181 ( .A(n16738), .B(p_input[281]), .Z(n19488) );
  XNOR U19182 ( .A(n19504), .B(n19503), .Z(n19486) );
  XNOR U19183 ( .A(n19522), .B(n19509), .Z(n19503) );
  XOR U19184 ( .A(p_input[2056]), .B(p_input[280]), .Z(n19509) );
  XOR U19185 ( .A(n19500), .B(n19508), .Z(n19522) );
  XOR U19186 ( .A(n19523), .B(n19505), .Z(n19508) );
  XOR U19187 ( .A(p_input[2054]), .B(p_input[278]), .Z(n19505) );
  XNOR U19188 ( .A(p_input[2055]), .B(p_input[279]), .Z(n19523) );
  XNOR U19189 ( .A(n16741), .B(p_input[274]), .Z(n19500) );
  XNOR U19190 ( .A(n19514), .B(n19513), .Z(n19504) );
  XOR U19191 ( .A(n19524), .B(n19510), .Z(n19513) );
  XOR U19192 ( .A(p_input[2051]), .B(p_input[275]), .Z(n19510) );
  XNOR U19193 ( .A(p_input[2052]), .B(p_input[276]), .Z(n19524) );
  XOR U19194 ( .A(p_input[2053]), .B(p_input[277]), .Z(n19514) );
  XNOR U19195 ( .A(n19525), .B(n19526), .Z(n19421) );
  AND U19196 ( .A(n226), .B(n19527), .Z(n19526) );
  XNOR U19197 ( .A(n19528), .B(n19529), .Z(n226) );
  AND U19198 ( .A(n19530), .B(n19531), .Z(n19529) );
  XOR U19199 ( .A(n19528), .B(n19431), .Z(n19531) );
  XNOR U19200 ( .A(n19528), .B(n19385), .Z(n19530) );
  XOR U19201 ( .A(n19532), .B(n19533), .Z(n19528) );
  AND U19202 ( .A(n19534), .B(n19535), .Z(n19533) );
  XOR U19203 ( .A(n19532), .B(n19395), .Z(n19534) );
  XOR U19204 ( .A(n19536), .B(n19537), .Z(n19374) );
  AND U19205 ( .A(n230), .B(n19527), .Z(n19537) );
  XNOR U19206 ( .A(n19525), .B(n19536), .Z(n19527) );
  XNOR U19207 ( .A(n19538), .B(n19539), .Z(n230) );
  AND U19208 ( .A(n19540), .B(n19541), .Z(n19539) );
  XNOR U19209 ( .A(n19542), .B(n19538), .Z(n19541) );
  IV U19210 ( .A(n19431), .Z(n19542) );
  XNOR U19211 ( .A(n19543), .B(n19544), .Z(n19431) );
  AND U19212 ( .A(n233), .B(n19545), .Z(n19544) );
  XNOR U19213 ( .A(n19543), .B(n19546), .Z(n19545) );
  XNOR U19214 ( .A(n19385), .B(n19538), .Z(n19540) );
  XOR U19215 ( .A(n19547), .B(n19548), .Z(n19385) );
  AND U19216 ( .A(n241), .B(n19549), .Z(n19548) );
  XOR U19217 ( .A(n19532), .B(n19550), .Z(n19538) );
  AND U19218 ( .A(n19551), .B(n19535), .Z(n19550) );
  XNOR U19219 ( .A(n19444), .B(n19532), .Z(n19535) );
  XNOR U19220 ( .A(n19552), .B(n19553), .Z(n19444) );
  AND U19221 ( .A(n233), .B(n19554), .Z(n19553) );
  XOR U19222 ( .A(n19555), .B(n19552), .Z(n19554) );
  XNOR U19223 ( .A(n19556), .B(n19532), .Z(n19551) );
  IV U19224 ( .A(n19395), .Z(n19556) );
  XOR U19225 ( .A(n19557), .B(n19558), .Z(n19395) );
  AND U19226 ( .A(n241), .B(n19559), .Z(n19558) );
  XOR U19227 ( .A(n19560), .B(n19561), .Z(n19532) );
  AND U19228 ( .A(n19562), .B(n19563), .Z(n19561) );
  XNOR U19229 ( .A(n19469), .B(n19560), .Z(n19563) );
  XNOR U19230 ( .A(n19564), .B(n19565), .Z(n19469) );
  AND U19231 ( .A(n233), .B(n19566), .Z(n19565) );
  XNOR U19232 ( .A(n19567), .B(n19564), .Z(n19566) );
  XOR U19233 ( .A(n19560), .B(n19406), .Z(n19562) );
  XOR U19234 ( .A(n19568), .B(n19569), .Z(n19406) );
  AND U19235 ( .A(n241), .B(n19570), .Z(n19569) );
  XOR U19236 ( .A(n19571), .B(n19572), .Z(n19560) );
  AND U19237 ( .A(n19573), .B(n19574), .Z(n19572) );
  XNOR U19238 ( .A(n19571), .B(n19515), .Z(n19574) );
  XNOR U19239 ( .A(n19575), .B(n19576), .Z(n19515) );
  AND U19240 ( .A(n233), .B(n19577), .Z(n19576) );
  XOR U19241 ( .A(n19578), .B(n19575), .Z(n19577) );
  XNOR U19242 ( .A(n19579), .B(n19571), .Z(n19573) );
  IV U19243 ( .A(n19418), .Z(n19579) );
  XOR U19244 ( .A(n19580), .B(n19581), .Z(n19418) );
  AND U19245 ( .A(n241), .B(n19582), .Z(n19581) );
  AND U19246 ( .A(n19536), .B(n19525), .Z(n19571) );
  XNOR U19247 ( .A(n19583), .B(n19584), .Z(n19525) );
  AND U19248 ( .A(n233), .B(n19585), .Z(n19584) );
  XNOR U19249 ( .A(n19586), .B(n19583), .Z(n19585) );
  XNOR U19250 ( .A(n19587), .B(n19588), .Z(n233) );
  AND U19251 ( .A(n19589), .B(n19590), .Z(n19588) );
  XOR U19252 ( .A(n19546), .B(n19587), .Z(n19590) );
  AND U19253 ( .A(n19591), .B(n19592), .Z(n19546) );
  XOR U19254 ( .A(n19587), .B(n19543), .Z(n19589) );
  XNOR U19255 ( .A(n19593), .B(n19594), .Z(n19543) );
  AND U19256 ( .A(n237), .B(n19549), .Z(n19594) );
  XOR U19257 ( .A(n19547), .B(n19593), .Z(n19549) );
  XOR U19258 ( .A(n19595), .B(n19596), .Z(n19587) );
  AND U19259 ( .A(n19597), .B(n19598), .Z(n19596) );
  XNOR U19260 ( .A(n19595), .B(n19591), .Z(n19598) );
  IV U19261 ( .A(n19555), .Z(n19591) );
  XOR U19262 ( .A(n19599), .B(n19600), .Z(n19555) );
  XOR U19263 ( .A(n19601), .B(n19592), .Z(n19600) );
  AND U19264 ( .A(n19567), .B(n19602), .Z(n19592) );
  AND U19265 ( .A(n19603), .B(n19604), .Z(n19601) );
  XOR U19266 ( .A(n19605), .B(n19599), .Z(n19603) );
  XNOR U19267 ( .A(n19552), .B(n19595), .Z(n19597) );
  XNOR U19268 ( .A(n19606), .B(n19607), .Z(n19552) );
  AND U19269 ( .A(n237), .B(n19559), .Z(n19607) );
  XOR U19270 ( .A(n19606), .B(n19557), .Z(n19559) );
  XOR U19271 ( .A(n19608), .B(n19609), .Z(n19595) );
  AND U19272 ( .A(n19610), .B(n19611), .Z(n19609) );
  XNOR U19273 ( .A(n19608), .B(n19567), .Z(n19611) );
  XOR U19274 ( .A(n19612), .B(n19604), .Z(n19567) );
  XNOR U19275 ( .A(n19613), .B(n19599), .Z(n19604) );
  XOR U19276 ( .A(n19614), .B(n19615), .Z(n19599) );
  AND U19277 ( .A(n19616), .B(n19617), .Z(n19615) );
  XOR U19278 ( .A(n19618), .B(n19614), .Z(n19616) );
  XNOR U19279 ( .A(n19619), .B(n19620), .Z(n19613) );
  AND U19280 ( .A(n19621), .B(n19622), .Z(n19620) );
  XOR U19281 ( .A(n19619), .B(n19623), .Z(n19621) );
  XNOR U19282 ( .A(n19605), .B(n19602), .Z(n19612) );
  AND U19283 ( .A(n19624), .B(n19625), .Z(n19602) );
  XOR U19284 ( .A(n19626), .B(n19627), .Z(n19605) );
  AND U19285 ( .A(n19628), .B(n19629), .Z(n19627) );
  XOR U19286 ( .A(n19626), .B(n19630), .Z(n19628) );
  XNOR U19287 ( .A(n19564), .B(n19608), .Z(n19610) );
  XNOR U19288 ( .A(n19631), .B(n19632), .Z(n19564) );
  AND U19289 ( .A(n237), .B(n19570), .Z(n19632) );
  XOR U19290 ( .A(n19631), .B(n19568), .Z(n19570) );
  XOR U19291 ( .A(n19633), .B(n19634), .Z(n19608) );
  AND U19292 ( .A(n19635), .B(n19636), .Z(n19634) );
  XNOR U19293 ( .A(n19633), .B(n19624), .Z(n19636) );
  IV U19294 ( .A(n19578), .Z(n19624) );
  XNOR U19295 ( .A(n19637), .B(n19617), .Z(n19578) );
  XNOR U19296 ( .A(n19638), .B(n19623), .Z(n19617) );
  XOR U19297 ( .A(n19639), .B(n19640), .Z(n19623) );
  NOR U19298 ( .A(n19641), .B(n19642), .Z(n19640) );
  XNOR U19299 ( .A(n19639), .B(n19643), .Z(n19641) );
  XNOR U19300 ( .A(n19622), .B(n19614), .Z(n19638) );
  XOR U19301 ( .A(n19644), .B(n19645), .Z(n19614) );
  AND U19302 ( .A(n19646), .B(n19647), .Z(n19645) );
  XNOR U19303 ( .A(n19644), .B(n19648), .Z(n19646) );
  XNOR U19304 ( .A(n19649), .B(n19619), .Z(n19622) );
  XOR U19305 ( .A(n19650), .B(n19651), .Z(n19619) );
  AND U19306 ( .A(n19652), .B(n19653), .Z(n19651) );
  XOR U19307 ( .A(n19650), .B(n19654), .Z(n19652) );
  XNOR U19308 ( .A(n19655), .B(n19656), .Z(n19649) );
  NOR U19309 ( .A(n19657), .B(n19658), .Z(n19656) );
  XOR U19310 ( .A(n19655), .B(n19659), .Z(n19657) );
  XNOR U19311 ( .A(n19618), .B(n19625), .Z(n19637) );
  NOR U19312 ( .A(n19586), .B(n19660), .Z(n19625) );
  XOR U19313 ( .A(n19630), .B(n19629), .Z(n19618) );
  XNOR U19314 ( .A(n19661), .B(n19626), .Z(n19629) );
  XOR U19315 ( .A(n19662), .B(n19663), .Z(n19626) );
  AND U19316 ( .A(n19664), .B(n19665), .Z(n19663) );
  XOR U19317 ( .A(n19662), .B(n19666), .Z(n19664) );
  XNOR U19318 ( .A(n19667), .B(n19668), .Z(n19661) );
  NOR U19319 ( .A(n19669), .B(n19670), .Z(n19668) );
  XNOR U19320 ( .A(n19667), .B(n19671), .Z(n19669) );
  XOR U19321 ( .A(n19672), .B(n19673), .Z(n19630) );
  NOR U19322 ( .A(n19674), .B(n19675), .Z(n19673) );
  XNOR U19323 ( .A(n19672), .B(n19676), .Z(n19674) );
  XNOR U19324 ( .A(n19575), .B(n19633), .Z(n19635) );
  XNOR U19325 ( .A(n19677), .B(n19678), .Z(n19575) );
  AND U19326 ( .A(n237), .B(n19582), .Z(n19678) );
  XOR U19327 ( .A(n19677), .B(n19580), .Z(n19582) );
  AND U19328 ( .A(n19583), .B(n19586), .Z(n19633) );
  XOR U19329 ( .A(n19679), .B(n19660), .Z(n19586) );
  XNOR U19330 ( .A(p_input[2048]), .B(p_input[288]), .Z(n19660) );
  XOR U19331 ( .A(n19648), .B(n19647), .Z(n19679) );
  XNOR U19332 ( .A(n19680), .B(n19654), .Z(n19647) );
  XNOR U19333 ( .A(n19643), .B(n19642), .Z(n19654) );
  XOR U19334 ( .A(n19681), .B(n19639), .Z(n19642) );
  XNOR U19335 ( .A(n16904), .B(p_input[298]), .Z(n19639) );
  XNOR U19336 ( .A(p_input[2059]), .B(p_input[299]), .Z(n19681) );
  XOR U19337 ( .A(p_input[2060]), .B(p_input[300]), .Z(n19643) );
  XNOR U19338 ( .A(n19653), .B(n19644), .Z(n19680) );
  XNOR U19339 ( .A(n17068), .B(p_input[289]), .Z(n19644) );
  XOR U19340 ( .A(n19682), .B(n19659), .Z(n19653) );
  XNOR U19341 ( .A(p_input[2063]), .B(p_input[303]), .Z(n19659) );
  XOR U19342 ( .A(n19650), .B(n19658), .Z(n19682) );
  XOR U19343 ( .A(n19683), .B(n19655), .Z(n19658) );
  XOR U19344 ( .A(p_input[2061]), .B(p_input[301]), .Z(n19655) );
  XNOR U19345 ( .A(p_input[2062]), .B(p_input[302]), .Z(n19683) );
  XNOR U19346 ( .A(n16738), .B(p_input[297]), .Z(n19650) );
  XNOR U19347 ( .A(n19666), .B(n19665), .Z(n19648) );
  XNOR U19348 ( .A(n19684), .B(n19671), .Z(n19665) );
  XOR U19349 ( .A(p_input[2056]), .B(p_input[296]), .Z(n19671) );
  XOR U19350 ( .A(n19662), .B(n19670), .Z(n19684) );
  XOR U19351 ( .A(n19685), .B(n19667), .Z(n19670) );
  XOR U19352 ( .A(p_input[2054]), .B(p_input[294]), .Z(n19667) );
  XNOR U19353 ( .A(p_input[2055]), .B(p_input[295]), .Z(n19685) );
  XNOR U19354 ( .A(n16741), .B(p_input[290]), .Z(n19662) );
  XNOR U19355 ( .A(n19676), .B(n19675), .Z(n19666) );
  XOR U19356 ( .A(n19686), .B(n19672), .Z(n19675) );
  XOR U19357 ( .A(p_input[2051]), .B(p_input[291]), .Z(n19672) );
  XNOR U19358 ( .A(p_input[2052]), .B(p_input[292]), .Z(n19686) );
  XOR U19359 ( .A(p_input[2053]), .B(p_input[293]), .Z(n19676) );
  XNOR U19360 ( .A(n19687), .B(n19688), .Z(n19583) );
  AND U19361 ( .A(n237), .B(n19689), .Z(n19688) );
  XNOR U19362 ( .A(n19690), .B(n19691), .Z(n237) );
  AND U19363 ( .A(n19692), .B(n19693), .Z(n19691) );
  XOR U19364 ( .A(n19690), .B(n19593), .Z(n19693) );
  XNOR U19365 ( .A(n19690), .B(n19547), .Z(n19692) );
  XOR U19366 ( .A(n19694), .B(n19695), .Z(n19690) );
  AND U19367 ( .A(n19696), .B(n19697), .Z(n19695) );
  XOR U19368 ( .A(n19694), .B(n19557), .Z(n19696) );
  XOR U19369 ( .A(n19698), .B(n19699), .Z(n19536) );
  AND U19370 ( .A(n241), .B(n19689), .Z(n19699) );
  XNOR U19371 ( .A(n19687), .B(n19698), .Z(n19689) );
  XNOR U19372 ( .A(n19700), .B(n19701), .Z(n241) );
  AND U19373 ( .A(n19702), .B(n19703), .Z(n19701) );
  XNOR U19374 ( .A(n19704), .B(n19700), .Z(n19703) );
  IV U19375 ( .A(n19593), .Z(n19704) );
  XNOR U19376 ( .A(n19705), .B(n19706), .Z(n19593) );
  AND U19377 ( .A(n244), .B(n19707), .Z(n19706) );
  XNOR U19378 ( .A(n19705), .B(n19708), .Z(n19707) );
  XNOR U19379 ( .A(n19547), .B(n19700), .Z(n19702) );
  XOR U19380 ( .A(n19709), .B(n19710), .Z(n19547) );
  AND U19381 ( .A(n252), .B(n19711), .Z(n19710) );
  XOR U19382 ( .A(n19694), .B(n19712), .Z(n19700) );
  AND U19383 ( .A(n19713), .B(n19697), .Z(n19712) );
  XNOR U19384 ( .A(n19606), .B(n19694), .Z(n19697) );
  XNOR U19385 ( .A(n19714), .B(n19715), .Z(n19606) );
  AND U19386 ( .A(n244), .B(n19716), .Z(n19715) );
  XOR U19387 ( .A(n19717), .B(n19714), .Z(n19716) );
  XNOR U19388 ( .A(n19718), .B(n19694), .Z(n19713) );
  IV U19389 ( .A(n19557), .Z(n19718) );
  XOR U19390 ( .A(n19719), .B(n19720), .Z(n19557) );
  AND U19391 ( .A(n252), .B(n19721), .Z(n19720) );
  XOR U19392 ( .A(n19722), .B(n19723), .Z(n19694) );
  AND U19393 ( .A(n19724), .B(n19725), .Z(n19723) );
  XNOR U19394 ( .A(n19631), .B(n19722), .Z(n19725) );
  XNOR U19395 ( .A(n19726), .B(n19727), .Z(n19631) );
  AND U19396 ( .A(n244), .B(n19728), .Z(n19727) );
  XNOR U19397 ( .A(n19729), .B(n19726), .Z(n19728) );
  XOR U19398 ( .A(n19722), .B(n19568), .Z(n19724) );
  XOR U19399 ( .A(n19730), .B(n19731), .Z(n19568) );
  AND U19400 ( .A(n252), .B(n19732), .Z(n19731) );
  XOR U19401 ( .A(n19733), .B(n19734), .Z(n19722) );
  AND U19402 ( .A(n19735), .B(n19736), .Z(n19734) );
  XNOR U19403 ( .A(n19733), .B(n19677), .Z(n19736) );
  XNOR U19404 ( .A(n19737), .B(n19738), .Z(n19677) );
  AND U19405 ( .A(n244), .B(n19739), .Z(n19738) );
  XOR U19406 ( .A(n19740), .B(n19737), .Z(n19739) );
  XNOR U19407 ( .A(n19741), .B(n19733), .Z(n19735) );
  IV U19408 ( .A(n19580), .Z(n19741) );
  XOR U19409 ( .A(n19742), .B(n19743), .Z(n19580) );
  AND U19410 ( .A(n252), .B(n19744), .Z(n19743) );
  AND U19411 ( .A(n19698), .B(n19687), .Z(n19733) );
  XNOR U19412 ( .A(n19745), .B(n19746), .Z(n19687) );
  AND U19413 ( .A(n244), .B(n19747), .Z(n19746) );
  XNOR U19414 ( .A(n19748), .B(n19745), .Z(n19747) );
  XNOR U19415 ( .A(n19749), .B(n19750), .Z(n244) );
  AND U19416 ( .A(n19751), .B(n19752), .Z(n19750) );
  XOR U19417 ( .A(n19708), .B(n19749), .Z(n19752) );
  AND U19418 ( .A(n19753), .B(n19754), .Z(n19708) );
  XOR U19419 ( .A(n19749), .B(n19705), .Z(n19751) );
  XNOR U19420 ( .A(n19755), .B(n19756), .Z(n19705) );
  AND U19421 ( .A(n248), .B(n19711), .Z(n19756) );
  XOR U19422 ( .A(n19709), .B(n19755), .Z(n19711) );
  XOR U19423 ( .A(n19757), .B(n19758), .Z(n19749) );
  AND U19424 ( .A(n19759), .B(n19760), .Z(n19758) );
  XNOR U19425 ( .A(n19757), .B(n19753), .Z(n19760) );
  IV U19426 ( .A(n19717), .Z(n19753) );
  XOR U19427 ( .A(n19761), .B(n19762), .Z(n19717) );
  XOR U19428 ( .A(n19763), .B(n19754), .Z(n19762) );
  AND U19429 ( .A(n19729), .B(n19764), .Z(n19754) );
  AND U19430 ( .A(n19765), .B(n19766), .Z(n19763) );
  XOR U19431 ( .A(n19767), .B(n19761), .Z(n19765) );
  XNOR U19432 ( .A(n19714), .B(n19757), .Z(n19759) );
  XNOR U19433 ( .A(n19768), .B(n19769), .Z(n19714) );
  AND U19434 ( .A(n248), .B(n19721), .Z(n19769) );
  XOR U19435 ( .A(n19768), .B(n19719), .Z(n19721) );
  XOR U19436 ( .A(n19770), .B(n19771), .Z(n19757) );
  AND U19437 ( .A(n19772), .B(n19773), .Z(n19771) );
  XNOR U19438 ( .A(n19770), .B(n19729), .Z(n19773) );
  XOR U19439 ( .A(n19774), .B(n19766), .Z(n19729) );
  XNOR U19440 ( .A(n19775), .B(n19761), .Z(n19766) );
  XOR U19441 ( .A(n19776), .B(n19777), .Z(n19761) );
  AND U19442 ( .A(n19778), .B(n19779), .Z(n19777) );
  XOR U19443 ( .A(n19780), .B(n19776), .Z(n19778) );
  XNOR U19444 ( .A(n19781), .B(n19782), .Z(n19775) );
  AND U19445 ( .A(n19783), .B(n19784), .Z(n19782) );
  XOR U19446 ( .A(n19781), .B(n19785), .Z(n19783) );
  XNOR U19447 ( .A(n19767), .B(n19764), .Z(n19774) );
  AND U19448 ( .A(n19786), .B(n19787), .Z(n19764) );
  XOR U19449 ( .A(n19788), .B(n19789), .Z(n19767) );
  AND U19450 ( .A(n19790), .B(n19791), .Z(n19789) );
  XOR U19451 ( .A(n19788), .B(n19792), .Z(n19790) );
  XNOR U19452 ( .A(n19726), .B(n19770), .Z(n19772) );
  XNOR U19453 ( .A(n19793), .B(n19794), .Z(n19726) );
  AND U19454 ( .A(n248), .B(n19732), .Z(n19794) );
  XOR U19455 ( .A(n19793), .B(n19730), .Z(n19732) );
  XOR U19456 ( .A(n19795), .B(n19796), .Z(n19770) );
  AND U19457 ( .A(n19797), .B(n19798), .Z(n19796) );
  XNOR U19458 ( .A(n19795), .B(n19786), .Z(n19798) );
  IV U19459 ( .A(n19740), .Z(n19786) );
  XNOR U19460 ( .A(n19799), .B(n19779), .Z(n19740) );
  XNOR U19461 ( .A(n19800), .B(n19785), .Z(n19779) );
  XOR U19462 ( .A(n19801), .B(n19802), .Z(n19785) );
  NOR U19463 ( .A(n19803), .B(n19804), .Z(n19802) );
  XNOR U19464 ( .A(n19801), .B(n19805), .Z(n19803) );
  XNOR U19465 ( .A(n19784), .B(n19776), .Z(n19800) );
  XOR U19466 ( .A(n19806), .B(n19807), .Z(n19776) );
  AND U19467 ( .A(n19808), .B(n19809), .Z(n19807) );
  XNOR U19468 ( .A(n19806), .B(n19810), .Z(n19808) );
  XNOR U19469 ( .A(n19811), .B(n19781), .Z(n19784) );
  XOR U19470 ( .A(n19812), .B(n19813), .Z(n19781) );
  AND U19471 ( .A(n19814), .B(n19815), .Z(n19813) );
  XOR U19472 ( .A(n19812), .B(n19816), .Z(n19814) );
  XNOR U19473 ( .A(n19817), .B(n19818), .Z(n19811) );
  NOR U19474 ( .A(n19819), .B(n19820), .Z(n19818) );
  XOR U19475 ( .A(n19817), .B(n19821), .Z(n19819) );
  XNOR U19476 ( .A(n19780), .B(n19787), .Z(n19799) );
  NOR U19477 ( .A(n19748), .B(n19822), .Z(n19787) );
  XOR U19478 ( .A(n19792), .B(n19791), .Z(n19780) );
  XNOR U19479 ( .A(n19823), .B(n19788), .Z(n19791) );
  XOR U19480 ( .A(n19824), .B(n19825), .Z(n19788) );
  AND U19481 ( .A(n19826), .B(n19827), .Z(n19825) );
  XOR U19482 ( .A(n19824), .B(n19828), .Z(n19826) );
  XNOR U19483 ( .A(n19829), .B(n19830), .Z(n19823) );
  NOR U19484 ( .A(n19831), .B(n19832), .Z(n19830) );
  XNOR U19485 ( .A(n19829), .B(n19833), .Z(n19831) );
  XOR U19486 ( .A(n19834), .B(n19835), .Z(n19792) );
  NOR U19487 ( .A(n19836), .B(n19837), .Z(n19835) );
  XNOR U19488 ( .A(n19834), .B(n19838), .Z(n19836) );
  XNOR U19489 ( .A(n19737), .B(n19795), .Z(n19797) );
  XNOR U19490 ( .A(n19839), .B(n19840), .Z(n19737) );
  AND U19491 ( .A(n248), .B(n19744), .Z(n19840) );
  XOR U19492 ( .A(n19839), .B(n19742), .Z(n19744) );
  AND U19493 ( .A(n19745), .B(n19748), .Z(n19795) );
  XOR U19494 ( .A(n19841), .B(n19822), .Z(n19748) );
  XNOR U19495 ( .A(p_input[2048]), .B(p_input[304]), .Z(n19822) );
  XOR U19496 ( .A(n19810), .B(n19809), .Z(n19841) );
  XNOR U19497 ( .A(n19842), .B(n19816), .Z(n19809) );
  XNOR U19498 ( .A(n19805), .B(n19804), .Z(n19816) );
  XOR U19499 ( .A(n19843), .B(n19801), .Z(n19804) );
  XNOR U19500 ( .A(n16904), .B(p_input[314]), .Z(n19801) );
  XNOR U19501 ( .A(p_input[2059]), .B(p_input[315]), .Z(n19843) );
  XOR U19502 ( .A(p_input[2060]), .B(p_input[316]), .Z(n19805) );
  XNOR U19503 ( .A(n19815), .B(n19806), .Z(n19842) );
  XNOR U19504 ( .A(n17068), .B(p_input[305]), .Z(n19806) );
  XOR U19505 ( .A(n19844), .B(n19821), .Z(n19815) );
  XNOR U19506 ( .A(p_input[2063]), .B(p_input[319]), .Z(n19821) );
  XOR U19507 ( .A(n19812), .B(n19820), .Z(n19844) );
  XOR U19508 ( .A(n19845), .B(n19817), .Z(n19820) );
  XOR U19509 ( .A(p_input[2061]), .B(p_input[317]), .Z(n19817) );
  XNOR U19510 ( .A(p_input[2062]), .B(p_input[318]), .Z(n19845) );
  XNOR U19511 ( .A(n16738), .B(p_input[313]), .Z(n19812) );
  XNOR U19512 ( .A(n19828), .B(n19827), .Z(n19810) );
  XNOR U19513 ( .A(n19846), .B(n19833), .Z(n19827) );
  XOR U19514 ( .A(p_input[2056]), .B(p_input[312]), .Z(n19833) );
  XOR U19515 ( .A(n19824), .B(n19832), .Z(n19846) );
  XOR U19516 ( .A(n19847), .B(n19829), .Z(n19832) );
  XOR U19517 ( .A(p_input[2054]), .B(p_input[310]), .Z(n19829) );
  XNOR U19518 ( .A(p_input[2055]), .B(p_input[311]), .Z(n19847) );
  XNOR U19519 ( .A(n16741), .B(p_input[306]), .Z(n19824) );
  XNOR U19520 ( .A(n19838), .B(n19837), .Z(n19828) );
  XOR U19521 ( .A(n19848), .B(n19834), .Z(n19837) );
  XOR U19522 ( .A(p_input[2051]), .B(p_input[307]), .Z(n19834) );
  XNOR U19523 ( .A(p_input[2052]), .B(p_input[308]), .Z(n19848) );
  XOR U19524 ( .A(p_input[2053]), .B(p_input[309]), .Z(n19838) );
  XNOR U19525 ( .A(n19849), .B(n19850), .Z(n19745) );
  AND U19526 ( .A(n248), .B(n19851), .Z(n19850) );
  XNOR U19527 ( .A(n19852), .B(n19853), .Z(n248) );
  AND U19528 ( .A(n19854), .B(n19855), .Z(n19853) );
  XOR U19529 ( .A(n19852), .B(n19755), .Z(n19855) );
  XNOR U19530 ( .A(n19852), .B(n19709), .Z(n19854) );
  XOR U19531 ( .A(n19856), .B(n19857), .Z(n19852) );
  AND U19532 ( .A(n19858), .B(n19859), .Z(n19857) );
  XOR U19533 ( .A(n19856), .B(n19719), .Z(n19858) );
  XOR U19534 ( .A(n19860), .B(n19861), .Z(n19698) );
  AND U19535 ( .A(n252), .B(n19851), .Z(n19861) );
  XNOR U19536 ( .A(n19849), .B(n19860), .Z(n19851) );
  XNOR U19537 ( .A(n19862), .B(n19863), .Z(n252) );
  AND U19538 ( .A(n19864), .B(n19865), .Z(n19863) );
  XNOR U19539 ( .A(n19866), .B(n19862), .Z(n19865) );
  IV U19540 ( .A(n19755), .Z(n19866) );
  XNOR U19541 ( .A(n19867), .B(n19868), .Z(n19755) );
  AND U19542 ( .A(n255), .B(n19869), .Z(n19868) );
  XNOR U19543 ( .A(n19867), .B(n19870), .Z(n19869) );
  XNOR U19544 ( .A(n19709), .B(n19862), .Z(n19864) );
  XOR U19545 ( .A(n19871), .B(n19872), .Z(n19709) );
  AND U19546 ( .A(n263), .B(n19873), .Z(n19872) );
  XOR U19547 ( .A(n19856), .B(n19874), .Z(n19862) );
  AND U19548 ( .A(n19875), .B(n19859), .Z(n19874) );
  XNOR U19549 ( .A(n19768), .B(n19856), .Z(n19859) );
  XNOR U19550 ( .A(n19876), .B(n19877), .Z(n19768) );
  AND U19551 ( .A(n255), .B(n19878), .Z(n19877) );
  XOR U19552 ( .A(n19879), .B(n19876), .Z(n19878) );
  XNOR U19553 ( .A(n19880), .B(n19856), .Z(n19875) );
  IV U19554 ( .A(n19719), .Z(n19880) );
  XOR U19555 ( .A(n19881), .B(n19882), .Z(n19719) );
  AND U19556 ( .A(n263), .B(n19883), .Z(n19882) );
  XOR U19557 ( .A(n19884), .B(n19885), .Z(n19856) );
  AND U19558 ( .A(n19886), .B(n19887), .Z(n19885) );
  XNOR U19559 ( .A(n19793), .B(n19884), .Z(n19887) );
  XNOR U19560 ( .A(n19888), .B(n19889), .Z(n19793) );
  AND U19561 ( .A(n255), .B(n19890), .Z(n19889) );
  XNOR U19562 ( .A(n19891), .B(n19888), .Z(n19890) );
  XOR U19563 ( .A(n19884), .B(n19730), .Z(n19886) );
  XOR U19564 ( .A(n19892), .B(n19893), .Z(n19730) );
  AND U19565 ( .A(n263), .B(n19894), .Z(n19893) );
  XOR U19566 ( .A(n19895), .B(n19896), .Z(n19884) );
  AND U19567 ( .A(n19897), .B(n19898), .Z(n19896) );
  XNOR U19568 ( .A(n19895), .B(n19839), .Z(n19898) );
  XNOR U19569 ( .A(n19899), .B(n19900), .Z(n19839) );
  AND U19570 ( .A(n255), .B(n19901), .Z(n19900) );
  XOR U19571 ( .A(n19902), .B(n19899), .Z(n19901) );
  XNOR U19572 ( .A(n19903), .B(n19895), .Z(n19897) );
  IV U19573 ( .A(n19742), .Z(n19903) );
  XOR U19574 ( .A(n19904), .B(n19905), .Z(n19742) );
  AND U19575 ( .A(n263), .B(n19906), .Z(n19905) );
  AND U19576 ( .A(n19860), .B(n19849), .Z(n19895) );
  XNOR U19577 ( .A(n19907), .B(n19908), .Z(n19849) );
  AND U19578 ( .A(n255), .B(n19909), .Z(n19908) );
  XNOR U19579 ( .A(n19910), .B(n19907), .Z(n19909) );
  XNOR U19580 ( .A(n19911), .B(n19912), .Z(n255) );
  AND U19581 ( .A(n19913), .B(n19914), .Z(n19912) );
  XOR U19582 ( .A(n19870), .B(n19911), .Z(n19914) );
  AND U19583 ( .A(n19915), .B(n19916), .Z(n19870) );
  XOR U19584 ( .A(n19911), .B(n19867), .Z(n19913) );
  XNOR U19585 ( .A(n19917), .B(n19918), .Z(n19867) );
  AND U19586 ( .A(n259), .B(n19873), .Z(n19918) );
  XOR U19587 ( .A(n19871), .B(n19917), .Z(n19873) );
  XOR U19588 ( .A(n19919), .B(n19920), .Z(n19911) );
  AND U19589 ( .A(n19921), .B(n19922), .Z(n19920) );
  XNOR U19590 ( .A(n19919), .B(n19915), .Z(n19922) );
  IV U19591 ( .A(n19879), .Z(n19915) );
  XOR U19592 ( .A(n19923), .B(n19924), .Z(n19879) );
  XOR U19593 ( .A(n19925), .B(n19916), .Z(n19924) );
  AND U19594 ( .A(n19891), .B(n19926), .Z(n19916) );
  AND U19595 ( .A(n19927), .B(n19928), .Z(n19925) );
  XOR U19596 ( .A(n19929), .B(n19923), .Z(n19927) );
  XNOR U19597 ( .A(n19876), .B(n19919), .Z(n19921) );
  XNOR U19598 ( .A(n19930), .B(n19931), .Z(n19876) );
  AND U19599 ( .A(n259), .B(n19883), .Z(n19931) );
  XOR U19600 ( .A(n19930), .B(n19881), .Z(n19883) );
  XOR U19601 ( .A(n19932), .B(n19933), .Z(n19919) );
  AND U19602 ( .A(n19934), .B(n19935), .Z(n19933) );
  XNOR U19603 ( .A(n19932), .B(n19891), .Z(n19935) );
  XOR U19604 ( .A(n19936), .B(n19928), .Z(n19891) );
  XNOR U19605 ( .A(n19937), .B(n19923), .Z(n19928) );
  XOR U19606 ( .A(n19938), .B(n19939), .Z(n19923) );
  AND U19607 ( .A(n19940), .B(n19941), .Z(n19939) );
  XOR U19608 ( .A(n19942), .B(n19938), .Z(n19940) );
  XNOR U19609 ( .A(n19943), .B(n19944), .Z(n19937) );
  AND U19610 ( .A(n19945), .B(n19946), .Z(n19944) );
  XOR U19611 ( .A(n19943), .B(n19947), .Z(n19945) );
  XNOR U19612 ( .A(n19929), .B(n19926), .Z(n19936) );
  AND U19613 ( .A(n19948), .B(n19949), .Z(n19926) );
  XOR U19614 ( .A(n19950), .B(n19951), .Z(n19929) );
  AND U19615 ( .A(n19952), .B(n19953), .Z(n19951) );
  XOR U19616 ( .A(n19950), .B(n19954), .Z(n19952) );
  XNOR U19617 ( .A(n19888), .B(n19932), .Z(n19934) );
  XNOR U19618 ( .A(n19955), .B(n19956), .Z(n19888) );
  AND U19619 ( .A(n259), .B(n19894), .Z(n19956) );
  XOR U19620 ( .A(n19955), .B(n19892), .Z(n19894) );
  XOR U19621 ( .A(n19957), .B(n19958), .Z(n19932) );
  AND U19622 ( .A(n19959), .B(n19960), .Z(n19958) );
  XNOR U19623 ( .A(n19957), .B(n19948), .Z(n19960) );
  IV U19624 ( .A(n19902), .Z(n19948) );
  XNOR U19625 ( .A(n19961), .B(n19941), .Z(n19902) );
  XNOR U19626 ( .A(n19962), .B(n19947), .Z(n19941) );
  XOR U19627 ( .A(n19963), .B(n19964), .Z(n19947) );
  NOR U19628 ( .A(n19965), .B(n19966), .Z(n19964) );
  XNOR U19629 ( .A(n19963), .B(n19967), .Z(n19965) );
  XNOR U19630 ( .A(n19946), .B(n19938), .Z(n19962) );
  XOR U19631 ( .A(n19968), .B(n19969), .Z(n19938) );
  AND U19632 ( .A(n19970), .B(n19971), .Z(n19969) );
  XNOR U19633 ( .A(n19968), .B(n19972), .Z(n19970) );
  XNOR U19634 ( .A(n19973), .B(n19943), .Z(n19946) );
  XOR U19635 ( .A(n19974), .B(n19975), .Z(n19943) );
  AND U19636 ( .A(n19976), .B(n19977), .Z(n19975) );
  XOR U19637 ( .A(n19974), .B(n19978), .Z(n19976) );
  XNOR U19638 ( .A(n19979), .B(n19980), .Z(n19973) );
  NOR U19639 ( .A(n19981), .B(n19982), .Z(n19980) );
  XOR U19640 ( .A(n19979), .B(n19983), .Z(n19981) );
  XNOR U19641 ( .A(n19942), .B(n19949), .Z(n19961) );
  NOR U19642 ( .A(n19910), .B(n19984), .Z(n19949) );
  XOR U19643 ( .A(n19954), .B(n19953), .Z(n19942) );
  XNOR U19644 ( .A(n19985), .B(n19950), .Z(n19953) );
  XOR U19645 ( .A(n19986), .B(n19987), .Z(n19950) );
  AND U19646 ( .A(n19988), .B(n19989), .Z(n19987) );
  XOR U19647 ( .A(n19986), .B(n19990), .Z(n19988) );
  XNOR U19648 ( .A(n19991), .B(n19992), .Z(n19985) );
  NOR U19649 ( .A(n19993), .B(n19994), .Z(n19992) );
  XNOR U19650 ( .A(n19991), .B(n19995), .Z(n19993) );
  XOR U19651 ( .A(n19996), .B(n19997), .Z(n19954) );
  NOR U19652 ( .A(n19998), .B(n19999), .Z(n19997) );
  XNOR U19653 ( .A(n19996), .B(n20000), .Z(n19998) );
  XNOR U19654 ( .A(n19899), .B(n19957), .Z(n19959) );
  XNOR U19655 ( .A(n20001), .B(n20002), .Z(n19899) );
  AND U19656 ( .A(n259), .B(n19906), .Z(n20002) );
  XOR U19657 ( .A(n20001), .B(n19904), .Z(n19906) );
  AND U19658 ( .A(n19907), .B(n19910), .Z(n19957) );
  XOR U19659 ( .A(n20003), .B(n19984), .Z(n19910) );
  XNOR U19660 ( .A(p_input[2048]), .B(p_input[320]), .Z(n19984) );
  XOR U19661 ( .A(n19972), .B(n19971), .Z(n20003) );
  XNOR U19662 ( .A(n20004), .B(n19978), .Z(n19971) );
  XNOR U19663 ( .A(n19967), .B(n19966), .Z(n19978) );
  XOR U19664 ( .A(n20005), .B(n19963), .Z(n19966) );
  XNOR U19665 ( .A(n16904), .B(p_input[330]), .Z(n19963) );
  XNOR U19666 ( .A(p_input[2059]), .B(p_input[331]), .Z(n20005) );
  XOR U19667 ( .A(p_input[2060]), .B(p_input[332]), .Z(n19967) );
  XNOR U19668 ( .A(n19977), .B(n19968), .Z(n20004) );
  XNOR U19669 ( .A(n17068), .B(p_input[321]), .Z(n19968) );
  XOR U19670 ( .A(n20006), .B(n19983), .Z(n19977) );
  XNOR U19671 ( .A(p_input[2063]), .B(p_input[335]), .Z(n19983) );
  XOR U19672 ( .A(n19974), .B(n19982), .Z(n20006) );
  XOR U19673 ( .A(n20007), .B(n19979), .Z(n19982) );
  XOR U19674 ( .A(p_input[2061]), .B(p_input[333]), .Z(n19979) );
  XNOR U19675 ( .A(p_input[2062]), .B(p_input[334]), .Z(n20007) );
  XNOR U19676 ( .A(n16738), .B(p_input[329]), .Z(n19974) );
  XNOR U19677 ( .A(n19990), .B(n19989), .Z(n19972) );
  XNOR U19678 ( .A(n20008), .B(n19995), .Z(n19989) );
  XOR U19679 ( .A(p_input[2056]), .B(p_input[328]), .Z(n19995) );
  XOR U19680 ( .A(n19986), .B(n19994), .Z(n20008) );
  XOR U19681 ( .A(n20009), .B(n19991), .Z(n19994) );
  XOR U19682 ( .A(p_input[2054]), .B(p_input[326]), .Z(n19991) );
  XNOR U19683 ( .A(p_input[2055]), .B(p_input[327]), .Z(n20009) );
  XNOR U19684 ( .A(n16741), .B(p_input[322]), .Z(n19986) );
  XNOR U19685 ( .A(n20000), .B(n19999), .Z(n19990) );
  XOR U19686 ( .A(n20010), .B(n19996), .Z(n19999) );
  XOR U19687 ( .A(p_input[2051]), .B(p_input[323]), .Z(n19996) );
  XNOR U19688 ( .A(p_input[2052]), .B(p_input[324]), .Z(n20010) );
  XOR U19689 ( .A(p_input[2053]), .B(p_input[325]), .Z(n20000) );
  XNOR U19690 ( .A(n20011), .B(n20012), .Z(n19907) );
  AND U19691 ( .A(n259), .B(n20013), .Z(n20012) );
  XNOR U19692 ( .A(n20014), .B(n20015), .Z(n259) );
  AND U19693 ( .A(n20016), .B(n20017), .Z(n20015) );
  XOR U19694 ( .A(n20014), .B(n19917), .Z(n20017) );
  XNOR U19695 ( .A(n20014), .B(n19871), .Z(n20016) );
  XOR U19696 ( .A(n20018), .B(n20019), .Z(n20014) );
  AND U19697 ( .A(n20020), .B(n20021), .Z(n20019) );
  XOR U19698 ( .A(n20018), .B(n19881), .Z(n20020) );
  XOR U19699 ( .A(n20022), .B(n20023), .Z(n19860) );
  AND U19700 ( .A(n263), .B(n20013), .Z(n20023) );
  XNOR U19701 ( .A(n20011), .B(n20022), .Z(n20013) );
  XNOR U19702 ( .A(n20024), .B(n20025), .Z(n263) );
  AND U19703 ( .A(n20026), .B(n20027), .Z(n20025) );
  XNOR U19704 ( .A(n20028), .B(n20024), .Z(n20027) );
  IV U19705 ( .A(n19917), .Z(n20028) );
  XNOR U19706 ( .A(n20029), .B(n20030), .Z(n19917) );
  AND U19707 ( .A(n266), .B(n20031), .Z(n20030) );
  XNOR U19708 ( .A(n20029), .B(n20032), .Z(n20031) );
  XNOR U19709 ( .A(n19871), .B(n20024), .Z(n20026) );
  XOR U19710 ( .A(n20033), .B(n20034), .Z(n19871) );
  AND U19711 ( .A(n274), .B(n20035), .Z(n20034) );
  XOR U19712 ( .A(n20018), .B(n20036), .Z(n20024) );
  AND U19713 ( .A(n20037), .B(n20021), .Z(n20036) );
  XNOR U19714 ( .A(n19930), .B(n20018), .Z(n20021) );
  XNOR U19715 ( .A(n20038), .B(n20039), .Z(n19930) );
  AND U19716 ( .A(n266), .B(n20040), .Z(n20039) );
  XOR U19717 ( .A(n20041), .B(n20038), .Z(n20040) );
  XNOR U19718 ( .A(n20042), .B(n20018), .Z(n20037) );
  IV U19719 ( .A(n19881), .Z(n20042) );
  XOR U19720 ( .A(n20043), .B(n20044), .Z(n19881) );
  AND U19721 ( .A(n274), .B(n20045), .Z(n20044) );
  XOR U19722 ( .A(n20046), .B(n20047), .Z(n20018) );
  AND U19723 ( .A(n20048), .B(n20049), .Z(n20047) );
  XNOR U19724 ( .A(n19955), .B(n20046), .Z(n20049) );
  XNOR U19725 ( .A(n20050), .B(n20051), .Z(n19955) );
  AND U19726 ( .A(n266), .B(n20052), .Z(n20051) );
  XNOR U19727 ( .A(n20053), .B(n20050), .Z(n20052) );
  XOR U19728 ( .A(n20046), .B(n19892), .Z(n20048) );
  XOR U19729 ( .A(n20054), .B(n20055), .Z(n19892) );
  AND U19730 ( .A(n274), .B(n20056), .Z(n20055) );
  XOR U19731 ( .A(n20057), .B(n20058), .Z(n20046) );
  AND U19732 ( .A(n20059), .B(n20060), .Z(n20058) );
  XNOR U19733 ( .A(n20057), .B(n20001), .Z(n20060) );
  XNOR U19734 ( .A(n20061), .B(n20062), .Z(n20001) );
  AND U19735 ( .A(n266), .B(n20063), .Z(n20062) );
  XOR U19736 ( .A(n20064), .B(n20061), .Z(n20063) );
  XNOR U19737 ( .A(n20065), .B(n20057), .Z(n20059) );
  IV U19738 ( .A(n19904), .Z(n20065) );
  XOR U19739 ( .A(n20066), .B(n20067), .Z(n19904) );
  AND U19740 ( .A(n274), .B(n20068), .Z(n20067) );
  AND U19741 ( .A(n20022), .B(n20011), .Z(n20057) );
  XNOR U19742 ( .A(n20069), .B(n20070), .Z(n20011) );
  AND U19743 ( .A(n266), .B(n20071), .Z(n20070) );
  XNOR U19744 ( .A(n20072), .B(n20069), .Z(n20071) );
  XNOR U19745 ( .A(n20073), .B(n20074), .Z(n266) );
  AND U19746 ( .A(n20075), .B(n20076), .Z(n20074) );
  XOR U19747 ( .A(n20032), .B(n20073), .Z(n20076) );
  AND U19748 ( .A(n20077), .B(n20078), .Z(n20032) );
  XOR U19749 ( .A(n20073), .B(n20029), .Z(n20075) );
  XNOR U19750 ( .A(n20079), .B(n20080), .Z(n20029) );
  AND U19751 ( .A(n270), .B(n20035), .Z(n20080) );
  XOR U19752 ( .A(n20033), .B(n20079), .Z(n20035) );
  XOR U19753 ( .A(n20081), .B(n20082), .Z(n20073) );
  AND U19754 ( .A(n20083), .B(n20084), .Z(n20082) );
  XNOR U19755 ( .A(n20081), .B(n20077), .Z(n20084) );
  IV U19756 ( .A(n20041), .Z(n20077) );
  XOR U19757 ( .A(n20085), .B(n20086), .Z(n20041) );
  XOR U19758 ( .A(n20087), .B(n20078), .Z(n20086) );
  AND U19759 ( .A(n20053), .B(n20088), .Z(n20078) );
  AND U19760 ( .A(n20089), .B(n20090), .Z(n20087) );
  XOR U19761 ( .A(n20091), .B(n20085), .Z(n20089) );
  XNOR U19762 ( .A(n20038), .B(n20081), .Z(n20083) );
  XNOR U19763 ( .A(n20092), .B(n20093), .Z(n20038) );
  AND U19764 ( .A(n270), .B(n20045), .Z(n20093) );
  XOR U19765 ( .A(n20092), .B(n20043), .Z(n20045) );
  XOR U19766 ( .A(n20094), .B(n20095), .Z(n20081) );
  AND U19767 ( .A(n20096), .B(n20097), .Z(n20095) );
  XNOR U19768 ( .A(n20094), .B(n20053), .Z(n20097) );
  XOR U19769 ( .A(n20098), .B(n20090), .Z(n20053) );
  XNOR U19770 ( .A(n20099), .B(n20085), .Z(n20090) );
  XOR U19771 ( .A(n20100), .B(n20101), .Z(n20085) );
  AND U19772 ( .A(n20102), .B(n20103), .Z(n20101) );
  XOR U19773 ( .A(n20104), .B(n20100), .Z(n20102) );
  XNOR U19774 ( .A(n20105), .B(n20106), .Z(n20099) );
  AND U19775 ( .A(n20107), .B(n20108), .Z(n20106) );
  XOR U19776 ( .A(n20105), .B(n20109), .Z(n20107) );
  XNOR U19777 ( .A(n20091), .B(n20088), .Z(n20098) );
  AND U19778 ( .A(n20110), .B(n20111), .Z(n20088) );
  XOR U19779 ( .A(n20112), .B(n20113), .Z(n20091) );
  AND U19780 ( .A(n20114), .B(n20115), .Z(n20113) );
  XOR U19781 ( .A(n20112), .B(n20116), .Z(n20114) );
  XNOR U19782 ( .A(n20050), .B(n20094), .Z(n20096) );
  XNOR U19783 ( .A(n20117), .B(n20118), .Z(n20050) );
  AND U19784 ( .A(n270), .B(n20056), .Z(n20118) );
  XOR U19785 ( .A(n20117), .B(n20054), .Z(n20056) );
  XOR U19786 ( .A(n20119), .B(n20120), .Z(n20094) );
  AND U19787 ( .A(n20121), .B(n20122), .Z(n20120) );
  XNOR U19788 ( .A(n20119), .B(n20110), .Z(n20122) );
  IV U19789 ( .A(n20064), .Z(n20110) );
  XNOR U19790 ( .A(n20123), .B(n20103), .Z(n20064) );
  XNOR U19791 ( .A(n20124), .B(n20109), .Z(n20103) );
  XOR U19792 ( .A(n20125), .B(n20126), .Z(n20109) );
  NOR U19793 ( .A(n20127), .B(n20128), .Z(n20126) );
  XNOR U19794 ( .A(n20125), .B(n20129), .Z(n20127) );
  XNOR U19795 ( .A(n20108), .B(n20100), .Z(n20124) );
  XOR U19796 ( .A(n20130), .B(n20131), .Z(n20100) );
  AND U19797 ( .A(n20132), .B(n20133), .Z(n20131) );
  XNOR U19798 ( .A(n20130), .B(n20134), .Z(n20132) );
  XNOR U19799 ( .A(n20135), .B(n20105), .Z(n20108) );
  XOR U19800 ( .A(n20136), .B(n20137), .Z(n20105) );
  AND U19801 ( .A(n20138), .B(n20139), .Z(n20137) );
  XOR U19802 ( .A(n20136), .B(n20140), .Z(n20138) );
  XNOR U19803 ( .A(n20141), .B(n20142), .Z(n20135) );
  NOR U19804 ( .A(n20143), .B(n20144), .Z(n20142) );
  XOR U19805 ( .A(n20141), .B(n20145), .Z(n20143) );
  XNOR U19806 ( .A(n20104), .B(n20111), .Z(n20123) );
  NOR U19807 ( .A(n20072), .B(n20146), .Z(n20111) );
  XOR U19808 ( .A(n20116), .B(n20115), .Z(n20104) );
  XNOR U19809 ( .A(n20147), .B(n20112), .Z(n20115) );
  XOR U19810 ( .A(n20148), .B(n20149), .Z(n20112) );
  AND U19811 ( .A(n20150), .B(n20151), .Z(n20149) );
  XOR U19812 ( .A(n20148), .B(n20152), .Z(n20150) );
  XNOR U19813 ( .A(n20153), .B(n20154), .Z(n20147) );
  NOR U19814 ( .A(n20155), .B(n20156), .Z(n20154) );
  XNOR U19815 ( .A(n20153), .B(n20157), .Z(n20155) );
  XOR U19816 ( .A(n20158), .B(n20159), .Z(n20116) );
  NOR U19817 ( .A(n20160), .B(n20161), .Z(n20159) );
  XNOR U19818 ( .A(n20158), .B(n20162), .Z(n20160) );
  XNOR U19819 ( .A(n20061), .B(n20119), .Z(n20121) );
  XNOR U19820 ( .A(n20163), .B(n20164), .Z(n20061) );
  AND U19821 ( .A(n270), .B(n20068), .Z(n20164) );
  XOR U19822 ( .A(n20163), .B(n20066), .Z(n20068) );
  AND U19823 ( .A(n20069), .B(n20072), .Z(n20119) );
  XOR U19824 ( .A(n20165), .B(n20146), .Z(n20072) );
  XNOR U19825 ( .A(p_input[2048]), .B(p_input[336]), .Z(n20146) );
  XOR U19826 ( .A(n20134), .B(n20133), .Z(n20165) );
  XNOR U19827 ( .A(n20166), .B(n20140), .Z(n20133) );
  XNOR U19828 ( .A(n20129), .B(n20128), .Z(n20140) );
  XOR U19829 ( .A(n20167), .B(n20125), .Z(n20128) );
  XNOR U19830 ( .A(n16904), .B(p_input[346]), .Z(n20125) );
  XNOR U19831 ( .A(p_input[2059]), .B(p_input[347]), .Z(n20167) );
  XOR U19832 ( .A(p_input[2060]), .B(p_input[348]), .Z(n20129) );
  XNOR U19833 ( .A(n20139), .B(n20130), .Z(n20166) );
  XNOR U19834 ( .A(n17068), .B(p_input[337]), .Z(n20130) );
  XOR U19835 ( .A(n20168), .B(n20145), .Z(n20139) );
  XNOR U19836 ( .A(p_input[2063]), .B(p_input[351]), .Z(n20145) );
  XOR U19837 ( .A(n20136), .B(n20144), .Z(n20168) );
  XOR U19838 ( .A(n20169), .B(n20141), .Z(n20144) );
  XOR U19839 ( .A(p_input[2061]), .B(p_input[349]), .Z(n20141) );
  XNOR U19840 ( .A(p_input[2062]), .B(p_input[350]), .Z(n20169) );
  XNOR U19841 ( .A(n16738), .B(p_input[345]), .Z(n20136) );
  XNOR U19842 ( .A(n20152), .B(n20151), .Z(n20134) );
  XNOR U19843 ( .A(n20170), .B(n20157), .Z(n20151) );
  XOR U19844 ( .A(p_input[2056]), .B(p_input[344]), .Z(n20157) );
  XOR U19845 ( .A(n20148), .B(n20156), .Z(n20170) );
  XOR U19846 ( .A(n20171), .B(n20153), .Z(n20156) );
  XOR U19847 ( .A(p_input[2054]), .B(p_input[342]), .Z(n20153) );
  XNOR U19848 ( .A(p_input[2055]), .B(p_input[343]), .Z(n20171) );
  XNOR U19849 ( .A(n16741), .B(p_input[338]), .Z(n20148) );
  XNOR U19850 ( .A(n20162), .B(n20161), .Z(n20152) );
  XOR U19851 ( .A(n20172), .B(n20158), .Z(n20161) );
  XOR U19852 ( .A(p_input[2051]), .B(p_input[339]), .Z(n20158) );
  XNOR U19853 ( .A(p_input[2052]), .B(p_input[340]), .Z(n20172) );
  XOR U19854 ( .A(p_input[2053]), .B(p_input[341]), .Z(n20162) );
  XNOR U19855 ( .A(n20173), .B(n20174), .Z(n20069) );
  AND U19856 ( .A(n270), .B(n20175), .Z(n20174) );
  XNOR U19857 ( .A(n20176), .B(n20177), .Z(n270) );
  AND U19858 ( .A(n20178), .B(n20179), .Z(n20177) );
  XOR U19859 ( .A(n20176), .B(n20079), .Z(n20179) );
  XNOR U19860 ( .A(n20176), .B(n20033), .Z(n20178) );
  XOR U19861 ( .A(n20180), .B(n20181), .Z(n20176) );
  AND U19862 ( .A(n20182), .B(n20183), .Z(n20181) );
  XOR U19863 ( .A(n20180), .B(n20043), .Z(n20182) );
  XOR U19864 ( .A(n20184), .B(n20185), .Z(n20022) );
  AND U19865 ( .A(n274), .B(n20175), .Z(n20185) );
  XNOR U19866 ( .A(n20173), .B(n20184), .Z(n20175) );
  XNOR U19867 ( .A(n20186), .B(n20187), .Z(n274) );
  AND U19868 ( .A(n20188), .B(n20189), .Z(n20187) );
  XNOR U19869 ( .A(n20190), .B(n20186), .Z(n20189) );
  IV U19870 ( .A(n20079), .Z(n20190) );
  XNOR U19871 ( .A(n20191), .B(n20192), .Z(n20079) );
  AND U19872 ( .A(n277), .B(n20193), .Z(n20192) );
  XNOR U19873 ( .A(n20191), .B(n20194), .Z(n20193) );
  XNOR U19874 ( .A(n20033), .B(n20186), .Z(n20188) );
  XOR U19875 ( .A(n20195), .B(n20196), .Z(n20033) );
  AND U19876 ( .A(n285), .B(n20197), .Z(n20196) );
  XOR U19877 ( .A(n20180), .B(n20198), .Z(n20186) );
  AND U19878 ( .A(n20199), .B(n20183), .Z(n20198) );
  XNOR U19879 ( .A(n20092), .B(n20180), .Z(n20183) );
  XNOR U19880 ( .A(n20200), .B(n20201), .Z(n20092) );
  AND U19881 ( .A(n277), .B(n20202), .Z(n20201) );
  XOR U19882 ( .A(n20203), .B(n20200), .Z(n20202) );
  XNOR U19883 ( .A(n20204), .B(n20180), .Z(n20199) );
  IV U19884 ( .A(n20043), .Z(n20204) );
  XOR U19885 ( .A(n20205), .B(n20206), .Z(n20043) );
  AND U19886 ( .A(n285), .B(n20207), .Z(n20206) );
  XOR U19887 ( .A(n20208), .B(n20209), .Z(n20180) );
  AND U19888 ( .A(n20210), .B(n20211), .Z(n20209) );
  XNOR U19889 ( .A(n20117), .B(n20208), .Z(n20211) );
  XNOR U19890 ( .A(n20212), .B(n20213), .Z(n20117) );
  AND U19891 ( .A(n277), .B(n20214), .Z(n20213) );
  XNOR U19892 ( .A(n20215), .B(n20212), .Z(n20214) );
  XOR U19893 ( .A(n20208), .B(n20054), .Z(n20210) );
  XOR U19894 ( .A(n20216), .B(n20217), .Z(n20054) );
  AND U19895 ( .A(n285), .B(n20218), .Z(n20217) );
  XOR U19896 ( .A(n20219), .B(n20220), .Z(n20208) );
  AND U19897 ( .A(n20221), .B(n20222), .Z(n20220) );
  XNOR U19898 ( .A(n20219), .B(n20163), .Z(n20222) );
  XNOR U19899 ( .A(n20223), .B(n20224), .Z(n20163) );
  AND U19900 ( .A(n277), .B(n20225), .Z(n20224) );
  XOR U19901 ( .A(n20226), .B(n20223), .Z(n20225) );
  XNOR U19902 ( .A(n20227), .B(n20219), .Z(n20221) );
  IV U19903 ( .A(n20066), .Z(n20227) );
  XOR U19904 ( .A(n20228), .B(n20229), .Z(n20066) );
  AND U19905 ( .A(n285), .B(n20230), .Z(n20229) );
  AND U19906 ( .A(n20184), .B(n20173), .Z(n20219) );
  XNOR U19907 ( .A(n20231), .B(n20232), .Z(n20173) );
  AND U19908 ( .A(n277), .B(n20233), .Z(n20232) );
  XNOR U19909 ( .A(n20234), .B(n20231), .Z(n20233) );
  XNOR U19910 ( .A(n20235), .B(n20236), .Z(n277) );
  AND U19911 ( .A(n20237), .B(n20238), .Z(n20236) );
  XOR U19912 ( .A(n20194), .B(n20235), .Z(n20238) );
  AND U19913 ( .A(n20239), .B(n20240), .Z(n20194) );
  XOR U19914 ( .A(n20235), .B(n20191), .Z(n20237) );
  XNOR U19915 ( .A(n20241), .B(n20242), .Z(n20191) );
  AND U19916 ( .A(n281), .B(n20197), .Z(n20242) );
  XOR U19917 ( .A(n20195), .B(n20241), .Z(n20197) );
  XOR U19918 ( .A(n20243), .B(n20244), .Z(n20235) );
  AND U19919 ( .A(n20245), .B(n20246), .Z(n20244) );
  XNOR U19920 ( .A(n20243), .B(n20239), .Z(n20246) );
  IV U19921 ( .A(n20203), .Z(n20239) );
  XOR U19922 ( .A(n20247), .B(n20248), .Z(n20203) );
  XOR U19923 ( .A(n20249), .B(n20240), .Z(n20248) );
  AND U19924 ( .A(n20215), .B(n20250), .Z(n20240) );
  AND U19925 ( .A(n20251), .B(n20252), .Z(n20249) );
  XOR U19926 ( .A(n20253), .B(n20247), .Z(n20251) );
  XNOR U19927 ( .A(n20200), .B(n20243), .Z(n20245) );
  XNOR U19928 ( .A(n20254), .B(n20255), .Z(n20200) );
  AND U19929 ( .A(n281), .B(n20207), .Z(n20255) );
  XOR U19930 ( .A(n20254), .B(n20205), .Z(n20207) );
  XOR U19931 ( .A(n20256), .B(n20257), .Z(n20243) );
  AND U19932 ( .A(n20258), .B(n20259), .Z(n20257) );
  XNOR U19933 ( .A(n20256), .B(n20215), .Z(n20259) );
  XOR U19934 ( .A(n20260), .B(n20252), .Z(n20215) );
  XNOR U19935 ( .A(n20261), .B(n20247), .Z(n20252) );
  XOR U19936 ( .A(n20262), .B(n20263), .Z(n20247) );
  AND U19937 ( .A(n20264), .B(n20265), .Z(n20263) );
  XOR U19938 ( .A(n20266), .B(n20262), .Z(n20264) );
  XNOR U19939 ( .A(n20267), .B(n20268), .Z(n20261) );
  AND U19940 ( .A(n20269), .B(n20270), .Z(n20268) );
  XOR U19941 ( .A(n20267), .B(n20271), .Z(n20269) );
  XNOR U19942 ( .A(n20253), .B(n20250), .Z(n20260) );
  AND U19943 ( .A(n20272), .B(n20273), .Z(n20250) );
  XOR U19944 ( .A(n20274), .B(n20275), .Z(n20253) );
  AND U19945 ( .A(n20276), .B(n20277), .Z(n20275) );
  XOR U19946 ( .A(n20274), .B(n20278), .Z(n20276) );
  XNOR U19947 ( .A(n20212), .B(n20256), .Z(n20258) );
  XNOR U19948 ( .A(n20279), .B(n20280), .Z(n20212) );
  AND U19949 ( .A(n281), .B(n20218), .Z(n20280) );
  XOR U19950 ( .A(n20279), .B(n20216), .Z(n20218) );
  XOR U19951 ( .A(n20281), .B(n20282), .Z(n20256) );
  AND U19952 ( .A(n20283), .B(n20284), .Z(n20282) );
  XNOR U19953 ( .A(n20281), .B(n20272), .Z(n20284) );
  IV U19954 ( .A(n20226), .Z(n20272) );
  XNOR U19955 ( .A(n20285), .B(n20265), .Z(n20226) );
  XNOR U19956 ( .A(n20286), .B(n20271), .Z(n20265) );
  XOR U19957 ( .A(n20287), .B(n20288), .Z(n20271) );
  NOR U19958 ( .A(n20289), .B(n20290), .Z(n20288) );
  XNOR U19959 ( .A(n20287), .B(n20291), .Z(n20289) );
  XNOR U19960 ( .A(n20270), .B(n20262), .Z(n20286) );
  XOR U19961 ( .A(n20292), .B(n20293), .Z(n20262) );
  AND U19962 ( .A(n20294), .B(n20295), .Z(n20293) );
  XNOR U19963 ( .A(n20292), .B(n20296), .Z(n20294) );
  XNOR U19964 ( .A(n20297), .B(n20267), .Z(n20270) );
  XOR U19965 ( .A(n20298), .B(n20299), .Z(n20267) );
  AND U19966 ( .A(n20300), .B(n20301), .Z(n20299) );
  XOR U19967 ( .A(n20298), .B(n20302), .Z(n20300) );
  XNOR U19968 ( .A(n20303), .B(n20304), .Z(n20297) );
  NOR U19969 ( .A(n20305), .B(n20306), .Z(n20304) );
  XOR U19970 ( .A(n20303), .B(n20307), .Z(n20305) );
  XNOR U19971 ( .A(n20266), .B(n20273), .Z(n20285) );
  NOR U19972 ( .A(n20234), .B(n20308), .Z(n20273) );
  XOR U19973 ( .A(n20278), .B(n20277), .Z(n20266) );
  XNOR U19974 ( .A(n20309), .B(n20274), .Z(n20277) );
  XOR U19975 ( .A(n20310), .B(n20311), .Z(n20274) );
  AND U19976 ( .A(n20312), .B(n20313), .Z(n20311) );
  XOR U19977 ( .A(n20310), .B(n20314), .Z(n20312) );
  XNOR U19978 ( .A(n20315), .B(n20316), .Z(n20309) );
  NOR U19979 ( .A(n20317), .B(n20318), .Z(n20316) );
  XNOR U19980 ( .A(n20315), .B(n20319), .Z(n20317) );
  XOR U19981 ( .A(n20320), .B(n20321), .Z(n20278) );
  NOR U19982 ( .A(n20322), .B(n20323), .Z(n20321) );
  XNOR U19983 ( .A(n20320), .B(n20324), .Z(n20322) );
  XNOR U19984 ( .A(n20223), .B(n20281), .Z(n20283) );
  XNOR U19985 ( .A(n20325), .B(n20326), .Z(n20223) );
  AND U19986 ( .A(n281), .B(n20230), .Z(n20326) );
  XOR U19987 ( .A(n20325), .B(n20228), .Z(n20230) );
  AND U19988 ( .A(n20231), .B(n20234), .Z(n20281) );
  XOR U19989 ( .A(n20327), .B(n20308), .Z(n20234) );
  XNOR U19990 ( .A(p_input[2048]), .B(p_input[352]), .Z(n20308) );
  XOR U19991 ( .A(n20296), .B(n20295), .Z(n20327) );
  XNOR U19992 ( .A(n20328), .B(n20302), .Z(n20295) );
  XNOR U19993 ( .A(n20291), .B(n20290), .Z(n20302) );
  XOR U19994 ( .A(n20329), .B(n20287), .Z(n20290) );
  XNOR U19995 ( .A(n16904), .B(p_input[362]), .Z(n20287) );
  XNOR U19996 ( .A(p_input[2059]), .B(p_input[363]), .Z(n20329) );
  XOR U19997 ( .A(p_input[2060]), .B(p_input[364]), .Z(n20291) );
  XNOR U19998 ( .A(n20301), .B(n20292), .Z(n20328) );
  XNOR U19999 ( .A(n17068), .B(p_input[353]), .Z(n20292) );
  XOR U20000 ( .A(n20330), .B(n20307), .Z(n20301) );
  XNOR U20001 ( .A(p_input[2063]), .B(p_input[367]), .Z(n20307) );
  XOR U20002 ( .A(n20298), .B(n20306), .Z(n20330) );
  XOR U20003 ( .A(n20331), .B(n20303), .Z(n20306) );
  XOR U20004 ( .A(p_input[2061]), .B(p_input[365]), .Z(n20303) );
  XNOR U20005 ( .A(p_input[2062]), .B(p_input[366]), .Z(n20331) );
  XNOR U20006 ( .A(n16738), .B(p_input[361]), .Z(n20298) );
  XNOR U20007 ( .A(n20314), .B(n20313), .Z(n20296) );
  XNOR U20008 ( .A(n20332), .B(n20319), .Z(n20313) );
  XOR U20009 ( .A(p_input[2056]), .B(p_input[360]), .Z(n20319) );
  XOR U20010 ( .A(n20310), .B(n20318), .Z(n20332) );
  XOR U20011 ( .A(n20333), .B(n20315), .Z(n20318) );
  XOR U20012 ( .A(p_input[2054]), .B(p_input[358]), .Z(n20315) );
  XNOR U20013 ( .A(p_input[2055]), .B(p_input[359]), .Z(n20333) );
  XNOR U20014 ( .A(n16741), .B(p_input[354]), .Z(n20310) );
  XNOR U20015 ( .A(n20324), .B(n20323), .Z(n20314) );
  XOR U20016 ( .A(n20334), .B(n20320), .Z(n20323) );
  XOR U20017 ( .A(p_input[2051]), .B(p_input[355]), .Z(n20320) );
  XNOR U20018 ( .A(p_input[2052]), .B(p_input[356]), .Z(n20334) );
  XOR U20019 ( .A(p_input[2053]), .B(p_input[357]), .Z(n20324) );
  XNOR U20020 ( .A(n20335), .B(n20336), .Z(n20231) );
  AND U20021 ( .A(n281), .B(n20337), .Z(n20336) );
  XNOR U20022 ( .A(n20338), .B(n20339), .Z(n281) );
  AND U20023 ( .A(n20340), .B(n20341), .Z(n20339) );
  XOR U20024 ( .A(n20338), .B(n20241), .Z(n20341) );
  XNOR U20025 ( .A(n20338), .B(n20195), .Z(n20340) );
  XOR U20026 ( .A(n20342), .B(n20343), .Z(n20338) );
  AND U20027 ( .A(n20344), .B(n20345), .Z(n20343) );
  XOR U20028 ( .A(n20342), .B(n20205), .Z(n20344) );
  XOR U20029 ( .A(n20346), .B(n20347), .Z(n20184) );
  AND U20030 ( .A(n285), .B(n20337), .Z(n20347) );
  XNOR U20031 ( .A(n20335), .B(n20346), .Z(n20337) );
  XNOR U20032 ( .A(n20348), .B(n20349), .Z(n285) );
  AND U20033 ( .A(n20350), .B(n20351), .Z(n20349) );
  XNOR U20034 ( .A(n20352), .B(n20348), .Z(n20351) );
  IV U20035 ( .A(n20241), .Z(n20352) );
  XNOR U20036 ( .A(n20353), .B(n20354), .Z(n20241) );
  AND U20037 ( .A(n288), .B(n20355), .Z(n20354) );
  XNOR U20038 ( .A(n20353), .B(n20356), .Z(n20355) );
  XNOR U20039 ( .A(n20195), .B(n20348), .Z(n20350) );
  XOR U20040 ( .A(n20357), .B(n20358), .Z(n20195) );
  AND U20041 ( .A(n296), .B(n20359), .Z(n20358) );
  XOR U20042 ( .A(n20342), .B(n20360), .Z(n20348) );
  AND U20043 ( .A(n20361), .B(n20345), .Z(n20360) );
  XNOR U20044 ( .A(n20254), .B(n20342), .Z(n20345) );
  XNOR U20045 ( .A(n20362), .B(n20363), .Z(n20254) );
  AND U20046 ( .A(n288), .B(n20364), .Z(n20363) );
  XOR U20047 ( .A(n20365), .B(n20362), .Z(n20364) );
  XNOR U20048 ( .A(n20366), .B(n20342), .Z(n20361) );
  IV U20049 ( .A(n20205), .Z(n20366) );
  XOR U20050 ( .A(n20367), .B(n20368), .Z(n20205) );
  AND U20051 ( .A(n296), .B(n20369), .Z(n20368) );
  XOR U20052 ( .A(n20370), .B(n20371), .Z(n20342) );
  AND U20053 ( .A(n20372), .B(n20373), .Z(n20371) );
  XNOR U20054 ( .A(n20279), .B(n20370), .Z(n20373) );
  XNOR U20055 ( .A(n20374), .B(n20375), .Z(n20279) );
  AND U20056 ( .A(n288), .B(n20376), .Z(n20375) );
  XNOR U20057 ( .A(n20377), .B(n20374), .Z(n20376) );
  XOR U20058 ( .A(n20370), .B(n20216), .Z(n20372) );
  XOR U20059 ( .A(n20378), .B(n20379), .Z(n20216) );
  AND U20060 ( .A(n296), .B(n20380), .Z(n20379) );
  XOR U20061 ( .A(n20381), .B(n20382), .Z(n20370) );
  AND U20062 ( .A(n20383), .B(n20384), .Z(n20382) );
  XNOR U20063 ( .A(n20381), .B(n20325), .Z(n20384) );
  XNOR U20064 ( .A(n20385), .B(n20386), .Z(n20325) );
  AND U20065 ( .A(n288), .B(n20387), .Z(n20386) );
  XOR U20066 ( .A(n20388), .B(n20385), .Z(n20387) );
  XNOR U20067 ( .A(n20389), .B(n20381), .Z(n20383) );
  IV U20068 ( .A(n20228), .Z(n20389) );
  XOR U20069 ( .A(n20390), .B(n20391), .Z(n20228) );
  AND U20070 ( .A(n296), .B(n20392), .Z(n20391) );
  AND U20071 ( .A(n20346), .B(n20335), .Z(n20381) );
  XNOR U20072 ( .A(n20393), .B(n20394), .Z(n20335) );
  AND U20073 ( .A(n288), .B(n20395), .Z(n20394) );
  XNOR U20074 ( .A(n20396), .B(n20393), .Z(n20395) );
  XNOR U20075 ( .A(n20397), .B(n20398), .Z(n288) );
  AND U20076 ( .A(n20399), .B(n20400), .Z(n20398) );
  XOR U20077 ( .A(n20356), .B(n20397), .Z(n20400) );
  AND U20078 ( .A(n20401), .B(n20402), .Z(n20356) );
  XOR U20079 ( .A(n20397), .B(n20353), .Z(n20399) );
  XNOR U20080 ( .A(n20403), .B(n20404), .Z(n20353) );
  AND U20081 ( .A(n292), .B(n20359), .Z(n20404) );
  XOR U20082 ( .A(n20357), .B(n20403), .Z(n20359) );
  XOR U20083 ( .A(n20405), .B(n20406), .Z(n20397) );
  AND U20084 ( .A(n20407), .B(n20408), .Z(n20406) );
  XNOR U20085 ( .A(n20405), .B(n20401), .Z(n20408) );
  IV U20086 ( .A(n20365), .Z(n20401) );
  XOR U20087 ( .A(n20409), .B(n20410), .Z(n20365) );
  XOR U20088 ( .A(n20411), .B(n20402), .Z(n20410) );
  AND U20089 ( .A(n20377), .B(n20412), .Z(n20402) );
  AND U20090 ( .A(n20413), .B(n20414), .Z(n20411) );
  XOR U20091 ( .A(n20415), .B(n20409), .Z(n20413) );
  XNOR U20092 ( .A(n20362), .B(n20405), .Z(n20407) );
  XNOR U20093 ( .A(n20416), .B(n20417), .Z(n20362) );
  AND U20094 ( .A(n292), .B(n20369), .Z(n20417) );
  XOR U20095 ( .A(n20416), .B(n20367), .Z(n20369) );
  XOR U20096 ( .A(n20418), .B(n20419), .Z(n20405) );
  AND U20097 ( .A(n20420), .B(n20421), .Z(n20419) );
  XNOR U20098 ( .A(n20418), .B(n20377), .Z(n20421) );
  XOR U20099 ( .A(n20422), .B(n20414), .Z(n20377) );
  XNOR U20100 ( .A(n20423), .B(n20409), .Z(n20414) );
  XOR U20101 ( .A(n20424), .B(n20425), .Z(n20409) );
  AND U20102 ( .A(n20426), .B(n20427), .Z(n20425) );
  XOR U20103 ( .A(n20428), .B(n20424), .Z(n20426) );
  XNOR U20104 ( .A(n20429), .B(n20430), .Z(n20423) );
  AND U20105 ( .A(n20431), .B(n20432), .Z(n20430) );
  XOR U20106 ( .A(n20429), .B(n20433), .Z(n20431) );
  XNOR U20107 ( .A(n20415), .B(n20412), .Z(n20422) );
  AND U20108 ( .A(n20434), .B(n20435), .Z(n20412) );
  XOR U20109 ( .A(n20436), .B(n20437), .Z(n20415) );
  AND U20110 ( .A(n20438), .B(n20439), .Z(n20437) );
  XOR U20111 ( .A(n20436), .B(n20440), .Z(n20438) );
  XNOR U20112 ( .A(n20374), .B(n20418), .Z(n20420) );
  XNOR U20113 ( .A(n20441), .B(n20442), .Z(n20374) );
  AND U20114 ( .A(n292), .B(n20380), .Z(n20442) );
  XOR U20115 ( .A(n20441), .B(n20378), .Z(n20380) );
  XOR U20116 ( .A(n20443), .B(n20444), .Z(n20418) );
  AND U20117 ( .A(n20445), .B(n20446), .Z(n20444) );
  XNOR U20118 ( .A(n20443), .B(n20434), .Z(n20446) );
  IV U20119 ( .A(n20388), .Z(n20434) );
  XNOR U20120 ( .A(n20447), .B(n20427), .Z(n20388) );
  XNOR U20121 ( .A(n20448), .B(n20433), .Z(n20427) );
  XOR U20122 ( .A(n20449), .B(n20450), .Z(n20433) );
  NOR U20123 ( .A(n20451), .B(n20452), .Z(n20450) );
  XNOR U20124 ( .A(n20449), .B(n20453), .Z(n20451) );
  XNOR U20125 ( .A(n20432), .B(n20424), .Z(n20448) );
  XOR U20126 ( .A(n20454), .B(n20455), .Z(n20424) );
  AND U20127 ( .A(n20456), .B(n20457), .Z(n20455) );
  XNOR U20128 ( .A(n20454), .B(n20458), .Z(n20456) );
  XNOR U20129 ( .A(n20459), .B(n20429), .Z(n20432) );
  XOR U20130 ( .A(n20460), .B(n20461), .Z(n20429) );
  AND U20131 ( .A(n20462), .B(n20463), .Z(n20461) );
  XOR U20132 ( .A(n20460), .B(n20464), .Z(n20462) );
  XNOR U20133 ( .A(n20465), .B(n20466), .Z(n20459) );
  NOR U20134 ( .A(n20467), .B(n20468), .Z(n20466) );
  XOR U20135 ( .A(n20465), .B(n20469), .Z(n20467) );
  XNOR U20136 ( .A(n20428), .B(n20435), .Z(n20447) );
  NOR U20137 ( .A(n20396), .B(n20470), .Z(n20435) );
  XOR U20138 ( .A(n20440), .B(n20439), .Z(n20428) );
  XNOR U20139 ( .A(n20471), .B(n20436), .Z(n20439) );
  XOR U20140 ( .A(n20472), .B(n20473), .Z(n20436) );
  AND U20141 ( .A(n20474), .B(n20475), .Z(n20473) );
  XOR U20142 ( .A(n20472), .B(n20476), .Z(n20474) );
  XNOR U20143 ( .A(n20477), .B(n20478), .Z(n20471) );
  NOR U20144 ( .A(n20479), .B(n20480), .Z(n20478) );
  XNOR U20145 ( .A(n20477), .B(n20481), .Z(n20479) );
  XOR U20146 ( .A(n20482), .B(n20483), .Z(n20440) );
  NOR U20147 ( .A(n20484), .B(n20485), .Z(n20483) );
  XNOR U20148 ( .A(n20482), .B(n20486), .Z(n20484) );
  XNOR U20149 ( .A(n20385), .B(n20443), .Z(n20445) );
  XNOR U20150 ( .A(n20487), .B(n20488), .Z(n20385) );
  AND U20151 ( .A(n292), .B(n20392), .Z(n20488) );
  XOR U20152 ( .A(n20487), .B(n20390), .Z(n20392) );
  AND U20153 ( .A(n20393), .B(n20396), .Z(n20443) );
  XOR U20154 ( .A(n20489), .B(n20470), .Z(n20396) );
  XNOR U20155 ( .A(p_input[2048]), .B(p_input[368]), .Z(n20470) );
  XOR U20156 ( .A(n20458), .B(n20457), .Z(n20489) );
  XNOR U20157 ( .A(n20490), .B(n20464), .Z(n20457) );
  XNOR U20158 ( .A(n20453), .B(n20452), .Z(n20464) );
  XOR U20159 ( .A(n20491), .B(n20449), .Z(n20452) );
  XNOR U20160 ( .A(n16904), .B(p_input[378]), .Z(n20449) );
  XNOR U20161 ( .A(p_input[2059]), .B(p_input[379]), .Z(n20491) );
  XOR U20162 ( .A(p_input[2060]), .B(p_input[380]), .Z(n20453) );
  XNOR U20163 ( .A(n20463), .B(n20454), .Z(n20490) );
  XNOR U20164 ( .A(n17068), .B(p_input[369]), .Z(n20454) );
  XOR U20165 ( .A(n20492), .B(n20469), .Z(n20463) );
  XNOR U20166 ( .A(p_input[2063]), .B(p_input[383]), .Z(n20469) );
  XOR U20167 ( .A(n20460), .B(n20468), .Z(n20492) );
  XOR U20168 ( .A(n20493), .B(n20465), .Z(n20468) );
  XOR U20169 ( .A(p_input[2061]), .B(p_input[381]), .Z(n20465) );
  XNOR U20170 ( .A(p_input[2062]), .B(p_input[382]), .Z(n20493) );
  XNOR U20171 ( .A(n16738), .B(p_input[377]), .Z(n20460) );
  XNOR U20172 ( .A(n20476), .B(n20475), .Z(n20458) );
  XNOR U20173 ( .A(n20494), .B(n20481), .Z(n20475) );
  XOR U20174 ( .A(p_input[2056]), .B(p_input[376]), .Z(n20481) );
  XOR U20175 ( .A(n20472), .B(n20480), .Z(n20494) );
  XOR U20176 ( .A(n20495), .B(n20477), .Z(n20480) );
  XOR U20177 ( .A(p_input[2054]), .B(p_input[374]), .Z(n20477) );
  XNOR U20178 ( .A(p_input[2055]), .B(p_input[375]), .Z(n20495) );
  XNOR U20179 ( .A(n16741), .B(p_input[370]), .Z(n20472) );
  XNOR U20180 ( .A(n20486), .B(n20485), .Z(n20476) );
  XOR U20181 ( .A(n20496), .B(n20482), .Z(n20485) );
  XOR U20182 ( .A(p_input[2051]), .B(p_input[371]), .Z(n20482) );
  XNOR U20183 ( .A(p_input[2052]), .B(p_input[372]), .Z(n20496) );
  XOR U20184 ( .A(p_input[2053]), .B(p_input[373]), .Z(n20486) );
  XNOR U20185 ( .A(n20497), .B(n20498), .Z(n20393) );
  AND U20186 ( .A(n292), .B(n20499), .Z(n20498) );
  XNOR U20187 ( .A(n20500), .B(n20501), .Z(n292) );
  AND U20188 ( .A(n20502), .B(n20503), .Z(n20501) );
  XOR U20189 ( .A(n20500), .B(n20403), .Z(n20503) );
  XNOR U20190 ( .A(n20500), .B(n20357), .Z(n20502) );
  XOR U20191 ( .A(n20504), .B(n20505), .Z(n20500) );
  AND U20192 ( .A(n20506), .B(n20507), .Z(n20505) );
  XOR U20193 ( .A(n20504), .B(n20367), .Z(n20506) );
  XOR U20194 ( .A(n20508), .B(n20509), .Z(n20346) );
  AND U20195 ( .A(n296), .B(n20499), .Z(n20509) );
  XNOR U20196 ( .A(n20497), .B(n20508), .Z(n20499) );
  XNOR U20197 ( .A(n20510), .B(n20511), .Z(n296) );
  AND U20198 ( .A(n20512), .B(n20513), .Z(n20511) );
  XNOR U20199 ( .A(n20514), .B(n20510), .Z(n20513) );
  IV U20200 ( .A(n20403), .Z(n20514) );
  XNOR U20201 ( .A(n20515), .B(n20516), .Z(n20403) );
  AND U20202 ( .A(n299), .B(n20517), .Z(n20516) );
  XNOR U20203 ( .A(n20515), .B(n20518), .Z(n20517) );
  XNOR U20204 ( .A(n20357), .B(n20510), .Z(n20512) );
  XOR U20205 ( .A(n20519), .B(n20520), .Z(n20357) );
  AND U20206 ( .A(n307), .B(n20521), .Z(n20520) );
  XOR U20207 ( .A(n20504), .B(n20522), .Z(n20510) );
  AND U20208 ( .A(n20523), .B(n20507), .Z(n20522) );
  XNOR U20209 ( .A(n20416), .B(n20504), .Z(n20507) );
  XNOR U20210 ( .A(n20524), .B(n20525), .Z(n20416) );
  AND U20211 ( .A(n299), .B(n20526), .Z(n20525) );
  XOR U20212 ( .A(n20527), .B(n20524), .Z(n20526) );
  XNOR U20213 ( .A(n20528), .B(n20504), .Z(n20523) );
  IV U20214 ( .A(n20367), .Z(n20528) );
  XOR U20215 ( .A(n20529), .B(n20530), .Z(n20367) );
  AND U20216 ( .A(n307), .B(n20531), .Z(n20530) );
  XOR U20217 ( .A(n20532), .B(n20533), .Z(n20504) );
  AND U20218 ( .A(n20534), .B(n20535), .Z(n20533) );
  XNOR U20219 ( .A(n20441), .B(n20532), .Z(n20535) );
  XNOR U20220 ( .A(n20536), .B(n20537), .Z(n20441) );
  AND U20221 ( .A(n299), .B(n20538), .Z(n20537) );
  XNOR U20222 ( .A(n20539), .B(n20536), .Z(n20538) );
  XOR U20223 ( .A(n20532), .B(n20378), .Z(n20534) );
  XOR U20224 ( .A(n20540), .B(n20541), .Z(n20378) );
  AND U20225 ( .A(n307), .B(n20542), .Z(n20541) );
  XOR U20226 ( .A(n20543), .B(n20544), .Z(n20532) );
  AND U20227 ( .A(n20545), .B(n20546), .Z(n20544) );
  XNOR U20228 ( .A(n20543), .B(n20487), .Z(n20546) );
  XNOR U20229 ( .A(n20547), .B(n20548), .Z(n20487) );
  AND U20230 ( .A(n299), .B(n20549), .Z(n20548) );
  XOR U20231 ( .A(n20550), .B(n20547), .Z(n20549) );
  XNOR U20232 ( .A(n20551), .B(n20543), .Z(n20545) );
  IV U20233 ( .A(n20390), .Z(n20551) );
  XOR U20234 ( .A(n20552), .B(n20553), .Z(n20390) );
  AND U20235 ( .A(n307), .B(n20554), .Z(n20553) );
  AND U20236 ( .A(n20508), .B(n20497), .Z(n20543) );
  XNOR U20237 ( .A(n20555), .B(n20556), .Z(n20497) );
  AND U20238 ( .A(n299), .B(n20557), .Z(n20556) );
  XNOR U20239 ( .A(n20558), .B(n20555), .Z(n20557) );
  XNOR U20240 ( .A(n20559), .B(n20560), .Z(n299) );
  AND U20241 ( .A(n20561), .B(n20562), .Z(n20560) );
  XOR U20242 ( .A(n20518), .B(n20559), .Z(n20562) );
  AND U20243 ( .A(n20563), .B(n20564), .Z(n20518) );
  XOR U20244 ( .A(n20559), .B(n20515), .Z(n20561) );
  XNOR U20245 ( .A(n20565), .B(n20566), .Z(n20515) );
  AND U20246 ( .A(n303), .B(n20521), .Z(n20566) );
  XOR U20247 ( .A(n20519), .B(n20565), .Z(n20521) );
  XOR U20248 ( .A(n20567), .B(n20568), .Z(n20559) );
  AND U20249 ( .A(n20569), .B(n20570), .Z(n20568) );
  XNOR U20250 ( .A(n20567), .B(n20563), .Z(n20570) );
  IV U20251 ( .A(n20527), .Z(n20563) );
  XOR U20252 ( .A(n20571), .B(n20572), .Z(n20527) );
  XOR U20253 ( .A(n20573), .B(n20564), .Z(n20572) );
  AND U20254 ( .A(n20539), .B(n20574), .Z(n20564) );
  AND U20255 ( .A(n20575), .B(n20576), .Z(n20573) );
  XOR U20256 ( .A(n20577), .B(n20571), .Z(n20575) );
  XNOR U20257 ( .A(n20524), .B(n20567), .Z(n20569) );
  XNOR U20258 ( .A(n20578), .B(n20579), .Z(n20524) );
  AND U20259 ( .A(n303), .B(n20531), .Z(n20579) );
  XOR U20260 ( .A(n20578), .B(n20529), .Z(n20531) );
  XOR U20261 ( .A(n20580), .B(n20581), .Z(n20567) );
  AND U20262 ( .A(n20582), .B(n20583), .Z(n20581) );
  XNOR U20263 ( .A(n20580), .B(n20539), .Z(n20583) );
  XOR U20264 ( .A(n20584), .B(n20576), .Z(n20539) );
  XNOR U20265 ( .A(n20585), .B(n20571), .Z(n20576) );
  XOR U20266 ( .A(n20586), .B(n20587), .Z(n20571) );
  AND U20267 ( .A(n20588), .B(n20589), .Z(n20587) );
  XOR U20268 ( .A(n20590), .B(n20586), .Z(n20588) );
  XNOR U20269 ( .A(n20591), .B(n20592), .Z(n20585) );
  AND U20270 ( .A(n20593), .B(n20594), .Z(n20592) );
  XOR U20271 ( .A(n20591), .B(n20595), .Z(n20593) );
  XNOR U20272 ( .A(n20577), .B(n20574), .Z(n20584) );
  AND U20273 ( .A(n20596), .B(n20597), .Z(n20574) );
  XOR U20274 ( .A(n20598), .B(n20599), .Z(n20577) );
  AND U20275 ( .A(n20600), .B(n20601), .Z(n20599) );
  XOR U20276 ( .A(n20598), .B(n20602), .Z(n20600) );
  XNOR U20277 ( .A(n20536), .B(n20580), .Z(n20582) );
  XNOR U20278 ( .A(n20603), .B(n20604), .Z(n20536) );
  AND U20279 ( .A(n303), .B(n20542), .Z(n20604) );
  XOR U20280 ( .A(n20603), .B(n20540), .Z(n20542) );
  XOR U20281 ( .A(n20605), .B(n20606), .Z(n20580) );
  AND U20282 ( .A(n20607), .B(n20608), .Z(n20606) );
  XNOR U20283 ( .A(n20605), .B(n20596), .Z(n20608) );
  IV U20284 ( .A(n20550), .Z(n20596) );
  XNOR U20285 ( .A(n20609), .B(n20589), .Z(n20550) );
  XNOR U20286 ( .A(n20610), .B(n20595), .Z(n20589) );
  XOR U20287 ( .A(n20611), .B(n20612), .Z(n20595) );
  NOR U20288 ( .A(n20613), .B(n20614), .Z(n20612) );
  XNOR U20289 ( .A(n20611), .B(n20615), .Z(n20613) );
  XNOR U20290 ( .A(n20594), .B(n20586), .Z(n20610) );
  XOR U20291 ( .A(n20616), .B(n20617), .Z(n20586) );
  AND U20292 ( .A(n20618), .B(n20619), .Z(n20617) );
  XNOR U20293 ( .A(n20616), .B(n20620), .Z(n20618) );
  XNOR U20294 ( .A(n20621), .B(n20591), .Z(n20594) );
  XOR U20295 ( .A(n20622), .B(n20623), .Z(n20591) );
  AND U20296 ( .A(n20624), .B(n20625), .Z(n20623) );
  XOR U20297 ( .A(n20622), .B(n20626), .Z(n20624) );
  XNOR U20298 ( .A(n20627), .B(n20628), .Z(n20621) );
  NOR U20299 ( .A(n20629), .B(n20630), .Z(n20628) );
  XOR U20300 ( .A(n20627), .B(n20631), .Z(n20629) );
  XNOR U20301 ( .A(n20590), .B(n20597), .Z(n20609) );
  NOR U20302 ( .A(n20558), .B(n20632), .Z(n20597) );
  XOR U20303 ( .A(n20602), .B(n20601), .Z(n20590) );
  XNOR U20304 ( .A(n20633), .B(n20598), .Z(n20601) );
  XOR U20305 ( .A(n20634), .B(n20635), .Z(n20598) );
  AND U20306 ( .A(n20636), .B(n20637), .Z(n20635) );
  XOR U20307 ( .A(n20634), .B(n20638), .Z(n20636) );
  XNOR U20308 ( .A(n20639), .B(n20640), .Z(n20633) );
  NOR U20309 ( .A(n20641), .B(n20642), .Z(n20640) );
  XNOR U20310 ( .A(n20639), .B(n20643), .Z(n20641) );
  XOR U20311 ( .A(n20644), .B(n20645), .Z(n20602) );
  NOR U20312 ( .A(n20646), .B(n20647), .Z(n20645) );
  XNOR U20313 ( .A(n20644), .B(n20648), .Z(n20646) );
  XNOR U20314 ( .A(n20547), .B(n20605), .Z(n20607) );
  XNOR U20315 ( .A(n20649), .B(n20650), .Z(n20547) );
  AND U20316 ( .A(n303), .B(n20554), .Z(n20650) );
  XOR U20317 ( .A(n20649), .B(n20552), .Z(n20554) );
  AND U20318 ( .A(n20555), .B(n20558), .Z(n20605) );
  XOR U20319 ( .A(n20651), .B(n20632), .Z(n20558) );
  XNOR U20320 ( .A(p_input[2048]), .B(p_input[384]), .Z(n20632) );
  XOR U20321 ( .A(n20620), .B(n20619), .Z(n20651) );
  XNOR U20322 ( .A(n20652), .B(n20626), .Z(n20619) );
  XNOR U20323 ( .A(n20615), .B(n20614), .Z(n20626) );
  XOR U20324 ( .A(n20653), .B(n20611), .Z(n20614) );
  XNOR U20325 ( .A(n16904), .B(p_input[394]), .Z(n20611) );
  XNOR U20326 ( .A(p_input[2059]), .B(p_input[395]), .Z(n20653) );
  XOR U20327 ( .A(p_input[2060]), .B(p_input[396]), .Z(n20615) );
  XNOR U20328 ( .A(n20625), .B(n20616), .Z(n20652) );
  XNOR U20329 ( .A(n17068), .B(p_input[385]), .Z(n20616) );
  XOR U20330 ( .A(n20654), .B(n20631), .Z(n20625) );
  XNOR U20331 ( .A(p_input[2063]), .B(p_input[399]), .Z(n20631) );
  XOR U20332 ( .A(n20622), .B(n20630), .Z(n20654) );
  XOR U20333 ( .A(n20655), .B(n20627), .Z(n20630) );
  XOR U20334 ( .A(p_input[2061]), .B(p_input[397]), .Z(n20627) );
  XNOR U20335 ( .A(p_input[2062]), .B(p_input[398]), .Z(n20655) );
  XNOR U20336 ( .A(n16738), .B(p_input[393]), .Z(n20622) );
  XNOR U20337 ( .A(n20638), .B(n20637), .Z(n20620) );
  XNOR U20338 ( .A(n20656), .B(n20643), .Z(n20637) );
  XOR U20339 ( .A(p_input[2056]), .B(p_input[392]), .Z(n20643) );
  XOR U20340 ( .A(n20634), .B(n20642), .Z(n20656) );
  XOR U20341 ( .A(n20657), .B(n20639), .Z(n20642) );
  XOR U20342 ( .A(p_input[2054]), .B(p_input[390]), .Z(n20639) );
  XNOR U20343 ( .A(p_input[2055]), .B(p_input[391]), .Z(n20657) );
  XNOR U20344 ( .A(n16741), .B(p_input[386]), .Z(n20634) );
  XNOR U20345 ( .A(n20648), .B(n20647), .Z(n20638) );
  XOR U20346 ( .A(n20658), .B(n20644), .Z(n20647) );
  XOR U20347 ( .A(p_input[2051]), .B(p_input[387]), .Z(n20644) );
  XNOR U20348 ( .A(p_input[2052]), .B(p_input[388]), .Z(n20658) );
  XOR U20349 ( .A(p_input[2053]), .B(p_input[389]), .Z(n20648) );
  XNOR U20350 ( .A(n20659), .B(n20660), .Z(n20555) );
  AND U20351 ( .A(n303), .B(n20661), .Z(n20660) );
  XNOR U20352 ( .A(n20662), .B(n20663), .Z(n303) );
  AND U20353 ( .A(n20664), .B(n20665), .Z(n20663) );
  XOR U20354 ( .A(n20662), .B(n20565), .Z(n20665) );
  XNOR U20355 ( .A(n20662), .B(n20519), .Z(n20664) );
  XOR U20356 ( .A(n20666), .B(n20667), .Z(n20662) );
  AND U20357 ( .A(n20668), .B(n20669), .Z(n20667) );
  XOR U20358 ( .A(n20666), .B(n20529), .Z(n20668) );
  XOR U20359 ( .A(n20670), .B(n20671), .Z(n20508) );
  AND U20360 ( .A(n307), .B(n20661), .Z(n20671) );
  XNOR U20361 ( .A(n20659), .B(n20670), .Z(n20661) );
  XNOR U20362 ( .A(n20672), .B(n20673), .Z(n307) );
  AND U20363 ( .A(n20674), .B(n20675), .Z(n20673) );
  XNOR U20364 ( .A(n20676), .B(n20672), .Z(n20675) );
  IV U20365 ( .A(n20565), .Z(n20676) );
  XNOR U20366 ( .A(n20677), .B(n20678), .Z(n20565) );
  AND U20367 ( .A(n310), .B(n20679), .Z(n20678) );
  XNOR U20368 ( .A(n20677), .B(n20680), .Z(n20679) );
  XNOR U20369 ( .A(n20519), .B(n20672), .Z(n20674) );
  XOR U20370 ( .A(n20681), .B(n20682), .Z(n20519) );
  AND U20371 ( .A(n318), .B(n20683), .Z(n20682) );
  XOR U20372 ( .A(n20666), .B(n20684), .Z(n20672) );
  AND U20373 ( .A(n20685), .B(n20669), .Z(n20684) );
  XNOR U20374 ( .A(n20578), .B(n20666), .Z(n20669) );
  XNOR U20375 ( .A(n20686), .B(n20687), .Z(n20578) );
  AND U20376 ( .A(n310), .B(n20688), .Z(n20687) );
  XOR U20377 ( .A(n20689), .B(n20686), .Z(n20688) );
  XNOR U20378 ( .A(n20690), .B(n20666), .Z(n20685) );
  IV U20379 ( .A(n20529), .Z(n20690) );
  XOR U20380 ( .A(n20691), .B(n20692), .Z(n20529) );
  AND U20381 ( .A(n318), .B(n20693), .Z(n20692) );
  XOR U20382 ( .A(n20694), .B(n20695), .Z(n20666) );
  AND U20383 ( .A(n20696), .B(n20697), .Z(n20695) );
  XNOR U20384 ( .A(n20603), .B(n20694), .Z(n20697) );
  XNOR U20385 ( .A(n20698), .B(n20699), .Z(n20603) );
  AND U20386 ( .A(n310), .B(n20700), .Z(n20699) );
  XNOR U20387 ( .A(n20701), .B(n20698), .Z(n20700) );
  XOR U20388 ( .A(n20694), .B(n20540), .Z(n20696) );
  XOR U20389 ( .A(n20702), .B(n20703), .Z(n20540) );
  AND U20390 ( .A(n318), .B(n20704), .Z(n20703) );
  XOR U20391 ( .A(n20705), .B(n20706), .Z(n20694) );
  AND U20392 ( .A(n20707), .B(n20708), .Z(n20706) );
  XNOR U20393 ( .A(n20705), .B(n20649), .Z(n20708) );
  XNOR U20394 ( .A(n20709), .B(n20710), .Z(n20649) );
  AND U20395 ( .A(n310), .B(n20711), .Z(n20710) );
  XOR U20396 ( .A(n20712), .B(n20709), .Z(n20711) );
  XNOR U20397 ( .A(n20713), .B(n20705), .Z(n20707) );
  IV U20398 ( .A(n20552), .Z(n20713) );
  XOR U20399 ( .A(n20714), .B(n20715), .Z(n20552) );
  AND U20400 ( .A(n318), .B(n20716), .Z(n20715) );
  AND U20401 ( .A(n20670), .B(n20659), .Z(n20705) );
  XNOR U20402 ( .A(n20717), .B(n20718), .Z(n20659) );
  AND U20403 ( .A(n310), .B(n20719), .Z(n20718) );
  XNOR U20404 ( .A(n20720), .B(n20717), .Z(n20719) );
  XNOR U20405 ( .A(n20721), .B(n20722), .Z(n310) );
  AND U20406 ( .A(n20723), .B(n20724), .Z(n20722) );
  XOR U20407 ( .A(n20680), .B(n20721), .Z(n20724) );
  AND U20408 ( .A(n20725), .B(n20726), .Z(n20680) );
  XOR U20409 ( .A(n20721), .B(n20677), .Z(n20723) );
  XNOR U20410 ( .A(n20727), .B(n20728), .Z(n20677) );
  AND U20411 ( .A(n314), .B(n20683), .Z(n20728) );
  XOR U20412 ( .A(n20681), .B(n20727), .Z(n20683) );
  XOR U20413 ( .A(n20729), .B(n20730), .Z(n20721) );
  AND U20414 ( .A(n20731), .B(n20732), .Z(n20730) );
  XNOR U20415 ( .A(n20729), .B(n20725), .Z(n20732) );
  IV U20416 ( .A(n20689), .Z(n20725) );
  XOR U20417 ( .A(n20733), .B(n20734), .Z(n20689) );
  XOR U20418 ( .A(n20735), .B(n20726), .Z(n20734) );
  AND U20419 ( .A(n20701), .B(n20736), .Z(n20726) );
  AND U20420 ( .A(n20737), .B(n20738), .Z(n20735) );
  XOR U20421 ( .A(n20739), .B(n20733), .Z(n20737) );
  XNOR U20422 ( .A(n20686), .B(n20729), .Z(n20731) );
  XNOR U20423 ( .A(n20740), .B(n20741), .Z(n20686) );
  AND U20424 ( .A(n314), .B(n20693), .Z(n20741) );
  XOR U20425 ( .A(n20740), .B(n20691), .Z(n20693) );
  XOR U20426 ( .A(n20742), .B(n20743), .Z(n20729) );
  AND U20427 ( .A(n20744), .B(n20745), .Z(n20743) );
  XNOR U20428 ( .A(n20742), .B(n20701), .Z(n20745) );
  XOR U20429 ( .A(n20746), .B(n20738), .Z(n20701) );
  XNOR U20430 ( .A(n20747), .B(n20733), .Z(n20738) );
  XOR U20431 ( .A(n20748), .B(n20749), .Z(n20733) );
  AND U20432 ( .A(n20750), .B(n20751), .Z(n20749) );
  XOR U20433 ( .A(n20752), .B(n20748), .Z(n20750) );
  XNOR U20434 ( .A(n20753), .B(n20754), .Z(n20747) );
  AND U20435 ( .A(n20755), .B(n20756), .Z(n20754) );
  XOR U20436 ( .A(n20753), .B(n20757), .Z(n20755) );
  XNOR U20437 ( .A(n20739), .B(n20736), .Z(n20746) );
  AND U20438 ( .A(n20758), .B(n20759), .Z(n20736) );
  XOR U20439 ( .A(n20760), .B(n20761), .Z(n20739) );
  AND U20440 ( .A(n20762), .B(n20763), .Z(n20761) );
  XOR U20441 ( .A(n20760), .B(n20764), .Z(n20762) );
  XNOR U20442 ( .A(n20698), .B(n20742), .Z(n20744) );
  XNOR U20443 ( .A(n20765), .B(n20766), .Z(n20698) );
  AND U20444 ( .A(n314), .B(n20704), .Z(n20766) );
  XOR U20445 ( .A(n20765), .B(n20702), .Z(n20704) );
  XOR U20446 ( .A(n20767), .B(n20768), .Z(n20742) );
  AND U20447 ( .A(n20769), .B(n20770), .Z(n20768) );
  XNOR U20448 ( .A(n20767), .B(n20758), .Z(n20770) );
  IV U20449 ( .A(n20712), .Z(n20758) );
  XNOR U20450 ( .A(n20771), .B(n20751), .Z(n20712) );
  XNOR U20451 ( .A(n20772), .B(n20757), .Z(n20751) );
  XOR U20452 ( .A(n20773), .B(n20774), .Z(n20757) );
  NOR U20453 ( .A(n20775), .B(n20776), .Z(n20774) );
  XNOR U20454 ( .A(n20773), .B(n20777), .Z(n20775) );
  XNOR U20455 ( .A(n20756), .B(n20748), .Z(n20772) );
  XOR U20456 ( .A(n20778), .B(n20779), .Z(n20748) );
  AND U20457 ( .A(n20780), .B(n20781), .Z(n20779) );
  XNOR U20458 ( .A(n20778), .B(n20782), .Z(n20780) );
  XNOR U20459 ( .A(n20783), .B(n20753), .Z(n20756) );
  XOR U20460 ( .A(n20784), .B(n20785), .Z(n20753) );
  AND U20461 ( .A(n20786), .B(n20787), .Z(n20785) );
  XOR U20462 ( .A(n20784), .B(n20788), .Z(n20786) );
  XNOR U20463 ( .A(n20789), .B(n20790), .Z(n20783) );
  NOR U20464 ( .A(n20791), .B(n20792), .Z(n20790) );
  XOR U20465 ( .A(n20789), .B(n20793), .Z(n20791) );
  XNOR U20466 ( .A(n20752), .B(n20759), .Z(n20771) );
  NOR U20467 ( .A(n20720), .B(n20794), .Z(n20759) );
  XOR U20468 ( .A(n20764), .B(n20763), .Z(n20752) );
  XNOR U20469 ( .A(n20795), .B(n20760), .Z(n20763) );
  XOR U20470 ( .A(n20796), .B(n20797), .Z(n20760) );
  AND U20471 ( .A(n20798), .B(n20799), .Z(n20797) );
  XOR U20472 ( .A(n20796), .B(n20800), .Z(n20798) );
  XNOR U20473 ( .A(n20801), .B(n20802), .Z(n20795) );
  NOR U20474 ( .A(n20803), .B(n20804), .Z(n20802) );
  XNOR U20475 ( .A(n20801), .B(n20805), .Z(n20803) );
  XOR U20476 ( .A(n20806), .B(n20807), .Z(n20764) );
  NOR U20477 ( .A(n20808), .B(n20809), .Z(n20807) );
  XNOR U20478 ( .A(n20806), .B(n20810), .Z(n20808) );
  XNOR U20479 ( .A(n20709), .B(n20767), .Z(n20769) );
  XNOR U20480 ( .A(n20811), .B(n20812), .Z(n20709) );
  AND U20481 ( .A(n314), .B(n20716), .Z(n20812) );
  XOR U20482 ( .A(n20811), .B(n20714), .Z(n20716) );
  AND U20483 ( .A(n20717), .B(n20720), .Z(n20767) );
  XOR U20484 ( .A(n20813), .B(n20794), .Z(n20720) );
  XNOR U20485 ( .A(p_input[2048]), .B(p_input[400]), .Z(n20794) );
  XOR U20486 ( .A(n20782), .B(n20781), .Z(n20813) );
  XNOR U20487 ( .A(n20814), .B(n20788), .Z(n20781) );
  XNOR U20488 ( .A(n20777), .B(n20776), .Z(n20788) );
  XOR U20489 ( .A(n20815), .B(n20773), .Z(n20776) );
  XNOR U20490 ( .A(n16904), .B(p_input[410]), .Z(n20773) );
  XNOR U20491 ( .A(p_input[2059]), .B(p_input[411]), .Z(n20815) );
  XOR U20492 ( .A(p_input[2060]), .B(p_input[412]), .Z(n20777) );
  XNOR U20493 ( .A(n20787), .B(n20778), .Z(n20814) );
  XNOR U20494 ( .A(n17068), .B(p_input[401]), .Z(n20778) );
  XOR U20495 ( .A(n20816), .B(n20793), .Z(n20787) );
  XNOR U20496 ( .A(p_input[2063]), .B(p_input[415]), .Z(n20793) );
  XOR U20497 ( .A(n20784), .B(n20792), .Z(n20816) );
  XOR U20498 ( .A(n20817), .B(n20789), .Z(n20792) );
  XOR U20499 ( .A(p_input[2061]), .B(p_input[413]), .Z(n20789) );
  XNOR U20500 ( .A(p_input[2062]), .B(p_input[414]), .Z(n20817) );
  XNOR U20501 ( .A(n16738), .B(p_input[409]), .Z(n20784) );
  XNOR U20502 ( .A(n20800), .B(n20799), .Z(n20782) );
  XNOR U20503 ( .A(n20818), .B(n20805), .Z(n20799) );
  XOR U20504 ( .A(p_input[2056]), .B(p_input[408]), .Z(n20805) );
  XOR U20505 ( .A(n20796), .B(n20804), .Z(n20818) );
  XOR U20506 ( .A(n20819), .B(n20801), .Z(n20804) );
  XOR U20507 ( .A(p_input[2054]), .B(p_input[406]), .Z(n20801) );
  XNOR U20508 ( .A(p_input[2055]), .B(p_input[407]), .Z(n20819) );
  XNOR U20509 ( .A(n16741), .B(p_input[402]), .Z(n20796) );
  XNOR U20510 ( .A(n20810), .B(n20809), .Z(n20800) );
  XOR U20511 ( .A(n20820), .B(n20806), .Z(n20809) );
  XOR U20512 ( .A(p_input[2051]), .B(p_input[403]), .Z(n20806) );
  XNOR U20513 ( .A(p_input[2052]), .B(p_input[404]), .Z(n20820) );
  XOR U20514 ( .A(p_input[2053]), .B(p_input[405]), .Z(n20810) );
  XNOR U20515 ( .A(n20821), .B(n20822), .Z(n20717) );
  AND U20516 ( .A(n314), .B(n20823), .Z(n20822) );
  XNOR U20517 ( .A(n20824), .B(n20825), .Z(n314) );
  AND U20518 ( .A(n20826), .B(n20827), .Z(n20825) );
  XOR U20519 ( .A(n20824), .B(n20727), .Z(n20827) );
  XNOR U20520 ( .A(n20824), .B(n20681), .Z(n20826) );
  XOR U20521 ( .A(n20828), .B(n20829), .Z(n20824) );
  AND U20522 ( .A(n20830), .B(n20831), .Z(n20829) );
  XOR U20523 ( .A(n20828), .B(n20691), .Z(n20830) );
  XOR U20524 ( .A(n20832), .B(n20833), .Z(n20670) );
  AND U20525 ( .A(n318), .B(n20823), .Z(n20833) );
  XNOR U20526 ( .A(n20821), .B(n20832), .Z(n20823) );
  XNOR U20527 ( .A(n20834), .B(n20835), .Z(n318) );
  AND U20528 ( .A(n20836), .B(n20837), .Z(n20835) );
  XNOR U20529 ( .A(n20838), .B(n20834), .Z(n20837) );
  IV U20530 ( .A(n20727), .Z(n20838) );
  XNOR U20531 ( .A(n20839), .B(n20840), .Z(n20727) );
  AND U20532 ( .A(n321), .B(n20841), .Z(n20840) );
  XNOR U20533 ( .A(n20839), .B(n20842), .Z(n20841) );
  XNOR U20534 ( .A(n20681), .B(n20834), .Z(n20836) );
  XOR U20535 ( .A(n20843), .B(n20844), .Z(n20681) );
  AND U20536 ( .A(n329), .B(n20845), .Z(n20844) );
  XOR U20537 ( .A(n20828), .B(n20846), .Z(n20834) );
  AND U20538 ( .A(n20847), .B(n20831), .Z(n20846) );
  XNOR U20539 ( .A(n20740), .B(n20828), .Z(n20831) );
  XNOR U20540 ( .A(n20848), .B(n20849), .Z(n20740) );
  AND U20541 ( .A(n321), .B(n20850), .Z(n20849) );
  XOR U20542 ( .A(n20851), .B(n20848), .Z(n20850) );
  XNOR U20543 ( .A(n20852), .B(n20828), .Z(n20847) );
  IV U20544 ( .A(n20691), .Z(n20852) );
  XOR U20545 ( .A(n20853), .B(n20854), .Z(n20691) );
  AND U20546 ( .A(n329), .B(n20855), .Z(n20854) );
  XOR U20547 ( .A(n20856), .B(n20857), .Z(n20828) );
  AND U20548 ( .A(n20858), .B(n20859), .Z(n20857) );
  XNOR U20549 ( .A(n20765), .B(n20856), .Z(n20859) );
  XNOR U20550 ( .A(n20860), .B(n20861), .Z(n20765) );
  AND U20551 ( .A(n321), .B(n20862), .Z(n20861) );
  XNOR U20552 ( .A(n20863), .B(n20860), .Z(n20862) );
  XOR U20553 ( .A(n20856), .B(n20702), .Z(n20858) );
  XOR U20554 ( .A(n20864), .B(n20865), .Z(n20702) );
  AND U20555 ( .A(n329), .B(n20866), .Z(n20865) );
  XOR U20556 ( .A(n20867), .B(n20868), .Z(n20856) );
  AND U20557 ( .A(n20869), .B(n20870), .Z(n20868) );
  XNOR U20558 ( .A(n20867), .B(n20811), .Z(n20870) );
  XNOR U20559 ( .A(n20871), .B(n20872), .Z(n20811) );
  AND U20560 ( .A(n321), .B(n20873), .Z(n20872) );
  XOR U20561 ( .A(n20874), .B(n20871), .Z(n20873) );
  XNOR U20562 ( .A(n20875), .B(n20867), .Z(n20869) );
  IV U20563 ( .A(n20714), .Z(n20875) );
  XOR U20564 ( .A(n20876), .B(n20877), .Z(n20714) );
  AND U20565 ( .A(n329), .B(n20878), .Z(n20877) );
  AND U20566 ( .A(n20832), .B(n20821), .Z(n20867) );
  XNOR U20567 ( .A(n20879), .B(n20880), .Z(n20821) );
  AND U20568 ( .A(n321), .B(n20881), .Z(n20880) );
  XNOR U20569 ( .A(n20882), .B(n20879), .Z(n20881) );
  XNOR U20570 ( .A(n20883), .B(n20884), .Z(n321) );
  AND U20571 ( .A(n20885), .B(n20886), .Z(n20884) );
  XOR U20572 ( .A(n20842), .B(n20883), .Z(n20886) );
  AND U20573 ( .A(n20887), .B(n20888), .Z(n20842) );
  XOR U20574 ( .A(n20883), .B(n20839), .Z(n20885) );
  XNOR U20575 ( .A(n20889), .B(n20890), .Z(n20839) );
  AND U20576 ( .A(n325), .B(n20845), .Z(n20890) );
  XOR U20577 ( .A(n20843), .B(n20889), .Z(n20845) );
  XOR U20578 ( .A(n20891), .B(n20892), .Z(n20883) );
  AND U20579 ( .A(n20893), .B(n20894), .Z(n20892) );
  XNOR U20580 ( .A(n20891), .B(n20887), .Z(n20894) );
  IV U20581 ( .A(n20851), .Z(n20887) );
  XOR U20582 ( .A(n20895), .B(n20896), .Z(n20851) );
  XOR U20583 ( .A(n20897), .B(n20888), .Z(n20896) );
  AND U20584 ( .A(n20863), .B(n20898), .Z(n20888) );
  AND U20585 ( .A(n20899), .B(n20900), .Z(n20897) );
  XOR U20586 ( .A(n20901), .B(n20895), .Z(n20899) );
  XNOR U20587 ( .A(n20848), .B(n20891), .Z(n20893) );
  XNOR U20588 ( .A(n20902), .B(n20903), .Z(n20848) );
  AND U20589 ( .A(n325), .B(n20855), .Z(n20903) );
  XOR U20590 ( .A(n20902), .B(n20853), .Z(n20855) );
  XOR U20591 ( .A(n20904), .B(n20905), .Z(n20891) );
  AND U20592 ( .A(n20906), .B(n20907), .Z(n20905) );
  XNOR U20593 ( .A(n20904), .B(n20863), .Z(n20907) );
  XOR U20594 ( .A(n20908), .B(n20900), .Z(n20863) );
  XNOR U20595 ( .A(n20909), .B(n20895), .Z(n20900) );
  XOR U20596 ( .A(n20910), .B(n20911), .Z(n20895) );
  AND U20597 ( .A(n20912), .B(n20913), .Z(n20911) );
  XOR U20598 ( .A(n20914), .B(n20910), .Z(n20912) );
  XNOR U20599 ( .A(n20915), .B(n20916), .Z(n20909) );
  AND U20600 ( .A(n20917), .B(n20918), .Z(n20916) );
  XOR U20601 ( .A(n20915), .B(n20919), .Z(n20917) );
  XNOR U20602 ( .A(n20901), .B(n20898), .Z(n20908) );
  AND U20603 ( .A(n20920), .B(n20921), .Z(n20898) );
  XOR U20604 ( .A(n20922), .B(n20923), .Z(n20901) );
  AND U20605 ( .A(n20924), .B(n20925), .Z(n20923) );
  XOR U20606 ( .A(n20922), .B(n20926), .Z(n20924) );
  XNOR U20607 ( .A(n20860), .B(n20904), .Z(n20906) );
  XNOR U20608 ( .A(n20927), .B(n20928), .Z(n20860) );
  AND U20609 ( .A(n325), .B(n20866), .Z(n20928) );
  XOR U20610 ( .A(n20927), .B(n20864), .Z(n20866) );
  XOR U20611 ( .A(n20929), .B(n20930), .Z(n20904) );
  AND U20612 ( .A(n20931), .B(n20932), .Z(n20930) );
  XNOR U20613 ( .A(n20929), .B(n20920), .Z(n20932) );
  IV U20614 ( .A(n20874), .Z(n20920) );
  XNOR U20615 ( .A(n20933), .B(n20913), .Z(n20874) );
  XNOR U20616 ( .A(n20934), .B(n20919), .Z(n20913) );
  XOR U20617 ( .A(n20935), .B(n20936), .Z(n20919) );
  NOR U20618 ( .A(n20937), .B(n20938), .Z(n20936) );
  XNOR U20619 ( .A(n20935), .B(n20939), .Z(n20937) );
  XNOR U20620 ( .A(n20918), .B(n20910), .Z(n20934) );
  XOR U20621 ( .A(n20940), .B(n20941), .Z(n20910) );
  AND U20622 ( .A(n20942), .B(n20943), .Z(n20941) );
  XNOR U20623 ( .A(n20940), .B(n20944), .Z(n20942) );
  XNOR U20624 ( .A(n20945), .B(n20915), .Z(n20918) );
  XOR U20625 ( .A(n20946), .B(n20947), .Z(n20915) );
  AND U20626 ( .A(n20948), .B(n20949), .Z(n20947) );
  XOR U20627 ( .A(n20946), .B(n20950), .Z(n20948) );
  XNOR U20628 ( .A(n20951), .B(n20952), .Z(n20945) );
  NOR U20629 ( .A(n20953), .B(n20954), .Z(n20952) );
  XOR U20630 ( .A(n20951), .B(n20955), .Z(n20953) );
  XNOR U20631 ( .A(n20914), .B(n20921), .Z(n20933) );
  NOR U20632 ( .A(n20882), .B(n20956), .Z(n20921) );
  XOR U20633 ( .A(n20926), .B(n20925), .Z(n20914) );
  XNOR U20634 ( .A(n20957), .B(n20922), .Z(n20925) );
  XOR U20635 ( .A(n20958), .B(n20959), .Z(n20922) );
  AND U20636 ( .A(n20960), .B(n20961), .Z(n20959) );
  XOR U20637 ( .A(n20958), .B(n20962), .Z(n20960) );
  XNOR U20638 ( .A(n20963), .B(n20964), .Z(n20957) );
  NOR U20639 ( .A(n20965), .B(n20966), .Z(n20964) );
  XNOR U20640 ( .A(n20963), .B(n20967), .Z(n20965) );
  XOR U20641 ( .A(n20968), .B(n20969), .Z(n20926) );
  NOR U20642 ( .A(n20970), .B(n20971), .Z(n20969) );
  XNOR U20643 ( .A(n20968), .B(n20972), .Z(n20970) );
  XNOR U20644 ( .A(n20871), .B(n20929), .Z(n20931) );
  XNOR U20645 ( .A(n20973), .B(n20974), .Z(n20871) );
  AND U20646 ( .A(n325), .B(n20878), .Z(n20974) );
  XOR U20647 ( .A(n20973), .B(n20876), .Z(n20878) );
  AND U20648 ( .A(n20879), .B(n20882), .Z(n20929) );
  XOR U20649 ( .A(n20975), .B(n20956), .Z(n20882) );
  XNOR U20650 ( .A(p_input[2048]), .B(p_input[416]), .Z(n20956) );
  XOR U20651 ( .A(n20944), .B(n20943), .Z(n20975) );
  XNOR U20652 ( .A(n20976), .B(n20950), .Z(n20943) );
  XNOR U20653 ( .A(n20939), .B(n20938), .Z(n20950) );
  XOR U20654 ( .A(n20977), .B(n20935), .Z(n20938) );
  XNOR U20655 ( .A(n16904), .B(p_input[426]), .Z(n20935) );
  XNOR U20656 ( .A(p_input[2059]), .B(p_input[427]), .Z(n20977) );
  XOR U20657 ( .A(p_input[2060]), .B(p_input[428]), .Z(n20939) );
  XNOR U20658 ( .A(n20949), .B(n20940), .Z(n20976) );
  XNOR U20659 ( .A(n17068), .B(p_input[417]), .Z(n20940) );
  XOR U20660 ( .A(n20978), .B(n20955), .Z(n20949) );
  XNOR U20661 ( .A(p_input[2063]), .B(p_input[431]), .Z(n20955) );
  XOR U20662 ( .A(n20946), .B(n20954), .Z(n20978) );
  XOR U20663 ( .A(n20979), .B(n20951), .Z(n20954) );
  XOR U20664 ( .A(p_input[2061]), .B(p_input[429]), .Z(n20951) );
  XNOR U20665 ( .A(p_input[2062]), .B(p_input[430]), .Z(n20979) );
  XNOR U20666 ( .A(n16738), .B(p_input[425]), .Z(n20946) );
  XNOR U20667 ( .A(n20962), .B(n20961), .Z(n20944) );
  XNOR U20668 ( .A(n20980), .B(n20967), .Z(n20961) );
  XOR U20669 ( .A(p_input[2056]), .B(p_input[424]), .Z(n20967) );
  XOR U20670 ( .A(n20958), .B(n20966), .Z(n20980) );
  XOR U20671 ( .A(n20981), .B(n20963), .Z(n20966) );
  XOR U20672 ( .A(p_input[2054]), .B(p_input[422]), .Z(n20963) );
  XNOR U20673 ( .A(p_input[2055]), .B(p_input[423]), .Z(n20981) );
  XNOR U20674 ( .A(n16741), .B(p_input[418]), .Z(n20958) );
  XNOR U20675 ( .A(n20972), .B(n20971), .Z(n20962) );
  XOR U20676 ( .A(n20982), .B(n20968), .Z(n20971) );
  XOR U20677 ( .A(p_input[2051]), .B(p_input[419]), .Z(n20968) );
  XNOR U20678 ( .A(p_input[2052]), .B(p_input[420]), .Z(n20982) );
  XOR U20679 ( .A(p_input[2053]), .B(p_input[421]), .Z(n20972) );
  XNOR U20680 ( .A(n20983), .B(n20984), .Z(n20879) );
  AND U20681 ( .A(n325), .B(n20985), .Z(n20984) );
  XNOR U20682 ( .A(n20986), .B(n20987), .Z(n325) );
  AND U20683 ( .A(n20988), .B(n20989), .Z(n20987) );
  XOR U20684 ( .A(n20986), .B(n20889), .Z(n20989) );
  XNOR U20685 ( .A(n20986), .B(n20843), .Z(n20988) );
  XOR U20686 ( .A(n20990), .B(n20991), .Z(n20986) );
  AND U20687 ( .A(n20992), .B(n20993), .Z(n20991) );
  XOR U20688 ( .A(n20990), .B(n20853), .Z(n20992) );
  XOR U20689 ( .A(n20994), .B(n20995), .Z(n20832) );
  AND U20690 ( .A(n329), .B(n20985), .Z(n20995) );
  XNOR U20691 ( .A(n20983), .B(n20994), .Z(n20985) );
  XNOR U20692 ( .A(n20996), .B(n20997), .Z(n329) );
  AND U20693 ( .A(n20998), .B(n20999), .Z(n20997) );
  XNOR U20694 ( .A(n21000), .B(n20996), .Z(n20999) );
  IV U20695 ( .A(n20889), .Z(n21000) );
  XNOR U20696 ( .A(n21001), .B(n21002), .Z(n20889) );
  AND U20697 ( .A(n332), .B(n21003), .Z(n21002) );
  XNOR U20698 ( .A(n21001), .B(n21004), .Z(n21003) );
  XNOR U20699 ( .A(n20843), .B(n20996), .Z(n20998) );
  XOR U20700 ( .A(n21005), .B(n21006), .Z(n20843) );
  AND U20701 ( .A(n340), .B(n21007), .Z(n21006) );
  XOR U20702 ( .A(n20990), .B(n21008), .Z(n20996) );
  AND U20703 ( .A(n21009), .B(n20993), .Z(n21008) );
  XNOR U20704 ( .A(n20902), .B(n20990), .Z(n20993) );
  XNOR U20705 ( .A(n21010), .B(n21011), .Z(n20902) );
  AND U20706 ( .A(n332), .B(n21012), .Z(n21011) );
  XOR U20707 ( .A(n21013), .B(n21010), .Z(n21012) );
  XNOR U20708 ( .A(n21014), .B(n20990), .Z(n21009) );
  IV U20709 ( .A(n20853), .Z(n21014) );
  XOR U20710 ( .A(n21015), .B(n21016), .Z(n20853) );
  AND U20711 ( .A(n340), .B(n21017), .Z(n21016) );
  XOR U20712 ( .A(n21018), .B(n21019), .Z(n20990) );
  AND U20713 ( .A(n21020), .B(n21021), .Z(n21019) );
  XNOR U20714 ( .A(n20927), .B(n21018), .Z(n21021) );
  XNOR U20715 ( .A(n21022), .B(n21023), .Z(n20927) );
  AND U20716 ( .A(n332), .B(n21024), .Z(n21023) );
  XNOR U20717 ( .A(n21025), .B(n21022), .Z(n21024) );
  XOR U20718 ( .A(n21018), .B(n20864), .Z(n21020) );
  XOR U20719 ( .A(n21026), .B(n21027), .Z(n20864) );
  AND U20720 ( .A(n340), .B(n21028), .Z(n21027) );
  XOR U20721 ( .A(n21029), .B(n21030), .Z(n21018) );
  AND U20722 ( .A(n21031), .B(n21032), .Z(n21030) );
  XNOR U20723 ( .A(n21029), .B(n20973), .Z(n21032) );
  XNOR U20724 ( .A(n21033), .B(n21034), .Z(n20973) );
  AND U20725 ( .A(n332), .B(n21035), .Z(n21034) );
  XOR U20726 ( .A(n21036), .B(n21033), .Z(n21035) );
  XNOR U20727 ( .A(n21037), .B(n21029), .Z(n21031) );
  IV U20728 ( .A(n20876), .Z(n21037) );
  XOR U20729 ( .A(n21038), .B(n21039), .Z(n20876) );
  AND U20730 ( .A(n340), .B(n21040), .Z(n21039) );
  AND U20731 ( .A(n20994), .B(n20983), .Z(n21029) );
  XNOR U20732 ( .A(n21041), .B(n21042), .Z(n20983) );
  AND U20733 ( .A(n332), .B(n21043), .Z(n21042) );
  XNOR U20734 ( .A(n21044), .B(n21041), .Z(n21043) );
  XNOR U20735 ( .A(n21045), .B(n21046), .Z(n332) );
  AND U20736 ( .A(n21047), .B(n21048), .Z(n21046) );
  XOR U20737 ( .A(n21004), .B(n21045), .Z(n21048) );
  AND U20738 ( .A(n21049), .B(n21050), .Z(n21004) );
  XOR U20739 ( .A(n21045), .B(n21001), .Z(n21047) );
  XNOR U20740 ( .A(n21051), .B(n21052), .Z(n21001) );
  AND U20741 ( .A(n336), .B(n21007), .Z(n21052) );
  XOR U20742 ( .A(n21005), .B(n21051), .Z(n21007) );
  XOR U20743 ( .A(n21053), .B(n21054), .Z(n21045) );
  AND U20744 ( .A(n21055), .B(n21056), .Z(n21054) );
  XNOR U20745 ( .A(n21053), .B(n21049), .Z(n21056) );
  IV U20746 ( .A(n21013), .Z(n21049) );
  XOR U20747 ( .A(n21057), .B(n21058), .Z(n21013) );
  XOR U20748 ( .A(n21059), .B(n21050), .Z(n21058) );
  AND U20749 ( .A(n21025), .B(n21060), .Z(n21050) );
  AND U20750 ( .A(n21061), .B(n21062), .Z(n21059) );
  XOR U20751 ( .A(n21063), .B(n21057), .Z(n21061) );
  XNOR U20752 ( .A(n21010), .B(n21053), .Z(n21055) );
  XNOR U20753 ( .A(n21064), .B(n21065), .Z(n21010) );
  AND U20754 ( .A(n336), .B(n21017), .Z(n21065) );
  XOR U20755 ( .A(n21064), .B(n21015), .Z(n21017) );
  XOR U20756 ( .A(n21066), .B(n21067), .Z(n21053) );
  AND U20757 ( .A(n21068), .B(n21069), .Z(n21067) );
  XNOR U20758 ( .A(n21066), .B(n21025), .Z(n21069) );
  XOR U20759 ( .A(n21070), .B(n21062), .Z(n21025) );
  XNOR U20760 ( .A(n21071), .B(n21057), .Z(n21062) );
  XOR U20761 ( .A(n21072), .B(n21073), .Z(n21057) );
  AND U20762 ( .A(n21074), .B(n21075), .Z(n21073) );
  XOR U20763 ( .A(n21076), .B(n21072), .Z(n21074) );
  XNOR U20764 ( .A(n21077), .B(n21078), .Z(n21071) );
  AND U20765 ( .A(n21079), .B(n21080), .Z(n21078) );
  XOR U20766 ( .A(n21077), .B(n21081), .Z(n21079) );
  XNOR U20767 ( .A(n21063), .B(n21060), .Z(n21070) );
  AND U20768 ( .A(n21082), .B(n21083), .Z(n21060) );
  XOR U20769 ( .A(n21084), .B(n21085), .Z(n21063) );
  AND U20770 ( .A(n21086), .B(n21087), .Z(n21085) );
  XOR U20771 ( .A(n21084), .B(n21088), .Z(n21086) );
  XNOR U20772 ( .A(n21022), .B(n21066), .Z(n21068) );
  XNOR U20773 ( .A(n21089), .B(n21090), .Z(n21022) );
  AND U20774 ( .A(n336), .B(n21028), .Z(n21090) );
  XOR U20775 ( .A(n21089), .B(n21026), .Z(n21028) );
  XOR U20776 ( .A(n21091), .B(n21092), .Z(n21066) );
  AND U20777 ( .A(n21093), .B(n21094), .Z(n21092) );
  XNOR U20778 ( .A(n21091), .B(n21082), .Z(n21094) );
  IV U20779 ( .A(n21036), .Z(n21082) );
  XNOR U20780 ( .A(n21095), .B(n21075), .Z(n21036) );
  XNOR U20781 ( .A(n21096), .B(n21081), .Z(n21075) );
  XOR U20782 ( .A(n21097), .B(n21098), .Z(n21081) );
  NOR U20783 ( .A(n21099), .B(n21100), .Z(n21098) );
  XNOR U20784 ( .A(n21097), .B(n21101), .Z(n21099) );
  XNOR U20785 ( .A(n21080), .B(n21072), .Z(n21096) );
  XOR U20786 ( .A(n21102), .B(n21103), .Z(n21072) );
  AND U20787 ( .A(n21104), .B(n21105), .Z(n21103) );
  XNOR U20788 ( .A(n21102), .B(n21106), .Z(n21104) );
  XNOR U20789 ( .A(n21107), .B(n21077), .Z(n21080) );
  XOR U20790 ( .A(n21108), .B(n21109), .Z(n21077) );
  AND U20791 ( .A(n21110), .B(n21111), .Z(n21109) );
  XOR U20792 ( .A(n21108), .B(n21112), .Z(n21110) );
  XNOR U20793 ( .A(n21113), .B(n21114), .Z(n21107) );
  NOR U20794 ( .A(n21115), .B(n21116), .Z(n21114) );
  XOR U20795 ( .A(n21113), .B(n21117), .Z(n21115) );
  XNOR U20796 ( .A(n21076), .B(n21083), .Z(n21095) );
  NOR U20797 ( .A(n21044), .B(n21118), .Z(n21083) );
  XOR U20798 ( .A(n21088), .B(n21087), .Z(n21076) );
  XNOR U20799 ( .A(n21119), .B(n21084), .Z(n21087) );
  XOR U20800 ( .A(n21120), .B(n21121), .Z(n21084) );
  AND U20801 ( .A(n21122), .B(n21123), .Z(n21121) );
  XOR U20802 ( .A(n21120), .B(n21124), .Z(n21122) );
  XNOR U20803 ( .A(n21125), .B(n21126), .Z(n21119) );
  NOR U20804 ( .A(n21127), .B(n21128), .Z(n21126) );
  XNOR U20805 ( .A(n21125), .B(n21129), .Z(n21127) );
  XOR U20806 ( .A(n21130), .B(n21131), .Z(n21088) );
  NOR U20807 ( .A(n21132), .B(n21133), .Z(n21131) );
  XNOR U20808 ( .A(n21130), .B(n21134), .Z(n21132) );
  XNOR U20809 ( .A(n21033), .B(n21091), .Z(n21093) );
  XNOR U20810 ( .A(n21135), .B(n21136), .Z(n21033) );
  AND U20811 ( .A(n336), .B(n21040), .Z(n21136) );
  XOR U20812 ( .A(n21135), .B(n21038), .Z(n21040) );
  AND U20813 ( .A(n21041), .B(n21044), .Z(n21091) );
  XOR U20814 ( .A(n21137), .B(n21118), .Z(n21044) );
  XNOR U20815 ( .A(p_input[2048]), .B(p_input[432]), .Z(n21118) );
  XOR U20816 ( .A(n21106), .B(n21105), .Z(n21137) );
  XNOR U20817 ( .A(n21138), .B(n21112), .Z(n21105) );
  XNOR U20818 ( .A(n21101), .B(n21100), .Z(n21112) );
  XOR U20819 ( .A(n21139), .B(n21097), .Z(n21100) );
  XNOR U20820 ( .A(n16904), .B(p_input[442]), .Z(n21097) );
  XNOR U20821 ( .A(p_input[2059]), .B(p_input[443]), .Z(n21139) );
  XOR U20822 ( .A(p_input[2060]), .B(p_input[444]), .Z(n21101) );
  XNOR U20823 ( .A(n21111), .B(n21102), .Z(n21138) );
  XNOR U20824 ( .A(n17068), .B(p_input[433]), .Z(n21102) );
  XOR U20825 ( .A(n21140), .B(n21117), .Z(n21111) );
  XNOR U20826 ( .A(p_input[2063]), .B(p_input[447]), .Z(n21117) );
  XOR U20827 ( .A(n21108), .B(n21116), .Z(n21140) );
  XOR U20828 ( .A(n21141), .B(n21113), .Z(n21116) );
  XOR U20829 ( .A(p_input[2061]), .B(p_input[445]), .Z(n21113) );
  XNOR U20830 ( .A(p_input[2062]), .B(p_input[446]), .Z(n21141) );
  XNOR U20831 ( .A(n16738), .B(p_input[441]), .Z(n21108) );
  XNOR U20832 ( .A(n21124), .B(n21123), .Z(n21106) );
  XNOR U20833 ( .A(n21142), .B(n21129), .Z(n21123) );
  XOR U20834 ( .A(p_input[2056]), .B(p_input[440]), .Z(n21129) );
  XOR U20835 ( .A(n21120), .B(n21128), .Z(n21142) );
  XOR U20836 ( .A(n21143), .B(n21125), .Z(n21128) );
  XOR U20837 ( .A(p_input[2054]), .B(p_input[438]), .Z(n21125) );
  XNOR U20838 ( .A(p_input[2055]), .B(p_input[439]), .Z(n21143) );
  XNOR U20839 ( .A(n16741), .B(p_input[434]), .Z(n21120) );
  XNOR U20840 ( .A(n21134), .B(n21133), .Z(n21124) );
  XOR U20841 ( .A(n21144), .B(n21130), .Z(n21133) );
  XOR U20842 ( .A(p_input[2051]), .B(p_input[435]), .Z(n21130) );
  XNOR U20843 ( .A(p_input[2052]), .B(p_input[436]), .Z(n21144) );
  XOR U20844 ( .A(p_input[2053]), .B(p_input[437]), .Z(n21134) );
  XNOR U20845 ( .A(n21145), .B(n21146), .Z(n21041) );
  AND U20846 ( .A(n336), .B(n21147), .Z(n21146) );
  XNOR U20847 ( .A(n21148), .B(n21149), .Z(n336) );
  AND U20848 ( .A(n21150), .B(n21151), .Z(n21149) );
  XOR U20849 ( .A(n21148), .B(n21051), .Z(n21151) );
  XNOR U20850 ( .A(n21148), .B(n21005), .Z(n21150) );
  XOR U20851 ( .A(n21152), .B(n21153), .Z(n21148) );
  AND U20852 ( .A(n21154), .B(n21155), .Z(n21153) );
  XOR U20853 ( .A(n21152), .B(n21015), .Z(n21154) );
  XOR U20854 ( .A(n21156), .B(n21157), .Z(n20994) );
  AND U20855 ( .A(n340), .B(n21147), .Z(n21157) );
  XNOR U20856 ( .A(n21145), .B(n21156), .Z(n21147) );
  XNOR U20857 ( .A(n21158), .B(n21159), .Z(n340) );
  AND U20858 ( .A(n21160), .B(n21161), .Z(n21159) );
  XNOR U20859 ( .A(n21162), .B(n21158), .Z(n21161) );
  IV U20860 ( .A(n21051), .Z(n21162) );
  XNOR U20861 ( .A(n21163), .B(n21164), .Z(n21051) );
  AND U20862 ( .A(n343), .B(n21165), .Z(n21164) );
  XNOR U20863 ( .A(n21163), .B(n21166), .Z(n21165) );
  XNOR U20864 ( .A(n21005), .B(n21158), .Z(n21160) );
  XOR U20865 ( .A(n21167), .B(n21168), .Z(n21005) );
  AND U20866 ( .A(n351), .B(n21169), .Z(n21168) );
  XOR U20867 ( .A(n21152), .B(n21170), .Z(n21158) );
  AND U20868 ( .A(n21171), .B(n21155), .Z(n21170) );
  XNOR U20869 ( .A(n21064), .B(n21152), .Z(n21155) );
  XNOR U20870 ( .A(n21172), .B(n21173), .Z(n21064) );
  AND U20871 ( .A(n343), .B(n21174), .Z(n21173) );
  XOR U20872 ( .A(n21175), .B(n21172), .Z(n21174) );
  XNOR U20873 ( .A(n21176), .B(n21152), .Z(n21171) );
  IV U20874 ( .A(n21015), .Z(n21176) );
  XOR U20875 ( .A(n21177), .B(n21178), .Z(n21015) );
  AND U20876 ( .A(n351), .B(n21179), .Z(n21178) );
  XOR U20877 ( .A(n21180), .B(n21181), .Z(n21152) );
  AND U20878 ( .A(n21182), .B(n21183), .Z(n21181) );
  XNOR U20879 ( .A(n21089), .B(n21180), .Z(n21183) );
  XNOR U20880 ( .A(n21184), .B(n21185), .Z(n21089) );
  AND U20881 ( .A(n343), .B(n21186), .Z(n21185) );
  XNOR U20882 ( .A(n21187), .B(n21184), .Z(n21186) );
  XOR U20883 ( .A(n21180), .B(n21026), .Z(n21182) );
  XOR U20884 ( .A(n21188), .B(n21189), .Z(n21026) );
  AND U20885 ( .A(n351), .B(n21190), .Z(n21189) );
  XOR U20886 ( .A(n21191), .B(n21192), .Z(n21180) );
  AND U20887 ( .A(n21193), .B(n21194), .Z(n21192) );
  XNOR U20888 ( .A(n21191), .B(n21135), .Z(n21194) );
  XNOR U20889 ( .A(n21195), .B(n21196), .Z(n21135) );
  AND U20890 ( .A(n343), .B(n21197), .Z(n21196) );
  XOR U20891 ( .A(n21198), .B(n21195), .Z(n21197) );
  XNOR U20892 ( .A(n21199), .B(n21191), .Z(n21193) );
  IV U20893 ( .A(n21038), .Z(n21199) );
  XOR U20894 ( .A(n21200), .B(n21201), .Z(n21038) );
  AND U20895 ( .A(n351), .B(n21202), .Z(n21201) );
  AND U20896 ( .A(n21156), .B(n21145), .Z(n21191) );
  XNOR U20897 ( .A(n21203), .B(n21204), .Z(n21145) );
  AND U20898 ( .A(n343), .B(n21205), .Z(n21204) );
  XNOR U20899 ( .A(n21206), .B(n21203), .Z(n21205) );
  XNOR U20900 ( .A(n21207), .B(n21208), .Z(n343) );
  AND U20901 ( .A(n21209), .B(n21210), .Z(n21208) );
  XOR U20902 ( .A(n21166), .B(n21207), .Z(n21210) );
  AND U20903 ( .A(n21211), .B(n21212), .Z(n21166) );
  XOR U20904 ( .A(n21207), .B(n21163), .Z(n21209) );
  XNOR U20905 ( .A(n21213), .B(n21214), .Z(n21163) );
  AND U20906 ( .A(n347), .B(n21169), .Z(n21214) );
  XOR U20907 ( .A(n21167), .B(n21213), .Z(n21169) );
  XOR U20908 ( .A(n21215), .B(n21216), .Z(n21207) );
  AND U20909 ( .A(n21217), .B(n21218), .Z(n21216) );
  XNOR U20910 ( .A(n21215), .B(n21211), .Z(n21218) );
  IV U20911 ( .A(n21175), .Z(n21211) );
  XOR U20912 ( .A(n21219), .B(n21220), .Z(n21175) );
  XOR U20913 ( .A(n21221), .B(n21212), .Z(n21220) );
  AND U20914 ( .A(n21187), .B(n21222), .Z(n21212) );
  AND U20915 ( .A(n21223), .B(n21224), .Z(n21221) );
  XOR U20916 ( .A(n21225), .B(n21219), .Z(n21223) );
  XNOR U20917 ( .A(n21172), .B(n21215), .Z(n21217) );
  XNOR U20918 ( .A(n21226), .B(n21227), .Z(n21172) );
  AND U20919 ( .A(n347), .B(n21179), .Z(n21227) );
  XOR U20920 ( .A(n21226), .B(n21177), .Z(n21179) );
  XOR U20921 ( .A(n21228), .B(n21229), .Z(n21215) );
  AND U20922 ( .A(n21230), .B(n21231), .Z(n21229) );
  XNOR U20923 ( .A(n21228), .B(n21187), .Z(n21231) );
  XOR U20924 ( .A(n21232), .B(n21224), .Z(n21187) );
  XNOR U20925 ( .A(n21233), .B(n21219), .Z(n21224) );
  XOR U20926 ( .A(n21234), .B(n21235), .Z(n21219) );
  AND U20927 ( .A(n21236), .B(n21237), .Z(n21235) );
  XOR U20928 ( .A(n21238), .B(n21234), .Z(n21236) );
  XNOR U20929 ( .A(n21239), .B(n21240), .Z(n21233) );
  AND U20930 ( .A(n21241), .B(n21242), .Z(n21240) );
  XOR U20931 ( .A(n21239), .B(n21243), .Z(n21241) );
  XNOR U20932 ( .A(n21225), .B(n21222), .Z(n21232) );
  AND U20933 ( .A(n21244), .B(n21245), .Z(n21222) );
  XOR U20934 ( .A(n21246), .B(n21247), .Z(n21225) );
  AND U20935 ( .A(n21248), .B(n21249), .Z(n21247) );
  XOR U20936 ( .A(n21246), .B(n21250), .Z(n21248) );
  XNOR U20937 ( .A(n21184), .B(n21228), .Z(n21230) );
  XNOR U20938 ( .A(n21251), .B(n21252), .Z(n21184) );
  AND U20939 ( .A(n347), .B(n21190), .Z(n21252) );
  XOR U20940 ( .A(n21251), .B(n21188), .Z(n21190) );
  XOR U20941 ( .A(n21253), .B(n21254), .Z(n21228) );
  AND U20942 ( .A(n21255), .B(n21256), .Z(n21254) );
  XNOR U20943 ( .A(n21253), .B(n21244), .Z(n21256) );
  IV U20944 ( .A(n21198), .Z(n21244) );
  XNOR U20945 ( .A(n21257), .B(n21237), .Z(n21198) );
  XNOR U20946 ( .A(n21258), .B(n21243), .Z(n21237) );
  XOR U20947 ( .A(n21259), .B(n21260), .Z(n21243) );
  NOR U20948 ( .A(n21261), .B(n21262), .Z(n21260) );
  XNOR U20949 ( .A(n21259), .B(n21263), .Z(n21261) );
  XNOR U20950 ( .A(n21242), .B(n21234), .Z(n21258) );
  XOR U20951 ( .A(n21264), .B(n21265), .Z(n21234) );
  AND U20952 ( .A(n21266), .B(n21267), .Z(n21265) );
  XNOR U20953 ( .A(n21264), .B(n21268), .Z(n21266) );
  XNOR U20954 ( .A(n21269), .B(n21239), .Z(n21242) );
  XOR U20955 ( .A(n21270), .B(n21271), .Z(n21239) );
  AND U20956 ( .A(n21272), .B(n21273), .Z(n21271) );
  XOR U20957 ( .A(n21270), .B(n21274), .Z(n21272) );
  XNOR U20958 ( .A(n21275), .B(n21276), .Z(n21269) );
  NOR U20959 ( .A(n21277), .B(n21278), .Z(n21276) );
  XOR U20960 ( .A(n21275), .B(n21279), .Z(n21277) );
  XNOR U20961 ( .A(n21238), .B(n21245), .Z(n21257) );
  NOR U20962 ( .A(n21206), .B(n21280), .Z(n21245) );
  XOR U20963 ( .A(n21250), .B(n21249), .Z(n21238) );
  XNOR U20964 ( .A(n21281), .B(n21246), .Z(n21249) );
  XOR U20965 ( .A(n21282), .B(n21283), .Z(n21246) );
  AND U20966 ( .A(n21284), .B(n21285), .Z(n21283) );
  XOR U20967 ( .A(n21282), .B(n21286), .Z(n21284) );
  XNOR U20968 ( .A(n21287), .B(n21288), .Z(n21281) );
  NOR U20969 ( .A(n21289), .B(n21290), .Z(n21288) );
  XNOR U20970 ( .A(n21287), .B(n21291), .Z(n21289) );
  XOR U20971 ( .A(n21292), .B(n21293), .Z(n21250) );
  NOR U20972 ( .A(n21294), .B(n21295), .Z(n21293) );
  XNOR U20973 ( .A(n21292), .B(n21296), .Z(n21294) );
  XNOR U20974 ( .A(n21195), .B(n21253), .Z(n21255) );
  XNOR U20975 ( .A(n21297), .B(n21298), .Z(n21195) );
  AND U20976 ( .A(n347), .B(n21202), .Z(n21298) );
  XOR U20977 ( .A(n21297), .B(n21200), .Z(n21202) );
  AND U20978 ( .A(n21203), .B(n21206), .Z(n21253) );
  XOR U20979 ( .A(n21299), .B(n21280), .Z(n21206) );
  XNOR U20980 ( .A(p_input[2048]), .B(p_input[448]), .Z(n21280) );
  XOR U20981 ( .A(n21268), .B(n21267), .Z(n21299) );
  XNOR U20982 ( .A(n21300), .B(n21274), .Z(n21267) );
  XNOR U20983 ( .A(n21263), .B(n21262), .Z(n21274) );
  XOR U20984 ( .A(n21301), .B(n21259), .Z(n21262) );
  XNOR U20985 ( .A(n16904), .B(p_input[458]), .Z(n21259) );
  XNOR U20986 ( .A(p_input[2059]), .B(p_input[459]), .Z(n21301) );
  XOR U20987 ( .A(p_input[2060]), .B(p_input[460]), .Z(n21263) );
  XNOR U20988 ( .A(n21273), .B(n21264), .Z(n21300) );
  XNOR U20989 ( .A(n17068), .B(p_input[449]), .Z(n21264) );
  XOR U20990 ( .A(n21302), .B(n21279), .Z(n21273) );
  XNOR U20991 ( .A(p_input[2063]), .B(p_input[463]), .Z(n21279) );
  XOR U20992 ( .A(n21270), .B(n21278), .Z(n21302) );
  XOR U20993 ( .A(n21303), .B(n21275), .Z(n21278) );
  XOR U20994 ( .A(p_input[2061]), .B(p_input[461]), .Z(n21275) );
  XNOR U20995 ( .A(p_input[2062]), .B(p_input[462]), .Z(n21303) );
  XNOR U20996 ( .A(n16738), .B(p_input[457]), .Z(n21270) );
  XNOR U20997 ( .A(n21286), .B(n21285), .Z(n21268) );
  XNOR U20998 ( .A(n21304), .B(n21291), .Z(n21285) );
  XOR U20999 ( .A(p_input[2056]), .B(p_input[456]), .Z(n21291) );
  XOR U21000 ( .A(n21282), .B(n21290), .Z(n21304) );
  XOR U21001 ( .A(n21305), .B(n21287), .Z(n21290) );
  XOR U21002 ( .A(p_input[2054]), .B(p_input[454]), .Z(n21287) );
  XNOR U21003 ( .A(p_input[2055]), .B(p_input[455]), .Z(n21305) );
  XNOR U21004 ( .A(n16741), .B(p_input[450]), .Z(n21282) );
  XNOR U21005 ( .A(n21296), .B(n21295), .Z(n21286) );
  XOR U21006 ( .A(n21306), .B(n21292), .Z(n21295) );
  XOR U21007 ( .A(p_input[2051]), .B(p_input[451]), .Z(n21292) );
  XNOR U21008 ( .A(p_input[2052]), .B(p_input[452]), .Z(n21306) );
  XOR U21009 ( .A(p_input[2053]), .B(p_input[453]), .Z(n21296) );
  XNOR U21010 ( .A(n21307), .B(n21308), .Z(n21203) );
  AND U21011 ( .A(n347), .B(n21309), .Z(n21308) );
  XNOR U21012 ( .A(n21310), .B(n21311), .Z(n347) );
  AND U21013 ( .A(n21312), .B(n21313), .Z(n21311) );
  XOR U21014 ( .A(n21310), .B(n21213), .Z(n21313) );
  XNOR U21015 ( .A(n21310), .B(n21167), .Z(n21312) );
  XOR U21016 ( .A(n21314), .B(n21315), .Z(n21310) );
  AND U21017 ( .A(n21316), .B(n21317), .Z(n21315) );
  XOR U21018 ( .A(n21314), .B(n21177), .Z(n21316) );
  XOR U21019 ( .A(n21318), .B(n21319), .Z(n21156) );
  AND U21020 ( .A(n351), .B(n21309), .Z(n21319) );
  XNOR U21021 ( .A(n21307), .B(n21318), .Z(n21309) );
  XNOR U21022 ( .A(n21320), .B(n21321), .Z(n351) );
  AND U21023 ( .A(n21322), .B(n21323), .Z(n21321) );
  XNOR U21024 ( .A(n21324), .B(n21320), .Z(n21323) );
  IV U21025 ( .A(n21213), .Z(n21324) );
  XNOR U21026 ( .A(n21325), .B(n21326), .Z(n21213) );
  AND U21027 ( .A(n354), .B(n21327), .Z(n21326) );
  XNOR U21028 ( .A(n21325), .B(n21328), .Z(n21327) );
  XNOR U21029 ( .A(n21167), .B(n21320), .Z(n21322) );
  XOR U21030 ( .A(n21329), .B(n21330), .Z(n21167) );
  AND U21031 ( .A(n362), .B(n21331), .Z(n21330) );
  XOR U21032 ( .A(n21314), .B(n21332), .Z(n21320) );
  AND U21033 ( .A(n21333), .B(n21317), .Z(n21332) );
  XNOR U21034 ( .A(n21226), .B(n21314), .Z(n21317) );
  XNOR U21035 ( .A(n21334), .B(n21335), .Z(n21226) );
  AND U21036 ( .A(n354), .B(n21336), .Z(n21335) );
  XOR U21037 ( .A(n21337), .B(n21334), .Z(n21336) );
  XNOR U21038 ( .A(n21338), .B(n21314), .Z(n21333) );
  IV U21039 ( .A(n21177), .Z(n21338) );
  XOR U21040 ( .A(n21339), .B(n21340), .Z(n21177) );
  AND U21041 ( .A(n362), .B(n21341), .Z(n21340) );
  XOR U21042 ( .A(n21342), .B(n21343), .Z(n21314) );
  AND U21043 ( .A(n21344), .B(n21345), .Z(n21343) );
  XNOR U21044 ( .A(n21251), .B(n21342), .Z(n21345) );
  XNOR U21045 ( .A(n21346), .B(n21347), .Z(n21251) );
  AND U21046 ( .A(n354), .B(n21348), .Z(n21347) );
  XNOR U21047 ( .A(n21349), .B(n21346), .Z(n21348) );
  XOR U21048 ( .A(n21342), .B(n21188), .Z(n21344) );
  XOR U21049 ( .A(n21350), .B(n21351), .Z(n21188) );
  AND U21050 ( .A(n362), .B(n21352), .Z(n21351) );
  XOR U21051 ( .A(n21353), .B(n21354), .Z(n21342) );
  AND U21052 ( .A(n21355), .B(n21356), .Z(n21354) );
  XNOR U21053 ( .A(n21353), .B(n21297), .Z(n21356) );
  XNOR U21054 ( .A(n21357), .B(n21358), .Z(n21297) );
  AND U21055 ( .A(n354), .B(n21359), .Z(n21358) );
  XOR U21056 ( .A(n21360), .B(n21357), .Z(n21359) );
  XNOR U21057 ( .A(n21361), .B(n21353), .Z(n21355) );
  IV U21058 ( .A(n21200), .Z(n21361) );
  XOR U21059 ( .A(n21362), .B(n21363), .Z(n21200) );
  AND U21060 ( .A(n362), .B(n21364), .Z(n21363) );
  AND U21061 ( .A(n21318), .B(n21307), .Z(n21353) );
  XNOR U21062 ( .A(n21365), .B(n21366), .Z(n21307) );
  AND U21063 ( .A(n354), .B(n21367), .Z(n21366) );
  XNOR U21064 ( .A(n21368), .B(n21365), .Z(n21367) );
  XNOR U21065 ( .A(n21369), .B(n21370), .Z(n354) );
  AND U21066 ( .A(n21371), .B(n21372), .Z(n21370) );
  XOR U21067 ( .A(n21328), .B(n21369), .Z(n21372) );
  AND U21068 ( .A(n21373), .B(n21374), .Z(n21328) );
  XOR U21069 ( .A(n21369), .B(n21325), .Z(n21371) );
  XNOR U21070 ( .A(n21375), .B(n21376), .Z(n21325) );
  AND U21071 ( .A(n358), .B(n21331), .Z(n21376) );
  XOR U21072 ( .A(n21329), .B(n21375), .Z(n21331) );
  XOR U21073 ( .A(n21377), .B(n21378), .Z(n21369) );
  AND U21074 ( .A(n21379), .B(n21380), .Z(n21378) );
  XNOR U21075 ( .A(n21377), .B(n21373), .Z(n21380) );
  IV U21076 ( .A(n21337), .Z(n21373) );
  XOR U21077 ( .A(n21381), .B(n21382), .Z(n21337) );
  XOR U21078 ( .A(n21383), .B(n21374), .Z(n21382) );
  AND U21079 ( .A(n21349), .B(n21384), .Z(n21374) );
  AND U21080 ( .A(n21385), .B(n21386), .Z(n21383) );
  XOR U21081 ( .A(n21387), .B(n21381), .Z(n21385) );
  XNOR U21082 ( .A(n21334), .B(n21377), .Z(n21379) );
  XNOR U21083 ( .A(n21388), .B(n21389), .Z(n21334) );
  AND U21084 ( .A(n358), .B(n21341), .Z(n21389) );
  XOR U21085 ( .A(n21388), .B(n21339), .Z(n21341) );
  XOR U21086 ( .A(n21390), .B(n21391), .Z(n21377) );
  AND U21087 ( .A(n21392), .B(n21393), .Z(n21391) );
  XNOR U21088 ( .A(n21390), .B(n21349), .Z(n21393) );
  XOR U21089 ( .A(n21394), .B(n21386), .Z(n21349) );
  XNOR U21090 ( .A(n21395), .B(n21381), .Z(n21386) );
  XOR U21091 ( .A(n21396), .B(n21397), .Z(n21381) );
  AND U21092 ( .A(n21398), .B(n21399), .Z(n21397) );
  XOR U21093 ( .A(n21400), .B(n21396), .Z(n21398) );
  XNOR U21094 ( .A(n21401), .B(n21402), .Z(n21395) );
  AND U21095 ( .A(n21403), .B(n21404), .Z(n21402) );
  XOR U21096 ( .A(n21401), .B(n21405), .Z(n21403) );
  XNOR U21097 ( .A(n21387), .B(n21384), .Z(n21394) );
  AND U21098 ( .A(n21406), .B(n21407), .Z(n21384) );
  XOR U21099 ( .A(n21408), .B(n21409), .Z(n21387) );
  AND U21100 ( .A(n21410), .B(n21411), .Z(n21409) );
  XOR U21101 ( .A(n21408), .B(n21412), .Z(n21410) );
  XNOR U21102 ( .A(n21346), .B(n21390), .Z(n21392) );
  XNOR U21103 ( .A(n21413), .B(n21414), .Z(n21346) );
  AND U21104 ( .A(n358), .B(n21352), .Z(n21414) );
  XOR U21105 ( .A(n21413), .B(n21350), .Z(n21352) );
  XOR U21106 ( .A(n21415), .B(n21416), .Z(n21390) );
  AND U21107 ( .A(n21417), .B(n21418), .Z(n21416) );
  XNOR U21108 ( .A(n21415), .B(n21406), .Z(n21418) );
  IV U21109 ( .A(n21360), .Z(n21406) );
  XNOR U21110 ( .A(n21419), .B(n21399), .Z(n21360) );
  XNOR U21111 ( .A(n21420), .B(n21405), .Z(n21399) );
  XOR U21112 ( .A(n21421), .B(n21422), .Z(n21405) );
  NOR U21113 ( .A(n21423), .B(n21424), .Z(n21422) );
  XNOR U21114 ( .A(n21421), .B(n21425), .Z(n21423) );
  XNOR U21115 ( .A(n21404), .B(n21396), .Z(n21420) );
  XOR U21116 ( .A(n21426), .B(n21427), .Z(n21396) );
  AND U21117 ( .A(n21428), .B(n21429), .Z(n21427) );
  XNOR U21118 ( .A(n21426), .B(n21430), .Z(n21428) );
  XNOR U21119 ( .A(n21431), .B(n21401), .Z(n21404) );
  XOR U21120 ( .A(n21432), .B(n21433), .Z(n21401) );
  AND U21121 ( .A(n21434), .B(n21435), .Z(n21433) );
  XOR U21122 ( .A(n21432), .B(n21436), .Z(n21434) );
  XNOR U21123 ( .A(n21437), .B(n21438), .Z(n21431) );
  NOR U21124 ( .A(n21439), .B(n21440), .Z(n21438) );
  XOR U21125 ( .A(n21437), .B(n21441), .Z(n21439) );
  XNOR U21126 ( .A(n21400), .B(n21407), .Z(n21419) );
  NOR U21127 ( .A(n21368), .B(n21442), .Z(n21407) );
  XOR U21128 ( .A(n21412), .B(n21411), .Z(n21400) );
  XNOR U21129 ( .A(n21443), .B(n21408), .Z(n21411) );
  XOR U21130 ( .A(n21444), .B(n21445), .Z(n21408) );
  AND U21131 ( .A(n21446), .B(n21447), .Z(n21445) );
  XOR U21132 ( .A(n21444), .B(n21448), .Z(n21446) );
  XNOR U21133 ( .A(n21449), .B(n21450), .Z(n21443) );
  NOR U21134 ( .A(n21451), .B(n21452), .Z(n21450) );
  XNOR U21135 ( .A(n21449), .B(n21453), .Z(n21451) );
  XOR U21136 ( .A(n21454), .B(n21455), .Z(n21412) );
  NOR U21137 ( .A(n21456), .B(n21457), .Z(n21455) );
  XNOR U21138 ( .A(n21454), .B(n21458), .Z(n21456) );
  XNOR U21139 ( .A(n21357), .B(n21415), .Z(n21417) );
  XNOR U21140 ( .A(n21459), .B(n21460), .Z(n21357) );
  AND U21141 ( .A(n358), .B(n21364), .Z(n21460) );
  XOR U21142 ( .A(n21459), .B(n21362), .Z(n21364) );
  AND U21143 ( .A(n21365), .B(n21368), .Z(n21415) );
  XOR U21144 ( .A(n21461), .B(n21442), .Z(n21368) );
  XNOR U21145 ( .A(p_input[2048]), .B(p_input[464]), .Z(n21442) );
  XOR U21146 ( .A(n21430), .B(n21429), .Z(n21461) );
  XNOR U21147 ( .A(n21462), .B(n21436), .Z(n21429) );
  XNOR U21148 ( .A(n21425), .B(n21424), .Z(n21436) );
  XOR U21149 ( .A(n21463), .B(n21421), .Z(n21424) );
  XNOR U21150 ( .A(n16904), .B(p_input[474]), .Z(n21421) );
  XNOR U21151 ( .A(p_input[2059]), .B(p_input[475]), .Z(n21463) );
  XOR U21152 ( .A(p_input[2060]), .B(p_input[476]), .Z(n21425) );
  XNOR U21153 ( .A(n21435), .B(n21426), .Z(n21462) );
  XNOR U21154 ( .A(n17068), .B(p_input[465]), .Z(n21426) );
  XOR U21155 ( .A(n21464), .B(n21441), .Z(n21435) );
  XNOR U21156 ( .A(p_input[2063]), .B(p_input[479]), .Z(n21441) );
  XOR U21157 ( .A(n21432), .B(n21440), .Z(n21464) );
  XOR U21158 ( .A(n21465), .B(n21437), .Z(n21440) );
  XOR U21159 ( .A(p_input[2061]), .B(p_input[477]), .Z(n21437) );
  XNOR U21160 ( .A(p_input[2062]), .B(p_input[478]), .Z(n21465) );
  XNOR U21161 ( .A(n16738), .B(p_input[473]), .Z(n21432) );
  XNOR U21162 ( .A(n21448), .B(n21447), .Z(n21430) );
  XNOR U21163 ( .A(n21466), .B(n21453), .Z(n21447) );
  XOR U21164 ( .A(p_input[2056]), .B(p_input[472]), .Z(n21453) );
  XOR U21165 ( .A(n21444), .B(n21452), .Z(n21466) );
  XOR U21166 ( .A(n21467), .B(n21449), .Z(n21452) );
  XOR U21167 ( .A(p_input[2054]), .B(p_input[470]), .Z(n21449) );
  XNOR U21168 ( .A(p_input[2055]), .B(p_input[471]), .Z(n21467) );
  XNOR U21169 ( .A(n16741), .B(p_input[466]), .Z(n21444) );
  XNOR U21170 ( .A(n21458), .B(n21457), .Z(n21448) );
  XOR U21171 ( .A(n21468), .B(n21454), .Z(n21457) );
  XOR U21172 ( .A(p_input[2051]), .B(p_input[467]), .Z(n21454) );
  XNOR U21173 ( .A(p_input[2052]), .B(p_input[468]), .Z(n21468) );
  XOR U21174 ( .A(p_input[2053]), .B(p_input[469]), .Z(n21458) );
  XNOR U21175 ( .A(n21469), .B(n21470), .Z(n21365) );
  AND U21176 ( .A(n358), .B(n21471), .Z(n21470) );
  XNOR U21177 ( .A(n21472), .B(n21473), .Z(n358) );
  AND U21178 ( .A(n21474), .B(n21475), .Z(n21473) );
  XOR U21179 ( .A(n21472), .B(n21375), .Z(n21475) );
  XNOR U21180 ( .A(n21472), .B(n21329), .Z(n21474) );
  XOR U21181 ( .A(n21476), .B(n21477), .Z(n21472) );
  AND U21182 ( .A(n21478), .B(n21479), .Z(n21477) );
  XOR U21183 ( .A(n21476), .B(n21339), .Z(n21478) );
  XOR U21184 ( .A(n21480), .B(n21481), .Z(n21318) );
  AND U21185 ( .A(n362), .B(n21471), .Z(n21481) );
  XNOR U21186 ( .A(n21469), .B(n21480), .Z(n21471) );
  XNOR U21187 ( .A(n21482), .B(n21483), .Z(n362) );
  AND U21188 ( .A(n21484), .B(n21485), .Z(n21483) );
  XNOR U21189 ( .A(n21486), .B(n21482), .Z(n21485) );
  IV U21190 ( .A(n21375), .Z(n21486) );
  XNOR U21191 ( .A(n21487), .B(n21488), .Z(n21375) );
  AND U21192 ( .A(n365), .B(n21489), .Z(n21488) );
  XNOR U21193 ( .A(n21487), .B(n21490), .Z(n21489) );
  XNOR U21194 ( .A(n21329), .B(n21482), .Z(n21484) );
  XOR U21195 ( .A(n21491), .B(n21492), .Z(n21329) );
  AND U21196 ( .A(n373), .B(n21493), .Z(n21492) );
  XOR U21197 ( .A(n21476), .B(n21494), .Z(n21482) );
  AND U21198 ( .A(n21495), .B(n21479), .Z(n21494) );
  XNOR U21199 ( .A(n21388), .B(n21476), .Z(n21479) );
  XNOR U21200 ( .A(n21496), .B(n21497), .Z(n21388) );
  AND U21201 ( .A(n365), .B(n21498), .Z(n21497) );
  XOR U21202 ( .A(n21499), .B(n21496), .Z(n21498) );
  XNOR U21203 ( .A(n21500), .B(n21476), .Z(n21495) );
  IV U21204 ( .A(n21339), .Z(n21500) );
  XOR U21205 ( .A(n21501), .B(n21502), .Z(n21339) );
  AND U21206 ( .A(n373), .B(n21503), .Z(n21502) );
  XOR U21207 ( .A(n21504), .B(n21505), .Z(n21476) );
  AND U21208 ( .A(n21506), .B(n21507), .Z(n21505) );
  XNOR U21209 ( .A(n21413), .B(n21504), .Z(n21507) );
  XNOR U21210 ( .A(n21508), .B(n21509), .Z(n21413) );
  AND U21211 ( .A(n365), .B(n21510), .Z(n21509) );
  XNOR U21212 ( .A(n21511), .B(n21508), .Z(n21510) );
  XOR U21213 ( .A(n21504), .B(n21350), .Z(n21506) );
  XOR U21214 ( .A(n21512), .B(n21513), .Z(n21350) );
  AND U21215 ( .A(n373), .B(n21514), .Z(n21513) );
  XOR U21216 ( .A(n21515), .B(n21516), .Z(n21504) );
  AND U21217 ( .A(n21517), .B(n21518), .Z(n21516) );
  XNOR U21218 ( .A(n21515), .B(n21459), .Z(n21518) );
  XNOR U21219 ( .A(n21519), .B(n21520), .Z(n21459) );
  AND U21220 ( .A(n365), .B(n21521), .Z(n21520) );
  XOR U21221 ( .A(n21522), .B(n21519), .Z(n21521) );
  XNOR U21222 ( .A(n21523), .B(n21515), .Z(n21517) );
  IV U21223 ( .A(n21362), .Z(n21523) );
  XOR U21224 ( .A(n21524), .B(n21525), .Z(n21362) );
  AND U21225 ( .A(n373), .B(n21526), .Z(n21525) );
  AND U21226 ( .A(n21480), .B(n21469), .Z(n21515) );
  XNOR U21227 ( .A(n21527), .B(n21528), .Z(n21469) );
  AND U21228 ( .A(n365), .B(n21529), .Z(n21528) );
  XNOR U21229 ( .A(n21530), .B(n21527), .Z(n21529) );
  XNOR U21230 ( .A(n21531), .B(n21532), .Z(n365) );
  AND U21231 ( .A(n21533), .B(n21534), .Z(n21532) );
  XOR U21232 ( .A(n21490), .B(n21531), .Z(n21534) );
  AND U21233 ( .A(n21535), .B(n21536), .Z(n21490) );
  XOR U21234 ( .A(n21531), .B(n21487), .Z(n21533) );
  XNOR U21235 ( .A(n21537), .B(n21538), .Z(n21487) );
  AND U21236 ( .A(n369), .B(n21493), .Z(n21538) );
  XOR U21237 ( .A(n21491), .B(n21537), .Z(n21493) );
  XOR U21238 ( .A(n21539), .B(n21540), .Z(n21531) );
  AND U21239 ( .A(n21541), .B(n21542), .Z(n21540) );
  XNOR U21240 ( .A(n21539), .B(n21535), .Z(n21542) );
  IV U21241 ( .A(n21499), .Z(n21535) );
  XOR U21242 ( .A(n21543), .B(n21544), .Z(n21499) );
  XOR U21243 ( .A(n21545), .B(n21536), .Z(n21544) );
  AND U21244 ( .A(n21511), .B(n21546), .Z(n21536) );
  AND U21245 ( .A(n21547), .B(n21548), .Z(n21545) );
  XOR U21246 ( .A(n21549), .B(n21543), .Z(n21547) );
  XNOR U21247 ( .A(n21496), .B(n21539), .Z(n21541) );
  XNOR U21248 ( .A(n21550), .B(n21551), .Z(n21496) );
  AND U21249 ( .A(n369), .B(n21503), .Z(n21551) );
  XOR U21250 ( .A(n21550), .B(n21501), .Z(n21503) );
  XOR U21251 ( .A(n21552), .B(n21553), .Z(n21539) );
  AND U21252 ( .A(n21554), .B(n21555), .Z(n21553) );
  XNOR U21253 ( .A(n21552), .B(n21511), .Z(n21555) );
  XOR U21254 ( .A(n21556), .B(n21548), .Z(n21511) );
  XNOR U21255 ( .A(n21557), .B(n21543), .Z(n21548) );
  XOR U21256 ( .A(n21558), .B(n21559), .Z(n21543) );
  AND U21257 ( .A(n21560), .B(n21561), .Z(n21559) );
  XOR U21258 ( .A(n21562), .B(n21558), .Z(n21560) );
  XNOR U21259 ( .A(n21563), .B(n21564), .Z(n21557) );
  AND U21260 ( .A(n21565), .B(n21566), .Z(n21564) );
  XOR U21261 ( .A(n21563), .B(n21567), .Z(n21565) );
  XNOR U21262 ( .A(n21549), .B(n21546), .Z(n21556) );
  AND U21263 ( .A(n21568), .B(n21569), .Z(n21546) );
  XOR U21264 ( .A(n21570), .B(n21571), .Z(n21549) );
  AND U21265 ( .A(n21572), .B(n21573), .Z(n21571) );
  XOR U21266 ( .A(n21570), .B(n21574), .Z(n21572) );
  XNOR U21267 ( .A(n21508), .B(n21552), .Z(n21554) );
  XNOR U21268 ( .A(n21575), .B(n21576), .Z(n21508) );
  AND U21269 ( .A(n369), .B(n21514), .Z(n21576) );
  XOR U21270 ( .A(n21575), .B(n21512), .Z(n21514) );
  XOR U21271 ( .A(n21577), .B(n21578), .Z(n21552) );
  AND U21272 ( .A(n21579), .B(n21580), .Z(n21578) );
  XNOR U21273 ( .A(n21577), .B(n21568), .Z(n21580) );
  IV U21274 ( .A(n21522), .Z(n21568) );
  XNOR U21275 ( .A(n21581), .B(n21561), .Z(n21522) );
  XNOR U21276 ( .A(n21582), .B(n21567), .Z(n21561) );
  XOR U21277 ( .A(n21583), .B(n21584), .Z(n21567) );
  NOR U21278 ( .A(n21585), .B(n21586), .Z(n21584) );
  XNOR U21279 ( .A(n21583), .B(n21587), .Z(n21585) );
  XNOR U21280 ( .A(n21566), .B(n21558), .Z(n21582) );
  XOR U21281 ( .A(n21588), .B(n21589), .Z(n21558) );
  AND U21282 ( .A(n21590), .B(n21591), .Z(n21589) );
  XNOR U21283 ( .A(n21588), .B(n21592), .Z(n21590) );
  XNOR U21284 ( .A(n21593), .B(n21563), .Z(n21566) );
  XOR U21285 ( .A(n21594), .B(n21595), .Z(n21563) );
  AND U21286 ( .A(n21596), .B(n21597), .Z(n21595) );
  XOR U21287 ( .A(n21594), .B(n21598), .Z(n21596) );
  XNOR U21288 ( .A(n21599), .B(n21600), .Z(n21593) );
  NOR U21289 ( .A(n21601), .B(n21602), .Z(n21600) );
  XOR U21290 ( .A(n21599), .B(n21603), .Z(n21601) );
  XNOR U21291 ( .A(n21562), .B(n21569), .Z(n21581) );
  NOR U21292 ( .A(n21530), .B(n21604), .Z(n21569) );
  XOR U21293 ( .A(n21574), .B(n21573), .Z(n21562) );
  XNOR U21294 ( .A(n21605), .B(n21570), .Z(n21573) );
  XOR U21295 ( .A(n21606), .B(n21607), .Z(n21570) );
  AND U21296 ( .A(n21608), .B(n21609), .Z(n21607) );
  XOR U21297 ( .A(n21606), .B(n21610), .Z(n21608) );
  XNOR U21298 ( .A(n21611), .B(n21612), .Z(n21605) );
  NOR U21299 ( .A(n21613), .B(n21614), .Z(n21612) );
  XNOR U21300 ( .A(n21611), .B(n21615), .Z(n21613) );
  XOR U21301 ( .A(n21616), .B(n21617), .Z(n21574) );
  NOR U21302 ( .A(n21618), .B(n21619), .Z(n21617) );
  XNOR U21303 ( .A(n21616), .B(n21620), .Z(n21618) );
  XNOR U21304 ( .A(n21519), .B(n21577), .Z(n21579) );
  XNOR U21305 ( .A(n21621), .B(n21622), .Z(n21519) );
  AND U21306 ( .A(n369), .B(n21526), .Z(n21622) );
  XOR U21307 ( .A(n21621), .B(n21524), .Z(n21526) );
  AND U21308 ( .A(n21527), .B(n21530), .Z(n21577) );
  XOR U21309 ( .A(n21623), .B(n21604), .Z(n21530) );
  XNOR U21310 ( .A(p_input[2048]), .B(p_input[480]), .Z(n21604) );
  XOR U21311 ( .A(n21592), .B(n21591), .Z(n21623) );
  XNOR U21312 ( .A(n21624), .B(n21598), .Z(n21591) );
  XNOR U21313 ( .A(n21587), .B(n21586), .Z(n21598) );
  XOR U21314 ( .A(n21625), .B(n21583), .Z(n21586) );
  XNOR U21315 ( .A(n16904), .B(p_input[490]), .Z(n21583) );
  XNOR U21316 ( .A(p_input[2059]), .B(p_input[491]), .Z(n21625) );
  XOR U21317 ( .A(p_input[2060]), .B(p_input[492]), .Z(n21587) );
  XNOR U21318 ( .A(n21597), .B(n21588), .Z(n21624) );
  XNOR U21319 ( .A(n17068), .B(p_input[481]), .Z(n21588) );
  XOR U21320 ( .A(n21626), .B(n21603), .Z(n21597) );
  XNOR U21321 ( .A(p_input[2063]), .B(p_input[495]), .Z(n21603) );
  XOR U21322 ( .A(n21594), .B(n21602), .Z(n21626) );
  XOR U21323 ( .A(n21627), .B(n21599), .Z(n21602) );
  XOR U21324 ( .A(p_input[2061]), .B(p_input[493]), .Z(n21599) );
  XNOR U21325 ( .A(p_input[2062]), .B(p_input[494]), .Z(n21627) );
  XNOR U21326 ( .A(n16738), .B(p_input[489]), .Z(n21594) );
  XNOR U21327 ( .A(n21610), .B(n21609), .Z(n21592) );
  XNOR U21328 ( .A(n21628), .B(n21615), .Z(n21609) );
  XOR U21329 ( .A(p_input[2056]), .B(p_input[488]), .Z(n21615) );
  XOR U21330 ( .A(n21606), .B(n21614), .Z(n21628) );
  XOR U21331 ( .A(n21629), .B(n21611), .Z(n21614) );
  XOR U21332 ( .A(p_input[2054]), .B(p_input[486]), .Z(n21611) );
  XNOR U21333 ( .A(p_input[2055]), .B(p_input[487]), .Z(n21629) );
  XNOR U21334 ( .A(n16741), .B(p_input[482]), .Z(n21606) );
  XNOR U21335 ( .A(n21620), .B(n21619), .Z(n21610) );
  XOR U21336 ( .A(n21630), .B(n21616), .Z(n21619) );
  XOR U21337 ( .A(p_input[2051]), .B(p_input[483]), .Z(n21616) );
  XNOR U21338 ( .A(p_input[2052]), .B(p_input[484]), .Z(n21630) );
  XOR U21339 ( .A(p_input[2053]), .B(p_input[485]), .Z(n21620) );
  XNOR U21340 ( .A(n21631), .B(n21632), .Z(n21527) );
  AND U21341 ( .A(n369), .B(n21633), .Z(n21632) );
  XNOR U21342 ( .A(n21634), .B(n21635), .Z(n369) );
  AND U21343 ( .A(n21636), .B(n21637), .Z(n21635) );
  XOR U21344 ( .A(n21634), .B(n21537), .Z(n21637) );
  XNOR U21345 ( .A(n21634), .B(n21491), .Z(n21636) );
  XOR U21346 ( .A(n21638), .B(n21639), .Z(n21634) );
  AND U21347 ( .A(n21640), .B(n21641), .Z(n21639) );
  XOR U21348 ( .A(n21638), .B(n21501), .Z(n21640) );
  XOR U21349 ( .A(n21642), .B(n21643), .Z(n21480) );
  AND U21350 ( .A(n373), .B(n21633), .Z(n21643) );
  XNOR U21351 ( .A(n21631), .B(n21642), .Z(n21633) );
  XNOR U21352 ( .A(n21644), .B(n21645), .Z(n373) );
  AND U21353 ( .A(n21646), .B(n21647), .Z(n21645) );
  XNOR U21354 ( .A(n21648), .B(n21644), .Z(n21647) );
  IV U21355 ( .A(n21537), .Z(n21648) );
  XNOR U21356 ( .A(n21649), .B(n21650), .Z(n21537) );
  AND U21357 ( .A(n376), .B(n21651), .Z(n21650) );
  XNOR U21358 ( .A(n21649), .B(n21652), .Z(n21651) );
  XNOR U21359 ( .A(n21491), .B(n21644), .Z(n21646) );
  XOR U21360 ( .A(n21653), .B(n21654), .Z(n21491) );
  AND U21361 ( .A(n384), .B(n21655), .Z(n21654) );
  XOR U21362 ( .A(n21638), .B(n21656), .Z(n21644) );
  AND U21363 ( .A(n21657), .B(n21641), .Z(n21656) );
  XNOR U21364 ( .A(n21550), .B(n21638), .Z(n21641) );
  XNOR U21365 ( .A(n21658), .B(n21659), .Z(n21550) );
  AND U21366 ( .A(n376), .B(n21660), .Z(n21659) );
  XOR U21367 ( .A(n21661), .B(n21658), .Z(n21660) );
  XNOR U21368 ( .A(n21662), .B(n21638), .Z(n21657) );
  IV U21369 ( .A(n21501), .Z(n21662) );
  XOR U21370 ( .A(n21663), .B(n21664), .Z(n21501) );
  AND U21371 ( .A(n384), .B(n21665), .Z(n21664) );
  XOR U21372 ( .A(n21666), .B(n21667), .Z(n21638) );
  AND U21373 ( .A(n21668), .B(n21669), .Z(n21667) );
  XNOR U21374 ( .A(n21575), .B(n21666), .Z(n21669) );
  XNOR U21375 ( .A(n21670), .B(n21671), .Z(n21575) );
  AND U21376 ( .A(n376), .B(n21672), .Z(n21671) );
  XNOR U21377 ( .A(n21673), .B(n21670), .Z(n21672) );
  XOR U21378 ( .A(n21666), .B(n21512), .Z(n21668) );
  XOR U21379 ( .A(n21674), .B(n21675), .Z(n21512) );
  AND U21380 ( .A(n384), .B(n21676), .Z(n21675) );
  XOR U21381 ( .A(n21677), .B(n21678), .Z(n21666) );
  AND U21382 ( .A(n21679), .B(n21680), .Z(n21678) );
  XNOR U21383 ( .A(n21677), .B(n21621), .Z(n21680) );
  XNOR U21384 ( .A(n21681), .B(n21682), .Z(n21621) );
  AND U21385 ( .A(n376), .B(n21683), .Z(n21682) );
  XOR U21386 ( .A(n21684), .B(n21681), .Z(n21683) );
  XNOR U21387 ( .A(n21685), .B(n21677), .Z(n21679) );
  IV U21388 ( .A(n21524), .Z(n21685) );
  XOR U21389 ( .A(n21686), .B(n21687), .Z(n21524) );
  AND U21390 ( .A(n384), .B(n21688), .Z(n21687) );
  AND U21391 ( .A(n21642), .B(n21631), .Z(n21677) );
  XNOR U21392 ( .A(n21689), .B(n21690), .Z(n21631) );
  AND U21393 ( .A(n376), .B(n21691), .Z(n21690) );
  XNOR U21394 ( .A(n21692), .B(n21689), .Z(n21691) );
  XNOR U21395 ( .A(n21693), .B(n21694), .Z(n376) );
  AND U21396 ( .A(n21695), .B(n21696), .Z(n21694) );
  XOR U21397 ( .A(n21652), .B(n21693), .Z(n21696) );
  AND U21398 ( .A(n21697), .B(n21698), .Z(n21652) );
  XOR U21399 ( .A(n21693), .B(n21649), .Z(n21695) );
  XNOR U21400 ( .A(n21699), .B(n21700), .Z(n21649) );
  AND U21401 ( .A(n380), .B(n21655), .Z(n21700) );
  XOR U21402 ( .A(n21653), .B(n21699), .Z(n21655) );
  XOR U21403 ( .A(n21701), .B(n21702), .Z(n21693) );
  AND U21404 ( .A(n21703), .B(n21704), .Z(n21702) );
  XNOR U21405 ( .A(n21701), .B(n21697), .Z(n21704) );
  IV U21406 ( .A(n21661), .Z(n21697) );
  XOR U21407 ( .A(n21705), .B(n21706), .Z(n21661) );
  XOR U21408 ( .A(n21707), .B(n21698), .Z(n21706) );
  AND U21409 ( .A(n21673), .B(n21708), .Z(n21698) );
  AND U21410 ( .A(n21709), .B(n21710), .Z(n21707) );
  XOR U21411 ( .A(n21711), .B(n21705), .Z(n21709) );
  XNOR U21412 ( .A(n21658), .B(n21701), .Z(n21703) );
  XNOR U21413 ( .A(n21712), .B(n21713), .Z(n21658) );
  AND U21414 ( .A(n380), .B(n21665), .Z(n21713) );
  XOR U21415 ( .A(n21712), .B(n21663), .Z(n21665) );
  XOR U21416 ( .A(n21714), .B(n21715), .Z(n21701) );
  AND U21417 ( .A(n21716), .B(n21717), .Z(n21715) );
  XNOR U21418 ( .A(n21714), .B(n21673), .Z(n21717) );
  XOR U21419 ( .A(n21718), .B(n21710), .Z(n21673) );
  XNOR U21420 ( .A(n21719), .B(n21705), .Z(n21710) );
  XOR U21421 ( .A(n21720), .B(n21721), .Z(n21705) );
  AND U21422 ( .A(n21722), .B(n21723), .Z(n21721) );
  XOR U21423 ( .A(n21724), .B(n21720), .Z(n21722) );
  XNOR U21424 ( .A(n21725), .B(n21726), .Z(n21719) );
  AND U21425 ( .A(n21727), .B(n21728), .Z(n21726) );
  XOR U21426 ( .A(n21725), .B(n21729), .Z(n21727) );
  XNOR U21427 ( .A(n21711), .B(n21708), .Z(n21718) );
  AND U21428 ( .A(n21730), .B(n21731), .Z(n21708) );
  XOR U21429 ( .A(n21732), .B(n21733), .Z(n21711) );
  AND U21430 ( .A(n21734), .B(n21735), .Z(n21733) );
  XOR U21431 ( .A(n21732), .B(n21736), .Z(n21734) );
  XNOR U21432 ( .A(n21670), .B(n21714), .Z(n21716) );
  XNOR U21433 ( .A(n21737), .B(n21738), .Z(n21670) );
  AND U21434 ( .A(n380), .B(n21676), .Z(n21738) );
  XOR U21435 ( .A(n21737), .B(n21674), .Z(n21676) );
  XOR U21436 ( .A(n21739), .B(n21740), .Z(n21714) );
  AND U21437 ( .A(n21741), .B(n21742), .Z(n21740) );
  XNOR U21438 ( .A(n21739), .B(n21730), .Z(n21742) );
  IV U21439 ( .A(n21684), .Z(n21730) );
  XNOR U21440 ( .A(n21743), .B(n21723), .Z(n21684) );
  XNOR U21441 ( .A(n21744), .B(n21729), .Z(n21723) );
  XOR U21442 ( .A(n21745), .B(n21746), .Z(n21729) );
  NOR U21443 ( .A(n21747), .B(n21748), .Z(n21746) );
  XNOR U21444 ( .A(n21745), .B(n21749), .Z(n21747) );
  XNOR U21445 ( .A(n21728), .B(n21720), .Z(n21744) );
  XOR U21446 ( .A(n21750), .B(n21751), .Z(n21720) );
  AND U21447 ( .A(n21752), .B(n21753), .Z(n21751) );
  XNOR U21448 ( .A(n21750), .B(n21754), .Z(n21752) );
  XNOR U21449 ( .A(n21755), .B(n21725), .Z(n21728) );
  XOR U21450 ( .A(n21756), .B(n21757), .Z(n21725) );
  AND U21451 ( .A(n21758), .B(n21759), .Z(n21757) );
  XOR U21452 ( .A(n21756), .B(n21760), .Z(n21758) );
  XNOR U21453 ( .A(n21761), .B(n21762), .Z(n21755) );
  NOR U21454 ( .A(n21763), .B(n21764), .Z(n21762) );
  XOR U21455 ( .A(n21761), .B(n21765), .Z(n21763) );
  XNOR U21456 ( .A(n21724), .B(n21731), .Z(n21743) );
  NOR U21457 ( .A(n21692), .B(n21766), .Z(n21731) );
  XOR U21458 ( .A(n21736), .B(n21735), .Z(n21724) );
  XNOR U21459 ( .A(n21767), .B(n21732), .Z(n21735) );
  XOR U21460 ( .A(n21768), .B(n21769), .Z(n21732) );
  AND U21461 ( .A(n21770), .B(n21771), .Z(n21769) );
  XOR U21462 ( .A(n21768), .B(n21772), .Z(n21770) );
  XNOR U21463 ( .A(n21773), .B(n21774), .Z(n21767) );
  NOR U21464 ( .A(n21775), .B(n21776), .Z(n21774) );
  XNOR U21465 ( .A(n21773), .B(n21777), .Z(n21775) );
  XOR U21466 ( .A(n21778), .B(n21779), .Z(n21736) );
  NOR U21467 ( .A(n21780), .B(n21781), .Z(n21779) );
  XNOR U21468 ( .A(n21778), .B(n21782), .Z(n21780) );
  XNOR U21469 ( .A(n21681), .B(n21739), .Z(n21741) );
  XNOR U21470 ( .A(n21783), .B(n21784), .Z(n21681) );
  AND U21471 ( .A(n380), .B(n21688), .Z(n21784) );
  XOR U21472 ( .A(n21783), .B(n21686), .Z(n21688) );
  AND U21473 ( .A(n21689), .B(n21692), .Z(n21739) );
  XOR U21474 ( .A(n21785), .B(n21766), .Z(n21692) );
  XNOR U21475 ( .A(p_input[2048]), .B(p_input[496]), .Z(n21766) );
  XOR U21476 ( .A(n21754), .B(n21753), .Z(n21785) );
  XNOR U21477 ( .A(n21786), .B(n21760), .Z(n21753) );
  XNOR U21478 ( .A(n21749), .B(n21748), .Z(n21760) );
  XOR U21479 ( .A(n21787), .B(n21745), .Z(n21748) );
  XNOR U21480 ( .A(n16904), .B(p_input[506]), .Z(n21745) );
  XNOR U21481 ( .A(p_input[2059]), .B(p_input[507]), .Z(n21787) );
  XOR U21482 ( .A(p_input[2060]), .B(p_input[508]), .Z(n21749) );
  XNOR U21483 ( .A(n21759), .B(n21750), .Z(n21786) );
  XNOR U21484 ( .A(n17068), .B(p_input[497]), .Z(n21750) );
  XOR U21485 ( .A(n21788), .B(n21765), .Z(n21759) );
  XNOR U21486 ( .A(p_input[2063]), .B(p_input[511]), .Z(n21765) );
  XOR U21487 ( .A(n21756), .B(n21764), .Z(n21788) );
  XOR U21488 ( .A(n21789), .B(n21761), .Z(n21764) );
  XOR U21489 ( .A(p_input[2061]), .B(p_input[509]), .Z(n21761) );
  XNOR U21490 ( .A(p_input[2062]), .B(p_input[510]), .Z(n21789) );
  XNOR U21491 ( .A(n16738), .B(p_input[505]), .Z(n21756) );
  XNOR U21492 ( .A(n21772), .B(n21771), .Z(n21754) );
  XNOR U21493 ( .A(n21790), .B(n21777), .Z(n21771) );
  XOR U21494 ( .A(p_input[2056]), .B(p_input[504]), .Z(n21777) );
  XOR U21495 ( .A(n21768), .B(n21776), .Z(n21790) );
  XOR U21496 ( .A(n21791), .B(n21773), .Z(n21776) );
  XOR U21497 ( .A(p_input[2054]), .B(p_input[502]), .Z(n21773) );
  XNOR U21498 ( .A(p_input[2055]), .B(p_input[503]), .Z(n21791) );
  XNOR U21499 ( .A(n16741), .B(p_input[498]), .Z(n21768) );
  XNOR U21500 ( .A(n21782), .B(n21781), .Z(n21772) );
  XOR U21501 ( .A(n21792), .B(n21778), .Z(n21781) );
  XOR U21502 ( .A(p_input[2051]), .B(p_input[499]), .Z(n21778) );
  XNOR U21503 ( .A(p_input[2052]), .B(p_input[500]), .Z(n21792) );
  XOR U21504 ( .A(p_input[2053]), .B(p_input[501]), .Z(n21782) );
  XNOR U21505 ( .A(n21793), .B(n21794), .Z(n21689) );
  AND U21506 ( .A(n380), .B(n21795), .Z(n21794) );
  XNOR U21507 ( .A(n21796), .B(n21797), .Z(n380) );
  AND U21508 ( .A(n21798), .B(n21799), .Z(n21797) );
  XOR U21509 ( .A(n21796), .B(n21699), .Z(n21799) );
  XNOR U21510 ( .A(n21796), .B(n21653), .Z(n21798) );
  XOR U21511 ( .A(n21800), .B(n21801), .Z(n21796) );
  AND U21512 ( .A(n21802), .B(n21803), .Z(n21801) );
  XOR U21513 ( .A(n21800), .B(n21663), .Z(n21802) );
  XOR U21514 ( .A(n21804), .B(n21805), .Z(n21642) );
  AND U21515 ( .A(n384), .B(n21795), .Z(n21805) );
  XNOR U21516 ( .A(n21793), .B(n21804), .Z(n21795) );
  XNOR U21517 ( .A(n21806), .B(n21807), .Z(n384) );
  AND U21518 ( .A(n21808), .B(n21809), .Z(n21807) );
  XNOR U21519 ( .A(n21810), .B(n21806), .Z(n21809) );
  IV U21520 ( .A(n21699), .Z(n21810) );
  XNOR U21521 ( .A(n21811), .B(n21812), .Z(n21699) );
  AND U21522 ( .A(n387), .B(n21813), .Z(n21812) );
  XNOR U21523 ( .A(n21811), .B(n21814), .Z(n21813) );
  XNOR U21524 ( .A(n21653), .B(n21806), .Z(n21808) );
  XOR U21525 ( .A(n21815), .B(n21816), .Z(n21653) );
  AND U21526 ( .A(n395), .B(n21817), .Z(n21816) );
  XOR U21527 ( .A(n21800), .B(n21818), .Z(n21806) );
  AND U21528 ( .A(n21819), .B(n21803), .Z(n21818) );
  XNOR U21529 ( .A(n21712), .B(n21800), .Z(n21803) );
  XNOR U21530 ( .A(n21820), .B(n21821), .Z(n21712) );
  AND U21531 ( .A(n387), .B(n21822), .Z(n21821) );
  XOR U21532 ( .A(n21823), .B(n21820), .Z(n21822) );
  XNOR U21533 ( .A(n21824), .B(n21800), .Z(n21819) );
  IV U21534 ( .A(n21663), .Z(n21824) );
  XOR U21535 ( .A(n21825), .B(n21826), .Z(n21663) );
  AND U21536 ( .A(n395), .B(n21827), .Z(n21826) );
  XOR U21537 ( .A(n21828), .B(n21829), .Z(n21800) );
  AND U21538 ( .A(n21830), .B(n21831), .Z(n21829) );
  XNOR U21539 ( .A(n21737), .B(n21828), .Z(n21831) );
  XNOR U21540 ( .A(n21832), .B(n21833), .Z(n21737) );
  AND U21541 ( .A(n387), .B(n21834), .Z(n21833) );
  XNOR U21542 ( .A(n21835), .B(n21832), .Z(n21834) );
  XOR U21543 ( .A(n21828), .B(n21674), .Z(n21830) );
  XOR U21544 ( .A(n21836), .B(n21837), .Z(n21674) );
  AND U21545 ( .A(n395), .B(n21838), .Z(n21837) );
  XOR U21546 ( .A(n21839), .B(n21840), .Z(n21828) );
  AND U21547 ( .A(n21841), .B(n21842), .Z(n21840) );
  XNOR U21548 ( .A(n21839), .B(n21783), .Z(n21842) );
  XNOR U21549 ( .A(n21843), .B(n21844), .Z(n21783) );
  AND U21550 ( .A(n387), .B(n21845), .Z(n21844) );
  XOR U21551 ( .A(n21846), .B(n21843), .Z(n21845) );
  XNOR U21552 ( .A(n21847), .B(n21839), .Z(n21841) );
  IV U21553 ( .A(n21686), .Z(n21847) );
  XOR U21554 ( .A(n21848), .B(n21849), .Z(n21686) );
  AND U21555 ( .A(n395), .B(n21850), .Z(n21849) );
  AND U21556 ( .A(n21804), .B(n21793), .Z(n21839) );
  XNOR U21557 ( .A(n21851), .B(n21852), .Z(n21793) );
  AND U21558 ( .A(n387), .B(n21853), .Z(n21852) );
  XNOR U21559 ( .A(n21854), .B(n21851), .Z(n21853) );
  XNOR U21560 ( .A(n21855), .B(n21856), .Z(n387) );
  AND U21561 ( .A(n21857), .B(n21858), .Z(n21856) );
  XOR U21562 ( .A(n21814), .B(n21855), .Z(n21858) );
  AND U21563 ( .A(n21859), .B(n21860), .Z(n21814) );
  XOR U21564 ( .A(n21855), .B(n21811), .Z(n21857) );
  XNOR U21565 ( .A(n21861), .B(n21862), .Z(n21811) );
  AND U21566 ( .A(n391), .B(n21817), .Z(n21862) );
  XOR U21567 ( .A(n21815), .B(n21861), .Z(n21817) );
  XOR U21568 ( .A(n21863), .B(n21864), .Z(n21855) );
  AND U21569 ( .A(n21865), .B(n21866), .Z(n21864) );
  XNOR U21570 ( .A(n21863), .B(n21859), .Z(n21866) );
  IV U21571 ( .A(n21823), .Z(n21859) );
  XOR U21572 ( .A(n21867), .B(n21868), .Z(n21823) );
  XOR U21573 ( .A(n21869), .B(n21860), .Z(n21868) );
  AND U21574 ( .A(n21835), .B(n21870), .Z(n21860) );
  AND U21575 ( .A(n21871), .B(n21872), .Z(n21869) );
  XOR U21576 ( .A(n21873), .B(n21867), .Z(n21871) );
  XNOR U21577 ( .A(n21820), .B(n21863), .Z(n21865) );
  XNOR U21578 ( .A(n21874), .B(n21875), .Z(n21820) );
  AND U21579 ( .A(n391), .B(n21827), .Z(n21875) );
  XOR U21580 ( .A(n21874), .B(n21825), .Z(n21827) );
  XOR U21581 ( .A(n21876), .B(n21877), .Z(n21863) );
  AND U21582 ( .A(n21878), .B(n21879), .Z(n21877) );
  XNOR U21583 ( .A(n21876), .B(n21835), .Z(n21879) );
  XOR U21584 ( .A(n21880), .B(n21872), .Z(n21835) );
  XNOR U21585 ( .A(n21881), .B(n21867), .Z(n21872) );
  XOR U21586 ( .A(n21882), .B(n21883), .Z(n21867) );
  AND U21587 ( .A(n21884), .B(n21885), .Z(n21883) );
  XOR U21588 ( .A(n21886), .B(n21882), .Z(n21884) );
  XNOR U21589 ( .A(n21887), .B(n21888), .Z(n21881) );
  AND U21590 ( .A(n21889), .B(n21890), .Z(n21888) );
  XOR U21591 ( .A(n21887), .B(n21891), .Z(n21889) );
  XNOR U21592 ( .A(n21873), .B(n21870), .Z(n21880) );
  AND U21593 ( .A(n21892), .B(n21893), .Z(n21870) );
  XOR U21594 ( .A(n21894), .B(n21895), .Z(n21873) );
  AND U21595 ( .A(n21896), .B(n21897), .Z(n21895) );
  XOR U21596 ( .A(n21894), .B(n21898), .Z(n21896) );
  XNOR U21597 ( .A(n21832), .B(n21876), .Z(n21878) );
  XNOR U21598 ( .A(n21899), .B(n21900), .Z(n21832) );
  AND U21599 ( .A(n391), .B(n21838), .Z(n21900) );
  XOR U21600 ( .A(n21899), .B(n21836), .Z(n21838) );
  XOR U21601 ( .A(n21901), .B(n21902), .Z(n21876) );
  AND U21602 ( .A(n21903), .B(n21904), .Z(n21902) );
  XNOR U21603 ( .A(n21901), .B(n21892), .Z(n21904) );
  IV U21604 ( .A(n21846), .Z(n21892) );
  XNOR U21605 ( .A(n21905), .B(n21885), .Z(n21846) );
  XNOR U21606 ( .A(n21906), .B(n21891), .Z(n21885) );
  XOR U21607 ( .A(n21907), .B(n21908), .Z(n21891) );
  NOR U21608 ( .A(n21909), .B(n21910), .Z(n21908) );
  XNOR U21609 ( .A(n21907), .B(n21911), .Z(n21909) );
  XNOR U21610 ( .A(n21890), .B(n21882), .Z(n21906) );
  XOR U21611 ( .A(n21912), .B(n21913), .Z(n21882) );
  AND U21612 ( .A(n21914), .B(n21915), .Z(n21913) );
  XNOR U21613 ( .A(n21912), .B(n21916), .Z(n21914) );
  XNOR U21614 ( .A(n21917), .B(n21887), .Z(n21890) );
  XOR U21615 ( .A(n21918), .B(n21919), .Z(n21887) );
  AND U21616 ( .A(n21920), .B(n21921), .Z(n21919) );
  XOR U21617 ( .A(n21918), .B(n21922), .Z(n21920) );
  XNOR U21618 ( .A(n21923), .B(n21924), .Z(n21917) );
  NOR U21619 ( .A(n21925), .B(n21926), .Z(n21924) );
  XOR U21620 ( .A(n21923), .B(n21927), .Z(n21925) );
  XNOR U21621 ( .A(n21886), .B(n21893), .Z(n21905) );
  NOR U21622 ( .A(n21854), .B(n21928), .Z(n21893) );
  XOR U21623 ( .A(n21898), .B(n21897), .Z(n21886) );
  XNOR U21624 ( .A(n21929), .B(n21894), .Z(n21897) );
  XOR U21625 ( .A(n21930), .B(n21931), .Z(n21894) );
  AND U21626 ( .A(n21932), .B(n21933), .Z(n21931) );
  XOR U21627 ( .A(n21930), .B(n21934), .Z(n21932) );
  XNOR U21628 ( .A(n21935), .B(n21936), .Z(n21929) );
  NOR U21629 ( .A(n21937), .B(n21938), .Z(n21936) );
  XNOR U21630 ( .A(n21935), .B(n21939), .Z(n21937) );
  XOR U21631 ( .A(n21940), .B(n21941), .Z(n21898) );
  NOR U21632 ( .A(n21942), .B(n21943), .Z(n21941) );
  XNOR U21633 ( .A(n21940), .B(n21944), .Z(n21942) );
  XNOR U21634 ( .A(n21843), .B(n21901), .Z(n21903) );
  XNOR U21635 ( .A(n21945), .B(n21946), .Z(n21843) );
  AND U21636 ( .A(n391), .B(n21850), .Z(n21946) );
  XOR U21637 ( .A(n21945), .B(n21848), .Z(n21850) );
  AND U21638 ( .A(n21851), .B(n21854), .Z(n21901) );
  XOR U21639 ( .A(n21947), .B(n21928), .Z(n21854) );
  XNOR U21640 ( .A(p_input[2048]), .B(p_input[512]), .Z(n21928) );
  XOR U21641 ( .A(n21916), .B(n21915), .Z(n21947) );
  XNOR U21642 ( .A(n21948), .B(n21922), .Z(n21915) );
  XNOR U21643 ( .A(n21911), .B(n21910), .Z(n21922) );
  XOR U21644 ( .A(n21949), .B(n21907), .Z(n21910) );
  XNOR U21645 ( .A(n16904), .B(p_input[522]), .Z(n21907) );
  XNOR U21646 ( .A(p_input[2059]), .B(p_input[523]), .Z(n21949) );
  XOR U21647 ( .A(p_input[2060]), .B(p_input[524]), .Z(n21911) );
  XNOR U21648 ( .A(n21921), .B(n21912), .Z(n21948) );
  XNOR U21649 ( .A(n17068), .B(p_input[513]), .Z(n21912) );
  XOR U21650 ( .A(n21950), .B(n21927), .Z(n21921) );
  XNOR U21651 ( .A(p_input[2063]), .B(p_input[527]), .Z(n21927) );
  XOR U21652 ( .A(n21918), .B(n21926), .Z(n21950) );
  XOR U21653 ( .A(n21951), .B(n21923), .Z(n21926) );
  XOR U21654 ( .A(p_input[2061]), .B(p_input[525]), .Z(n21923) );
  XNOR U21655 ( .A(p_input[2062]), .B(p_input[526]), .Z(n21951) );
  XNOR U21656 ( .A(n16738), .B(p_input[521]), .Z(n21918) );
  XNOR U21657 ( .A(n21934), .B(n21933), .Z(n21916) );
  XNOR U21658 ( .A(n21952), .B(n21939), .Z(n21933) );
  XOR U21659 ( .A(p_input[2056]), .B(p_input[520]), .Z(n21939) );
  XOR U21660 ( .A(n21930), .B(n21938), .Z(n21952) );
  XOR U21661 ( .A(n21953), .B(n21935), .Z(n21938) );
  XOR U21662 ( .A(p_input[2054]), .B(p_input[518]), .Z(n21935) );
  XNOR U21663 ( .A(p_input[2055]), .B(p_input[519]), .Z(n21953) );
  XNOR U21664 ( .A(n16741), .B(p_input[514]), .Z(n21930) );
  XNOR U21665 ( .A(n21944), .B(n21943), .Z(n21934) );
  XOR U21666 ( .A(n21954), .B(n21940), .Z(n21943) );
  XOR U21667 ( .A(p_input[2051]), .B(p_input[515]), .Z(n21940) );
  XNOR U21668 ( .A(p_input[2052]), .B(p_input[516]), .Z(n21954) );
  XOR U21669 ( .A(p_input[2053]), .B(p_input[517]), .Z(n21944) );
  XNOR U21670 ( .A(n21955), .B(n21956), .Z(n21851) );
  AND U21671 ( .A(n391), .B(n21957), .Z(n21956) );
  XNOR U21672 ( .A(n21958), .B(n21959), .Z(n391) );
  AND U21673 ( .A(n21960), .B(n21961), .Z(n21959) );
  XOR U21674 ( .A(n21958), .B(n21861), .Z(n21961) );
  XNOR U21675 ( .A(n21958), .B(n21815), .Z(n21960) );
  XOR U21676 ( .A(n21962), .B(n21963), .Z(n21958) );
  AND U21677 ( .A(n21964), .B(n21965), .Z(n21963) );
  XOR U21678 ( .A(n21962), .B(n21825), .Z(n21964) );
  XOR U21679 ( .A(n21966), .B(n21967), .Z(n21804) );
  AND U21680 ( .A(n395), .B(n21957), .Z(n21967) );
  XNOR U21681 ( .A(n21955), .B(n21966), .Z(n21957) );
  XNOR U21682 ( .A(n21968), .B(n21969), .Z(n395) );
  AND U21683 ( .A(n21970), .B(n21971), .Z(n21969) );
  XNOR U21684 ( .A(n21972), .B(n21968), .Z(n21971) );
  IV U21685 ( .A(n21861), .Z(n21972) );
  XNOR U21686 ( .A(n21973), .B(n21974), .Z(n21861) );
  AND U21687 ( .A(n398), .B(n21975), .Z(n21974) );
  XNOR U21688 ( .A(n21973), .B(n21976), .Z(n21975) );
  XNOR U21689 ( .A(n21815), .B(n21968), .Z(n21970) );
  XOR U21690 ( .A(n21977), .B(n21978), .Z(n21815) );
  AND U21691 ( .A(n406), .B(n21979), .Z(n21978) );
  XOR U21692 ( .A(n21962), .B(n21980), .Z(n21968) );
  AND U21693 ( .A(n21981), .B(n21965), .Z(n21980) );
  XNOR U21694 ( .A(n21874), .B(n21962), .Z(n21965) );
  XNOR U21695 ( .A(n21982), .B(n21983), .Z(n21874) );
  AND U21696 ( .A(n398), .B(n21984), .Z(n21983) );
  XOR U21697 ( .A(n21985), .B(n21982), .Z(n21984) );
  XNOR U21698 ( .A(n21986), .B(n21962), .Z(n21981) );
  IV U21699 ( .A(n21825), .Z(n21986) );
  XOR U21700 ( .A(n21987), .B(n21988), .Z(n21825) );
  AND U21701 ( .A(n406), .B(n21989), .Z(n21988) );
  XOR U21702 ( .A(n21990), .B(n21991), .Z(n21962) );
  AND U21703 ( .A(n21992), .B(n21993), .Z(n21991) );
  XNOR U21704 ( .A(n21899), .B(n21990), .Z(n21993) );
  XNOR U21705 ( .A(n21994), .B(n21995), .Z(n21899) );
  AND U21706 ( .A(n398), .B(n21996), .Z(n21995) );
  XNOR U21707 ( .A(n21997), .B(n21994), .Z(n21996) );
  XOR U21708 ( .A(n21990), .B(n21836), .Z(n21992) );
  XOR U21709 ( .A(n21998), .B(n21999), .Z(n21836) );
  AND U21710 ( .A(n406), .B(n22000), .Z(n21999) );
  XOR U21711 ( .A(n22001), .B(n22002), .Z(n21990) );
  AND U21712 ( .A(n22003), .B(n22004), .Z(n22002) );
  XNOR U21713 ( .A(n22001), .B(n21945), .Z(n22004) );
  XNOR U21714 ( .A(n22005), .B(n22006), .Z(n21945) );
  AND U21715 ( .A(n398), .B(n22007), .Z(n22006) );
  XOR U21716 ( .A(n22008), .B(n22005), .Z(n22007) );
  XNOR U21717 ( .A(n22009), .B(n22001), .Z(n22003) );
  IV U21718 ( .A(n21848), .Z(n22009) );
  XOR U21719 ( .A(n22010), .B(n22011), .Z(n21848) );
  AND U21720 ( .A(n406), .B(n22012), .Z(n22011) );
  AND U21721 ( .A(n21966), .B(n21955), .Z(n22001) );
  XNOR U21722 ( .A(n22013), .B(n22014), .Z(n21955) );
  AND U21723 ( .A(n398), .B(n22015), .Z(n22014) );
  XNOR U21724 ( .A(n22016), .B(n22013), .Z(n22015) );
  XNOR U21725 ( .A(n22017), .B(n22018), .Z(n398) );
  AND U21726 ( .A(n22019), .B(n22020), .Z(n22018) );
  XOR U21727 ( .A(n21976), .B(n22017), .Z(n22020) );
  AND U21728 ( .A(n22021), .B(n22022), .Z(n21976) );
  XOR U21729 ( .A(n22017), .B(n21973), .Z(n22019) );
  XNOR U21730 ( .A(n22023), .B(n22024), .Z(n21973) );
  AND U21731 ( .A(n402), .B(n21979), .Z(n22024) );
  XOR U21732 ( .A(n21977), .B(n22023), .Z(n21979) );
  XOR U21733 ( .A(n22025), .B(n22026), .Z(n22017) );
  AND U21734 ( .A(n22027), .B(n22028), .Z(n22026) );
  XNOR U21735 ( .A(n22025), .B(n22021), .Z(n22028) );
  IV U21736 ( .A(n21985), .Z(n22021) );
  XOR U21737 ( .A(n22029), .B(n22030), .Z(n21985) );
  XOR U21738 ( .A(n22031), .B(n22022), .Z(n22030) );
  AND U21739 ( .A(n21997), .B(n22032), .Z(n22022) );
  AND U21740 ( .A(n22033), .B(n22034), .Z(n22031) );
  XOR U21741 ( .A(n22035), .B(n22029), .Z(n22033) );
  XNOR U21742 ( .A(n21982), .B(n22025), .Z(n22027) );
  XNOR U21743 ( .A(n22036), .B(n22037), .Z(n21982) );
  AND U21744 ( .A(n402), .B(n21989), .Z(n22037) );
  XOR U21745 ( .A(n22036), .B(n21987), .Z(n21989) );
  XOR U21746 ( .A(n22038), .B(n22039), .Z(n22025) );
  AND U21747 ( .A(n22040), .B(n22041), .Z(n22039) );
  XNOR U21748 ( .A(n22038), .B(n21997), .Z(n22041) );
  XOR U21749 ( .A(n22042), .B(n22034), .Z(n21997) );
  XNOR U21750 ( .A(n22043), .B(n22029), .Z(n22034) );
  XOR U21751 ( .A(n22044), .B(n22045), .Z(n22029) );
  AND U21752 ( .A(n22046), .B(n22047), .Z(n22045) );
  XOR U21753 ( .A(n22048), .B(n22044), .Z(n22046) );
  XNOR U21754 ( .A(n22049), .B(n22050), .Z(n22043) );
  AND U21755 ( .A(n22051), .B(n22052), .Z(n22050) );
  XOR U21756 ( .A(n22049), .B(n22053), .Z(n22051) );
  XNOR U21757 ( .A(n22035), .B(n22032), .Z(n22042) );
  AND U21758 ( .A(n22054), .B(n22055), .Z(n22032) );
  XOR U21759 ( .A(n22056), .B(n22057), .Z(n22035) );
  AND U21760 ( .A(n22058), .B(n22059), .Z(n22057) );
  XOR U21761 ( .A(n22056), .B(n22060), .Z(n22058) );
  XNOR U21762 ( .A(n21994), .B(n22038), .Z(n22040) );
  XNOR U21763 ( .A(n22061), .B(n22062), .Z(n21994) );
  AND U21764 ( .A(n402), .B(n22000), .Z(n22062) );
  XOR U21765 ( .A(n22061), .B(n21998), .Z(n22000) );
  XOR U21766 ( .A(n22063), .B(n22064), .Z(n22038) );
  AND U21767 ( .A(n22065), .B(n22066), .Z(n22064) );
  XNOR U21768 ( .A(n22063), .B(n22054), .Z(n22066) );
  IV U21769 ( .A(n22008), .Z(n22054) );
  XNOR U21770 ( .A(n22067), .B(n22047), .Z(n22008) );
  XNOR U21771 ( .A(n22068), .B(n22053), .Z(n22047) );
  XOR U21772 ( .A(n22069), .B(n22070), .Z(n22053) );
  NOR U21773 ( .A(n22071), .B(n22072), .Z(n22070) );
  XNOR U21774 ( .A(n22069), .B(n22073), .Z(n22071) );
  XNOR U21775 ( .A(n22052), .B(n22044), .Z(n22068) );
  XOR U21776 ( .A(n22074), .B(n22075), .Z(n22044) );
  AND U21777 ( .A(n22076), .B(n22077), .Z(n22075) );
  XNOR U21778 ( .A(n22074), .B(n22078), .Z(n22076) );
  XNOR U21779 ( .A(n22079), .B(n22049), .Z(n22052) );
  XOR U21780 ( .A(n22080), .B(n22081), .Z(n22049) );
  AND U21781 ( .A(n22082), .B(n22083), .Z(n22081) );
  XOR U21782 ( .A(n22080), .B(n22084), .Z(n22082) );
  XNOR U21783 ( .A(n22085), .B(n22086), .Z(n22079) );
  NOR U21784 ( .A(n22087), .B(n22088), .Z(n22086) );
  XOR U21785 ( .A(n22085), .B(n22089), .Z(n22087) );
  XNOR U21786 ( .A(n22048), .B(n22055), .Z(n22067) );
  NOR U21787 ( .A(n22016), .B(n22090), .Z(n22055) );
  XOR U21788 ( .A(n22060), .B(n22059), .Z(n22048) );
  XNOR U21789 ( .A(n22091), .B(n22056), .Z(n22059) );
  XOR U21790 ( .A(n22092), .B(n22093), .Z(n22056) );
  AND U21791 ( .A(n22094), .B(n22095), .Z(n22093) );
  XOR U21792 ( .A(n22092), .B(n22096), .Z(n22094) );
  XNOR U21793 ( .A(n22097), .B(n22098), .Z(n22091) );
  NOR U21794 ( .A(n22099), .B(n22100), .Z(n22098) );
  XNOR U21795 ( .A(n22097), .B(n22101), .Z(n22099) );
  XOR U21796 ( .A(n22102), .B(n22103), .Z(n22060) );
  NOR U21797 ( .A(n22104), .B(n22105), .Z(n22103) );
  XNOR U21798 ( .A(n22102), .B(n22106), .Z(n22104) );
  XNOR U21799 ( .A(n22005), .B(n22063), .Z(n22065) );
  XNOR U21800 ( .A(n22107), .B(n22108), .Z(n22005) );
  AND U21801 ( .A(n402), .B(n22012), .Z(n22108) );
  XOR U21802 ( .A(n22107), .B(n22010), .Z(n22012) );
  AND U21803 ( .A(n22013), .B(n22016), .Z(n22063) );
  XOR U21804 ( .A(n22109), .B(n22090), .Z(n22016) );
  XNOR U21805 ( .A(p_input[2048]), .B(p_input[528]), .Z(n22090) );
  XOR U21806 ( .A(n22078), .B(n22077), .Z(n22109) );
  XNOR U21807 ( .A(n22110), .B(n22084), .Z(n22077) );
  XNOR U21808 ( .A(n22073), .B(n22072), .Z(n22084) );
  XOR U21809 ( .A(n22111), .B(n22069), .Z(n22072) );
  XNOR U21810 ( .A(n16904), .B(p_input[538]), .Z(n22069) );
  XNOR U21811 ( .A(p_input[2059]), .B(p_input[539]), .Z(n22111) );
  XOR U21812 ( .A(p_input[2060]), .B(p_input[540]), .Z(n22073) );
  XNOR U21813 ( .A(n22083), .B(n22074), .Z(n22110) );
  XNOR U21814 ( .A(n17068), .B(p_input[529]), .Z(n22074) );
  XOR U21815 ( .A(n22112), .B(n22089), .Z(n22083) );
  XNOR U21816 ( .A(p_input[2063]), .B(p_input[543]), .Z(n22089) );
  XOR U21817 ( .A(n22080), .B(n22088), .Z(n22112) );
  XOR U21818 ( .A(n22113), .B(n22085), .Z(n22088) );
  XOR U21819 ( .A(p_input[2061]), .B(p_input[541]), .Z(n22085) );
  XNOR U21820 ( .A(p_input[2062]), .B(p_input[542]), .Z(n22113) );
  XNOR U21821 ( .A(n16738), .B(p_input[537]), .Z(n22080) );
  XNOR U21822 ( .A(n22096), .B(n22095), .Z(n22078) );
  XNOR U21823 ( .A(n22114), .B(n22101), .Z(n22095) );
  XOR U21824 ( .A(p_input[2056]), .B(p_input[536]), .Z(n22101) );
  XOR U21825 ( .A(n22092), .B(n22100), .Z(n22114) );
  XOR U21826 ( .A(n22115), .B(n22097), .Z(n22100) );
  XOR U21827 ( .A(p_input[2054]), .B(p_input[534]), .Z(n22097) );
  XNOR U21828 ( .A(p_input[2055]), .B(p_input[535]), .Z(n22115) );
  XNOR U21829 ( .A(n16741), .B(p_input[530]), .Z(n22092) );
  XNOR U21830 ( .A(n22106), .B(n22105), .Z(n22096) );
  XOR U21831 ( .A(n22116), .B(n22102), .Z(n22105) );
  XOR U21832 ( .A(p_input[2051]), .B(p_input[531]), .Z(n22102) );
  XNOR U21833 ( .A(p_input[2052]), .B(p_input[532]), .Z(n22116) );
  XOR U21834 ( .A(p_input[2053]), .B(p_input[533]), .Z(n22106) );
  XNOR U21835 ( .A(n22117), .B(n22118), .Z(n22013) );
  AND U21836 ( .A(n402), .B(n22119), .Z(n22118) );
  XNOR U21837 ( .A(n22120), .B(n22121), .Z(n402) );
  AND U21838 ( .A(n22122), .B(n22123), .Z(n22121) );
  XOR U21839 ( .A(n22120), .B(n22023), .Z(n22123) );
  XNOR U21840 ( .A(n22120), .B(n21977), .Z(n22122) );
  XOR U21841 ( .A(n22124), .B(n22125), .Z(n22120) );
  AND U21842 ( .A(n22126), .B(n22127), .Z(n22125) );
  XOR U21843 ( .A(n22124), .B(n21987), .Z(n22126) );
  XOR U21844 ( .A(n22128), .B(n22129), .Z(n21966) );
  AND U21845 ( .A(n406), .B(n22119), .Z(n22129) );
  XNOR U21846 ( .A(n22117), .B(n22128), .Z(n22119) );
  XNOR U21847 ( .A(n22130), .B(n22131), .Z(n406) );
  AND U21848 ( .A(n22132), .B(n22133), .Z(n22131) );
  XNOR U21849 ( .A(n22134), .B(n22130), .Z(n22133) );
  IV U21850 ( .A(n22023), .Z(n22134) );
  XNOR U21851 ( .A(n22135), .B(n22136), .Z(n22023) );
  AND U21852 ( .A(n409), .B(n22137), .Z(n22136) );
  XNOR U21853 ( .A(n22135), .B(n22138), .Z(n22137) );
  XNOR U21854 ( .A(n21977), .B(n22130), .Z(n22132) );
  XOR U21855 ( .A(n22139), .B(n22140), .Z(n21977) );
  AND U21856 ( .A(n417), .B(n22141), .Z(n22140) );
  XOR U21857 ( .A(n22124), .B(n22142), .Z(n22130) );
  AND U21858 ( .A(n22143), .B(n22127), .Z(n22142) );
  XNOR U21859 ( .A(n22036), .B(n22124), .Z(n22127) );
  XNOR U21860 ( .A(n22144), .B(n22145), .Z(n22036) );
  AND U21861 ( .A(n409), .B(n22146), .Z(n22145) );
  XOR U21862 ( .A(n22147), .B(n22144), .Z(n22146) );
  XNOR U21863 ( .A(n22148), .B(n22124), .Z(n22143) );
  IV U21864 ( .A(n21987), .Z(n22148) );
  XOR U21865 ( .A(n22149), .B(n22150), .Z(n21987) );
  AND U21866 ( .A(n417), .B(n22151), .Z(n22150) );
  XOR U21867 ( .A(n22152), .B(n22153), .Z(n22124) );
  AND U21868 ( .A(n22154), .B(n22155), .Z(n22153) );
  XNOR U21869 ( .A(n22061), .B(n22152), .Z(n22155) );
  XNOR U21870 ( .A(n22156), .B(n22157), .Z(n22061) );
  AND U21871 ( .A(n409), .B(n22158), .Z(n22157) );
  XNOR U21872 ( .A(n22159), .B(n22156), .Z(n22158) );
  XOR U21873 ( .A(n22152), .B(n21998), .Z(n22154) );
  XOR U21874 ( .A(n22160), .B(n22161), .Z(n21998) );
  AND U21875 ( .A(n417), .B(n22162), .Z(n22161) );
  XOR U21876 ( .A(n22163), .B(n22164), .Z(n22152) );
  AND U21877 ( .A(n22165), .B(n22166), .Z(n22164) );
  XNOR U21878 ( .A(n22163), .B(n22107), .Z(n22166) );
  XNOR U21879 ( .A(n22167), .B(n22168), .Z(n22107) );
  AND U21880 ( .A(n409), .B(n22169), .Z(n22168) );
  XOR U21881 ( .A(n22170), .B(n22167), .Z(n22169) );
  XNOR U21882 ( .A(n22171), .B(n22163), .Z(n22165) );
  IV U21883 ( .A(n22010), .Z(n22171) );
  XOR U21884 ( .A(n22172), .B(n22173), .Z(n22010) );
  AND U21885 ( .A(n417), .B(n22174), .Z(n22173) );
  AND U21886 ( .A(n22128), .B(n22117), .Z(n22163) );
  XNOR U21887 ( .A(n22175), .B(n22176), .Z(n22117) );
  AND U21888 ( .A(n409), .B(n22177), .Z(n22176) );
  XNOR U21889 ( .A(n22178), .B(n22175), .Z(n22177) );
  XNOR U21890 ( .A(n22179), .B(n22180), .Z(n409) );
  AND U21891 ( .A(n22181), .B(n22182), .Z(n22180) );
  XOR U21892 ( .A(n22138), .B(n22179), .Z(n22182) );
  AND U21893 ( .A(n22183), .B(n22184), .Z(n22138) );
  XOR U21894 ( .A(n22179), .B(n22135), .Z(n22181) );
  XNOR U21895 ( .A(n22185), .B(n22186), .Z(n22135) );
  AND U21896 ( .A(n413), .B(n22141), .Z(n22186) );
  XOR U21897 ( .A(n22139), .B(n22185), .Z(n22141) );
  XOR U21898 ( .A(n22187), .B(n22188), .Z(n22179) );
  AND U21899 ( .A(n22189), .B(n22190), .Z(n22188) );
  XNOR U21900 ( .A(n22187), .B(n22183), .Z(n22190) );
  IV U21901 ( .A(n22147), .Z(n22183) );
  XOR U21902 ( .A(n22191), .B(n22192), .Z(n22147) );
  XOR U21903 ( .A(n22193), .B(n22184), .Z(n22192) );
  AND U21904 ( .A(n22159), .B(n22194), .Z(n22184) );
  AND U21905 ( .A(n22195), .B(n22196), .Z(n22193) );
  XOR U21906 ( .A(n22197), .B(n22191), .Z(n22195) );
  XNOR U21907 ( .A(n22144), .B(n22187), .Z(n22189) );
  XNOR U21908 ( .A(n22198), .B(n22199), .Z(n22144) );
  AND U21909 ( .A(n413), .B(n22151), .Z(n22199) );
  XOR U21910 ( .A(n22198), .B(n22149), .Z(n22151) );
  XOR U21911 ( .A(n22200), .B(n22201), .Z(n22187) );
  AND U21912 ( .A(n22202), .B(n22203), .Z(n22201) );
  XNOR U21913 ( .A(n22200), .B(n22159), .Z(n22203) );
  XOR U21914 ( .A(n22204), .B(n22196), .Z(n22159) );
  XNOR U21915 ( .A(n22205), .B(n22191), .Z(n22196) );
  XOR U21916 ( .A(n22206), .B(n22207), .Z(n22191) );
  AND U21917 ( .A(n22208), .B(n22209), .Z(n22207) );
  XOR U21918 ( .A(n22210), .B(n22206), .Z(n22208) );
  XNOR U21919 ( .A(n22211), .B(n22212), .Z(n22205) );
  AND U21920 ( .A(n22213), .B(n22214), .Z(n22212) );
  XOR U21921 ( .A(n22211), .B(n22215), .Z(n22213) );
  XNOR U21922 ( .A(n22197), .B(n22194), .Z(n22204) );
  AND U21923 ( .A(n22216), .B(n22217), .Z(n22194) );
  XOR U21924 ( .A(n22218), .B(n22219), .Z(n22197) );
  AND U21925 ( .A(n22220), .B(n22221), .Z(n22219) );
  XOR U21926 ( .A(n22218), .B(n22222), .Z(n22220) );
  XNOR U21927 ( .A(n22156), .B(n22200), .Z(n22202) );
  XNOR U21928 ( .A(n22223), .B(n22224), .Z(n22156) );
  AND U21929 ( .A(n413), .B(n22162), .Z(n22224) );
  XOR U21930 ( .A(n22223), .B(n22160), .Z(n22162) );
  XOR U21931 ( .A(n22225), .B(n22226), .Z(n22200) );
  AND U21932 ( .A(n22227), .B(n22228), .Z(n22226) );
  XNOR U21933 ( .A(n22225), .B(n22216), .Z(n22228) );
  IV U21934 ( .A(n22170), .Z(n22216) );
  XNOR U21935 ( .A(n22229), .B(n22209), .Z(n22170) );
  XNOR U21936 ( .A(n22230), .B(n22215), .Z(n22209) );
  XOR U21937 ( .A(n22231), .B(n22232), .Z(n22215) );
  NOR U21938 ( .A(n22233), .B(n22234), .Z(n22232) );
  XNOR U21939 ( .A(n22231), .B(n22235), .Z(n22233) );
  XNOR U21940 ( .A(n22214), .B(n22206), .Z(n22230) );
  XOR U21941 ( .A(n22236), .B(n22237), .Z(n22206) );
  AND U21942 ( .A(n22238), .B(n22239), .Z(n22237) );
  XNOR U21943 ( .A(n22236), .B(n22240), .Z(n22238) );
  XNOR U21944 ( .A(n22241), .B(n22211), .Z(n22214) );
  XOR U21945 ( .A(n22242), .B(n22243), .Z(n22211) );
  AND U21946 ( .A(n22244), .B(n22245), .Z(n22243) );
  XOR U21947 ( .A(n22242), .B(n22246), .Z(n22244) );
  XNOR U21948 ( .A(n22247), .B(n22248), .Z(n22241) );
  NOR U21949 ( .A(n22249), .B(n22250), .Z(n22248) );
  XOR U21950 ( .A(n22247), .B(n22251), .Z(n22249) );
  XNOR U21951 ( .A(n22210), .B(n22217), .Z(n22229) );
  NOR U21952 ( .A(n22178), .B(n22252), .Z(n22217) );
  XOR U21953 ( .A(n22222), .B(n22221), .Z(n22210) );
  XNOR U21954 ( .A(n22253), .B(n22218), .Z(n22221) );
  XOR U21955 ( .A(n22254), .B(n22255), .Z(n22218) );
  AND U21956 ( .A(n22256), .B(n22257), .Z(n22255) );
  XOR U21957 ( .A(n22254), .B(n22258), .Z(n22256) );
  XNOR U21958 ( .A(n22259), .B(n22260), .Z(n22253) );
  NOR U21959 ( .A(n22261), .B(n22262), .Z(n22260) );
  XNOR U21960 ( .A(n22259), .B(n22263), .Z(n22261) );
  XOR U21961 ( .A(n22264), .B(n22265), .Z(n22222) );
  NOR U21962 ( .A(n22266), .B(n22267), .Z(n22265) );
  XNOR U21963 ( .A(n22264), .B(n22268), .Z(n22266) );
  XNOR U21964 ( .A(n22167), .B(n22225), .Z(n22227) );
  XNOR U21965 ( .A(n22269), .B(n22270), .Z(n22167) );
  AND U21966 ( .A(n413), .B(n22174), .Z(n22270) );
  XOR U21967 ( .A(n22269), .B(n22172), .Z(n22174) );
  AND U21968 ( .A(n22175), .B(n22178), .Z(n22225) );
  XOR U21969 ( .A(n22271), .B(n22252), .Z(n22178) );
  XNOR U21970 ( .A(p_input[2048]), .B(p_input[544]), .Z(n22252) );
  XOR U21971 ( .A(n22240), .B(n22239), .Z(n22271) );
  XNOR U21972 ( .A(n22272), .B(n22246), .Z(n22239) );
  XNOR U21973 ( .A(n22235), .B(n22234), .Z(n22246) );
  XOR U21974 ( .A(n22273), .B(n22231), .Z(n22234) );
  XNOR U21975 ( .A(n16904), .B(p_input[554]), .Z(n22231) );
  XNOR U21976 ( .A(p_input[2059]), .B(p_input[555]), .Z(n22273) );
  XOR U21977 ( .A(p_input[2060]), .B(p_input[556]), .Z(n22235) );
  XNOR U21978 ( .A(n22245), .B(n22236), .Z(n22272) );
  XNOR U21979 ( .A(n17068), .B(p_input[545]), .Z(n22236) );
  XOR U21980 ( .A(n22274), .B(n22251), .Z(n22245) );
  XNOR U21981 ( .A(p_input[2063]), .B(p_input[559]), .Z(n22251) );
  XOR U21982 ( .A(n22242), .B(n22250), .Z(n22274) );
  XOR U21983 ( .A(n22275), .B(n22247), .Z(n22250) );
  XOR U21984 ( .A(p_input[2061]), .B(p_input[557]), .Z(n22247) );
  XNOR U21985 ( .A(p_input[2062]), .B(p_input[558]), .Z(n22275) );
  XNOR U21986 ( .A(n16738), .B(p_input[553]), .Z(n22242) );
  XNOR U21987 ( .A(n22258), .B(n22257), .Z(n22240) );
  XNOR U21988 ( .A(n22276), .B(n22263), .Z(n22257) );
  XOR U21989 ( .A(p_input[2056]), .B(p_input[552]), .Z(n22263) );
  XOR U21990 ( .A(n22254), .B(n22262), .Z(n22276) );
  XOR U21991 ( .A(n22277), .B(n22259), .Z(n22262) );
  XOR U21992 ( .A(p_input[2054]), .B(p_input[550]), .Z(n22259) );
  XNOR U21993 ( .A(p_input[2055]), .B(p_input[551]), .Z(n22277) );
  XNOR U21994 ( .A(n16741), .B(p_input[546]), .Z(n22254) );
  XNOR U21995 ( .A(n22268), .B(n22267), .Z(n22258) );
  XOR U21996 ( .A(n22278), .B(n22264), .Z(n22267) );
  XOR U21997 ( .A(p_input[2051]), .B(p_input[547]), .Z(n22264) );
  XNOR U21998 ( .A(p_input[2052]), .B(p_input[548]), .Z(n22278) );
  XOR U21999 ( .A(p_input[2053]), .B(p_input[549]), .Z(n22268) );
  XNOR U22000 ( .A(n22279), .B(n22280), .Z(n22175) );
  AND U22001 ( .A(n413), .B(n22281), .Z(n22280) );
  XNOR U22002 ( .A(n22282), .B(n22283), .Z(n413) );
  AND U22003 ( .A(n22284), .B(n22285), .Z(n22283) );
  XOR U22004 ( .A(n22282), .B(n22185), .Z(n22285) );
  XNOR U22005 ( .A(n22282), .B(n22139), .Z(n22284) );
  XOR U22006 ( .A(n22286), .B(n22287), .Z(n22282) );
  AND U22007 ( .A(n22288), .B(n22289), .Z(n22287) );
  XOR U22008 ( .A(n22286), .B(n22149), .Z(n22288) );
  XOR U22009 ( .A(n22290), .B(n22291), .Z(n22128) );
  AND U22010 ( .A(n417), .B(n22281), .Z(n22291) );
  XNOR U22011 ( .A(n22279), .B(n22290), .Z(n22281) );
  XNOR U22012 ( .A(n22292), .B(n22293), .Z(n417) );
  AND U22013 ( .A(n22294), .B(n22295), .Z(n22293) );
  XNOR U22014 ( .A(n22296), .B(n22292), .Z(n22295) );
  IV U22015 ( .A(n22185), .Z(n22296) );
  XNOR U22016 ( .A(n22297), .B(n22298), .Z(n22185) );
  AND U22017 ( .A(n420), .B(n22299), .Z(n22298) );
  XNOR U22018 ( .A(n22297), .B(n22300), .Z(n22299) );
  XNOR U22019 ( .A(n22139), .B(n22292), .Z(n22294) );
  XOR U22020 ( .A(n22301), .B(n22302), .Z(n22139) );
  AND U22021 ( .A(n428), .B(n22303), .Z(n22302) );
  XOR U22022 ( .A(n22286), .B(n22304), .Z(n22292) );
  AND U22023 ( .A(n22305), .B(n22289), .Z(n22304) );
  XNOR U22024 ( .A(n22198), .B(n22286), .Z(n22289) );
  XNOR U22025 ( .A(n22306), .B(n22307), .Z(n22198) );
  AND U22026 ( .A(n420), .B(n22308), .Z(n22307) );
  XOR U22027 ( .A(n22309), .B(n22306), .Z(n22308) );
  XNOR U22028 ( .A(n22310), .B(n22286), .Z(n22305) );
  IV U22029 ( .A(n22149), .Z(n22310) );
  XOR U22030 ( .A(n22311), .B(n22312), .Z(n22149) );
  AND U22031 ( .A(n428), .B(n22313), .Z(n22312) );
  XOR U22032 ( .A(n22314), .B(n22315), .Z(n22286) );
  AND U22033 ( .A(n22316), .B(n22317), .Z(n22315) );
  XNOR U22034 ( .A(n22223), .B(n22314), .Z(n22317) );
  XNOR U22035 ( .A(n22318), .B(n22319), .Z(n22223) );
  AND U22036 ( .A(n420), .B(n22320), .Z(n22319) );
  XNOR U22037 ( .A(n22321), .B(n22318), .Z(n22320) );
  XOR U22038 ( .A(n22314), .B(n22160), .Z(n22316) );
  XOR U22039 ( .A(n22322), .B(n22323), .Z(n22160) );
  AND U22040 ( .A(n428), .B(n22324), .Z(n22323) );
  XOR U22041 ( .A(n22325), .B(n22326), .Z(n22314) );
  AND U22042 ( .A(n22327), .B(n22328), .Z(n22326) );
  XNOR U22043 ( .A(n22325), .B(n22269), .Z(n22328) );
  XNOR U22044 ( .A(n22329), .B(n22330), .Z(n22269) );
  AND U22045 ( .A(n420), .B(n22331), .Z(n22330) );
  XOR U22046 ( .A(n22332), .B(n22329), .Z(n22331) );
  XNOR U22047 ( .A(n22333), .B(n22325), .Z(n22327) );
  IV U22048 ( .A(n22172), .Z(n22333) );
  XOR U22049 ( .A(n22334), .B(n22335), .Z(n22172) );
  AND U22050 ( .A(n428), .B(n22336), .Z(n22335) );
  AND U22051 ( .A(n22290), .B(n22279), .Z(n22325) );
  XNOR U22052 ( .A(n22337), .B(n22338), .Z(n22279) );
  AND U22053 ( .A(n420), .B(n22339), .Z(n22338) );
  XNOR U22054 ( .A(n22340), .B(n22337), .Z(n22339) );
  XNOR U22055 ( .A(n22341), .B(n22342), .Z(n420) );
  AND U22056 ( .A(n22343), .B(n22344), .Z(n22342) );
  XOR U22057 ( .A(n22300), .B(n22341), .Z(n22344) );
  AND U22058 ( .A(n22345), .B(n22346), .Z(n22300) );
  XOR U22059 ( .A(n22341), .B(n22297), .Z(n22343) );
  XNOR U22060 ( .A(n22347), .B(n22348), .Z(n22297) );
  AND U22061 ( .A(n424), .B(n22303), .Z(n22348) );
  XOR U22062 ( .A(n22301), .B(n22347), .Z(n22303) );
  XOR U22063 ( .A(n22349), .B(n22350), .Z(n22341) );
  AND U22064 ( .A(n22351), .B(n22352), .Z(n22350) );
  XNOR U22065 ( .A(n22349), .B(n22345), .Z(n22352) );
  IV U22066 ( .A(n22309), .Z(n22345) );
  XOR U22067 ( .A(n22353), .B(n22354), .Z(n22309) );
  XOR U22068 ( .A(n22355), .B(n22346), .Z(n22354) );
  AND U22069 ( .A(n22321), .B(n22356), .Z(n22346) );
  AND U22070 ( .A(n22357), .B(n22358), .Z(n22355) );
  XOR U22071 ( .A(n22359), .B(n22353), .Z(n22357) );
  XNOR U22072 ( .A(n22306), .B(n22349), .Z(n22351) );
  XNOR U22073 ( .A(n22360), .B(n22361), .Z(n22306) );
  AND U22074 ( .A(n424), .B(n22313), .Z(n22361) );
  XOR U22075 ( .A(n22360), .B(n22311), .Z(n22313) );
  XOR U22076 ( .A(n22362), .B(n22363), .Z(n22349) );
  AND U22077 ( .A(n22364), .B(n22365), .Z(n22363) );
  XNOR U22078 ( .A(n22362), .B(n22321), .Z(n22365) );
  XOR U22079 ( .A(n22366), .B(n22358), .Z(n22321) );
  XNOR U22080 ( .A(n22367), .B(n22353), .Z(n22358) );
  XOR U22081 ( .A(n22368), .B(n22369), .Z(n22353) );
  AND U22082 ( .A(n22370), .B(n22371), .Z(n22369) );
  XOR U22083 ( .A(n22372), .B(n22368), .Z(n22370) );
  XNOR U22084 ( .A(n22373), .B(n22374), .Z(n22367) );
  AND U22085 ( .A(n22375), .B(n22376), .Z(n22374) );
  XOR U22086 ( .A(n22373), .B(n22377), .Z(n22375) );
  XNOR U22087 ( .A(n22359), .B(n22356), .Z(n22366) );
  AND U22088 ( .A(n22378), .B(n22379), .Z(n22356) );
  XOR U22089 ( .A(n22380), .B(n22381), .Z(n22359) );
  AND U22090 ( .A(n22382), .B(n22383), .Z(n22381) );
  XOR U22091 ( .A(n22380), .B(n22384), .Z(n22382) );
  XNOR U22092 ( .A(n22318), .B(n22362), .Z(n22364) );
  XNOR U22093 ( .A(n22385), .B(n22386), .Z(n22318) );
  AND U22094 ( .A(n424), .B(n22324), .Z(n22386) );
  XOR U22095 ( .A(n22385), .B(n22322), .Z(n22324) );
  XOR U22096 ( .A(n22387), .B(n22388), .Z(n22362) );
  AND U22097 ( .A(n22389), .B(n22390), .Z(n22388) );
  XNOR U22098 ( .A(n22387), .B(n22378), .Z(n22390) );
  IV U22099 ( .A(n22332), .Z(n22378) );
  XNOR U22100 ( .A(n22391), .B(n22371), .Z(n22332) );
  XNOR U22101 ( .A(n22392), .B(n22377), .Z(n22371) );
  XOR U22102 ( .A(n22393), .B(n22394), .Z(n22377) );
  NOR U22103 ( .A(n22395), .B(n22396), .Z(n22394) );
  XNOR U22104 ( .A(n22393), .B(n22397), .Z(n22395) );
  XNOR U22105 ( .A(n22376), .B(n22368), .Z(n22392) );
  XOR U22106 ( .A(n22398), .B(n22399), .Z(n22368) );
  AND U22107 ( .A(n22400), .B(n22401), .Z(n22399) );
  XNOR U22108 ( .A(n22398), .B(n22402), .Z(n22400) );
  XNOR U22109 ( .A(n22403), .B(n22373), .Z(n22376) );
  XOR U22110 ( .A(n22404), .B(n22405), .Z(n22373) );
  AND U22111 ( .A(n22406), .B(n22407), .Z(n22405) );
  XOR U22112 ( .A(n22404), .B(n22408), .Z(n22406) );
  XNOR U22113 ( .A(n22409), .B(n22410), .Z(n22403) );
  NOR U22114 ( .A(n22411), .B(n22412), .Z(n22410) );
  XOR U22115 ( .A(n22409), .B(n22413), .Z(n22411) );
  XNOR U22116 ( .A(n22372), .B(n22379), .Z(n22391) );
  NOR U22117 ( .A(n22340), .B(n22414), .Z(n22379) );
  XOR U22118 ( .A(n22384), .B(n22383), .Z(n22372) );
  XNOR U22119 ( .A(n22415), .B(n22380), .Z(n22383) );
  XOR U22120 ( .A(n22416), .B(n22417), .Z(n22380) );
  AND U22121 ( .A(n22418), .B(n22419), .Z(n22417) );
  XOR U22122 ( .A(n22416), .B(n22420), .Z(n22418) );
  XNOR U22123 ( .A(n22421), .B(n22422), .Z(n22415) );
  NOR U22124 ( .A(n22423), .B(n22424), .Z(n22422) );
  XNOR U22125 ( .A(n22421), .B(n22425), .Z(n22423) );
  XOR U22126 ( .A(n22426), .B(n22427), .Z(n22384) );
  NOR U22127 ( .A(n22428), .B(n22429), .Z(n22427) );
  XNOR U22128 ( .A(n22426), .B(n22430), .Z(n22428) );
  XNOR U22129 ( .A(n22329), .B(n22387), .Z(n22389) );
  XNOR U22130 ( .A(n22431), .B(n22432), .Z(n22329) );
  AND U22131 ( .A(n424), .B(n22336), .Z(n22432) );
  XOR U22132 ( .A(n22431), .B(n22334), .Z(n22336) );
  AND U22133 ( .A(n22337), .B(n22340), .Z(n22387) );
  XOR U22134 ( .A(n22433), .B(n22414), .Z(n22340) );
  XNOR U22135 ( .A(p_input[2048]), .B(p_input[560]), .Z(n22414) );
  XOR U22136 ( .A(n22402), .B(n22401), .Z(n22433) );
  XNOR U22137 ( .A(n22434), .B(n22408), .Z(n22401) );
  XNOR U22138 ( .A(n22397), .B(n22396), .Z(n22408) );
  XOR U22139 ( .A(n22435), .B(n22393), .Z(n22396) );
  XNOR U22140 ( .A(n16904), .B(p_input[570]), .Z(n22393) );
  XNOR U22141 ( .A(p_input[2059]), .B(p_input[571]), .Z(n22435) );
  XOR U22142 ( .A(p_input[2060]), .B(p_input[572]), .Z(n22397) );
  XNOR U22143 ( .A(n22407), .B(n22398), .Z(n22434) );
  XNOR U22144 ( .A(n17068), .B(p_input[561]), .Z(n22398) );
  XOR U22145 ( .A(n22436), .B(n22413), .Z(n22407) );
  XNOR U22146 ( .A(p_input[2063]), .B(p_input[575]), .Z(n22413) );
  XOR U22147 ( .A(n22404), .B(n22412), .Z(n22436) );
  XOR U22148 ( .A(n22437), .B(n22409), .Z(n22412) );
  XOR U22149 ( .A(p_input[2061]), .B(p_input[573]), .Z(n22409) );
  XNOR U22150 ( .A(p_input[2062]), .B(p_input[574]), .Z(n22437) );
  XNOR U22151 ( .A(n16738), .B(p_input[569]), .Z(n22404) );
  XNOR U22152 ( .A(n22420), .B(n22419), .Z(n22402) );
  XNOR U22153 ( .A(n22438), .B(n22425), .Z(n22419) );
  XOR U22154 ( .A(p_input[2056]), .B(p_input[568]), .Z(n22425) );
  XOR U22155 ( .A(n22416), .B(n22424), .Z(n22438) );
  XOR U22156 ( .A(n22439), .B(n22421), .Z(n22424) );
  XOR U22157 ( .A(p_input[2054]), .B(p_input[566]), .Z(n22421) );
  XNOR U22158 ( .A(p_input[2055]), .B(p_input[567]), .Z(n22439) );
  XNOR U22159 ( .A(n16741), .B(p_input[562]), .Z(n22416) );
  XNOR U22160 ( .A(n22430), .B(n22429), .Z(n22420) );
  XOR U22161 ( .A(n22440), .B(n22426), .Z(n22429) );
  XOR U22162 ( .A(p_input[2051]), .B(p_input[563]), .Z(n22426) );
  XNOR U22163 ( .A(p_input[2052]), .B(p_input[564]), .Z(n22440) );
  XOR U22164 ( .A(p_input[2053]), .B(p_input[565]), .Z(n22430) );
  XNOR U22165 ( .A(n22441), .B(n22442), .Z(n22337) );
  AND U22166 ( .A(n424), .B(n22443), .Z(n22442) );
  XNOR U22167 ( .A(n22444), .B(n22445), .Z(n424) );
  AND U22168 ( .A(n22446), .B(n22447), .Z(n22445) );
  XOR U22169 ( .A(n22444), .B(n22347), .Z(n22447) );
  XNOR U22170 ( .A(n22444), .B(n22301), .Z(n22446) );
  XOR U22171 ( .A(n22448), .B(n22449), .Z(n22444) );
  AND U22172 ( .A(n22450), .B(n22451), .Z(n22449) );
  XOR U22173 ( .A(n22448), .B(n22311), .Z(n22450) );
  XOR U22174 ( .A(n22452), .B(n22453), .Z(n22290) );
  AND U22175 ( .A(n428), .B(n22443), .Z(n22453) );
  XNOR U22176 ( .A(n22441), .B(n22452), .Z(n22443) );
  XNOR U22177 ( .A(n22454), .B(n22455), .Z(n428) );
  AND U22178 ( .A(n22456), .B(n22457), .Z(n22455) );
  XNOR U22179 ( .A(n22458), .B(n22454), .Z(n22457) );
  IV U22180 ( .A(n22347), .Z(n22458) );
  XNOR U22181 ( .A(n22459), .B(n22460), .Z(n22347) );
  AND U22182 ( .A(n431), .B(n22461), .Z(n22460) );
  XNOR U22183 ( .A(n22459), .B(n22462), .Z(n22461) );
  XNOR U22184 ( .A(n22301), .B(n22454), .Z(n22456) );
  XOR U22185 ( .A(n22463), .B(n22464), .Z(n22301) );
  AND U22186 ( .A(n439), .B(n22465), .Z(n22464) );
  XOR U22187 ( .A(n22448), .B(n22466), .Z(n22454) );
  AND U22188 ( .A(n22467), .B(n22451), .Z(n22466) );
  XNOR U22189 ( .A(n22360), .B(n22448), .Z(n22451) );
  XNOR U22190 ( .A(n22468), .B(n22469), .Z(n22360) );
  AND U22191 ( .A(n431), .B(n22470), .Z(n22469) );
  XOR U22192 ( .A(n22471), .B(n22468), .Z(n22470) );
  XNOR U22193 ( .A(n22472), .B(n22448), .Z(n22467) );
  IV U22194 ( .A(n22311), .Z(n22472) );
  XOR U22195 ( .A(n22473), .B(n22474), .Z(n22311) );
  AND U22196 ( .A(n439), .B(n22475), .Z(n22474) );
  XOR U22197 ( .A(n22476), .B(n22477), .Z(n22448) );
  AND U22198 ( .A(n22478), .B(n22479), .Z(n22477) );
  XNOR U22199 ( .A(n22385), .B(n22476), .Z(n22479) );
  XNOR U22200 ( .A(n22480), .B(n22481), .Z(n22385) );
  AND U22201 ( .A(n431), .B(n22482), .Z(n22481) );
  XNOR U22202 ( .A(n22483), .B(n22480), .Z(n22482) );
  XOR U22203 ( .A(n22476), .B(n22322), .Z(n22478) );
  XOR U22204 ( .A(n22484), .B(n22485), .Z(n22322) );
  AND U22205 ( .A(n439), .B(n22486), .Z(n22485) );
  XOR U22206 ( .A(n22487), .B(n22488), .Z(n22476) );
  AND U22207 ( .A(n22489), .B(n22490), .Z(n22488) );
  XNOR U22208 ( .A(n22487), .B(n22431), .Z(n22490) );
  XNOR U22209 ( .A(n22491), .B(n22492), .Z(n22431) );
  AND U22210 ( .A(n431), .B(n22493), .Z(n22492) );
  XOR U22211 ( .A(n22494), .B(n22491), .Z(n22493) );
  XNOR U22212 ( .A(n22495), .B(n22487), .Z(n22489) );
  IV U22213 ( .A(n22334), .Z(n22495) );
  XOR U22214 ( .A(n22496), .B(n22497), .Z(n22334) );
  AND U22215 ( .A(n439), .B(n22498), .Z(n22497) );
  AND U22216 ( .A(n22452), .B(n22441), .Z(n22487) );
  XNOR U22217 ( .A(n22499), .B(n22500), .Z(n22441) );
  AND U22218 ( .A(n431), .B(n22501), .Z(n22500) );
  XNOR U22219 ( .A(n22502), .B(n22499), .Z(n22501) );
  XNOR U22220 ( .A(n22503), .B(n22504), .Z(n431) );
  AND U22221 ( .A(n22505), .B(n22506), .Z(n22504) );
  XOR U22222 ( .A(n22462), .B(n22503), .Z(n22506) );
  AND U22223 ( .A(n22507), .B(n22508), .Z(n22462) );
  XOR U22224 ( .A(n22503), .B(n22459), .Z(n22505) );
  XNOR U22225 ( .A(n22509), .B(n22510), .Z(n22459) );
  AND U22226 ( .A(n435), .B(n22465), .Z(n22510) );
  XOR U22227 ( .A(n22463), .B(n22509), .Z(n22465) );
  XOR U22228 ( .A(n22511), .B(n22512), .Z(n22503) );
  AND U22229 ( .A(n22513), .B(n22514), .Z(n22512) );
  XNOR U22230 ( .A(n22511), .B(n22507), .Z(n22514) );
  IV U22231 ( .A(n22471), .Z(n22507) );
  XOR U22232 ( .A(n22515), .B(n22516), .Z(n22471) );
  XOR U22233 ( .A(n22517), .B(n22508), .Z(n22516) );
  AND U22234 ( .A(n22483), .B(n22518), .Z(n22508) );
  AND U22235 ( .A(n22519), .B(n22520), .Z(n22517) );
  XOR U22236 ( .A(n22521), .B(n22515), .Z(n22519) );
  XNOR U22237 ( .A(n22468), .B(n22511), .Z(n22513) );
  XNOR U22238 ( .A(n22522), .B(n22523), .Z(n22468) );
  AND U22239 ( .A(n435), .B(n22475), .Z(n22523) );
  XOR U22240 ( .A(n22522), .B(n22473), .Z(n22475) );
  XOR U22241 ( .A(n22524), .B(n22525), .Z(n22511) );
  AND U22242 ( .A(n22526), .B(n22527), .Z(n22525) );
  XNOR U22243 ( .A(n22524), .B(n22483), .Z(n22527) );
  XOR U22244 ( .A(n22528), .B(n22520), .Z(n22483) );
  XNOR U22245 ( .A(n22529), .B(n22515), .Z(n22520) );
  XOR U22246 ( .A(n22530), .B(n22531), .Z(n22515) );
  AND U22247 ( .A(n22532), .B(n22533), .Z(n22531) );
  XOR U22248 ( .A(n22534), .B(n22530), .Z(n22532) );
  XNOR U22249 ( .A(n22535), .B(n22536), .Z(n22529) );
  AND U22250 ( .A(n22537), .B(n22538), .Z(n22536) );
  XOR U22251 ( .A(n22535), .B(n22539), .Z(n22537) );
  XNOR U22252 ( .A(n22521), .B(n22518), .Z(n22528) );
  AND U22253 ( .A(n22540), .B(n22541), .Z(n22518) );
  XOR U22254 ( .A(n22542), .B(n22543), .Z(n22521) );
  AND U22255 ( .A(n22544), .B(n22545), .Z(n22543) );
  XOR U22256 ( .A(n22542), .B(n22546), .Z(n22544) );
  XNOR U22257 ( .A(n22480), .B(n22524), .Z(n22526) );
  XNOR U22258 ( .A(n22547), .B(n22548), .Z(n22480) );
  AND U22259 ( .A(n435), .B(n22486), .Z(n22548) );
  XOR U22260 ( .A(n22547), .B(n22484), .Z(n22486) );
  XOR U22261 ( .A(n22549), .B(n22550), .Z(n22524) );
  AND U22262 ( .A(n22551), .B(n22552), .Z(n22550) );
  XNOR U22263 ( .A(n22549), .B(n22540), .Z(n22552) );
  IV U22264 ( .A(n22494), .Z(n22540) );
  XNOR U22265 ( .A(n22553), .B(n22533), .Z(n22494) );
  XNOR U22266 ( .A(n22554), .B(n22539), .Z(n22533) );
  XOR U22267 ( .A(n22555), .B(n22556), .Z(n22539) );
  NOR U22268 ( .A(n22557), .B(n22558), .Z(n22556) );
  XNOR U22269 ( .A(n22555), .B(n22559), .Z(n22557) );
  XNOR U22270 ( .A(n22538), .B(n22530), .Z(n22554) );
  XOR U22271 ( .A(n22560), .B(n22561), .Z(n22530) );
  AND U22272 ( .A(n22562), .B(n22563), .Z(n22561) );
  XNOR U22273 ( .A(n22560), .B(n22564), .Z(n22562) );
  XNOR U22274 ( .A(n22565), .B(n22535), .Z(n22538) );
  XOR U22275 ( .A(n22566), .B(n22567), .Z(n22535) );
  AND U22276 ( .A(n22568), .B(n22569), .Z(n22567) );
  XOR U22277 ( .A(n22566), .B(n22570), .Z(n22568) );
  XNOR U22278 ( .A(n22571), .B(n22572), .Z(n22565) );
  NOR U22279 ( .A(n22573), .B(n22574), .Z(n22572) );
  XOR U22280 ( .A(n22571), .B(n22575), .Z(n22573) );
  XNOR U22281 ( .A(n22534), .B(n22541), .Z(n22553) );
  NOR U22282 ( .A(n22502), .B(n22576), .Z(n22541) );
  XOR U22283 ( .A(n22546), .B(n22545), .Z(n22534) );
  XNOR U22284 ( .A(n22577), .B(n22542), .Z(n22545) );
  XOR U22285 ( .A(n22578), .B(n22579), .Z(n22542) );
  AND U22286 ( .A(n22580), .B(n22581), .Z(n22579) );
  XOR U22287 ( .A(n22578), .B(n22582), .Z(n22580) );
  XNOR U22288 ( .A(n22583), .B(n22584), .Z(n22577) );
  NOR U22289 ( .A(n22585), .B(n22586), .Z(n22584) );
  XNOR U22290 ( .A(n22583), .B(n22587), .Z(n22585) );
  XOR U22291 ( .A(n22588), .B(n22589), .Z(n22546) );
  NOR U22292 ( .A(n22590), .B(n22591), .Z(n22589) );
  XNOR U22293 ( .A(n22588), .B(n22592), .Z(n22590) );
  XNOR U22294 ( .A(n22491), .B(n22549), .Z(n22551) );
  XNOR U22295 ( .A(n22593), .B(n22594), .Z(n22491) );
  AND U22296 ( .A(n435), .B(n22498), .Z(n22594) );
  XOR U22297 ( .A(n22593), .B(n22496), .Z(n22498) );
  AND U22298 ( .A(n22499), .B(n22502), .Z(n22549) );
  XOR U22299 ( .A(n22595), .B(n22576), .Z(n22502) );
  XNOR U22300 ( .A(p_input[2048]), .B(p_input[576]), .Z(n22576) );
  XOR U22301 ( .A(n22564), .B(n22563), .Z(n22595) );
  XNOR U22302 ( .A(n22596), .B(n22570), .Z(n22563) );
  XNOR U22303 ( .A(n22559), .B(n22558), .Z(n22570) );
  XOR U22304 ( .A(n22597), .B(n22555), .Z(n22558) );
  XNOR U22305 ( .A(n16904), .B(p_input[586]), .Z(n22555) );
  XNOR U22306 ( .A(p_input[2059]), .B(p_input[587]), .Z(n22597) );
  XOR U22307 ( .A(p_input[2060]), .B(p_input[588]), .Z(n22559) );
  XNOR U22308 ( .A(n22569), .B(n22560), .Z(n22596) );
  XNOR U22309 ( .A(n17068), .B(p_input[577]), .Z(n22560) );
  XOR U22310 ( .A(n22598), .B(n22575), .Z(n22569) );
  XNOR U22311 ( .A(p_input[2063]), .B(p_input[591]), .Z(n22575) );
  XOR U22312 ( .A(n22566), .B(n22574), .Z(n22598) );
  XOR U22313 ( .A(n22599), .B(n22571), .Z(n22574) );
  XOR U22314 ( .A(p_input[2061]), .B(p_input[589]), .Z(n22571) );
  XNOR U22315 ( .A(p_input[2062]), .B(p_input[590]), .Z(n22599) );
  XNOR U22316 ( .A(n16738), .B(p_input[585]), .Z(n22566) );
  XNOR U22317 ( .A(n22582), .B(n22581), .Z(n22564) );
  XNOR U22318 ( .A(n22600), .B(n22587), .Z(n22581) );
  XOR U22319 ( .A(p_input[2056]), .B(p_input[584]), .Z(n22587) );
  XOR U22320 ( .A(n22578), .B(n22586), .Z(n22600) );
  XOR U22321 ( .A(n22601), .B(n22583), .Z(n22586) );
  XOR U22322 ( .A(p_input[2054]), .B(p_input[582]), .Z(n22583) );
  XNOR U22323 ( .A(p_input[2055]), .B(p_input[583]), .Z(n22601) );
  XNOR U22324 ( .A(n16741), .B(p_input[578]), .Z(n22578) );
  XNOR U22325 ( .A(n22592), .B(n22591), .Z(n22582) );
  XOR U22326 ( .A(n22602), .B(n22588), .Z(n22591) );
  XOR U22327 ( .A(p_input[2051]), .B(p_input[579]), .Z(n22588) );
  XNOR U22328 ( .A(p_input[2052]), .B(p_input[580]), .Z(n22602) );
  XOR U22329 ( .A(p_input[2053]), .B(p_input[581]), .Z(n22592) );
  XNOR U22330 ( .A(n22603), .B(n22604), .Z(n22499) );
  AND U22331 ( .A(n435), .B(n22605), .Z(n22604) );
  XNOR U22332 ( .A(n22606), .B(n22607), .Z(n435) );
  AND U22333 ( .A(n22608), .B(n22609), .Z(n22607) );
  XOR U22334 ( .A(n22606), .B(n22509), .Z(n22609) );
  XNOR U22335 ( .A(n22606), .B(n22463), .Z(n22608) );
  XOR U22336 ( .A(n22610), .B(n22611), .Z(n22606) );
  AND U22337 ( .A(n22612), .B(n22613), .Z(n22611) );
  XOR U22338 ( .A(n22610), .B(n22473), .Z(n22612) );
  XOR U22339 ( .A(n22614), .B(n22615), .Z(n22452) );
  AND U22340 ( .A(n439), .B(n22605), .Z(n22615) );
  XNOR U22341 ( .A(n22603), .B(n22614), .Z(n22605) );
  XNOR U22342 ( .A(n22616), .B(n22617), .Z(n439) );
  AND U22343 ( .A(n22618), .B(n22619), .Z(n22617) );
  XNOR U22344 ( .A(n22620), .B(n22616), .Z(n22619) );
  IV U22345 ( .A(n22509), .Z(n22620) );
  XNOR U22346 ( .A(n22621), .B(n22622), .Z(n22509) );
  AND U22347 ( .A(n442), .B(n22623), .Z(n22622) );
  XNOR U22348 ( .A(n22621), .B(n22624), .Z(n22623) );
  XNOR U22349 ( .A(n22463), .B(n22616), .Z(n22618) );
  XOR U22350 ( .A(n22625), .B(n22626), .Z(n22463) );
  AND U22351 ( .A(n450), .B(n22627), .Z(n22626) );
  XOR U22352 ( .A(n22610), .B(n22628), .Z(n22616) );
  AND U22353 ( .A(n22629), .B(n22613), .Z(n22628) );
  XNOR U22354 ( .A(n22522), .B(n22610), .Z(n22613) );
  XNOR U22355 ( .A(n22630), .B(n22631), .Z(n22522) );
  AND U22356 ( .A(n442), .B(n22632), .Z(n22631) );
  XOR U22357 ( .A(n22633), .B(n22630), .Z(n22632) );
  XNOR U22358 ( .A(n22634), .B(n22610), .Z(n22629) );
  IV U22359 ( .A(n22473), .Z(n22634) );
  XOR U22360 ( .A(n22635), .B(n22636), .Z(n22473) );
  AND U22361 ( .A(n450), .B(n22637), .Z(n22636) );
  XOR U22362 ( .A(n22638), .B(n22639), .Z(n22610) );
  AND U22363 ( .A(n22640), .B(n22641), .Z(n22639) );
  XNOR U22364 ( .A(n22547), .B(n22638), .Z(n22641) );
  XNOR U22365 ( .A(n22642), .B(n22643), .Z(n22547) );
  AND U22366 ( .A(n442), .B(n22644), .Z(n22643) );
  XNOR U22367 ( .A(n22645), .B(n22642), .Z(n22644) );
  XOR U22368 ( .A(n22638), .B(n22484), .Z(n22640) );
  XOR U22369 ( .A(n22646), .B(n22647), .Z(n22484) );
  AND U22370 ( .A(n450), .B(n22648), .Z(n22647) );
  XOR U22371 ( .A(n22649), .B(n22650), .Z(n22638) );
  AND U22372 ( .A(n22651), .B(n22652), .Z(n22650) );
  XNOR U22373 ( .A(n22649), .B(n22593), .Z(n22652) );
  XNOR U22374 ( .A(n22653), .B(n22654), .Z(n22593) );
  AND U22375 ( .A(n442), .B(n22655), .Z(n22654) );
  XOR U22376 ( .A(n22656), .B(n22653), .Z(n22655) );
  XNOR U22377 ( .A(n22657), .B(n22649), .Z(n22651) );
  IV U22378 ( .A(n22496), .Z(n22657) );
  XOR U22379 ( .A(n22658), .B(n22659), .Z(n22496) );
  AND U22380 ( .A(n450), .B(n22660), .Z(n22659) );
  AND U22381 ( .A(n22614), .B(n22603), .Z(n22649) );
  XNOR U22382 ( .A(n22661), .B(n22662), .Z(n22603) );
  AND U22383 ( .A(n442), .B(n22663), .Z(n22662) );
  XNOR U22384 ( .A(n22664), .B(n22661), .Z(n22663) );
  XNOR U22385 ( .A(n22665), .B(n22666), .Z(n442) );
  AND U22386 ( .A(n22667), .B(n22668), .Z(n22666) );
  XOR U22387 ( .A(n22624), .B(n22665), .Z(n22668) );
  AND U22388 ( .A(n22669), .B(n22670), .Z(n22624) );
  XOR U22389 ( .A(n22665), .B(n22621), .Z(n22667) );
  XNOR U22390 ( .A(n22671), .B(n22672), .Z(n22621) );
  AND U22391 ( .A(n446), .B(n22627), .Z(n22672) );
  XOR U22392 ( .A(n22625), .B(n22671), .Z(n22627) );
  XOR U22393 ( .A(n22673), .B(n22674), .Z(n22665) );
  AND U22394 ( .A(n22675), .B(n22676), .Z(n22674) );
  XNOR U22395 ( .A(n22673), .B(n22669), .Z(n22676) );
  IV U22396 ( .A(n22633), .Z(n22669) );
  XOR U22397 ( .A(n22677), .B(n22678), .Z(n22633) );
  XOR U22398 ( .A(n22679), .B(n22670), .Z(n22678) );
  AND U22399 ( .A(n22645), .B(n22680), .Z(n22670) );
  AND U22400 ( .A(n22681), .B(n22682), .Z(n22679) );
  XOR U22401 ( .A(n22683), .B(n22677), .Z(n22681) );
  XNOR U22402 ( .A(n22630), .B(n22673), .Z(n22675) );
  XNOR U22403 ( .A(n22684), .B(n22685), .Z(n22630) );
  AND U22404 ( .A(n446), .B(n22637), .Z(n22685) );
  XOR U22405 ( .A(n22684), .B(n22635), .Z(n22637) );
  XOR U22406 ( .A(n22686), .B(n22687), .Z(n22673) );
  AND U22407 ( .A(n22688), .B(n22689), .Z(n22687) );
  XNOR U22408 ( .A(n22686), .B(n22645), .Z(n22689) );
  XOR U22409 ( .A(n22690), .B(n22682), .Z(n22645) );
  XNOR U22410 ( .A(n22691), .B(n22677), .Z(n22682) );
  XOR U22411 ( .A(n22692), .B(n22693), .Z(n22677) );
  AND U22412 ( .A(n22694), .B(n22695), .Z(n22693) );
  XOR U22413 ( .A(n22696), .B(n22692), .Z(n22694) );
  XNOR U22414 ( .A(n22697), .B(n22698), .Z(n22691) );
  AND U22415 ( .A(n22699), .B(n22700), .Z(n22698) );
  XOR U22416 ( .A(n22697), .B(n22701), .Z(n22699) );
  XNOR U22417 ( .A(n22683), .B(n22680), .Z(n22690) );
  AND U22418 ( .A(n22702), .B(n22703), .Z(n22680) );
  XOR U22419 ( .A(n22704), .B(n22705), .Z(n22683) );
  AND U22420 ( .A(n22706), .B(n22707), .Z(n22705) );
  XOR U22421 ( .A(n22704), .B(n22708), .Z(n22706) );
  XNOR U22422 ( .A(n22642), .B(n22686), .Z(n22688) );
  XNOR U22423 ( .A(n22709), .B(n22710), .Z(n22642) );
  AND U22424 ( .A(n446), .B(n22648), .Z(n22710) );
  XOR U22425 ( .A(n22709), .B(n22646), .Z(n22648) );
  XOR U22426 ( .A(n22711), .B(n22712), .Z(n22686) );
  AND U22427 ( .A(n22713), .B(n22714), .Z(n22712) );
  XNOR U22428 ( .A(n22711), .B(n22702), .Z(n22714) );
  IV U22429 ( .A(n22656), .Z(n22702) );
  XNOR U22430 ( .A(n22715), .B(n22695), .Z(n22656) );
  XNOR U22431 ( .A(n22716), .B(n22701), .Z(n22695) );
  XOR U22432 ( .A(n22717), .B(n22718), .Z(n22701) );
  NOR U22433 ( .A(n22719), .B(n22720), .Z(n22718) );
  XNOR U22434 ( .A(n22717), .B(n22721), .Z(n22719) );
  XNOR U22435 ( .A(n22700), .B(n22692), .Z(n22716) );
  XOR U22436 ( .A(n22722), .B(n22723), .Z(n22692) );
  AND U22437 ( .A(n22724), .B(n22725), .Z(n22723) );
  XNOR U22438 ( .A(n22722), .B(n22726), .Z(n22724) );
  XNOR U22439 ( .A(n22727), .B(n22697), .Z(n22700) );
  XOR U22440 ( .A(n22728), .B(n22729), .Z(n22697) );
  AND U22441 ( .A(n22730), .B(n22731), .Z(n22729) );
  XOR U22442 ( .A(n22728), .B(n22732), .Z(n22730) );
  XNOR U22443 ( .A(n22733), .B(n22734), .Z(n22727) );
  NOR U22444 ( .A(n22735), .B(n22736), .Z(n22734) );
  XOR U22445 ( .A(n22733), .B(n22737), .Z(n22735) );
  XNOR U22446 ( .A(n22696), .B(n22703), .Z(n22715) );
  NOR U22447 ( .A(n22664), .B(n22738), .Z(n22703) );
  XOR U22448 ( .A(n22708), .B(n22707), .Z(n22696) );
  XNOR U22449 ( .A(n22739), .B(n22704), .Z(n22707) );
  XOR U22450 ( .A(n22740), .B(n22741), .Z(n22704) );
  AND U22451 ( .A(n22742), .B(n22743), .Z(n22741) );
  XOR U22452 ( .A(n22740), .B(n22744), .Z(n22742) );
  XNOR U22453 ( .A(n22745), .B(n22746), .Z(n22739) );
  NOR U22454 ( .A(n22747), .B(n22748), .Z(n22746) );
  XNOR U22455 ( .A(n22745), .B(n22749), .Z(n22747) );
  XOR U22456 ( .A(n22750), .B(n22751), .Z(n22708) );
  NOR U22457 ( .A(n22752), .B(n22753), .Z(n22751) );
  XNOR U22458 ( .A(n22750), .B(n22754), .Z(n22752) );
  XNOR U22459 ( .A(n22653), .B(n22711), .Z(n22713) );
  XNOR U22460 ( .A(n22755), .B(n22756), .Z(n22653) );
  AND U22461 ( .A(n446), .B(n22660), .Z(n22756) );
  XOR U22462 ( .A(n22755), .B(n22658), .Z(n22660) );
  AND U22463 ( .A(n22661), .B(n22664), .Z(n22711) );
  XOR U22464 ( .A(n22757), .B(n22738), .Z(n22664) );
  XNOR U22465 ( .A(p_input[2048]), .B(p_input[592]), .Z(n22738) );
  XOR U22466 ( .A(n22726), .B(n22725), .Z(n22757) );
  XNOR U22467 ( .A(n22758), .B(n22732), .Z(n22725) );
  XNOR U22468 ( .A(n22721), .B(n22720), .Z(n22732) );
  XOR U22469 ( .A(n22759), .B(n22717), .Z(n22720) );
  XNOR U22470 ( .A(n16904), .B(p_input[602]), .Z(n22717) );
  XNOR U22471 ( .A(p_input[2059]), .B(p_input[603]), .Z(n22759) );
  XOR U22472 ( .A(p_input[2060]), .B(p_input[604]), .Z(n22721) );
  XNOR U22473 ( .A(n22731), .B(n22722), .Z(n22758) );
  XNOR U22474 ( .A(n17068), .B(p_input[593]), .Z(n22722) );
  XOR U22475 ( .A(n22760), .B(n22737), .Z(n22731) );
  XNOR U22476 ( .A(p_input[2063]), .B(p_input[607]), .Z(n22737) );
  XOR U22477 ( .A(n22728), .B(n22736), .Z(n22760) );
  XOR U22478 ( .A(n22761), .B(n22733), .Z(n22736) );
  XOR U22479 ( .A(p_input[2061]), .B(p_input[605]), .Z(n22733) );
  XNOR U22480 ( .A(p_input[2062]), .B(p_input[606]), .Z(n22761) );
  XNOR U22481 ( .A(n16738), .B(p_input[601]), .Z(n22728) );
  XNOR U22482 ( .A(n22744), .B(n22743), .Z(n22726) );
  XNOR U22483 ( .A(n22762), .B(n22749), .Z(n22743) );
  XOR U22484 ( .A(p_input[2056]), .B(p_input[600]), .Z(n22749) );
  XOR U22485 ( .A(n22740), .B(n22748), .Z(n22762) );
  XOR U22486 ( .A(n22763), .B(n22745), .Z(n22748) );
  XOR U22487 ( .A(p_input[2054]), .B(p_input[598]), .Z(n22745) );
  XNOR U22488 ( .A(p_input[2055]), .B(p_input[599]), .Z(n22763) );
  XNOR U22489 ( .A(n16741), .B(p_input[594]), .Z(n22740) );
  XNOR U22490 ( .A(n22754), .B(n22753), .Z(n22744) );
  XOR U22491 ( .A(n22764), .B(n22750), .Z(n22753) );
  XOR U22492 ( .A(p_input[2051]), .B(p_input[595]), .Z(n22750) );
  XNOR U22493 ( .A(p_input[2052]), .B(p_input[596]), .Z(n22764) );
  XOR U22494 ( .A(p_input[2053]), .B(p_input[597]), .Z(n22754) );
  XNOR U22495 ( .A(n22765), .B(n22766), .Z(n22661) );
  AND U22496 ( .A(n446), .B(n22767), .Z(n22766) );
  XNOR U22497 ( .A(n22768), .B(n22769), .Z(n446) );
  AND U22498 ( .A(n22770), .B(n22771), .Z(n22769) );
  XOR U22499 ( .A(n22768), .B(n22671), .Z(n22771) );
  XNOR U22500 ( .A(n22768), .B(n22625), .Z(n22770) );
  XOR U22501 ( .A(n22772), .B(n22773), .Z(n22768) );
  AND U22502 ( .A(n22774), .B(n22775), .Z(n22773) );
  XOR U22503 ( .A(n22772), .B(n22635), .Z(n22774) );
  XOR U22504 ( .A(n22776), .B(n22777), .Z(n22614) );
  AND U22505 ( .A(n450), .B(n22767), .Z(n22777) );
  XNOR U22506 ( .A(n22765), .B(n22776), .Z(n22767) );
  XNOR U22507 ( .A(n22778), .B(n22779), .Z(n450) );
  AND U22508 ( .A(n22780), .B(n22781), .Z(n22779) );
  XNOR U22509 ( .A(n22782), .B(n22778), .Z(n22781) );
  IV U22510 ( .A(n22671), .Z(n22782) );
  XNOR U22511 ( .A(n22783), .B(n22784), .Z(n22671) );
  AND U22512 ( .A(n453), .B(n22785), .Z(n22784) );
  XNOR U22513 ( .A(n22783), .B(n22786), .Z(n22785) );
  XNOR U22514 ( .A(n22625), .B(n22778), .Z(n22780) );
  XOR U22515 ( .A(n22787), .B(n22788), .Z(n22625) );
  AND U22516 ( .A(n461), .B(n22789), .Z(n22788) );
  XOR U22517 ( .A(n22772), .B(n22790), .Z(n22778) );
  AND U22518 ( .A(n22791), .B(n22775), .Z(n22790) );
  XNOR U22519 ( .A(n22684), .B(n22772), .Z(n22775) );
  XNOR U22520 ( .A(n22792), .B(n22793), .Z(n22684) );
  AND U22521 ( .A(n453), .B(n22794), .Z(n22793) );
  XOR U22522 ( .A(n22795), .B(n22792), .Z(n22794) );
  XNOR U22523 ( .A(n22796), .B(n22772), .Z(n22791) );
  IV U22524 ( .A(n22635), .Z(n22796) );
  XOR U22525 ( .A(n22797), .B(n22798), .Z(n22635) );
  AND U22526 ( .A(n461), .B(n22799), .Z(n22798) );
  XOR U22527 ( .A(n22800), .B(n22801), .Z(n22772) );
  AND U22528 ( .A(n22802), .B(n22803), .Z(n22801) );
  XNOR U22529 ( .A(n22709), .B(n22800), .Z(n22803) );
  XNOR U22530 ( .A(n22804), .B(n22805), .Z(n22709) );
  AND U22531 ( .A(n453), .B(n22806), .Z(n22805) );
  XNOR U22532 ( .A(n22807), .B(n22804), .Z(n22806) );
  XOR U22533 ( .A(n22800), .B(n22646), .Z(n22802) );
  XOR U22534 ( .A(n22808), .B(n22809), .Z(n22646) );
  AND U22535 ( .A(n461), .B(n22810), .Z(n22809) );
  XOR U22536 ( .A(n22811), .B(n22812), .Z(n22800) );
  AND U22537 ( .A(n22813), .B(n22814), .Z(n22812) );
  XNOR U22538 ( .A(n22811), .B(n22755), .Z(n22814) );
  XNOR U22539 ( .A(n22815), .B(n22816), .Z(n22755) );
  AND U22540 ( .A(n453), .B(n22817), .Z(n22816) );
  XOR U22541 ( .A(n22818), .B(n22815), .Z(n22817) );
  XNOR U22542 ( .A(n22819), .B(n22811), .Z(n22813) );
  IV U22543 ( .A(n22658), .Z(n22819) );
  XOR U22544 ( .A(n22820), .B(n22821), .Z(n22658) );
  AND U22545 ( .A(n461), .B(n22822), .Z(n22821) );
  AND U22546 ( .A(n22776), .B(n22765), .Z(n22811) );
  XNOR U22547 ( .A(n22823), .B(n22824), .Z(n22765) );
  AND U22548 ( .A(n453), .B(n22825), .Z(n22824) );
  XNOR U22549 ( .A(n22826), .B(n22823), .Z(n22825) );
  XNOR U22550 ( .A(n22827), .B(n22828), .Z(n453) );
  AND U22551 ( .A(n22829), .B(n22830), .Z(n22828) );
  XOR U22552 ( .A(n22786), .B(n22827), .Z(n22830) );
  AND U22553 ( .A(n22831), .B(n22832), .Z(n22786) );
  XOR U22554 ( .A(n22827), .B(n22783), .Z(n22829) );
  XNOR U22555 ( .A(n22833), .B(n22834), .Z(n22783) );
  AND U22556 ( .A(n457), .B(n22789), .Z(n22834) );
  XOR U22557 ( .A(n22787), .B(n22833), .Z(n22789) );
  XOR U22558 ( .A(n22835), .B(n22836), .Z(n22827) );
  AND U22559 ( .A(n22837), .B(n22838), .Z(n22836) );
  XNOR U22560 ( .A(n22835), .B(n22831), .Z(n22838) );
  IV U22561 ( .A(n22795), .Z(n22831) );
  XOR U22562 ( .A(n22839), .B(n22840), .Z(n22795) );
  XOR U22563 ( .A(n22841), .B(n22832), .Z(n22840) );
  AND U22564 ( .A(n22807), .B(n22842), .Z(n22832) );
  AND U22565 ( .A(n22843), .B(n22844), .Z(n22841) );
  XOR U22566 ( .A(n22845), .B(n22839), .Z(n22843) );
  XNOR U22567 ( .A(n22792), .B(n22835), .Z(n22837) );
  XNOR U22568 ( .A(n22846), .B(n22847), .Z(n22792) );
  AND U22569 ( .A(n457), .B(n22799), .Z(n22847) );
  XOR U22570 ( .A(n22846), .B(n22797), .Z(n22799) );
  XOR U22571 ( .A(n22848), .B(n22849), .Z(n22835) );
  AND U22572 ( .A(n22850), .B(n22851), .Z(n22849) );
  XNOR U22573 ( .A(n22848), .B(n22807), .Z(n22851) );
  XOR U22574 ( .A(n22852), .B(n22844), .Z(n22807) );
  XNOR U22575 ( .A(n22853), .B(n22839), .Z(n22844) );
  XOR U22576 ( .A(n22854), .B(n22855), .Z(n22839) );
  AND U22577 ( .A(n22856), .B(n22857), .Z(n22855) );
  XOR U22578 ( .A(n22858), .B(n22854), .Z(n22856) );
  XNOR U22579 ( .A(n22859), .B(n22860), .Z(n22853) );
  AND U22580 ( .A(n22861), .B(n22862), .Z(n22860) );
  XOR U22581 ( .A(n22859), .B(n22863), .Z(n22861) );
  XNOR U22582 ( .A(n22845), .B(n22842), .Z(n22852) );
  AND U22583 ( .A(n22864), .B(n22865), .Z(n22842) );
  XOR U22584 ( .A(n22866), .B(n22867), .Z(n22845) );
  AND U22585 ( .A(n22868), .B(n22869), .Z(n22867) );
  XOR U22586 ( .A(n22866), .B(n22870), .Z(n22868) );
  XNOR U22587 ( .A(n22804), .B(n22848), .Z(n22850) );
  XNOR U22588 ( .A(n22871), .B(n22872), .Z(n22804) );
  AND U22589 ( .A(n457), .B(n22810), .Z(n22872) );
  XOR U22590 ( .A(n22871), .B(n22808), .Z(n22810) );
  XOR U22591 ( .A(n22873), .B(n22874), .Z(n22848) );
  AND U22592 ( .A(n22875), .B(n22876), .Z(n22874) );
  XNOR U22593 ( .A(n22873), .B(n22864), .Z(n22876) );
  IV U22594 ( .A(n22818), .Z(n22864) );
  XNOR U22595 ( .A(n22877), .B(n22857), .Z(n22818) );
  XNOR U22596 ( .A(n22878), .B(n22863), .Z(n22857) );
  XOR U22597 ( .A(n22879), .B(n22880), .Z(n22863) );
  NOR U22598 ( .A(n22881), .B(n22882), .Z(n22880) );
  XNOR U22599 ( .A(n22879), .B(n22883), .Z(n22881) );
  XNOR U22600 ( .A(n22862), .B(n22854), .Z(n22878) );
  XOR U22601 ( .A(n22884), .B(n22885), .Z(n22854) );
  AND U22602 ( .A(n22886), .B(n22887), .Z(n22885) );
  XNOR U22603 ( .A(n22884), .B(n22888), .Z(n22886) );
  XNOR U22604 ( .A(n22889), .B(n22859), .Z(n22862) );
  XOR U22605 ( .A(n22890), .B(n22891), .Z(n22859) );
  AND U22606 ( .A(n22892), .B(n22893), .Z(n22891) );
  XOR U22607 ( .A(n22890), .B(n22894), .Z(n22892) );
  XNOR U22608 ( .A(n22895), .B(n22896), .Z(n22889) );
  NOR U22609 ( .A(n22897), .B(n22898), .Z(n22896) );
  XOR U22610 ( .A(n22895), .B(n22899), .Z(n22897) );
  XNOR U22611 ( .A(n22858), .B(n22865), .Z(n22877) );
  NOR U22612 ( .A(n22826), .B(n22900), .Z(n22865) );
  XOR U22613 ( .A(n22870), .B(n22869), .Z(n22858) );
  XNOR U22614 ( .A(n22901), .B(n22866), .Z(n22869) );
  XOR U22615 ( .A(n22902), .B(n22903), .Z(n22866) );
  AND U22616 ( .A(n22904), .B(n22905), .Z(n22903) );
  XOR U22617 ( .A(n22902), .B(n22906), .Z(n22904) );
  XNOR U22618 ( .A(n22907), .B(n22908), .Z(n22901) );
  NOR U22619 ( .A(n22909), .B(n22910), .Z(n22908) );
  XNOR U22620 ( .A(n22907), .B(n22911), .Z(n22909) );
  XOR U22621 ( .A(n22912), .B(n22913), .Z(n22870) );
  NOR U22622 ( .A(n22914), .B(n22915), .Z(n22913) );
  XNOR U22623 ( .A(n22912), .B(n22916), .Z(n22914) );
  XNOR U22624 ( .A(n22815), .B(n22873), .Z(n22875) );
  XNOR U22625 ( .A(n22917), .B(n22918), .Z(n22815) );
  AND U22626 ( .A(n457), .B(n22822), .Z(n22918) );
  XOR U22627 ( .A(n22917), .B(n22820), .Z(n22822) );
  AND U22628 ( .A(n22823), .B(n22826), .Z(n22873) );
  XOR U22629 ( .A(n22919), .B(n22900), .Z(n22826) );
  XNOR U22630 ( .A(p_input[2048]), .B(p_input[608]), .Z(n22900) );
  XOR U22631 ( .A(n22888), .B(n22887), .Z(n22919) );
  XNOR U22632 ( .A(n22920), .B(n22894), .Z(n22887) );
  XNOR U22633 ( .A(n22883), .B(n22882), .Z(n22894) );
  XOR U22634 ( .A(n22921), .B(n22879), .Z(n22882) );
  XNOR U22635 ( .A(n16904), .B(p_input[618]), .Z(n22879) );
  XNOR U22636 ( .A(p_input[2059]), .B(p_input[619]), .Z(n22921) );
  XOR U22637 ( .A(p_input[2060]), .B(p_input[620]), .Z(n22883) );
  XNOR U22638 ( .A(n22893), .B(n22884), .Z(n22920) );
  XNOR U22639 ( .A(n17068), .B(p_input[609]), .Z(n22884) );
  XOR U22640 ( .A(n22922), .B(n22899), .Z(n22893) );
  XNOR U22641 ( .A(p_input[2063]), .B(p_input[623]), .Z(n22899) );
  XOR U22642 ( .A(n22890), .B(n22898), .Z(n22922) );
  XOR U22643 ( .A(n22923), .B(n22895), .Z(n22898) );
  XOR U22644 ( .A(p_input[2061]), .B(p_input[621]), .Z(n22895) );
  XNOR U22645 ( .A(p_input[2062]), .B(p_input[622]), .Z(n22923) );
  XNOR U22646 ( .A(n16738), .B(p_input[617]), .Z(n22890) );
  XNOR U22647 ( .A(n22906), .B(n22905), .Z(n22888) );
  XNOR U22648 ( .A(n22924), .B(n22911), .Z(n22905) );
  XOR U22649 ( .A(p_input[2056]), .B(p_input[616]), .Z(n22911) );
  XOR U22650 ( .A(n22902), .B(n22910), .Z(n22924) );
  XOR U22651 ( .A(n22925), .B(n22907), .Z(n22910) );
  XOR U22652 ( .A(p_input[2054]), .B(p_input[614]), .Z(n22907) );
  XNOR U22653 ( .A(p_input[2055]), .B(p_input[615]), .Z(n22925) );
  XNOR U22654 ( .A(n16741), .B(p_input[610]), .Z(n22902) );
  XNOR U22655 ( .A(n22916), .B(n22915), .Z(n22906) );
  XOR U22656 ( .A(n22926), .B(n22912), .Z(n22915) );
  XOR U22657 ( .A(p_input[2051]), .B(p_input[611]), .Z(n22912) );
  XNOR U22658 ( .A(p_input[2052]), .B(p_input[612]), .Z(n22926) );
  XOR U22659 ( .A(p_input[2053]), .B(p_input[613]), .Z(n22916) );
  XNOR U22660 ( .A(n22927), .B(n22928), .Z(n22823) );
  AND U22661 ( .A(n457), .B(n22929), .Z(n22928) );
  XNOR U22662 ( .A(n22930), .B(n22931), .Z(n457) );
  AND U22663 ( .A(n22932), .B(n22933), .Z(n22931) );
  XOR U22664 ( .A(n22930), .B(n22833), .Z(n22933) );
  XNOR U22665 ( .A(n22930), .B(n22787), .Z(n22932) );
  XOR U22666 ( .A(n22934), .B(n22935), .Z(n22930) );
  AND U22667 ( .A(n22936), .B(n22937), .Z(n22935) );
  XOR U22668 ( .A(n22934), .B(n22797), .Z(n22936) );
  XOR U22669 ( .A(n22938), .B(n22939), .Z(n22776) );
  AND U22670 ( .A(n461), .B(n22929), .Z(n22939) );
  XNOR U22671 ( .A(n22927), .B(n22938), .Z(n22929) );
  XNOR U22672 ( .A(n22940), .B(n22941), .Z(n461) );
  AND U22673 ( .A(n22942), .B(n22943), .Z(n22941) );
  XNOR U22674 ( .A(n22944), .B(n22940), .Z(n22943) );
  IV U22675 ( .A(n22833), .Z(n22944) );
  XNOR U22676 ( .A(n22945), .B(n22946), .Z(n22833) );
  AND U22677 ( .A(n464), .B(n22947), .Z(n22946) );
  XNOR U22678 ( .A(n22945), .B(n22948), .Z(n22947) );
  XNOR U22679 ( .A(n22787), .B(n22940), .Z(n22942) );
  XOR U22680 ( .A(n22949), .B(n22950), .Z(n22787) );
  AND U22681 ( .A(n472), .B(n22951), .Z(n22950) );
  XOR U22682 ( .A(n22934), .B(n22952), .Z(n22940) );
  AND U22683 ( .A(n22953), .B(n22937), .Z(n22952) );
  XNOR U22684 ( .A(n22846), .B(n22934), .Z(n22937) );
  XNOR U22685 ( .A(n22954), .B(n22955), .Z(n22846) );
  AND U22686 ( .A(n464), .B(n22956), .Z(n22955) );
  XOR U22687 ( .A(n22957), .B(n22954), .Z(n22956) );
  XNOR U22688 ( .A(n22958), .B(n22934), .Z(n22953) );
  IV U22689 ( .A(n22797), .Z(n22958) );
  XOR U22690 ( .A(n22959), .B(n22960), .Z(n22797) );
  AND U22691 ( .A(n472), .B(n22961), .Z(n22960) );
  XOR U22692 ( .A(n22962), .B(n22963), .Z(n22934) );
  AND U22693 ( .A(n22964), .B(n22965), .Z(n22963) );
  XNOR U22694 ( .A(n22871), .B(n22962), .Z(n22965) );
  XNOR U22695 ( .A(n22966), .B(n22967), .Z(n22871) );
  AND U22696 ( .A(n464), .B(n22968), .Z(n22967) );
  XNOR U22697 ( .A(n22969), .B(n22966), .Z(n22968) );
  XOR U22698 ( .A(n22962), .B(n22808), .Z(n22964) );
  XOR U22699 ( .A(n22970), .B(n22971), .Z(n22808) );
  AND U22700 ( .A(n472), .B(n22972), .Z(n22971) );
  XOR U22701 ( .A(n22973), .B(n22974), .Z(n22962) );
  AND U22702 ( .A(n22975), .B(n22976), .Z(n22974) );
  XNOR U22703 ( .A(n22973), .B(n22917), .Z(n22976) );
  XNOR U22704 ( .A(n22977), .B(n22978), .Z(n22917) );
  AND U22705 ( .A(n464), .B(n22979), .Z(n22978) );
  XOR U22706 ( .A(n22980), .B(n22977), .Z(n22979) );
  XNOR U22707 ( .A(n22981), .B(n22973), .Z(n22975) );
  IV U22708 ( .A(n22820), .Z(n22981) );
  XOR U22709 ( .A(n22982), .B(n22983), .Z(n22820) );
  AND U22710 ( .A(n472), .B(n22984), .Z(n22983) );
  AND U22711 ( .A(n22938), .B(n22927), .Z(n22973) );
  XNOR U22712 ( .A(n22985), .B(n22986), .Z(n22927) );
  AND U22713 ( .A(n464), .B(n22987), .Z(n22986) );
  XNOR U22714 ( .A(n22988), .B(n22985), .Z(n22987) );
  XNOR U22715 ( .A(n22989), .B(n22990), .Z(n464) );
  AND U22716 ( .A(n22991), .B(n22992), .Z(n22990) );
  XOR U22717 ( .A(n22948), .B(n22989), .Z(n22992) );
  AND U22718 ( .A(n22993), .B(n22994), .Z(n22948) );
  XOR U22719 ( .A(n22989), .B(n22945), .Z(n22991) );
  XNOR U22720 ( .A(n22995), .B(n22996), .Z(n22945) );
  AND U22721 ( .A(n468), .B(n22951), .Z(n22996) );
  XOR U22722 ( .A(n22949), .B(n22995), .Z(n22951) );
  XOR U22723 ( .A(n22997), .B(n22998), .Z(n22989) );
  AND U22724 ( .A(n22999), .B(n23000), .Z(n22998) );
  XNOR U22725 ( .A(n22997), .B(n22993), .Z(n23000) );
  IV U22726 ( .A(n22957), .Z(n22993) );
  XOR U22727 ( .A(n23001), .B(n23002), .Z(n22957) );
  XOR U22728 ( .A(n23003), .B(n22994), .Z(n23002) );
  AND U22729 ( .A(n22969), .B(n23004), .Z(n22994) );
  AND U22730 ( .A(n23005), .B(n23006), .Z(n23003) );
  XOR U22731 ( .A(n23007), .B(n23001), .Z(n23005) );
  XNOR U22732 ( .A(n22954), .B(n22997), .Z(n22999) );
  XNOR U22733 ( .A(n23008), .B(n23009), .Z(n22954) );
  AND U22734 ( .A(n468), .B(n22961), .Z(n23009) );
  XOR U22735 ( .A(n23008), .B(n22959), .Z(n22961) );
  XOR U22736 ( .A(n23010), .B(n23011), .Z(n22997) );
  AND U22737 ( .A(n23012), .B(n23013), .Z(n23011) );
  XNOR U22738 ( .A(n23010), .B(n22969), .Z(n23013) );
  XOR U22739 ( .A(n23014), .B(n23006), .Z(n22969) );
  XNOR U22740 ( .A(n23015), .B(n23001), .Z(n23006) );
  XOR U22741 ( .A(n23016), .B(n23017), .Z(n23001) );
  AND U22742 ( .A(n23018), .B(n23019), .Z(n23017) );
  XOR U22743 ( .A(n23020), .B(n23016), .Z(n23018) );
  XNOR U22744 ( .A(n23021), .B(n23022), .Z(n23015) );
  AND U22745 ( .A(n23023), .B(n23024), .Z(n23022) );
  XOR U22746 ( .A(n23021), .B(n23025), .Z(n23023) );
  XNOR U22747 ( .A(n23007), .B(n23004), .Z(n23014) );
  AND U22748 ( .A(n23026), .B(n23027), .Z(n23004) );
  XOR U22749 ( .A(n23028), .B(n23029), .Z(n23007) );
  AND U22750 ( .A(n23030), .B(n23031), .Z(n23029) );
  XOR U22751 ( .A(n23028), .B(n23032), .Z(n23030) );
  XNOR U22752 ( .A(n22966), .B(n23010), .Z(n23012) );
  XNOR U22753 ( .A(n23033), .B(n23034), .Z(n22966) );
  AND U22754 ( .A(n468), .B(n22972), .Z(n23034) );
  XOR U22755 ( .A(n23033), .B(n22970), .Z(n22972) );
  XOR U22756 ( .A(n23035), .B(n23036), .Z(n23010) );
  AND U22757 ( .A(n23037), .B(n23038), .Z(n23036) );
  XNOR U22758 ( .A(n23035), .B(n23026), .Z(n23038) );
  IV U22759 ( .A(n22980), .Z(n23026) );
  XNOR U22760 ( .A(n23039), .B(n23019), .Z(n22980) );
  XNOR U22761 ( .A(n23040), .B(n23025), .Z(n23019) );
  XOR U22762 ( .A(n23041), .B(n23042), .Z(n23025) );
  NOR U22763 ( .A(n23043), .B(n23044), .Z(n23042) );
  XNOR U22764 ( .A(n23041), .B(n23045), .Z(n23043) );
  XNOR U22765 ( .A(n23024), .B(n23016), .Z(n23040) );
  XOR U22766 ( .A(n23046), .B(n23047), .Z(n23016) );
  AND U22767 ( .A(n23048), .B(n23049), .Z(n23047) );
  XNOR U22768 ( .A(n23046), .B(n23050), .Z(n23048) );
  XNOR U22769 ( .A(n23051), .B(n23021), .Z(n23024) );
  XOR U22770 ( .A(n23052), .B(n23053), .Z(n23021) );
  AND U22771 ( .A(n23054), .B(n23055), .Z(n23053) );
  XOR U22772 ( .A(n23052), .B(n23056), .Z(n23054) );
  XNOR U22773 ( .A(n23057), .B(n23058), .Z(n23051) );
  NOR U22774 ( .A(n23059), .B(n23060), .Z(n23058) );
  XOR U22775 ( .A(n23057), .B(n23061), .Z(n23059) );
  XNOR U22776 ( .A(n23020), .B(n23027), .Z(n23039) );
  NOR U22777 ( .A(n22988), .B(n23062), .Z(n23027) );
  XOR U22778 ( .A(n23032), .B(n23031), .Z(n23020) );
  XNOR U22779 ( .A(n23063), .B(n23028), .Z(n23031) );
  XOR U22780 ( .A(n23064), .B(n23065), .Z(n23028) );
  AND U22781 ( .A(n23066), .B(n23067), .Z(n23065) );
  XOR U22782 ( .A(n23064), .B(n23068), .Z(n23066) );
  XNOR U22783 ( .A(n23069), .B(n23070), .Z(n23063) );
  NOR U22784 ( .A(n23071), .B(n23072), .Z(n23070) );
  XNOR U22785 ( .A(n23069), .B(n23073), .Z(n23071) );
  XOR U22786 ( .A(n23074), .B(n23075), .Z(n23032) );
  NOR U22787 ( .A(n23076), .B(n23077), .Z(n23075) );
  XNOR U22788 ( .A(n23074), .B(n23078), .Z(n23076) );
  XNOR U22789 ( .A(n22977), .B(n23035), .Z(n23037) );
  XNOR U22790 ( .A(n23079), .B(n23080), .Z(n22977) );
  AND U22791 ( .A(n468), .B(n22984), .Z(n23080) );
  XOR U22792 ( .A(n23079), .B(n22982), .Z(n22984) );
  AND U22793 ( .A(n22985), .B(n22988), .Z(n23035) );
  XOR U22794 ( .A(n23081), .B(n23062), .Z(n22988) );
  XNOR U22795 ( .A(p_input[2048]), .B(p_input[624]), .Z(n23062) );
  XOR U22796 ( .A(n23050), .B(n23049), .Z(n23081) );
  XNOR U22797 ( .A(n23082), .B(n23056), .Z(n23049) );
  XNOR U22798 ( .A(n23045), .B(n23044), .Z(n23056) );
  XOR U22799 ( .A(n23083), .B(n23041), .Z(n23044) );
  XNOR U22800 ( .A(n16904), .B(p_input[634]), .Z(n23041) );
  XNOR U22801 ( .A(p_input[2059]), .B(p_input[635]), .Z(n23083) );
  XOR U22802 ( .A(p_input[2060]), .B(p_input[636]), .Z(n23045) );
  XNOR U22803 ( .A(n23055), .B(n23046), .Z(n23082) );
  XNOR U22804 ( .A(n17068), .B(p_input[625]), .Z(n23046) );
  XOR U22805 ( .A(n23084), .B(n23061), .Z(n23055) );
  XNOR U22806 ( .A(p_input[2063]), .B(p_input[639]), .Z(n23061) );
  XOR U22807 ( .A(n23052), .B(n23060), .Z(n23084) );
  XOR U22808 ( .A(n23085), .B(n23057), .Z(n23060) );
  XOR U22809 ( .A(p_input[2061]), .B(p_input[637]), .Z(n23057) );
  XNOR U22810 ( .A(p_input[2062]), .B(p_input[638]), .Z(n23085) );
  XNOR U22811 ( .A(n16738), .B(p_input[633]), .Z(n23052) );
  XNOR U22812 ( .A(n23068), .B(n23067), .Z(n23050) );
  XNOR U22813 ( .A(n23086), .B(n23073), .Z(n23067) );
  XOR U22814 ( .A(p_input[2056]), .B(p_input[632]), .Z(n23073) );
  XOR U22815 ( .A(n23064), .B(n23072), .Z(n23086) );
  XOR U22816 ( .A(n23087), .B(n23069), .Z(n23072) );
  XOR U22817 ( .A(p_input[2054]), .B(p_input[630]), .Z(n23069) );
  XNOR U22818 ( .A(p_input[2055]), .B(p_input[631]), .Z(n23087) );
  XNOR U22819 ( .A(n16741), .B(p_input[626]), .Z(n23064) );
  XNOR U22820 ( .A(n23078), .B(n23077), .Z(n23068) );
  XOR U22821 ( .A(n23088), .B(n23074), .Z(n23077) );
  XOR U22822 ( .A(p_input[2051]), .B(p_input[627]), .Z(n23074) );
  XNOR U22823 ( .A(p_input[2052]), .B(p_input[628]), .Z(n23088) );
  XOR U22824 ( .A(p_input[2053]), .B(p_input[629]), .Z(n23078) );
  XNOR U22825 ( .A(n23089), .B(n23090), .Z(n22985) );
  AND U22826 ( .A(n468), .B(n23091), .Z(n23090) );
  XNOR U22827 ( .A(n23092), .B(n23093), .Z(n468) );
  AND U22828 ( .A(n23094), .B(n23095), .Z(n23093) );
  XOR U22829 ( .A(n23092), .B(n22995), .Z(n23095) );
  XNOR U22830 ( .A(n23092), .B(n22949), .Z(n23094) );
  XOR U22831 ( .A(n23096), .B(n23097), .Z(n23092) );
  AND U22832 ( .A(n23098), .B(n23099), .Z(n23097) );
  XOR U22833 ( .A(n23096), .B(n22959), .Z(n23098) );
  XOR U22834 ( .A(n23100), .B(n23101), .Z(n22938) );
  AND U22835 ( .A(n472), .B(n23091), .Z(n23101) );
  XNOR U22836 ( .A(n23089), .B(n23100), .Z(n23091) );
  XNOR U22837 ( .A(n23102), .B(n23103), .Z(n472) );
  AND U22838 ( .A(n23104), .B(n23105), .Z(n23103) );
  XNOR U22839 ( .A(n23106), .B(n23102), .Z(n23105) );
  IV U22840 ( .A(n22995), .Z(n23106) );
  XNOR U22841 ( .A(n23107), .B(n23108), .Z(n22995) );
  AND U22842 ( .A(n475), .B(n23109), .Z(n23108) );
  XNOR U22843 ( .A(n23107), .B(n23110), .Z(n23109) );
  XNOR U22844 ( .A(n22949), .B(n23102), .Z(n23104) );
  XOR U22845 ( .A(n23111), .B(n23112), .Z(n22949) );
  AND U22846 ( .A(n483), .B(n23113), .Z(n23112) );
  XOR U22847 ( .A(n23096), .B(n23114), .Z(n23102) );
  AND U22848 ( .A(n23115), .B(n23099), .Z(n23114) );
  XNOR U22849 ( .A(n23008), .B(n23096), .Z(n23099) );
  XNOR U22850 ( .A(n23116), .B(n23117), .Z(n23008) );
  AND U22851 ( .A(n475), .B(n23118), .Z(n23117) );
  XOR U22852 ( .A(n23119), .B(n23116), .Z(n23118) );
  XNOR U22853 ( .A(n23120), .B(n23096), .Z(n23115) );
  IV U22854 ( .A(n22959), .Z(n23120) );
  XOR U22855 ( .A(n23121), .B(n23122), .Z(n22959) );
  AND U22856 ( .A(n483), .B(n23123), .Z(n23122) );
  XOR U22857 ( .A(n23124), .B(n23125), .Z(n23096) );
  AND U22858 ( .A(n23126), .B(n23127), .Z(n23125) );
  XNOR U22859 ( .A(n23033), .B(n23124), .Z(n23127) );
  XNOR U22860 ( .A(n23128), .B(n23129), .Z(n23033) );
  AND U22861 ( .A(n475), .B(n23130), .Z(n23129) );
  XNOR U22862 ( .A(n23131), .B(n23128), .Z(n23130) );
  XOR U22863 ( .A(n23124), .B(n22970), .Z(n23126) );
  XOR U22864 ( .A(n23132), .B(n23133), .Z(n22970) );
  AND U22865 ( .A(n483), .B(n23134), .Z(n23133) );
  XOR U22866 ( .A(n23135), .B(n23136), .Z(n23124) );
  AND U22867 ( .A(n23137), .B(n23138), .Z(n23136) );
  XNOR U22868 ( .A(n23135), .B(n23079), .Z(n23138) );
  XNOR U22869 ( .A(n23139), .B(n23140), .Z(n23079) );
  AND U22870 ( .A(n475), .B(n23141), .Z(n23140) );
  XOR U22871 ( .A(n23142), .B(n23139), .Z(n23141) );
  XNOR U22872 ( .A(n23143), .B(n23135), .Z(n23137) );
  IV U22873 ( .A(n22982), .Z(n23143) );
  XOR U22874 ( .A(n23144), .B(n23145), .Z(n22982) );
  AND U22875 ( .A(n483), .B(n23146), .Z(n23145) );
  AND U22876 ( .A(n23100), .B(n23089), .Z(n23135) );
  XNOR U22877 ( .A(n23147), .B(n23148), .Z(n23089) );
  AND U22878 ( .A(n475), .B(n23149), .Z(n23148) );
  XNOR U22879 ( .A(n23150), .B(n23147), .Z(n23149) );
  XNOR U22880 ( .A(n23151), .B(n23152), .Z(n475) );
  AND U22881 ( .A(n23153), .B(n23154), .Z(n23152) );
  XOR U22882 ( .A(n23110), .B(n23151), .Z(n23154) );
  AND U22883 ( .A(n23155), .B(n23156), .Z(n23110) );
  XOR U22884 ( .A(n23151), .B(n23107), .Z(n23153) );
  XNOR U22885 ( .A(n23157), .B(n23158), .Z(n23107) );
  AND U22886 ( .A(n479), .B(n23113), .Z(n23158) );
  XOR U22887 ( .A(n23111), .B(n23157), .Z(n23113) );
  XOR U22888 ( .A(n23159), .B(n23160), .Z(n23151) );
  AND U22889 ( .A(n23161), .B(n23162), .Z(n23160) );
  XNOR U22890 ( .A(n23159), .B(n23155), .Z(n23162) );
  IV U22891 ( .A(n23119), .Z(n23155) );
  XOR U22892 ( .A(n23163), .B(n23164), .Z(n23119) );
  XOR U22893 ( .A(n23165), .B(n23156), .Z(n23164) );
  AND U22894 ( .A(n23131), .B(n23166), .Z(n23156) );
  AND U22895 ( .A(n23167), .B(n23168), .Z(n23165) );
  XOR U22896 ( .A(n23169), .B(n23163), .Z(n23167) );
  XNOR U22897 ( .A(n23116), .B(n23159), .Z(n23161) );
  XNOR U22898 ( .A(n23170), .B(n23171), .Z(n23116) );
  AND U22899 ( .A(n479), .B(n23123), .Z(n23171) );
  XOR U22900 ( .A(n23170), .B(n23121), .Z(n23123) );
  XOR U22901 ( .A(n23172), .B(n23173), .Z(n23159) );
  AND U22902 ( .A(n23174), .B(n23175), .Z(n23173) );
  XNOR U22903 ( .A(n23172), .B(n23131), .Z(n23175) );
  XOR U22904 ( .A(n23176), .B(n23168), .Z(n23131) );
  XNOR U22905 ( .A(n23177), .B(n23163), .Z(n23168) );
  XOR U22906 ( .A(n23178), .B(n23179), .Z(n23163) );
  AND U22907 ( .A(n23180), .B(n23181), .Z(n23179) );
  XOR U22908 ( .A(n23182), .B(n23178), .Z(n23180) );
  XNOR U22909 ( .A(n23183), .B(n23184), .Z(n23177) );
  AND U22910 ( .A(n23185), .B(n23186), .Z(n23184) );
  XOR U22911 ( .A(n23183), .B(n23187), .Z(n23185) );
  XNOR U22912 ( .A(n23169), .B(n23166), .Z(n23176) );
  AND U22913 ( .A(n23188), .B(n23189), .Z(n23166) );
  XOR U22914 ( .A(n23190), .B(n23191), .Z(n23169) );
  AND U22915 ( .A(n23192), .B(n23193), .Z(n23191) );
  XOR U22916 ( .A(n23190), .B(n23194), .Z(n23192) );
  XNOR U22917 ( .A(n23128), .B(n23172), .Z(n23174) );
  XNOR U22918 ( .A(n23195), .B(n23196), .Z(n23128) );
  AND U22919 ( .A(n479), .B(n23134), .Z(n23196) );
  XOR U22920 ( .A(n23195), .B(n23132), .Z(n23134) );
  XOR U22921 ( .A(n23197), .B(n23198), .Z(n23172) );
  AND U22922 ( .A(n23199), .B(n23200), .Z(n23198) );
  XNOR U22923 ( .A(n23197), .B(n23188), .Z(n23200) );
  IV U22924 ( .A(n23142), .Z(n23188) );
  XNOR U22925 ( .A(n23201), .B(n23181), .Z(n23142) );
  XNOR U22926 ( .A(n23202), .B(n23187), .Z(n23181) );
  XOR U22927 ( .A(n23203), .B(n23204), .Z(n23187) );
  NOR U22928 ( .A(n23205), .B(n23206), .Z(n23204) );
  XNOR U22929 ( .A(n23203), .B(n23207), .Z(n23205) );
  XNOR U22930 ( .A(n23186), .B(n23178), .Z(n23202) );
  XOR U22931 ( .A(n23208), .B(n23209), .Z(n23178) );
  AND U22932 ( .A(n23210), .B(n23211), .Z(n23209) );
  XNOR U22933 ( .A(n23208), .B(n23212), .Z(n23210) );
  XNOR U22934 ( .A(n23213), .B(n23183), .Z(n23186) );
  XOR U22935 ( .A(n23214), .B(n23215), .Z(n23183) );
  AND U22936 ( .A(n23216), .B(n23217), .Z(n23215) );
  XOR U22937 ( .A(n23214), .B(n23218), .Z(n23216) );
  XNOR U22938 ( .A(n23219), .B(n23220), .Z(n23213) );
  NOR U22939 ( .A(n23221), .B(n23222), .Z(n23220) );
  XOR U22940 ( .A(n23219), .B(n23223), .Z(n23221) );
  XNOR U22941 ( .A(n23182), .B(n23189), .Z(n23201) );
  NOR U22942 ( .A(n23150), .B(n23224), .Z(n23189) );
  XOR U22943 ( .A(n23194), .B(n23193), .Z(n23182) );
  XNOR U22944 ( .A(n23225), .B(n23190), .Z(n23193) );
  XOR U22945 ( .A(n23226), .B(n23227), .Z(n23190) );
  AND U22946 ( .A(n23228), .B(n23229), .Z(n23227) );
  XOR U22947 ( .A(n23226), .B(n23230), .Z(n23228) );
  XNOR U22948 ( .A(n23231), .B(n23232), .Z(n23225) );
  NOR U22949 ( .A(n23233), .B(n23234), .Z(n23232) );
  XNOR U22950 ( .A(n23231), .B(n23235), .Z(n23233) );
  XOR U22951 ( .A(n23236), .B(n23237), .Z(n23194) );
  NOR U22952 ( .A(n23238), .B(n23239), .Z(n23237) );
  XNOR U22953 ( .A(n23236), .B(n23240), .Z(n23238) );
  XNOR U22954 ( .A(n23139), .B(n23197), .Z(n23199) );
  XNOR U22955 ( .A(n23241), .B(n23242), .Z(n23139) );
  AND U22956 ( .A(n479), .B(n23146), .Z(n23242) );
  XOR U22957 ( .A(n23241), .B(n23144), .Z(n23146) );
  AND U22958 ( .A(n23147), .B(n23150), .Z(n23197) );
  XOR U22959 ( .A(n23243), .B(n23224), .Z(n23150) );
  XNOR U22960 ( .A(p_input[2048]), .B(p_input[640]), .Z(n23224) );
  XOR U22961 ( .A(n23212), .B(n23211), .Z(n23243) );
  XNOR U22962 ( .A(n23244), .B(n23218), .Z(n23211) );
  XNOR U22963 ( .A(n23207), .B(n23206), .Z(n23218) );
  XOR U22964 ( .A(n23245), .B(n23203), .Z(n23206) );
  XNOR U22965 ( .A(n16904), .B(p_input[650]), .Z(n23203) );
  XNOR U22966 ( .A(p_input[2059]), .B(p_input[651]), .Z(n23245) );
  XOR U22967 ( .A(p_input[2060]), .B(p_input[652]), .Z(n23207) );
  XNOR U22968 ( .A(n23217), .B(n23208), .Z(n23244) );
  XNOR U22969 ( .A(n17068), .B(p_input[641]), .Z(n23208) );
  XOR U22970 ( .A(n23246), .B(n23223), .Z(n23217) );
  XNOR U22971 ( .A(p_input[2063]), .B(p_input[655]), .Z(n23223) );
  XOR U22972 ( .A(n23214), .B(n23222), .Z(n23246) );
  XOR U22973 ( .A(n23247), .B(n23219), .Z(n23222) );
  XOR U22974 ( .A(p_input[2061]), .B(p_input[653]), .Z(n23219) );
  XNOR U22975 ( .A(p_input[2062]), .B(p_input[654]), .Z(n23247) );
  XNOR U22976 ( .A(n16738), .B(p_input[649]), .Z(n23214) );
  XNOR U22977 ( .A(n23230), .B(n23229), .Z(n23212) );
  XNOR U22978 ( .A(n23248), .B(n23235), .Z(n23229) );
  XOR U22979 ( .A(p_input[2056]), .B(p_input[648]), .Z(n23235) );
  XOR U22980 ( .A(n23226), .B(n23234), .Z(n23248) );
  XOR U22981 ( .A(n23249), .B(n23231), .Z(n23234) );
  XOR U22982 ( .A(p_input[2054]), .B(p_input[646]), .Z(n23231) );
  XNOR U22983 ( .A(p_input[2055]), .B(p_input[647]), .Z(n23249) );
  XNOR U22984 ( .A(n16741), .B(p_input[642]), .Z(n23226) );
  XNOR U22985 ( .A(n23240), .B(n23239), .Z(n23230) );
  XOR U22986 ( .A(n23250), .B(n23236), .Z(n23239) );
  XOR U22987 ( .A(p_input[2051]), .B(p_input[643]), .Z(n23236) );
  XNOR U22988 ( .A(p_input[2052]), .B(p_input[644]), .Z(n23250) );
  XOR U22989 ( .A(p_input[2053]), .B(p_input[645]), .Z(n23240) );
  XNOR U22990 ( .A(n23251), .B(n23252), .Z(n23147) );
  AND U22991 ( .A(n479), .B(n23253), .Z(n23252) );
  XNOR U22992 ( .A(n23254), .B(n23255), .Z(n479) );
  AND U22993 ( .A(n23256), .B(n23257), .Z(n23255) );
  XOR U22994 ( .A(n23254), .B(n23157), .Z(n23257) );
  XNOR U22995 ( .A(n23254), .B(n23111), .Z(n23256) );
  XOR U22996 ( .A(n23258), .B(n23259), .Z(n23254) );
  AND U22997 ( .A(n23260), .B(n23261), .Z(n23259) );
  XOR U22998 ( .A(n23258), .B(n23121), .Z(n23260) );
  XOR U22999 ( .A(n23262), .B(n23263), .Z(n23100) );
  AND U23000 ( .A(n483), .B(n23253), .Z(n23263) );
  XNOR U23001 ( .A(n23251), .B(n23262), .Z(n23253) );
  XNOR U23002 ( .A(n23264), .B(n23265), .Z(n483) );
  AND U23003 ( .A(n23266), .B(n23267), .Z(n23265) );
  XNOR U23004 ( .A(n23268), .B(n23264), .Z(n23267) );
  IV U23005 ( .A(n23157), .Z(n23268) );
  XNOR U23006 ( .A(n23269), .B(n23270), .Z(n23157) );
  AND U23007 ( .A(n486), .B(n23271), .Z(n23270) );
  XNOR U23008 ( .A(n23269), .B(n23272), .Z(n23271) );
  XNOR U23009 ( .A(n23111), .B(n23264), .Z(n23266) );
  XOR U23010 ( .A(n23273), .B(n23274), .Z(n23111) );
  AND U23011 ( .A(n494), .B(n23275), .Z(n23274) );
  XOR U23012 ( .A(n23258), .B(n23276), .Z(n23264) );
  AND U23013 ( .A(n23277), .B(n23261), .Z(n23276) );
  XNOR U23014 ( .A(n23170), .B(n23258), .Z(n23261) );
  XNOR U23015 ( .A(n23278), .B(n23279), .Z(n23170) );
  AND U23016 ( .A(n486), .B(n23280), .Z(n23279) );
  XOR U23017 ( .A(n23281), .B(n23278), .Z(n23280) );
  XNOR U23018 ( .A(n23282), .B(n23258), .Z(n23277) );
  IV U23019 ( .A(n23121), .Z(n23282) );
  XOR U23020 ( .A(n23283), .B(n23284), .Z(n23121) );
  AND U23021 ( .A(n494), .B(n23285), .Z(n23284) );
  XOR U23022 ( .A(n23286), .B(n23287), .Z(n23258) );
  AND U23023 ( .A(n23288), .B(n23289), .Z(n23287) );
  XNOR U23024 ( .A(n23195), .B(n23286), .Z(n23289) );
  XNOR U23025 ( .A(n23290), .B(n23291), .Z(n23195) );
  AND U23026 ( .A(n486), .B(n23292), .Z(n23291) );
  XNOR U23027 ( .A(n23293), .B(n23290), .Z(n23292) );
  XOR U23028 ( .A(n23286), .B(n23132), .Z(n23288) );
  XOR U23029 ( .A(n23294), .B(n23295), .Z(n23132) );
  AND U23030 ( .A(n494), .B(n23296), .Z(n23295) );
  XOR U23031 ( .A(n23297), .B(n23298), .Z(n23286) );
  AND U23032 ( .A(n23299), .B(n23300), .Z(n23298) );
  XNOR U23033 ( .A(n23297), .B(n23241), .Z(n23300) );
  XNOR U23034 ( .A(n23301), .B(n23302), .Z(n23241) );
  AND U23035 ( .A(n486), .B(n23303), .Z(n23302) );
  XOR U23036 ( .A(n23304), .B(n23301), .Z(n23303) );
  XNOR U23037 ( .A(n23305), .B(n23297), .Z(n23299) );
  IV U23038 ( .A(n23144), .Z(n23305) );
  XOR U23039 ( .A(n23306), .B(n23307), .Z(n23144) );
  AND U23040 ( .A(n494), .B(n23308), .Z(n23307) );
  AND U23041 ( .A(n23262), .B(n23251), .Z(n23297) );
  XNOR U23042 ( .A(n23309), .B(n23310), .Z(n23251) );
  AND U23043 ( .A(n486), .B(n23311), .Z(n23310) );
  XNOR U23044 ( .A(n23312), .B(n23309), .Z(n23311) );
  XNOR U23045 ( .A(n23313), .B(n23314), .Z(n486) );
  AND U23046 ( .A(n23315), .B(n23316), .Z(n23314) );
  XOR U23047 ( .A(n23272), .B(n23313), .Z(n23316) );
  AND U23048 ( .A(n23317), .B(n23318), .Z(n23272) );
  XOR U23049 ( .A(n23313), .B(n23269), .Z(n23315) );
  XNOR U23050 ( .A(n23319), .B(n23320), .Z(n23269) );
  AND U23051 ( .A(n490), .B(n23275), .Z(n23320) );
  XOR U23052 ( .A(n23273), .B(n23319), .Z(n23275) );
  XOR U23053 ( .A(n23321), .B(n23322), .Z(n23313) );
  AND U23054 ( .A(n23323), .B(n23324), .Z(n23322) );
  XNOR U23055 ( .A(n23321), .B(n23317), .Z(n23324) );
  IV U23056 ( .A(n23281), .Z(n23317) );
  XOR U23057 ( .A(n23325), .B(n23326), .Z(n23281) );
  XOR U23058 ( .A(n23327), .B(n23318), .Z(n23326) );
  AND U23059 ( .A(n23293), .B(n23328), .Z(n23318) );
  AND U23060 ( .A(n23329), .B(n23330), .Z(n23327) );
  XOR U23061 ( .A(n23331), .B(n23325), .Z(n23329) );
  XNOR U23062 ( .A(n23278), .B(n23321), .Z(n23323) );
  XNOR U23063 ( .A(n23332), .B(n23333), .Z(n23278) );
  AND U23064 ( .A(n490), .B(n23285), .Z(n23333) );
  XOR U23065 ( .A(n23332), .B(n23283), .Z(n23285) );
  XOR U23066 ( .A(n23334), .B(n23335), .Z(n23321) );
  AND U23067 ( .A(n23336), .B(n23337), .Z(n23335) );
  XNOR U23068 ( .A(n23334), .B(n23293), .Z(n23337) );
  XOR U23069 ( .A(n23338), .B(n23330), .Z(n23293) );
  XNOR U23070 ( .A(n23339), .B(n23325), .Z(n23330) );
  XOR U23071 ( .A(n23340), .B(n23341), .Z(n23325) );
  AND U23072 ( .A(n23342), .B(n23343), .Z(n23341) );
  XOR U23073 ( .A(n23344), .B(n23340), .Z(n23342) );
  XNOR U23074 ( .A(n23345), .B(n23346), .Z(n23339) );
  AND U23075 ( .A(n23347), .B(n23348), .Z(n23346) );
  XOR U23076 ( .A(n23345), .B(n23349), .Z(n23347) );
  XNOR U23077 ( .A(n23331), .B(n23328), .Z(n23338) );
  AND U23078 ( .A(n23350), .B(n23351), .Z(n23328) );
  XOR U23079 ( .A(n23352), .B(n23353), .Z(n23331) );
  AND U23080 ( .A(n23354), .B(n23355), .Z(n23353) );
  XOR U23081 ( .A(n23352), .B(n23356), .Z(n23354) );
  XNOR U23082 ( .A(n23290), .B(n23334), .Z(n23336) );
  XNOR U23083 ( .A(n23357), .B(n23358), .Z(n23290) );
  AND U23084 ( .A(n490), .B(n23296), .Z(n23358) );
  XOR U23085 ( .A(n23357), .B(n23294), .Z(n23296) );
  XOR U23086 ( .A(n23359), .B(n23360), .Z(n23334) );
  AND U23087 ( .A(n23361), .B(n23362), .Z(n23360) );
  XNOR U23088 ( .A(n23359), .B(n23350), .Z(n23362) );
  IV U23089 ( .A(n23304), .Z(n23350) );
  XNOR U23090 ( .A(n23363), .B(n23343), .Z(n23304) );
  XNOR U23091 ( .A(n23364), .B(n23349), .Z(n23343) );
  XOR U23092 ( .A(n23365), .B(n23366), .Z(n23349) );
  NOR U23093 ( .A(n23367), .B(n23368), .Z(n23366) );
  XNOR U23094 ( .A(n23365), .B(n23369), .Z(n23367) );
  XNOR U23095 ( .A(n23348), .B(n23340), .Z(n23364) );
  XOR U23096 ( .A(n23370), .B(n23371), .Z(n23340) );
  AND U23097 ( .A(n23372), .B(n23373), .Z(n23371) );
  XNOR U23098 ( .A(n23370), .B(n23374), .Z(n23372) );
  XNOR U23099 ( .A(n23375), .B(n23345), .Z(n23348) );
  XOR U23100 ( .A(n23376), .B(n23377), .Z(n23345) );
  AND U23101 ( .A(n23378), .B(n23379), .Z(n23377) );
  XOR U23102 ( .A(n23376), .B(n23380), .Z(n23378) );
  XNOR U23103 ( .A(n23381), .B(n23382), .Z(n23375) );
  NOR U23104 ( .A(n23383), .B(n23384), .Z(n23382) );
  XOR U23105 ( .A(n23381), .B(n23385), .Z(n23383) );
  XNOR U23106 ( .A(n23344), .B(n23351), .Z(n23363) );
  NOR U23107 ( .A(n23312), .B(n23386), .Z(n23351) );
  XOR U23108 ( .A(n23356), .B(n23355), .Z(n23344) );
  XNOR U23109 ( .A(n23387), .B(n23352), .Z(n23355) );
  XOR U23110 ( .A(n23388), .B(n23389), .Z(n23352) );
  AND U23111 ( .A(n23390), .B(n23391), .Z(n23389) );
  XOR U23112 ( .A(n23388), .B(n23392), .Z(n23390) );
  XNOR U23113 ( .A(n23393), .B(n23394), .Z(n23387) );
  NOR U23114 ( .A(n23395), .B(n23396), .Z(n23394) );
  XNOR U23115 ( .A(n23393), .B(n23397), .Z(n23395) );
  XOR U23116 ( .A(n23398), .B(n23399), .Z(n23356) );
  NOR U23117 ( .A(n23400), .B(n23401), .Z(n23399) );
  XNOR U23118 ( .A(n23398), .B(n23402), .Z(n23400) );
  XNOR U23119 ( .A(n23301), .B(n23359), .Z(n23361) );
  XNOR U23120 ( .A(n23403), .B(n23404), .Z(n23301) );
  AND U23121 ( .A(n490), .B(n23308), .Z(n23404) );
  XOR U23122 ( .A(n23403), .B(n23306), .Z(n23308) );
  AND U23123 ( .A(n23309), .B(n23312), .Z(n23359) );
  XOR U23124 ( .A(n23405), .B(n23386), .Z(n23312) );
  XNOR U23125 ( .A(p_input[2048]), .B(p_input[656]), .Z(n23386) );
  XOR U23126 ( .A(n23374), .B(n23373), .Z(n23405) );
  XNOR U23127 ( .A(n23406), .B(n23380), .Z(n23373) );
  XNOR U23128 ( .A(n23369), .B(n23368), .Z(n23380) );
  XOR U23129 ( .A(n23407), .B(n23365), .Z(n23368) );
  XNOR U23130 ( .A(n16904), .B(p_input[666]), .Z(n23365) );
  XNOR U23131 ( .A(p_input[2059]), .B(p_input[667]), .Z(n23407) );
  XOR U23132 ( .A(p_input[2060]), .B(p_input[668]), .Z(n23369) );
  XNOR U23133 ( .A(n23379), .B(n23370), .Z(n23406) );
  XNOR U23134 ( .A(n17068), .B(p_input[657]), .Z(n23370) );
  XOR U23135 ( .A(n23408), .B(n23385), .Z(n23379) );
  XNOR U23136 ( .A(p_input[2063]), .B(p_input[671]), .Z(n23385) );
  XOR U23137 ( .A(n23376), .B(n23384), .Z(n23408) );
  XOR U23138 ( .A(n23409), .B(n23381), .Z(n23384) );
  XOR U23139 ( .A(p_input[2061]), .B(p_input[669]), .Z(n23381) );
  XNOR U23140 ( .A(p_input[2062]), .B(p_input[670]), .Z(n23409) );
  XNOR U23141 ( .A(n16738), .B(p_input[665]), .Z(n23376) );
  XNOR U23142 ( .A(n23392), .B(n23391), .Z(n23374) );
  XNOR U23143 ( .A(n23410), .B(n23397), .Z(n23391) );
  XOR U23144 ( .A(p_input[2056]), .B(p_input[664]), .Z(n23397) );
  XOR U23145 ( .A(n23388), .B(n23396), .Z(n23410) );
  XOR U23146 ( .A(n23411), .B(n23393), .Z(n23396) );
  XOR U23147 ( .A(p_input[2054]), .B(p_input[662]), .Z(n23393) );
  XNOR U23148 ( .A(p_input[2055]), .B(p_input[663]), .Z(n23411) );
  XNOR U23149 ( .A(n16741), .B(p_input[658]), .Z(n23388) );
  XNOR U23150 ( .A(n23402), .B(n23401), .Z(n23392) );
  XOR U23151 ( .A(n23412), .B(n23398), .Z(n23401) );
  XOR U23152 ( .A(p_input[2051]), .B(p_input[659]), .Z(n23398) );
  XNOR U23153 ( .A(p_input[2052]), .B(p_input[660]), .Z(n23412) );
  XOR U23154 ( .A(p_input[2053]), .B(p_input[661]), .Z(n23402) );
  XNOR U23155 ( .A(n23413), .B(n23414), .Z(n23309) );
  AND U23156 ( .A(n490), .B(n23415), .Z(n23414) );
  XNOR U23157 ( .A(n23416), .B(n23417), .Z(n490) );
  AND U23158 ( .A(n23418), .B(n23419), .Z(n23417) );
  XOR U23159 ( .A(n23416), .B(n23319), .Z(n23419) );
  XNOR U23160 ( .A(n23416), .B(n23273), .Z(n23418) );
  XOR U23161 ( .A(n23420), .B(n23421), .Z(n23416) );
  AND U23162 ( .A(n23422), .B(n23423), .Z(n23421) );
  XOR U23163 ( .A(n23420), .B(n23283), .Z(n23422) );
  XOR U23164 ( .A(n23424), .B(n23425), .Z(n23262) );
  AND U23165 ( .A(n494), .B(n23415), .Z(n23425) );
  XNOR U23166 ( .A(n23413), .B(n23424), .Z(n23415) );
  XNOR U23167 ( .A(n23426), .B(n23427), .Z(n494) );
  AND U23168 ( .A(n23428), .B(n23429), .Z(n23427) );
  XNOR U23169 ( .A(n23430), .B(n23426), .Z(n23429) );
  IV U23170 ( .A(n23319), .Z(n23430) );
  XNOR U23171 ( .A(n23431), .B(n23432), .Z(n23319) );
  AND U23172 ( .A(n497), .B(n23433), .Z(n23432) );
  XNOR U23173 ( .A(n23431), .B(n23434), .Z(n23433) );
  XNOR U23174 ( .A(n23273), .B(n23426), .Z(n23428) );
  XOR U23175 ( .A(n23435), .B(n23436), .Z(n23273) );
  AND U23176 ( .A(n505), .B(n23437), .Z(n23436) );
  XOR U23177 ( .A(n23420), .B(n23438), .Z(n23426) );
  AND U23178 ( .A(n23439), .B(n23423), .Z(n23438) );
  XNOR U23179 ( .A(n23332), .B(n23420), .Z(n23423) );
  XNOR U23180 ( .A(n23440), .B(n23441), .Z(n23332) );
  AND U23181 ( .A(n497), .B(n23442), .Z(n23441) );
  XOR U23182 ( .A(n23443), .B(n23440), .Z(n23442) );
  XNOR U23183 ( .A(n23444), .B(n23420), .Z(n23439) );
  IV U23184 ( .A(n23283), .Z(n23444) );
  XOR U23185 ( .A(n23445), .B(n23446), .Z(n23283) );
  AND U23186 ( .A(n505), .B(n23447), .Z(n23446) );
  XOR U23187 ( .A(n23448), .B(n23449), .Z(n23420) );
  AND U23188 ( .A(n23450), .B(n23451), .Z(n23449) );
  XNOR U23189 ( .A(n23357), .B(n23448), .Z(n23451) );
  XNOR U23190 ( .A(n23452), .B(n23453), .Z(n23357) );
  AND U23191 ( .A(n497), .B(n23454), .Z(n23453) );
  XNOR U23192 ( .A(n23455), .B(n23452), .Z(n23454) );
  XOR U23193 ( .A(n23448), .B(n23294), .Z(n23450) );
  XOR U23194 ( .A(n23456), .B(n23457), .Z(n23294) );
  AND U23195 ( .A(n505), .B(n23458), .Z(n23457) );
  XOR U23196 ( .A(n23459), .B(n23460), .Z(n23448) );
  AND U23197 ( .A(n23461), .B(n23462), .Z(n23460) );
  XNOR U23198 ( .A(n23459), .B(n23403), .Z(n23462) );
  XNOR U23199 ( .A(n23463), .B(n23464), .Z(n23403) );
  AND U23200 ( .A(n497), .B(n23465), .Z(n23464) );
  XOR U23201 ( .A(n23466), .B(n23463), .Z(n23465) );
  XNOR U23202 ( .A(n23467), .B(n23459), .Z(n23461) );
  IV U23203 ( .A(n23306), .Z(n23467) );
  XOR U23204 ( .A(n23468), .B(n23469), .Z(n23306) );
  AND U23205 ( .A(n505), .B(n23470), .Z(n23469) );
  AND U23206 ( .A(n23424), .B(n23413), .Z(n23459) );
  XNOR U23207 ( .A(n23471), .B(n23472), .Z(n23413) );
  AND U23208 ( .A(n497), .B(n23473), .Z(n23472) );
  XNOR U23209 ( .A(n23474), .B(n23471), .Z(n23473) );
  XNOR U23210 ( .A(n23475), .B(n23476), .Z(n497) );
  AND U23211 ( .A(n23477), .B(n23478), .Z(n23476) );
  XOR U23212 ( .A(n23434), .B(n23475), .Z(n23478) );
  AND U23213 ( .A(n23479), .B(n23480), .Z(n23434) );
  XOR U23214 ( .A(n23475), .B(n23431), .Z(n23477) );
  XNOR U23215 ( .A(n23481), .B(n23482), .Z(n23431) );
  AND U23216 ( .A(n501), .B(n23437), .Z(n23482) );
  XOR U23217 ( .A(n23435), .B(n23481), .Z(n23437) );
  XOR U23218 ( .A(n23483), .B(n23484), .Z(n23475) );
  AND U23219 ( .A(n23485), .B(n23486), .Z(n23484) );
  XNOR U23220 ( .A(n23483), .B(n23479), .Z(n23486) );
  IV U23221 ( .A(n23443), .Z(n23479) );
  XOR U23222 ( .A(n23487), .B(n23488), .Z(n23443) );
  XOR U23223 ( .A(n23489), .B(n23480), .Z(n23488) );
  AND U23224 ( .A(n23455), .B(n23490), .Z(n23480) );
  AND U23225 ( .A(n23491), .B(n23492), .Z(n23489) );
  XOR U23226 ( .A(n23493), .B(n23487), .Z(n23491) );
  XNOR U23227 ( .A(n23440), .B(n23483), .Z(n23485) );
  XNOR U23228 ( .A(n23494), .B(n23495), .Z(n23440) );
  AND U23229 ( .A(n501), .B(n23447), .Z(n23495) );
  XOR U23230 ( .A(n23494), .B(n23445), .Z(n23447) );
  XOR U23231 ( .A(n23496), .B(n23497), .Z(n23483) );
  AND U23232 ( .A(n23498), .B(n23499), .Z(n23497) );
  XNOR U23233 ( .A(n23496), .B(n23455), .Z(n23499) );
  XOR U23234 ( .A(n23500), .B(n23492), .Z(n23455) );
  XNOR U23235 ( .A(n23501), .B(n23487), .Z(n23492) );
  XOR U23236 ( .A(n23502), .B(n23503), .Z(n23487) );
  AND U23237 ( .A(n23504), .B(n23505), .Z(n23503) );
  XOR U23238 ( .A(n23506), .B(n23502), .Z(n23504) );
  XNOR U23239 ( .A(n23507), .B(n23508), .Z(n23501) );
  AND U23240 ( .A(n23509), .B(n23510), .Z(n23508) );
  XOR U23241 ( .A(n23507), .B(n23511), .Z(n23509) );
  XNOR U23242 ( .A(n23493), .B(n23490), .Z(n23500) );
  AND U23243 ( .A(n23512), .B(n23513), .Z(n23490) );
  XOR U23244 ( .A(n23514), .B(n23515), .Z(n23493) );
  AND U23245 ( .A(n23516), .B(n23517), .Z(n23515) );
  XOR U23246 ( .A(n23514), .B(n23518), .Z(n23516) );
  XNOR U23247 ( .A(n23452), .B(n23496), .Z(n23498) );
  XNOR U23248 ( .A(n23519), .B(n23520), .Z(n23452) );
  AND U23249 ( .A(n501), .B(n23458), .Z(n23520) );
  XOR U23250 ( .A(n23519), .B(n23456), .Z(n23458) );
  XOR U23251 ( .A(n23521), .B(n23522), .Z(n23496) );
  AND U23252 ( .A(n23523), .B(n23524), .Z(n23522) );
  XNOR U23253 ( .A(n23521), .B(n23512), .Z(n23524) );
  IV U23254 ( .A(n23466), .Z(n23512) );
  XNOR U23255 ( .A(n23525), .B(n23505), .Z(n23466) );
  XNOR U23256 ( .A(n23526), .B(n23511), .Z(n23505) );
  XOR U23257 ( .A(n23527), .B(n23528), .Z(n23511) );
  NOR U23258 ( .A(n23529), .B(n23530), .Z(n23528) );
  XNOR U23259 ( .A(n23527), .B(n23531), .Z(n23529) );
  XNOR U23260 ( .A(n23510), .B(n23502), .Z(n23526) );
  XOR U23261 ( .A(n23532), .B(n23533), .Z(n23502) );
  AND U23262 ( .A(n23534), .B(n23535), .Z(n23533) );
  XNOR U23263 ( .A(n23532), .B(n23536), .Z(n23534) );
  XNOR U23264 ( .A(n23537), .B(n23507), .Z(n23510) );
  XOR U23265 ( .A(n23538), .B(n23539), .Z(n23507) );
  AND U23266 ( .A(n23540), .B(n23541), .Z(n23539) );
  XOR U23267 ( .A(n23538), .B(n23542), .Z(n23540) );
  XNOR U23268 ( .A(n23543), .B(n23544), .Z(n23537) );
  NOR U23269 ( .A(n23545), .B(n23546), .Z(n23544) );
  XOR U23270 ( .A(n23543), .B(n23547), .Z(n23545) );
  XNOR U23271 ( .A(n23506), .B(n23513), .Z(n23525) );
  NOR U23272 ( .A(n23474), .B(n23548), .Z(n23513) );
  XOR U23273 ( .A(n23518), .B(n23517), .Z(n23506) );
  XNOR U23274 ( .A(n23549), .B(n23514), .Z(n23517) );
  XOR U23275 ( .A(n23550), .B(n23551), .Z(n23514) );
  AND U23276 ( .A(n23552), .B(n23553), .Z(n23551) );
  XOR U23277 ( .A(n23550), .B(n23554), .Z(n23552) );
  XNOR U23278 ( .A(n23555), .B(n23556), .Z(n23549) );
  NOR U23279 ( .A(n23557), .B(n23558), .Z(n23556) );
  XNOR U23280 ( .A(n23555), .B(n23559), .Z(n23557) );
  XOR U23281 ( .A(n23560), .B(n23561), .Z(n23518) );
  NOR U23282 ( .A(n23562), .B(n23563), .Z(n23561) );
  XNOR U23283 ( .A(n23560), .B(n23564), .Z(n23562) );
  XNOR U23284 ( .A(n23463), .B(n23521), .Z(n23523) );
  XNOR U23285 ( .A(n23565), .B(n23566), .Z(n23463) );
  AND U23286 ( .A(n501), .B(n23470), .Z(n23566) );
  XOR U23287 ( .A(n23565), .B(n23468), .Z(n23470) );
  AND U23288 ( .A(n23471), .B(n23474), .Z(n23521) );
  XOR U23289 ( .A(n23567), .B(n23548), .Z(n23474) );
  XNOR U23290 ( .A(p_input[2048]), .B(p_input[672]), .Z(n23548) );
  XOR U23291 ( .A(n23536), .B(n23535), .Z(n23567) );
  XNOR U23292 ( .A(n23568), .B(n23542), .Z(n23535) );
  XNOR U23293 ( .A(n23531), .B(n23530), .Z(n23542) );
  XOR U23294 ( .A(n23569), .B(n23527), .Z(n23530) );
  XNOR U23295 ( .A(n16904), .B(p_input[682]), .Z(n23527) );
  XNOR U23296 ( .A(p_input[2059]), .B(p_input[683]), .Z(n23569) );
  XOR U23297 ( .A(p_input[2060]), .B(p_input[684]), .Z(n23531) );
  XNOR U23298 ( .A(n23541), .B(n23532), .Z(n23568) );
  XNOR U23299 ( .A(n17068), .B(p_input[673]), .Z(n23532) );
  XOR U23300 ( .A(n23570), .B(n23547), .Z(n23541) );
  XNOR U23301 ( .A(p_input[2063]), .B(p_input[687]), .Z(n23547) );
  XOR U23302 ( .A(n23538), .B(n23546), .Z(n23570) );
  XOR U23303 ( .A(n23571), .B(n23543), .Z(n23546) );
  XOR U23304 ( .A(p_input[2061]), .B(p_input[685]), .Z(n23543) );
  XNOR U23305 ( .A(p_input[2062]), .B(p_input[686]), .Z(n23571) );
  XNOR U23306 ( .A(n16738), .B(p_input[681]), .Z(n23538) );
  XNOR U23307 ( .A(n23554), .B(n23553), .Z(n23536) );
  XNOR U23308 ( .A(n23572), .B(n23559), .Z(n23553) );
  XOR U23309 ( .A(p_input[2056]), .B(p_input[680]), .Z(n23559) );
  XOR U23310 ( .A(n23550), .B(n23558), .Z(n23572) );
  XOR U23311 ( .A(n23573), .B(n23555), .Z(n23558) );
  XOR U23312 ( .A(p_input[2054]), .B(p_input[678]), .Z(n23555) );
  XNOR U23313 ( .A(p_input[2055]), .B(p_input[679]), .Z(n23573) );
  XNOR U23314 ( .A(n16741), .B(p_input[674]), .Z(n23550) );
  XNOR U23315 ( .A(n23564), .B(n23563), .Z(n23554) );
  XOR U23316 ( .A(n23574), .B(n23560), .Z(n23563) );
  XOR U23317 ( .A(p_input[2051]), .B(p_input[675]), .Z(n23560) );
  XNOR U23318 ( .A(p_input[2052]), .B(p_input[676]), .Z(n23574) );
  XOR U23319 ( .A(p_input[2053]), .B(p_input[677]), .Z(n23564) );
  XNOR U23320 ( .A(n23575), .B(n23576), .Z(n23471) );
  AND U23321 ( .A(n501), .B(n23577), .Z(n23576) );
  XNOR U23322 ( .A(n23578), .B(n23579), .Z(n501) );
  AND U23323 ( .A(n23580), .B(n23581), .Z(n23579) );
  XOR U23324 ( .A(n23578), .B(n23481), .Z(n23581) );
  XNOR U23325 ( .A(n23578), .B(n23435), .Z(n23580) );
  XOR U23326 ( .A(n23582), .B(n23583), .Z(n23578) );
  AND U23327 ( .A(n23584), .B(n23585), .Z(n23583) );
  XOR U23328 ( .A(n23582), .B(n23445), .Z(n23584) );
  XOR U23329 ( .A(n23586), .B(n23587), .Z(n23424) );
  AND U23330 ( .A(n505), .B(n23577), .Z(n23587) );
  XNOR U23331 ( .A(n23575), .B(n23586), .Z(n23577) );
  XNOR U23332 ( .A(n23588), .B(n23589), .Z(n505) );
  AND U23333 ( .A(n23590), .B(n23591), .Z(n23589) );
  XNOR U23334 ( .A(n23592), .B(n23588), .Z(n23591) );
  IV U23335 ( .A(n23481), .Z(n23592) );
  XNOR U23336 ( .A(n23593), .B(n23594), .Z(n23481) );
  AND U23337 ( .A(n508), .B(n23595), .Z(n23594) );
  XNOR U23338 ( .A(n23593), .B(n23596), .Z(n23595) );
  XNOR U23339 ( .A(n23435), .B(n23588), .Z(n23590) );
  XOR U23340 ( .A(n23597), .B(n23598), .Z(n23435) );
  AND U23341 ( .A(n516), .B(n23599), .Z(n23598) );
  XOR U23342 ( .A(n23582), .B(n23600), .Z(n23588) );
  AND U23343 ( .A(n23601), .B(n23585), .Z(n23600) );
  XNOR U23344 ( .A(n23494), .B(n23582), .Z(n23585) );
  XNOR U23345 ( .A(n23602), .B(n23603), .Z(n23494) );
  AND U23346 ( .A(n508), .B(n23604), .Z(n23603) );
  XOR U23347 ( .A(n23605), .B(n23602), .Z(n23604) );
  XNOR U23348 ( .A(n23606), .B(n23582), .Z(n23601) );
  IV U23349 ( .A(n23445), .Z(n23606) );
  XOR U23350 ( .A(n23607), .B(n23608), .Z(n23445) );
  AND U23351 ( .A(n516), .B(n23609), .Z(n23608) );
  XOR U23352 ( .A(n23610), .B(n23611), .Z(n23582) );
  AND U23353 ( .A(n23612), .B(n23613), .Z(n23611) );
  XNOR U23354 ( .A(n23519), .B(n23610), .Z(n23613) );
  XNOR U23355 ( .A(n23614), .B(n23615), .Z(n23519) );
  AND U23356 ( .A(n508), .B(n23616), .Z(n23615) );
  XNOR U23357 ( .A(n23617), .B(n23614), .Z(n23616) );
  XOR U23358 ( .A(n23610), .B(n23456), .Z(n23612) );
  XOR U23359 ( .A(n23618), .B(n23619), .Z(n23456) );
  AND U23360 ( .A(n516), .B(n23620), .Z(n23619) );
  XOR U23361 ( .A(n23621), .B(n23622), .Z(n23610) );
  AND U23362 ( .A(n23623), .B(n23624), .Z(n23622) );
  XNOR U23363 ( .A(n23621), .B(n23565), .Z(n23624) );
  XNOR U23364 ( .A(n23625), .B(n23626), .Z(n23565) );
  AND U23365 ( .A(n508), .B(n23627), .Z(n23626) );
  XOR U23366 ( .A(n23628), .B(n23625), .Z(n23627) );
  XNOR U23367 ( .A(n23629), .B(n23621), .Z(n23623) );
  IV U23368 ( .A(n23468), .Z(n23629) );
  XOR U23369 ( .A(n23630), .B(n23631), .Z(n23468) );
  AND U23370 ( .A(n516), .B(n23632), .Z(n23631) );
  AND U23371 ( .A(n23586), .B(n23575), .Z(n23621) );
  XNOR U23372 ( .A(n23633), .B(n23634), .Z(n23575) );
  AND U23373 ( .A(n508), .B(n23635), .Z(n23634) );
  XNOR U23374 ( .A(n23636), .B(n23633), .Z(n23635) );
  XNOR U23375 ( .A(n23637), .B(n23638), .Z(n508) );
  AND U23376 ( .A(n23639), .B(n23640), .Z(n23638) );
  XOR U23377 ( .A(n23596), .B(n23637), .Z(n23640) );
  AND U23378 ( .A(n23641), .B(n23642), .Z(n23596) );
  XOR U23379 ( .A(n23637), .B(n23593), .Z(n23639) );
  XNOR U23380 ( .A(n23643), .B(n23644), .Z(n23593) );
  AND U23381 ( .A(n512), .B(n23599), .Z(n23644) );
  XOR U23382 ( .A(n23597), .B(n23643), .Z(n23599) );
  XOR U23383 ( .A(n23645), .B(n23646), .Z(n23637) );
  AND U23384 ( .A(n23647), .B(n23648), .Z(n23646) );
  XNOR U23385 ( .A(n23645), .B(n23641), .Z(n23648) );
  IV U23386 ( .A(n23605), .Z(n23641) );
  XOR U23387 ( .A(n23649), .B(n23650), .Z(n23605) );
  XOR U23388 ( .A(n23651), .B(n23642), .Z(n23650) );
  AND U23389 ( .A(n23617), .B(n23652), .Z(n23642) );
  AND U23390 ( .A(n23653), .B(n23654), .Z(n23651) );
  XOR U23391 ( .A(n23655), .B(n23649), .Z(n23653) );
  XNOR U23392 ( .A(n23602), .B(n23645), .Z(n23647) );
  XNOR U23393 ( .A(n23656), .B(n23657), .Z(n23602) );
  AND U23394 ( .A(n512), .B(n23609), .Z(n23657) );
  XOR U23395 ( .A(n23656), .B(n23607), .Z(n23609) );
  XOR U23396 ( .A(n23658), .B(n23659), .Z(n23645) );
  AND U23397 ( .A(n23660), .B(n23661), .Z(n23659) );
  XNOR U23398 ( .A(n23658), .B(n23617), .Z(n23661) );
  XOR U23399 ( .A(n23662), .B(n23654), .Z(n23617) );
  XNOR U23400 ( .A(n23663), .B(n23649), .Z(n23654) );
  XOR U23401 ( .A(n23664), .B(n23665), .Z(n23649) );
  AND U23402 ( .A(n23666), .B(n23667), .Z(n23665) );
  XOR U23403 ( .A(n23668), .B(n23664), .Z(n23666) );
  XNOR U23404 ( .A(n23669), .B(n23670), .Z(n23663) );
  AND U23405 ( .A(n23671), .B(n23672), .Z(n23670) );
  XOR U23406 ( .A(n23669), .B(n23673), .Z(n23671) );
  XNOR U23407 ( .A(n23655), .B(n23652), .Z(n23662) );
  AND U23408 ( .A(n23674), .B(n23675), .Z(n23652) );
  XOR U23409 ( .A(n23676), .B(n23677), .Z(n23655) );
  AND U23410 ( .A(n23678), .B(n23679), .Z(n23677) );
  XOR U23411 ( .A(n23676), .B(n23680), .Z(n23678) );
  XNOR U23412 ( .A(n23614), .B(n23658), .Z(n23660) );
  XNOR U23413 ( .A(n23681), .B(n23682), .Z(n23614) );
  AND U23414 ( .A(n512), .B(n23620), .Z(n23682) );
  XOR U23415 ( .A(n23681), .B(n23618), .Z(n23620) );
  XOR U23416 ( .A(n23683), .B(n23684), .Z(n23658) );
  AND U23417 ( .A(n23685), .B(n23686), .Z(n23684) );
  XNOR U23418 ( .A(n23683), .B(n23674), .Z(n23686) );
  IV U23419 ( .A(n23628), .Z(n23674) );
  XNOR U23420 ( .A(n23687), .B(n23667), .Z(n23628) );
  XNOR U23421 ( .A(n23688), .B(n23673), .Z(n23667) );
  XOR U23422 ( .A(n23689), .B(n23690), .Z(n23673) );
  NOR U23423 ( .A(n23691), .B(n23692), .Z(n23690) );
  XNOR U23424 ( .A(n23689), .B(n23693), .Z(n23691) );
  XNOR U23425 ( .A(n23672), .B(n23664), .Z(n23688) );
  XOR U23426 ( .A(n23694), .B(n23695), .Z(n23664) );
  AND U23427 ( .A(n23696), .B(n23697), .Z(n23695) );
  XNOR U23428 ( .A(n23694), .B(n23698), .Z(n23696) );
  XNOR U23429 ( .A(n23699), .B(n23669), .Z(n23672) );
  XOR U23430 ( .A(n23700), .B(n23701), .Z(n23669) );
  AND U23431 ( .A(n23702), .B(n23703), .Z(n23701) );
  XOR U23432 ( .A(n23700), .B(n23704), .Z(n23702) );
  XNOR U23433 ( .A(n23705), .B(n23706), .Z(n23699) );
  NOR U23434 ( .A(n23707), .B(n23708), .Z(n23706) );
  XOR U23435 ( .A(n23705), .B(n23709), .Z(n23707) );
  XNOR U23436 ( .A(n23668), .B(n23675), .Z(n23687) );
  NOR U23437 ( .A(n23636), .B(n23710), .Z(n23675) );
  XOR U23438 ( .A(n23680), .B(n23679), .Z(n23668) );
  XNOR U23439 ( .A(n23711), .B(n23676), .Z(n23679) );
  XOR U23440 ( .A(n23712), .B(n23713), .Z(n23676) );
  AND U23441 ( .A(n23714), .B(n23715), .Z(n23713) );
  XOR U23442 ( .A(n23712), .B(n23716), .Z(n23714) );
  XNOR U23443 ( .A(n23717), .B(n23718), .Z(n23711) );
  NOR U23444 ( .A(n23719), .B(n23720), .Z(n23718) );
  XNOR U23445 ( .A(n23717), .B(n23721), .Z(n23719) );
  XOR U23446 ( .A(n23722), .B(n23723), .Z(n23680) );
  NOR U23447 ( .A(n23724), .B(n23725), .Z(n23723) );
  XNOR U23448 ( .A(n23722), .B(n23726), .Z(n23724) );
  XNOR U23449 ( .A(n23625), .B(n23683), .Z(n23685) );
  XNOR U23450 ( .A(n23727), .B(n23728), .Z(n23625) );
  AND U23451 ( .A(n512), .B(n23632), .Z(n23728) );
  XOR U23452 ( .A(n23727), .B(n23630), .Z(n23632) );
  AND U23453 ( .A(n23633), .B(n23636), .Z(n23683) );
  XOR U23454 ( .A(n23729), .B(n23710), .Z(n23636) );
  XNOR U23455 ( .A(p_input[2048]), .B(p_input[688]), .Z(n23710) );
  XOR U23456 ( .A(n23698), .B(n23697), .Z(n23729) );
  XNOR U23457 ( .A(n23730), .B(n23704), .Z(n23697) );
  XNOR U23458 ( .A(n23693), .B(n23692), .Z(n23704) );
  XOR U23459 ( .A(n23731), .B(n23689), .Z(n23692) );
  XNOR U23460 ( .A(n16904), .B(p_input[698]), .Z(n23689) );
  XNOR U23461 ( .A(p_input[2059]), .B(p_input[699]), .Z(n23731) );
  XOR U23462 ( .A(p_input[2060]), .B(p_input[700]), .Z(n23693) );
  XNOR U23463 ( .A(n23703), .B(n23694), .Z(n23730) );
  XNOR U23464 ( .A(n17068), .B(p_input[689]), .Z(n23694) );
  XOR U23465 ( .A(n23732), .B(n23709), .Z(n23703) );
  XNOR U23466 ( .A(p_input[2063]), .B(p_input[703]), .Z(n23709) );
  XOR U23467 ( .A(n23700), .B(n23708), .Z(n23732) );
  XOR U23468 ( .A(n23733), .B(n23705), .Z(n23708) );
  XOR U23469 ( .A(p_input[2061]), .B(p_input[701]), .Z(n23705) );
  XNOR U23470 ( .A(p_input[2062]), .B(p_input[702]), .Z(n23733) );
  XNOR U23471 ( .A(n16738), .B(p_input[697]), .Z(n23700) );
  XNOR U23472 ( .A(n23716), .B(n23715), .Z(n23698) );
  XNOR U23473 ( .A(n23734), .B(n23721), .Z(n23715) );
  XOR U23474 ( .A(p_input[2056]), .B(p_input[696]), .Z(n23721) );
  XOR U23475 ( .A(n23712), .B(n23720), .Z(n23734) );
  XOR U23476 ( .A(n23735), .B(n23717), .Z(n23720) );
  XOR U23477 ( .A(p_input[2054]), .B(p_input[694]), .Z(n23717) );
  XNOR U23478 ( .A(p_input[2055]), .B(p_input[695]), .Z(n23735) );
  XNOR U23479 ( .A(n16741), .B(p_input[690]), .Z(n23712) );
  XNOR U23480 ( .A(n23726), .B(n23725), .Z(n23716) );
  XOR U23481 ( .A(n23736), .B(n23722), .Z(n23725) );
  XOR U23482 ( .A(p_input[2051]), .B(p_input[691]), .Z(n23722) );
  XNOR U23483 ( .A(p_input[2052]), .B(p_input[692]), .Z(n23736) );
  XOR U23484 ( .A(p_input[2053]), .B(p_input[693]), .Z(n23726) );
  XNOR U23485 ( .A(n23737), .B(n23738), .Z(n23633) );
  AND U23486 ( .A(n512), .B(n23739), .Z(n23738) );
  XNOR U23487 ( .A(n23740), .B(n23741), .Z(n512) );
  AND U23488 ( .A(n23742), .B(n23743), .Z(n23741) );
  XOR U23489 ( .A(n23740), .B(n23643), .Z(n23743) );
  XNOR U23490 ( .A(n23740), .B(n23597), .Z(n23742) );
  XOR U23491 ( .A(n23744), .B(n23745), .Z(n23740) );
  AND U23492 ( .A(n23746), .B(n23747), .Z(n23745) );
  XOR U23493 ( .A(n23744), .B(n23607), .Z(n23746) );
  XOR U23494 ( .A(n23748), .B(n23749), .Z(n23586) );
  AND U23495 ( .A(n516), .B(n23739), .Z(n23749) );
  XNOR U23496 ( .A(n23737), .B(n23748), .Z(n23739) );
  XNOR U23497 ( .A(n23750), .B(n23751), .Z(n516) );
  AND U23498 ( .A(n23752), .B(n23753), .Z(n23751) );
  XNOR U23499 ( .A(n23754), .B(n23750), .Z(n23753) );
  IV U23500 ( .A(n23643), .Z(n23754) );
  XNOR U23501 ( .A(n23755), .B(n23756), .Z(n23643) );
  AND U23502 ( .A(n519), .B(n23757), .Z(n23756) );
  XNOR U23503 ( .A(n23755), .B(n23758), .Z(n23757) );
  XNOR U23504 ( .A(n23597), .B(n23750), .Z(n23752) );
  XOR U23505 ( .A(n23759), .B(n23760), .Z(n23597) );
  AND U23506 ( .A(n527), .B(n23761), .Z(n23760) );
  XOR U23507 ( .A(n23744), .B(n23762), .Z(n23750) );
  AND U23508 ( .A(n23763), .B(n23747), .Z(n23762) );
  XNOR U23509 ( .A(n23656), .B(n23744), .Z(n23747) );
  XNOR U23510 ( .A(n23764), .B(n23765), .Z(n23656) );
  AND U23511 ( .A(n519), .B(n23766), .Z(n23765) );
  XOR U23512 ( .A(n23767), .B(n23764), .Z(n23766) );
  XNOR U23513 ( .A(n23768), .B(n23744), .Z(n23763) );
  IV U23514 ( .A(n23607), .Z(n23768) );
  XOR U23515 ( .A(n23769), .B(n23770), .Z(n23607) );
  AND U23516 ( .A(n527), .B(n23771), .Z(n23770) );
  XOR U23517 ( .A(n23772), .B(n23773), .Z(n23744) );
  AND U23518 ( .A(n23774), .B(n23775), .Z(n23773) );
  XNOR U23519 ( .A(n23681), .B(n23772), .Z(n23775) );
  XNOR U23520 ( .A(n23776), .B(n23777), .Z(n23681) );
  AND U23521 ( .A(n519), .B(n23778), .Z(n23777) );
  XNOR U23522 ( .A(n23779), .B(n23776), .Z(n23778) );
  XOR U23523 ( .A(n23772), .B(n23618), .Z(n23774) );
  XOR U23524 ( .A(n23780), .B(n23781), .Z(n23618) );
  AND U23525 ( .A(n527), .B(n23782), .Z(n23781) );
  XOR U23526 ( .A(n23783), .B(n23784), .Z(n23772) );
  AND U23527 ( .A(n23785), .B(n23786), .Z(n23784) );
  XNOR U23528 ( .A(n23783), .B(n23727), .Z(n23786) );
  XNOR U23529 ( .A(n23787), .B(n23788), .Z(n23727) );
  AND U23530 ( .A(n519), .B(n23789), .Z(n23788) );
  XOR U23531 ( .A(n23790), .B(n23787), .Z(n23789) );
  XNOR U23532 ( .A(n23791), .B(n23783), .Z(n23785) );
  IV U23533 ( .A(n23630), .Z(n23791) );
  XOR U23534 ( .A(n23792), .B(n23793), .Z(n23630) );
  AND U23535 ( .A(n527), .B(n23794), .Z(n23793) );
  AND U23536 ( .A(n23748), .B(n23737), .Z(n23783) );
  XNOR U23537 ( .A(n23795), .B(n23796), .Z(n23737) );
  AND U23538 ( .A(n519), .B(n23797), .Z(n23796) );
  XNOR U23539 ( .A(n23798), .B(n23795), .Z(n23797) );
  XNOR U23540 ( .A(n23799), .B(n23800), .Z(n519) );
  AND U23541 ( .A(n23801), .B(n23802), .Z(n23800) );
  XOR U23542 ( .A(n23758), .B(n23799), .Z(n23802) );
  AND U23543 ( .A(n23803), .B(n23804), .Z(n23758) );
  XOR U23544 ( .A(n23799), .B(n23755), .Z(n23801) );
  XNOR U23545 ( .A(n23805), .B(n23806), .Z(n23755) );
  AND U23546 ( .A(n523), .B(n23761), .Z(n23806) );
  XOR U23547 ( .A(n23759), .B(n23805), .Z(n23761) );
  XOR U23548 ( .A(n23807), .B(n23808), .Z(n23799) );
  AND U23549 ( .A(n23809), .B(n23810), .Z(n23808) );
  XNOR U23550 ( .A(n23807), .B(n23803), .Z(n23810) );
  IV U23551 ( .A(n23767), .Z(n23803) );
  XOR U23552 ( .A(n23811), .B(n23812), .Z(n23767) );
  XOR U23553 ( .A(n23813), .B(n23804), .Z(n23812) );
  AND U23554 ( .A(n23779), .B(n23814), .Z(n23804) );
  AND U23555 ( .A(n23815), .B(n23816), .Z(n23813) );
  XOR U23556 ( .A(n23817), .B(n23811), .Z(n23815) );
  XNOR U23557 ( .A(n23764), .B(n23807), .Z(n23809) );
  XNOR U23558 ( .A(n23818), .B(n23819), .Z(n23764) );
  AND U23559 ( .A(n523), .B(n23771), .Z(n23819) );
  XOR U23560 ( .A(n23818), .B(n23769), .Z(n23771) );
  XOR U23561 ( .A(n23820), .B(n23821), .Z(n23807) );
  AND U23562 ( .A(n23822), .B(n23823), .Z(n23821) );
  XNOR U23563 ( .A(n23820), .B(n23779), .Z(n23823) );
  XOR U23564 ( .A(n23824), .B(n23816), .Z(n23779) );
  XNOR U23565 ( .A(n23825), .B(n23811), .Z(n23816) );
  XOR U23566 ( .A(n23826), .B(n23827), .Z(n23811) );
  AND U23567 ( .A(n23828), .B(n23829), .Z(n23827) );
  XOR U23568 ( .A(n23830), .B(n23826), .Z(n23828) );
  XNOR U23569 ( .A(n23831), .B(n23832), .Z(n23825) );
  AND U23570 ( .A(n23833), .B(n23834), .Z(n23832) );
  XOR U23571 ( .A(n23831), .B(n23835), .Z(n23833) );
  XNOR U23572 ( .A(n23817), .B(n23814), .Z(n23824) );
  AND U23573 ( .A(n23836), .B(n23837), .Z(n23814) );
  XOR U23574 ( .A(n23838), .B(n23839), .Z(n23817) );
  AND U23575 ( .A(n23840), .B(n23841), .Z(n23839) );
  XOR U23576 ( .A(n23838), .B(n23842), .Z(n23840) );
  XNOR U23577 ( .A(n23776), .B(n23820), .Z(n23822) );
  XNOR U23578 ( .A(n23843), .B(n23844), .Z(n23776) );
  AND U23579 ( .A(n523), .B(n23782), .Z(n23844) );
  XOR U23580 ( .A(n23843), .B(n23780), .Z(n23782) );
  XOR U23581 ( .A(n23845), .B(n23846), .Z(n23820) );
  AND U23582 ( .A(n23847), .B(n23848), .Z(n23846) );
  XNOR U23583 ( .A(n23845), .B(n23836), .Z(n23848) );
  IV U23584 ( .A(n23790), .Z(n23836) );
  XNOR U23585 ( .A(n23849), .B(n23829), .Z(n23790) );
  XNOR U23586 ( .A(n23850), .B(n23835), .Z(n23829) );
  XOR U23587 ( .A(n23851), .B(n23852), .Z(n23835) );
  NOR U23588 ( .A(n23853), .B(n23854), .Z(n23852) );
  XNOR U23589 ( .A(n23851), .B(n23855), .Z(n23853) );
  XNOR U23590 ( .A(n23834), .B(n23826), .Z(n23850) );
  XOR U23591 ( .A(n23856), .B(n23857), .Z(n23826) );
  AND U23592 ( .A(n23858), .B(n23859), .Z(n23857) );
  XNOR U23593 ( .A(n23856), .B(n23860), .Z(n23858) );
  XNOR U23594 ( .A(n23861), .B(n23831), .Z(n23834) );
  XOR U23595 ( .A(n23862), .B(n23863), .Z(n23831) );
  AND U23596 ( .A(n23864), .B(n23865), .Z(n23863) );
  XOR U23597 ( .A(n23862), .B(n23866), .Z(n23864) );
  XNOR U23598 ( .A(n23867), .B(n23868), .Z(n23861) );
  NOR U23599 ( .A(n23869), .B(n23870), .Z(n23868) );
  XOR U23600 ( .A(n23867), .B(n23871), .Z(n23869) );
  XNOR U23601 ( .A(n23830), .B(n23837), .Z(n23849) );
  NOR U23602 ( .A(n23798), .B(n23872), .Z(n23837) );
  XOR U23603 ( .A(n23842), .B(n23841), .Z(n23830) );
  XNOR U23604 ( .A(n23873), .B(n23838), .Z(n23841) );
  XOR U23605 ( .A(n23874), .B(n23875), .Z(n23838) );
  AND U23606 ( .A(n23876), .B(n23877), .Z(n23875) );
  XOR U23607 ( .A(n23874), .B(n23878), .Z(n23876) );
  XNOR U23608 ( .A(n23879), .B(n23880), .Z(n23873) );
  NOR U23609 ( .A(n23881), .B(n23882), .Z(n23880) );
  XNOR U23610 ( .A(n23879), .B(n23883), .Z(n23881) );
  XOR U23611 ( .A(n23884), .B(n23885), .Z(n23842) );
  NOR U23612 ( .A(n23886), .B(n23887), .Z(n23885) );
  XNOR U23613 ( .A(n23884), .B(n23888), .Z(n23886) );
  XNOR U23614 ( .A(n23787), .B(n23845), .Z(n23847) );
  XNOR U23615 ( .A(n23889), .B(n23890), .Z(n23787) );
  AND U23616 ( .A(n523), .B(n23794), .Z(n23890) );
  XOR U23617 ( .A(n23889), .B(n23792), .Z(n23794) );
  AND U23618 ( .A(n23795), .B(n23798), .Z(n23845) );
  XOR U23619 ( .A(n23891), .B(n23872), .Z(n23798) );
  XNOR U23620 ( .A(p_input[2048]), .B(p_input[704]), .Z(n23872) );
  XOR U23621 ( .A(n23860), .B(n23859), .Z(n23891) );
  XNOR U23622 ( .A(n23892), .B(n23866), .Z(n23859) );
  XNOR U23623 ( .A(n23855), .B(n23854), .Z(n23866) );
  XOR U23624 ( .A(n23893), .B(n23851), .Z(n23854) );
  XNOR U23625 ( .A(n16904), .B(p_input[714]), .Z(n23851) );
  XNOR U23626 ( .A(p_input[2059]), .B(p_input[715]), .Z(n23893) );
  XOR U23627 ( .A(p_input[2060]), .B(p_input[716]), .Z(n23855) );
  XNOR U23628 ( .A(n23865), .B(n23856), .Z(n23892) );
  XNOR U23629 ( .A(n17068), .B(p_input[705]), .Z(n23856) );
  XOR U23630 ( .A(n23894), .B(n23871), .Z(n23865) );
  XNOR U23631 ( .A(p_input[2063]), .B(p_input[719]), .Z(n23871) );
  XOR U23632 ( .A(n23862), .B(n23870), .Z(n23894) );
  XOR U23633 ( .A(n23895), .B(n23867), .Z(n23870) );
  XOR U23634 ( .A(p_input[2061]), .B(p_input[717]), .Z(n23867) );
  XNOR U23635 ( .A(p_input[2062]), .B(p_input[718]), .Z(n23895) );
  XNOR U23636 ( .A(n16738), .B(p_input[713]), .Z(n23862) );
  XNOR U23637 ( .A(n23878), .B(n23877), .Z(n23860) );
  XNOR U23638 ( .A(n23896), .B(n23883), .Z(n23877) );
  XOR U23639 ( .A(p_input[2056]), .B(p_input[712]), .Z(n23883) );
  XOR U23640 ( .A(n23874), .B(n23882), .Z(n23896) );
  XOR U23641 ( .A(n23897), .B(n23879), .Z(n23882) );
  XOR U23642 ( .A(p_input[2054]), .B(p_input[710]), .Z(n23879) );
  XNOR U23643 ( .A(p_input[2055]), .B(p_input[711]), .Z(n23897) );
  XNOR U23644 ( .A(n16741), .B(p_input[706]), .Z(n23874) );
  XNOR U23645 ( .A(n23888), .B(n23887), .Z(n23878) );
  XOR U23646 ( .A(n23898), .B(n23884), .Z(n23887) );
  XOR U23647 ( .A(p_input[2051]), .B(p_input[707]), .Z(n23884) );
  XNOR U23648 ( .A(p_input[2052]), .B(p_input[708]), .Z(n23898) );
  XOR U23649 ( .A(p_input[2053]), .B(p_input[709]), .Z(n23888) );
  XNOR U23650 ( .A(n23899), .B(n23900), .Z(n23795) );
  AND U23651 ( .A(n523), .B(n23901), .Z(n23900) );
  XNOR U23652 ( .A(n23902), .B(n23903), .Z(n523) );
  AND U23653 ( .A(n23904), .B(n23905), .Z(n23903) );
  XOR U23654 ( .A(n23902), .B(n23805), .Z(n23905) );
  XNOR U23655 ( .A(n23902), .B(n23759), .Z(n23904) );
  XOR U23656 ( .A(n23906), .B(n23907), .Z(n23902) );
  AND U23657 ( .A(n23908), .B(n23909), .Z(n23907) );
  XOR U23658 ( .A(n23906), .B(n23769), .Z(n23908) );
  XOR U23659 ( .A(n23910), .B(n23911), .Z(n23748) );
  AND U23660 ( .A(n527), .B(n23901), .Z(n23911) );
  XNOR U23661 ( .A(n23899), .B(n23910), .Z(n23901) );
  XNOR U23662 ( .A(n23912), .B(n23913), .Z(n527) );
  AND U23663 ( .A(n23914), .B(n23915), .Z(n23913) );
  XNOR U23664 ( .A(n23916), .B(n23912), .Z(n23915) );
  IV U23665 ( .A(n23805), .Z(n23916) );
  XNOR U23666 ( .A(n23917), .B(n23918), .Z(n23805) );
  AND U23667 ( .A(n530), .B(n23919), .Z(n23918) );
  XNOR U23668 ( .A(n23917), .B(n23920), .Z(n23919) );
  XNOR U23669 ( .A(n23759), .B(n23912), .Z(n23914) );
  XOR U23670 ( .A(n23921), .B(n23922), .Z(n23759) );
  AND U23671 ( .A(n538), .B(n23923), .Z(n23922) );
  XOR U23672 ( .A(n23906), .B(n23924), .Z(n23912) );
  AND U23673 ( .A(n23925), .B(n23909), .Z(n23924) );
  XNOR U23674 ( .A(n23818), .B(n23906), .Z(n23909) );
  XNOR U23675 ( .A(n23926), .B(n23927), .Z(n23818) );
  AND U23676 ( .A(n530), .B(n23928), .Z(n23927) );
  XOR U23677 ( .A(n23929), .B(n23926), .Z(n23928) );
  XNOR U23678 ( .A(n23930), .B(n23906), .Z(n23925) );
  IV U23679 ( .A(n23769), .Z(n23930) );
  XOR U23680 ( .A(n23931), .B(n23932), .Z(n23769) );
  AND U23681 ( .A(n538), .B(n23933), .Z(n23932) );
  XOR U23682 ( .A(n23934), .B(n23935), .Z(n23906) );
  AND U23683 ( .A(n23936), .B(n23937), .Z(n23935) );
  XNOR U23684 ( .A(n23843), .B(n23934), .Z(n23937) );
  XNOR U23685 ( .A(n23938), .B(n23939), .Z(n23843) );
  AND U23686 ( .A(n530), .B(n23940), .Z(n23939) );
  XNOR U23687 ( .A(n23941), .B(n23938), .Z(n23940) );
  XOR U23688 ( .A(n23934), .B(n23780), .Z(n23936) );
  XOR U23689 ( .A(n23942), .B(n23943), .Z(n23780) );
  AND U23690 ( .A(n538), .B(n23944), .Z(n23943) );
  XOR U23691 ( .A(n23945), .B(n23946), .Z(n23934) );
  AND U23692 ( .A(n23947), .B(n23948), .Z(n23946) );
  XNOR U23693 ( .A(n23945), .B(n23889), .Z(n23948) );
  XNOR U23694 ( .A(n23949), .B(n23950), .Z(n23889) );
  AND U23695 ( .A(n530), .B(n23951), .Z(n23950) );
  XOR U23696 ( .A(n23952), .B(n23949), .Z(n23951) );
  XNOR U23697 ( .A(n23953), .B(n23945), .Z(n23947) );
  IV U23698 ( .A(n23792), .Z(n23953) );
  XOR U23699 ( .A(n23954), .B(n23955), .Z(n23792) );
  AND U23700 ( .A(n538), .B(n23956), .Z(n23955) );
  AND U23701 ( .A(n23910), .B(n23899), .Z(n23945) );
  XNOR U23702 ( .A(n23957), .B(n23958), .Z(n23899) );
  AND U23703 ( .A(n530), .B(n23959), .Z(n23958) );
  XNOR U23704 ( .A(n23960), .B(n23957), .Z(n23959) );
  XNOR U23705 ( .A(n23961), .B(n23962), .Z(n530) );
  AND U23706 ( .A(n23963), .B(n23964), .Z(n23962) );
  XOR U23707 ( .A(n23920), .B(n23961), .Z(n23964) );
  AND U23708 ( .A(n23965), .B(n23966), .Z(n23920) );
  XOR U23709 ( .A(n23961), .B(n23917), .Z(n23963) );
  XNOR U23710 ( .A(n23967), .B(n23968), .Z(n23917) );
  AND U23711 ( .A(n534), .B(n23923), .Z(n23968) );
  XOR U23712 ( .A(n23921), .B(n23967), .Z(n23923) );
  XOR U23713 ( .A(n23969), .B(n23970), .Z(n23961) );
  AND U23714 ( .A(n23971), .B(n23972), .Z(n23970) );
  XNOR U23715 ( .A(n23969), .B(n23965), .Z(n23972) );
  IV U23716 ( .A(n23929), .Z(n23965) );
  XOR U23717 ( .A(n23973), .B(n23974), .Z(n23929) );
  XOR U23718 ( .A(n23975), .B(n23966), .Z(n23974) );
  AND U23719 ( .A(n23941), .B(n23976), .Z(n23966) );
  AND U23720 ( .A(n23977), .B(n23978), .Z(n23975) );
  XOR U23721 ( .A(n23979), .B(n23973), .Z(n23977) );
  XNOR U23722 ( .A(n23926), .B(n23969), .Z(n23971) );
  XNOR U23723 ( .A(n23980), .B(n23981), .Z(n23926) );
  AND U23724 ( .A(n534), .B(n23933), .Z(n23981) );
  XOR U23725 ( .A(n23980), .B(n23931), .Z(n23933) );
  XOR U23726 ( .A(n23982), .B(n23983), .Z(n23969) );
  AND U23727 ( .A(n23984), .B(n23985), .Z(n23983) );
  XNOR U23728 ( .A(n23982), .B(n23941), .Z(n23985) );
  XOR U23729 ( .A(n23986), .B(n23978), .Z(n23941) );
  XNOR U23730 ( .A(n23987), .B(n23973), .Z(n23978) );
  XOR U23731 ( .A(n23988), .B(n23989), .Z(n23973) );
  AND U23732 ( .A(n23990), .B(n23991), .Z(n23989) );
  XOR U23733 ( .A(n23992), .B(n23988), .Z(n23990) );
  XNOR U23734 ( .A(n23993), .B(n23994), .Z(n23987) );
  AND U23735 ( .A(n23995), .B(n23996), .Z(n23994) );
  XOR U23736 ( .A(n23993), .B(n23997), .Z(n23995) );
  XNOR U23737 ( .A(n23979), .B(n23976), .Z(n23986) );
  AND U23738 ( .A(n23998), .B(n23999), .Z(n23976) );
  XOR U23739 ( .A(n24000), .B(n24001), .Z(n23979) );
  AND U23740 ( .A(n24002), .B(n24003), .Z(n24001) );
  XOR U23741 ( .A(n24000), .B(n24004), .Z(n24002) );
  XNOR U23742 ( .A(n23938), .B(n23982), .Z(n23984) );
  XNOR U23743 ( .A(n24005), .B(n24006), .Z(n23938) );
  AND U23744 ( .A(n534), .B(n23944), .Z(n24006) );
  XOR U23745 ( .A(n24005), .B(n23942), .Z(n23944) );
  XOR U23746 ( .A(n24007), .B(n24008), .Z(n23982) );
  AND U23747 ( .A(n24009), .B(n24010), .Z(n24008) );
  XNOR U23748 ( .A(n24007), .B(n23998), .Z(n24010) );
  IV U23749 ( .A(n23952), .Z(n23998) );
  XNOR U23750 ( .A(n24011), .B(n23991), .Z(n23952) );
  XNOR U23751 ( .A(n24012), .B(n23997), .Z(n23991) );
  XOR U23752 ( .A(n24013), .B(n24014), .Z(n23997) );
  NOR U23753 ( .A(n24015), .B(n24016), .Z(n24014) );
  XNOR U23754 ( .A(n24013), .B(n24017), .Z(n24015) );
  XNOR U23755 ( .A(n23996), .B(n23988), .Z(n24012) );
  XOR U23756 ( .A(n24018), .B(n24019), .Z(n23988) );
  AND U23757 ( .A(n24020), .B(n24021), .Z(n24019) );
  XNOR U23758 ( .A(n24018), .B(n24022), .Z(n24020) );
  XNOR U23759 ( .A(n24023), .B(n23993), .Z(n23996) );
  XOR U23760 ( .A(n24024), .B(n24025), .Z(n23993) );
  AND U23761 ( .A(n24026), .B(n24027), .Z(n24025) );
  XOR U23762 ( .A(n24024), .B(n24028), .Z(n24026) );
  XNOR U23763 ( .A(n24029), .B(n24030), .Z(n24023) );
  NOR U23764 ( .A(n24031), .B(n24032), .Z(n24030) );
  XOR U23765 ( .A(n24029), .B(n24033), .Z(n24031) );
  XNOR U23766 ( .A(n23992), .B(n23999), .Z(n24011) );
  NOR U23767 ( .A(n23960), .B(n24034), .Z(n23999) );
  XOR U23768 ( .A(n24004), .B(n24003), .Z(n23992) );
  XNOR U23769 ( .A(n24035), .B(n24000), .Z(n24003) );
  XOR U23770 ( .A(n24036), .B(n24037), .Z(n24000) );
  AND U23771 ( .A(n24038), .B(n24039), .Z(n24037) );
  XOR U23772 ( .A(n24036), .B(n24040), .Z(n24038) );
  XNOR U23773 ( .A(n24041), .B(n24042), .Z(n24035) );
  NOR U23774 ( .A(n24043), .B(n24044), .Z(n24042) );
  XNOR U23775 ( .A(n24041), .B(n24045), .Z(n24043) );
  XOR U23776 ( .A(n24046), .B(n24047), .Z(n24004) );
  NOR U23777 ( .A(n24048), .B(n24049), .Z(n24047) );
  XNOR U23778 ( .A(n24046), .B(n24050), .Z(n24048) );
  XNOR U23779 ( .A(n23949), .B(n24007), .Z(n24009) );
  XNOR U23780 ( .A(n24051), .B(n24052), .Z(n23949) );
  AND U23781 ( .A(n534), .B(n23956), .Z(n24052) );
  XOR U23782 ( .A(n24051), .B(n23954), .Z(n23956) );
  AND U23783 ( .A(n23957), .B(n23960), .Z(n24007) );
  XOR U23784 ( .A(n24053), .B(n24034), .Z(n23960) );
  XNOR U23785 ( .A(p_input[2048]), .B(p_input[720]), .Z(n24034) );
  XOR U23786 ( .A(n24022), .B(n24021), .Z(n24053) );
  XNOR U23787 ( .A(n24054), .B(n24028), .Z(n24021) );
  XNOR U23788 ( .A(n24017), .B(n24016), .Z(n24028) );
  XOR U23789 ( .A(n24055), .B(n24013), .Z(n24016) );
  XNOR U23790 ( .A(n16904), .B(p_input[730]), .Z(n24013) );
  XNOR U23791 ( .A(p_input[2059]), .B(p_input[731]), .Z(n24055) );
  XOR U23792 ( .A(p_input[2060]), .B(p_input[732]), .Z(n24017) );
  XNOR U23793 ( .A(n24027), .B(n24018), .Z(n24054) );
  XNOR U23794 ( .A(n17068), .B(p_input[721]), .Z(n24018) );
  XOR U23795 ( .A(n24056), .B(n24033), .Z(n24027) );
  XNOR U23796 ( .A(p_input[2063]), .B(p_input[735]), .Z(n24033) );
  XOR U23797 ( .A(n24024), .B(n24032), .Z(n24056) );
  XOR U23798 ( .A(n24057), .B(n24029), .Z(n24032) );
  XOR U23799 ( .A(p_input[2061]), .B(p_input[733]), .Z(n24029) );
  XNOR U23800 ( .A(p_input[2062]), .B(p_input[734]), .Z(n24057) );
  XNOR U23801 ( .A(n16738), .B(p_input[729]), .Z(n24024) );
  XNOR U23802 ( .A(n24040), .B(n24039), .Z(n24022) );
  XNOR U23803 ( .A(n24058), .B(n24045), .Z(n24039) );
  XOR U23804 ( .A(p_input[2056]), .B(p_input[728]), .Z(n24045) );
  XOR U23805 ( .A(n24036), .B(n24044), .Z(n24058) );
  XOR U23806 ( .A(n24059), .B(n24041), .Z(n24044) );
  XOR U23807 ( .A(p_input[2054]), .B(p_input[726]), .Z(n24041) );
  XNOR U23808 ( .A(p_input[2055]), .B(p_input[727]), .Z(n24059) );
  XNOR U23809 ( .A(n16741), .B(p_input[722]), .Z(n24036) );
  XNOR U23810 ( .A(n24050), .B(n24049), .Z(n24040) );
  XOR U23811 ( .A(n24060), .B(n24046), .Z(n24049) );
  XOR U23812 ( .A(p_input[2051]), .B(p_input[723]), .Z(n24046) );
  XNOR U23813 ( .A(p_input[2052]), .B(p_input[724]), .Z(n24060) );
  XOR U23814 ( .A(p_input[2053]), .B(p_input[725]), .Z(n24050) );
  XNOR U23815 ( .A(n24061), .B(n24062), .Z(n23957) );
  AND U23816 ( .A(n534), .B(n24063), .Z(n24062) );
  XNOR U23817 ( .A(n24064), .B(n24065), .Z(n534) );
  AND U23818 ( .A(n24066), .B(n24067), .Z(n24065) );
  XOR U23819 ( .A(n24064), .B(n23967), .Z(n24067) );
  XNOR U23820 ( .A(n24064), .B(n23921), .Z(n24066) );
  XOR U23821 ( .A(n24068), .B(n24069), .Z(n24064) );
  AND U23822 ( .A(n24070), .B(n24071), .Z(n24069) );
  XOR U23823 ( .A(n24068), .B(n23931), .Z(n24070) );
  XOR U23824 ( .A(n24072), .B(n24073), .Z(n23910) );
  AND U23825 ( .A(n538), .B(n24063), .Z(n24073) );
  XNOR U23826 ( .A(n24061), .B(n24072), .Z(n24063) );
  XNOR U23827 ( .A(n24074), .B(n24075), .Z(n538) );
  AND U23828 ( .A(n24076), .B(n24077), .Z(n24075) );
  XNOR U23829 ( .A(n24078), .B(n24074), .Z(n24077) );
  IV U23830 ( .A(n23967), .Z(n24078) );
  XNOR U23831 ( .A(n24079), .B(n24080), .Z(n23967) );
  AND U23832 ( .A(n541), .B(n24081), .Z(n24080) );
  XNOR U23833 ( .A(n24079), .B(n24082), .Z(n24081) );
  XNOR U23834 ( .A(n23921), .B(n24074), .Z(n24076) );
  XOR U23835 ( .A(n24083), .B(n24084), .Z(n23921) );
  AND U23836 ( .A(n549), .B(n24085), .Z(n24084) );
  XOR U23837 ( .A(n24068), .B(n24086), .Z(n24074) );
  AND U23838 ( .A(n24087), .B(n24071), .Z(n24086) );
  XNOR U23839 ( .A(n23980), .B(n24068), .Z(n24071) );
  XNOR U23840 ( .A(n24088), .B(n24089), .Z(n23980) );
  AND U23841 ( .A(n541), .B(n24090), .Z(n24089) );
  XOR U23842 ( .A(n24091), .B(n24088), .Z(n24090) );
  XNOR U23843 ( .A(n24092), .B(n24068), .Z(n24087) );
  IV U23844 ( .A(n23931), .Z(n24092) );
  XOR U23845 ( .A(n24093), .B(n24094), .Z(n23931) );
  AND U23846 ( .A(n549), .B(n24095), .Z(n24094) );
  XOR U23847 ( .A(n24096), .B(n24097), .Z(n24068) );
  AND U23848 ( .A(n24098), .B(n24099), .Z(n24097) );
  XNOR U23849 ( .A(n24005), .B(n24096), .Z(n24099) );
  XNOR U23850 ( .A(n24100), .B(n24101), .Z(n24005) );
  AND U23851 ( .A(n541), .B(n24102), .Z(n24101) );
  XNOR U23852 ( .A(n24103), .B(n24100), .Z(n24102) );
  XOR U23853 ( .A(n24096), .B(n23942), .Z(n24098) );
  XOR U23854 ( .A(n24104), .B(n24105), .Z(n23942) );
  AND U23855 ( .A(n549), .B(n24106), .Z(n24105) );
  XOR U23856 ( .A(n24107), .B(n24108), .Z(n24096) );
  AND U23857 ( .A(n24109), .B(n24110), .Z(n24108) );
  XNOR U23858 ( .A(n24107), .B(n24051), .Z(n24110) );
  XNOR U23859 ( .A(n24111), .B(n24112), .Z(n24051) );
  AND U23860 ( .A(n541), .B(n24113), .Z(n24112) );
  XOR U23861 ( .A(n24114), .B(n24111), .Z(n24113) );
  XNOR U23862 ( .A(n24115), .B(n24107), .Z(n24109) );
  IV U23863 ( .A(n23954), .Z(n24115) );
  XOR U23864 ( .A(n24116), .B(n24117), .Z(n23954) );
  AND U23865 ( .A(n549), .B(n24118), .Z(n24117) );
  AND U23866 ( .A(n24072), .B(n24061), .Z(n24107) );
  XNOR U23867 ( .A(n24119), .B(n24120), .Z(n24061) );
  AND U23868 ( .A(n541), .B(n24121), .Z(n24120) );
  XNOR U23869 ( .A(n24122), .B(n24119), .Z(n24121) );
  XNOR U23870 ( .A(n24123), .B(n24124), .Z(n541) );
  AND U23871 ( .A(n24125), .B(n24126), .Z(n24124) );
  XOR U23872 ( .A(n24082), .B(n24123), .Z(n24126) );
  AND U23873 ( .A(n24127), .B(n24128), .Z(n24082) );
  XOR U23874 ( .A(n24123), .B(n24079), .Z(n24125) );
  XNOR U23875 ( .A(n24129), .B(n24130), .Z(n24079) );
  AND U23876 ( .A(n545), .B(n24085), .Z(n24130) );
  XOR U23877 ( .A(n24083), .B(n24129), .Z(n24085) );
  XOR U23878 ( .A(n24131), .B(n24132), .Z(n24123) );
  AND U23879 ( .A(n24133), .B(n24134), .Z(n24132) );
  XNOR U23880 ( .A(n24131), .B(n24127), .Z(n24134) );
  IV U23881 ( .A(n24091), .Z(n24127) );
  XOR U23882 ( .A(n24135), .B(n24136), .Z(n24091) );
  XOR U23883 ( .A(n24137), .B(n24128), .Z(n24136) );
  AND U23884 ( .A(n24103), .B(n24138), .Z(n24128) );
  AND U23885 ( .A(n24139), .B(n24140), .Z(n24137) );
  XOR U23886 ( .A(n24141), .B(n24135), .Z(n24139) );
  XNOR U23887 ( .A(n24088), .B(n24131), .Z(n24133) );
  XNOR U23888 ( .A(n24142), .B(n24143), .Z(n24088) );
  AND U23889 ( .A(n545), .B(n24095), .Z(n24143) );
  XOR U23890 ( .A(n24142), .B(n24093), .Z(n24095) );
  XOR U23891 ( .A(n24144), .B(n24145), .Z(n24131) );
  AND U23892 ( .A(n24146), .B(n24147), .Z(n24145) );
  XNOR U23893 ( .A(n24144), .B(n24103), .Z(n24147) );
  XOR U23894 ( .A(n24148), .B(n24140), .Z(n24103) );
  XNOR U23895 ( .A(n24149), .B(n24135), .Z(n24140) );
  XOR U23896 ( .A(n24150), .B(n24151), .Z(n24135) );
  AND U23897 ( .A(n24152), .B(n24153), .Z(n24151) );
  XOR U23898 ( .A(n24154), .B(n24150), .Z(n24152) );
  XNOR U23899 ( .A(n24155), .B(n24156), .Z(n24149) );
  AND U23900 ( .A(n24157), .B(n24158), .Z(n24156) );
  XOR U23901 ( .A(n24155), .B(n24159), .Z(n24157) );
  XNOR U23902 ( .A(n24141), .B(n24138), .Z(n24148) );
  AND U23903 ( .A(n24160), .B(n24161), .Z(n24138) );
  XOR U23904 ( .A(n24162), .B(n24163), .Z(n24141) );
  AND U23905 ( .A(n24164), .B(n24165), .Z(n24163) );
  XOR U23906 ( .A(n24162), .B(n24166), .Z(n24164) );
  XNOR U23907 ( .A(n24100), .B(n24144), .Z(n24146) );
  XNOR U23908 ( .A(n24167), .B(n24168), .Z(n24100) );
  AND U23909 ( .A(n545), .B(n24106), .Z(n24168) );
  XOR U23910 ( .A(n24167), .B(n24104), .Z(n24106) );
  XOR U23911 ( .A(n24169), .B(n24170), .Z(n24144) );
  AND U23912 ( .A(n24171), .B(n24172), .Z(n24170) );
  XNOR U23913 ( .A(n24169), .B(n24160), .Z(n24172) );
  IV U23914 ( .A(n24114), .Z(n24160) );
  XNOR U23915 ( .A(n24173), .B(n24153), .Z(n24114) );
  XNOR U23916 ( .A(n24174), .B(n24159), .Z(n24153) );
  XOR U23917 ( .A(n24175), .B(n24176), .Z(n24159) );
  NOR U23918 ( .A(n24177), .B(n24178), .Z(n24176) );
  XNOR U23919 ( .A(n24175), .B(n24179), .Z(n24177) );
  XNOR U23920 ( .A(n24158), .B(n24150), .Z(n24174) );
  XOR U23921 ( .A(n24180), .B(n24181), .Z(n24150) );
  AND U23922 ( .A(n24182), .B(n24183), .Z(n24181) );
  XNOR U23923 ( .A(n24180), .B(n24184), .Z(n24182) );
  XNOR U23924 ( .A(n24185), .B(n24155), .Z(n24158) );
  XOR U23925 ( .A(n24186), .B(n24187), .Z(n24155) );
  AND U23926 ( .A(n24188), .B(n24189), .Z(n24187) );
  XOR U23927 ( .A(n24186), .B(n24190), .Z(n24188) );
  XNOR U23928 ( .A(n24191), .B(n24192), .Z(n24185) );
  NOR U23929 ( .A(n24193), .B(n24194), .Z(n24192) );
  XOR U23930 ( .A(n24191), .B(n24195), .Z(n24193) );
  XNOR U23931 ( .A(n24154), .B(n24161), .Z(n24173) );
  NOR U23932 ( .A(n24122), .B(n24196), .Z(n24161) );
  XOR U23933 ( .A(n24166), .B(n24165), .Z(n24154) );
  XNOR U23934 ( .A(n24197), .B(n24162), .Z(n24165) );
  XOR U23935 ( .A(n24198), .B(n24199), .Z(n24162) );
  AND U23936 ( .A(n24200), .B(n24201), .Z(n24199) );
  XOR U23937 ( .A(n24198), .B(n24202), .Z(n24200) );
  XNOR U23938 ( .A(n24203), .B(n24204), .Z(n24197) );
  NOR U23939 ( .A(n24205), .B(n24206), .Z(n24204) );
  XNOR U23940 ( .A(n24203), .B(n24207), .Z(n24205) );
  XOR U23941 ( .A(n24208), .B(n24209), .Z(n24166) );
  NOR U23942 ( .A(n24210), .B(n24211), .Z(n24209) );
  XNOR U23943 ( .A(n24208), .B(n24212), .Z(n24210) );
  XNOR U23944 ( .A(n24111), .B(n24169), .Z(n24171) );
  XNOR U23945 ( .A(n24213), .B(n24214), .Z(n24111) );
  AND U23946 ( .A(n545), .B(n24118), .Z(n24214) );
  XOR U23947 ( .A(n24213), .B(n24116), .Z(n24118) );
  AND U23948 ( .A(n24119), .B(n24122), .Z(n24169) );
  XOR U23949 ( .A(n24215), .B(n24196), .Z(n24122) );
  XNOR U23950 ( .A(p_input[2048]), .B(p_input[736]), .Z(n24196) );
  XOR U23951 ( .A(n24184), .B(n24183), .Z(n24215) );
  XNOR U23952 ( .A(n24216), .B(n24190), .Z(n24183) );
  XNOR U23953 ( .A(n24179), .B(n24178), .Z(n24190) );
  XOR U23954 ( .A(n24217), .B(n24175), .Z(n24178) );
  XNOR U23955 ( .A(n16904), .B(p_input[746]), .Z(n24175) );
  XNOR U23956 ( .A(p_input[2059]), .B(p_input[747]), .Z(n24217) );
  XOR U23957 ( .A(p_input[2060]), .B(p_input[748]), .Z(n24179) );
  XNOR U23958 ( .A(n24189), .B(n24180), .Z(n24216) );
  XNOR U23959 ( .A(n17068), .B(p_input[737]), .Z(n24180) );
  XOR U23960 ( .A(n24218), .B(n24195), .Z(n24189) );
  XNOR U23961 ( .A(p_input[2063]), .B(p_input[751]), .Z(n24195) );
  XOR U23962 ( .A(n24186), .B(n24194), .Z(n24218) );
  XOR U23963 ( .A(n24219), .B(n24191), .Z(n24194) );
  XOR U23964 ( .A(p_input[2061]), .B(p_input[749]), .Z(n24191) );
  XNOR U23965 ( .A(p_input[2062]), .B(p_input[750]), .Z(n24219) );
  XNOR U23966 ( .A(n16738), .B(p_input[745]), .Z(n24186) );
  XNOR U23967 ( .A(n24202), .B(n24201), .Z(n24184) );
  XNOR U23968 ( .A(n24220), .B(n24207), .Z(n24201) );
  XOR U23969 ( .A(p_input[2056]), .B(p_input[744]), .Z(n24207) );
  XOR U23970 ( .A(n24198), .B(n24206), .Z(n24220) );
  XOR U23971 ( .A(n24221), .B(n24203), .Z(n24206) );
  XOR U23972 ( .A(p_input[2054]), .B(p_input[742]), .Z(n24203) );
  XNOR U23973 ( .A(p_input[2055]), .B(p_input[743]), .Z(n24221) );
  XNOR U23974 ( .A(n16741), .B(p_input[738]), .Z(n24198) );
  XNOR U23975 ( .A(n24212), .B(n24211), .Z(n24202) );
  XOR U23976 ( .A(n24222), .B(n24208), .Z(n24211) );
  XOR U23977 ( .A(p_input[2051]), .B(p_input[739]), .Z(n24208) );
  XNOR U23978 ( .A(p_input[2052]), .B(p_input[740]), .Z(n24222) );
  XOR U23979 ( .A(p_input[2053]), .B(p_input[741]), .Z(n24212) );
  XNOR U23980 ( .A(n24223), .B(n24224), .Z(n24119) );
  AND U23981 ( .A(n545), .B(n24225), .Z(n24224) );
  XNOR U23982 ( .A(n24226), .B(n24227), .Z(n545) );
  AND U23983 ( .A(n24228), .B(n24229), .Z(n24227) );
  XOR U23984 ( .A(n24226), .B(n24129), .Z(n24229) );
  XNOR U23985 ( .A(n24226), .B(n24083), .Z(n24228) );
  XOR U23986 ( .A(n24230), .B(n24231), .Z(n24226) );
  AND U23987 ( .A(n24232), .B(n24233), .Z(n24231) );
  XOR U23988 ( .A(n24230), .B(n24093), .Z(n24232) );
  XOR U23989 ( .A(n24234), .B(n24235), .Z(n24072) );
  AND U23990 ( .A(n549), .B(n24225), .Z(n24235) );
  XNOR U23991 ( .A(n24223), .B(n24234), .Z(n24225) );
  XNOR U23992 ( .A(n24236), .B(n24237), .Z(n549) );
  AND U23993 ( .A(n24238), .B(n24239), .Z(n24237) );
  XNOR U23994 ( .A(n24240), .B(n24236), .Z(n24239) );
  IV U23995 ( .A(n24129), .Z(n24240) );
  XNOR U23996 ( .A(n24241), .B(n24242), .Z(n24129) );
  AND U23997 ( .A(n552), .B(n24243), .Z(n24242) );
  XNOR U23998 ( .A(n24241), .B(n24244), .Z(n24243) );
  XNOR U23999 ( .A(n24083), .B(n24236), .Z(n24238) );
  XOR U24000 ( .A(n24245), .B(n24246), .Z(n24083) );
  AND U24001 ( .A(n560), .B(n24247), .Z(n24246) );
  XOR U24002 ( .A(n24230), .B(n24248), .Z(n24236) );
  AND U24003 ( .A(n24249), .B(n24233), .Z(n24248) );
  XNOR U24004 ( .A(n24142), .B(n24230), .Z(n24233) );
  XNOR U24005 ( .A(n24250), .B(n24251), .Z(n24142) );
  AND U24006 ( .A(n552), .B(n24252), .Z(n24251) );
  XOR U24007 ( .A(n24253), .B(n24250), .Z(n24252) );
  XNOR U24008 ( .A(n24254), .B(n24230), .Z(n24249) );
  IV U24009 ( .A(n24093), .Z(n24254) );
  XOR U24010 ( .A(n24255), .B(n24256), .Z(n24093) );
  AND U24011 ( .A(n560), .B(n24257), .Z(n24256) );
  XOR U24012 ( .A(n24258), .B(n24259), .Z(n24230) );
  AND U24013 ( .A(n24260), .B(n24261), .Z(n24259) );
  XNOR U24014 ( .A(n24167), .B(n24258), .Z(n24261) );
  XNOR U24015 ( .A(n24262), .B(n24263), .Z(n24167) );
  AND U24016 ( .A(n552), .B(n24264), .Z(n24263) );
  XNOR U24017 ( .A(n24265), .B(n24262), .Z(n24264) );
  XOR U24018 ( .A(n24258), .B(n24104), .Z(n24260) );
  XOR U24019 ( .A(n24266), .B(n24267), .Z(n24104) );
  AND U24020 ( .A(n560), .B(n24268), .Z(n24267) );
  XOR U24021 ( .A(n24269), .B(n24270), .Z(n24258) );
  AND U24022 ( .A(n24271), .B(n24272), .Z(n24270) );
  XNOR U24023 ( .A(n24269), .B(n24213), .Z(n24272) );
  XNOR U24024 ( .A(n24273), .B(n24274), .Z(n24213) );
  AND U24025 ( .A(n552), .B(n24275), .Z(n24274) );
  XOR U24026 ( .A(n24276), .B(n24273), .Z(n24275) );
  XNOR U24027 ( .A(n24277), .B(n24269), .Z(n24271) );
  IV U24028 ( .A(n24116), .Z(n24277) );
  XOR U24029 ( .A(n24278), .B(n24279), .Z(n24116) );
  AND U24030 ( .A(n560), .B(n24280), .Z(n24279) );
  AND U24031 ( .A(n24234), .B(n24223), .Z(n24269) );
  XNOR U24032 ( .A(n24281), .B(n24282), .Z(n24223) );
  AND U24033 ( .A(n552), .B(n24283), .Z(n24282) );
  XNOR U24034 ( .A(n24284), .B(n24281), .Z(n24283) );
  XNOR U24035 ( .A(n24285), .B(n24286), .Z(n552) );
  AND U24036 ( .A(n24287), .B(n24288), .Z(n24286) );
  XOR U24037 ( .A(n24244), .B(n24285), .Z(n24288) );
  AND U24038 ( .A(n24289), .B(n24290), .Z(n24244) );
  XOR U24039 ( .A(n24285), .B(n24241), .Z(n24287) );
  XNOR U24040 ( .A(n24291), .B(n24292), .Z(n24241) );
  AND U24041 ( .A(n556), .B(n24247), .Z(n24292) );
  XOR U24042 ( .A(n24245), .B(n24291), .Z(n24247) );
  XOR U24043 ( .A(n24293), .B(n24294), .Z(n24285) );
  AND U24044 ( .A(n24295), .B(n24296), .Z(n24294) );
  XNOR U24045 ( .A(n24293), .B(n24289), .Z(n24296) );
  IV U24046 ( .A(n24253), .Z(n24289) );
  XOR U24047 ( .A(n24297), .B(n24298), .Z(n24253) );
  XOR U24048 ( .A(n24299), .B(n24290), .Z(n24298) );
  AND U24049 ( .A(n24265), .B(n24300), .Z(n24290) );
  AND U24050 ( .A(n24301), .B(n24302), .Z(n24299) );
  XOR U24051 ( .A(n24303), .B(n24297), .Z(n24301) );
  XNOR U24052 ( .A(n24250), .B(n24293), .Z(n24295) );
  XNOR U24053 ( .A(n24304), .B(n24305), .Z(n24250) );
  AND U24054 ( .A(n556), .B(n24257), .Z(n24305) );
  XOR U24055 ( .A(n24304), .B(n24255), .Z(n24257) );
  XOR U24056 ( .A(n24306), .B(n24307), .Z(n24293) );
  AND U24057 ( .A(n24308), .B(n24309), .Z(n24307) );
  XNOR U24058 ( .A(n24306), .B(n24265), .Z(n24309) );
  XOR U24059 ( .A(n24310), .B(n24302), .Z(n24265) );
  XNOR U24060 ( .A(n24311), .B(n24297), .Z(n24302) );
  XOR U24061 ( .A(n24312), .B(n24313), .Z(n24297) );
  AND U24062 ( .A(n24314), .B(n24315), .Z(n24313) );
  XOR U24063 ( .A(n24316), .B(n24312), .Z(n24314) );
  XNOR U24064 ( .A(n24317), .B(n24318), .Z(n24311) );
  AND U24065 ( .A(n24319), .B(n24320), .Z(n24318) );
  XOR U24066 ( .A(n24317), .B(n24321), .Z(n24319) );
  XNOR U24067 ( .A(n24303), .B(n24300), .Z(n24310) );
  AND U24068 ( .A(n24322), .B(n24323), .Z(n24300) );
  XOR U24069 ( .A(n24324), .B(n24325), .Z(n24303) );
  AND U24070 ( .A(n24326), .B(n24327), .Z(n24325) );
  XOR U24071 ( .A(n24324), .B(n24328), .Z(n24326) );
  XNOR U24072 ( .A(n24262), .B(n24306), .Z(n24308) );
  XNOR U24073 ( .A(n24329), .B(n24330), .Z(n24262) );
  AND U24074 ( .A(n556), .B(n24268), .Z(n24330) );
  XOR U24075 ( .A(n24329), .B(n24266), .Z(n24268) );
  XOR U24076 ( .A(n24331), .B(n24332), .Z(n24306) );
  AND U24077 ( .A(n24333), .B(n24334), .Z(n24332) );
  XNOR U24078 ( .A(n24331), .B(n24322), .Z(n24334) );
  IV U24079 ( .A(n24276), .Z(n24322) );
  XNOR U24080 ( .A(n24335), .B(n24315), .Z(n24276) );
  XNOR U24081 ( .A(n24336), .B(n24321), .Z(n24315) );
  XOR U24082 ( .A(n24337), .B(n24338), .Z(n24321) );
  NOR U24083 ( .A(n24339), .B(n24340), .Z(n24338) );
  XNOR U24084 ( .A(n24337), .B(n24341), .Z(n24339) );
  XNOR U24085 ( .A(n24320), .B(n24312), .Z(n24336) );
  XOR U24086 ( .A(n24342), .B(n24343), .Z(n24312) );
  AND U24087 ( .A(n24344), .B(n24345), .Z(n24343) );
  XNOR U24088 ( .A(n24342), .B(n24346), .Z(n24344) );
  XNOR U24089 ( .A(n24347), .B(n24317), .Z(n24320) );
  XOR U24090 ( .A(n24348), .B(n24349), .Z(n24317) );
  AND U24091 ( .A(n24350), .B(n24351), .Z(n24349) );
  XOR U24092 ( .A(n24348), .B(n24352), .Z(n24350) );
  XNOR U24093 ( .A(n24353), .B(n24354), .Z(n24347) );
  NOR U24094 ( .A(n24355), .B(n24356), .Z(n24354) );
  XOR U24095 ( .A(n24353), .B(n24357), .Z(n24355) );
  XNOR U24096 ( .A(n24316), .B(n24323), .Z(n24335) );
  NOR U24097 ( .A(n24284), .B(n24358), .Z(n24323) );
  XOR U24098 ( .A(n24328), .B(n24327), .Z(n24316) );
  XNOR U24099 ( .A(n24359), .B(n24324), .Z(n24327) );
  XOR U24100 ( .A(n24360), .B(n24361), .Z(n24324) );
  AND U24101 ( .A(n24362), .B(n24363), .Z(n24361) );
  XOR U24102 ( .A(n24360), .B(n24364), .Z(n24362) );
  XNOR U24103 ( .A(n24365), .B(n24366), .Z(n24359) );
  NOR U24104 ( .A(n24367), .B(n24368), .Z(n24366) );
  XNOR U24105 ( .A(n24365), .B(n24369), .Z(n24367) );
  XOR U24106 ( .A(n24370), .B(n24371), .Z(n24328) );
  NOR U24107 ( .A(n24372), .B(n24373), .Z(n24371) );
  XNOR U24108 ( .A(n24370), .B(n24374), .Z(n24372) );
  XNOR U24109 ( .A(n24273), .B(n24331), .Z(n24333) );
  XNOR U24110 ( .A(n24375), .B(n24376), .Z(n24273) );
  AND U24111 ( .A(n556), .B(n24280), .Z(n24376) );
  XOR U24112 ( .A(n24375), .B(n24278), .Z(n24280) );
  AND U24113 ( .A(n24281), .B(n24284), .Z(n24331) );
  XOR U24114 ( .A(n24377), .B(n24358), .Z(n24284) );
  XNOR U24115 ( .A(p_input[2048]), .B(p_input[752]), .Z(n24358) );
  XOR U24116 ( .A(n24346), .B(n24345), .Z(n24377) );
  XNOR U24117 ( .A(n24378), .B(n24352), .Z(n24345) );
  XNOR U24118 ( .A(n24341), .B(n24340), .Z(n24352) );
  XOR U24119 ( .A(n24379), .B(n24337), .Z(n24340) );
  XNOR U24120 ( .A(n16904), .B(p_input[762]), .Z(n24337) );
  XNOR U24121 ( .A(p_input[2059]), .B(p_input[763]), .Z(n24379) );
  XOR U24122 ( .A(p_input[2060]), .B(p_input[764]), .Z(n24341) );
  XNOR U24123 ( .A(n24351), .B(n24342), .Z(n24378) );
  XNOR U24124 ( .A(n17068), .B(p_input[753]), .Z(n24342) );
  XOR U24125 ( .A(n24380), .B(n24357), .Z(n24351) );
  XNOR U24126 ( .A(p_input[2063]), .B(p_input[767]), .Z(n24357) );
  XOR U24127 ( .A(n24348), .B(n24356), .Z(n24380) );
  XOR U24128 ( .A(n24381), .B(n24353), .Z(n24356) );
  XOR U24129 ( .A(p_input[2061]), .B(p_input[765]), .Z(n24353) );
  XNOR U24130 ( .A(p_input[2062]), .B(p_input[766]), .Z(n24381) );
  XNOR U24131 ( .A(n16738), .B(p_input[761]), .Z(n24348) );
  XNOR U24132 ( .A(n24364), .B(n24363), .Z(n24346) );
  XNOR U24133 ( .A(n24382), .B(n24369), .Z(n24363) );
  XOR U24134 ( .A(p_input[2056]), .B(p_input[760]), .Z(n24369) );
  XOR U24135 ( .A(n24360), .B(n24368), .Z(n24382) );
  XOR U24136 ( .A(n24383), .B(n24365), .Z(n24368) );
  XOR U24137 ( .A(p_input[2054]), .B(p_input[758]), .Z(n24365) );
  XNOR U24138 ( .A(p_input[2055]), .B(p_input[759]), .Z(n24383) );
  XNOR U24139 ( .A(n16741), .B(p_input[754]), .Z(n24360) );
  XNOR U24140 ( .A(n24374), .B(n24373), .Z(n24364) );
  XOR U24141 ( .A(n24384), .B(n24370), .Z(n24373) );
  XOR U24142 ( .A(p_input[2051]), .B(p_input[755]), .Z(n24370) );
  XNOR U24143 ( .A(p_input[2052]), .B(p_input[756]), .Z(n24384) );
  XOR U24144 ( .A(p_input[2053]), .B(p_input[757]), .Z(n24374) );
  XNOR U24145 ( .A(n24385), .B(n24386), .Z(n24281) );
  AND U24146 ( .A(n556), .B(n24387), .Z(n24386) );
  XNOR U24147 ( .A(n24388), .B(n24389), .Z(n556) );
  AND U24148 ( .A(n24390), .B(n24391), .Z(n24389) );
  XOR U24149 ( .A(n24388), .B(n24291), .Z(n24391) );
  XNOR U24150 ( .A(n24388), .B(n24245), .Z(n24390) );
  XOR U24151 ( .A(n24392), .B(n24393), .Z(n24388) );
  AND U24152 ( .A(n24394), .B(n24395), .Z(n24393) );
  XOR U24153 ( .A(n24392), .B(n24255), .Z(n24394) );
  XOR U24154 ( .A(n24396), .B(n24397), .Z(n24234) );
  AND U24155 ( .A(n560), .B(n24387), .Z(n24397) );
  XNOR U24156 ( .A(n24385), .B(n24396), .Z(n24387) );
  XNOR U24157 ( .A(n24398), .B(n24399), .Z(n560) );
  AND U24158 ( .A(n24400), .B(n24401), .Z(n24399) );
  XNOR U24159 ( .A(n24402), .B(n24398), .Z(n24401) );
  IV U24160 ( .A(n24291), .Z(n24402) );
  XNOR U24161 ( .A(n24403), .B(n24404), .Z(n24291) );
  AND U24162 ( .A(n563), .B(n24405), .Z(n24404) );
  XNOR U24163 ( .A(n24403), .B(n24406), .Z(n24405) );
  XNOR U24164 ( .A(n24245), .B(n24398), .Z(n24400) );
  XOR U24165 ( .A(n24407), .B(n24408), .Z(n24245) );
  AND U24166 ( .A(n571), .B(n24409), .Z(n24408) );
  XOR U24167 ( .A(n24392), .B(n24410), .Z(n24398) );
  AND U24168 ( .A(n24411), .B(n24395), .Z(n24410) );
  XNOR U24169 ( .A(n24304), .B(n24392), .Z(n24395) );
  XNOR U24170 ( .A(n24412), .B(n24413), .Z(n24304) );
  AND U24171 ( .A(n563), .B(n24414), .Z(n24413) );
  XOR U24172 ( .A(n24415), .B(n24412), .Z(n24414) );
  XNOR U24173 ( .A(n24416), .B(n24392), .Z(n24411) );
  IV U24174 ( .A(n24255), .Z(n24416) );
  XOR U24175 ( .A(n24417), .B(n24418), .Z(n24255) );
  AND U24176 ( .A(n571), .B(n24419), .Z(n24418) );
  XOR U24177 ( .A(n24420), .B(n24421), .Z(n24392) );
  AND U24178 ( .A(n24422), .B(n24423), .Z(n24421) );
  XNOR U24179 ( .A(n24329), .B(n24420), .Z(n24423) );
  XNOR U24180 ( .A(n24424), .B(n24425), .Z(n24329) );
  AND U24181 ( .A(n563), .B(n24426), .Z(n24425) );
  XNOR U24182 ( .A(n24427), .B(n24424), .Z(n24426) );
  XOR U24183 ( .A(n24420), .B(n24266), .Z(n24422) );
  XOR U24184 ( .A(n24428), .B(n24429), .Z(n24266) );
  AND U24185 ( .A(n571), .B(n24430), .Z(n24429) );
  XOR U24186 ( .A(n24431), .B(n24432), .Z(n24420) );
  AND U24187 ( .A(n24433), .B(n24434), .Z(n24432) );
  XNOR U24188 ( .A(n24431), .B(n24375), .Z(n24434) );
  XNOR U24189 ( .A(n24435), .B(n24436), .Z(n24375) );
  AND U24190 ( .A(n563), .B(n24437), .Z(n24436) );
  XOR U24191 ( .A(n24438), .B(n24435), .Z(n24437) );
  XNOR U24192 ( .A(n24439), .B(n24431), .Z(n24433) );
  IV U24193 ( .A(n24278), .Z(n24439) );
  XOR U24194 ( .A(n24440), .B(n24441), .Z(n24278) );
  AND U24195 ( .A(n571), .B(n24442), .Z(n24441) );
  AND U24196 ( .A(n24396), .B(n24385), .Z(n24431) );
  XNOR U24197 ( .A(n24443), .B(n24444), .Z(n24385) );
  AND U24198 ( .A(n563), .B(n24445), .Z(n24444) );
  XNOR U24199 ( .A(n24446), .B(n24443), .Z(n24445) );
  XNOR U24200 ( .A(n24447), .B(n24448), .Z(n563) );
  AND U24201 ( .A(n24449), .B(n24450), .Z(n24448) );
  XOR U24202 ( .A(n24406), .B(n24447), .Z(n24450) );
  AND U24203 ( .A(n24451), .B(n24452), .Z(n24406) );
  XOR U24204 ( .A(n24447), .B(n24403), .Z(n24449) );
  XNOR U24205 ( .A(n24453), .B(n24454), .Z(n24403) );
  AND U24206 ( .A(n567), .B(n24409), .Z(n24454) );
  XOR U24207 ( .A(n24407), .B(n24453), .Z(n24409) );
  XOR U24208 ( .A(n24455), .B(n24456), .Z(n24447) );
  AND U24209 ( .A(n24457), .B(n24458), .Z(n24456) );
  XNOR U24210 ( .A(n24455), .B(n24451), .Z(n24458) );
  IV U24211 ( .A(n24415), .Z(n24451) );
  XOR U24212 ( .A(n24459), .B(n24460), .Z(n24415) );
  XOR U24213 ( .A(n24461), .B(n24452), .Z(n24460) );
  AND U24214 ( .A(n24427), .B(n24462), .Z(n24452) );
  AND U24215 ( .A(n24463), .B(n24464), .Z(n24461) );
  XOR U24216 ( .A(n24465), .B(n24459), .Z(n24463) );
  XNOR U24217 ( .A(n24412), .B(n24455), .Z(n24457) );
  XNOR U24218 ( .A(n24466), .B(n24467), .Z(n24412) );
  AND U24219 ( .A(n567), .B(n24419), .Z(n24467) );
  XOR U24220 ( .A(n24466), .B(n24417), .Z(n24419) );
  XOR U24221 ( .A(n24468), .B(n24469), .Z(n24455) );
  AND U24222 ( .A(n24470), .B(n24471), .Z(n24469) );
  XNOR U24223 ( .A(n24468), .B(n24427), .Z(n24471) );
  XOR U24224 ( .A(n24472), .B(n24464), .Z(n24427) );
  XNOR U24225 ( .A(n24473), .B(n24459), .Z(n24464) );
  XOR U24226 ( .A(n24474), .B(n24475), .Z(n24459) );
  AND U24227 ( .A(n24476), .B(n24477), .Z(n24475) );
  XOR U24228 ( .A(n24478), .B(n24474), .Z(n24476) );
  XNOR U24229 ( .A(n24479), .B(n24480), .Z(n24473) );
  AND U24230 ( .A(n24481), .B(n24482), .Z(n24480) );
  XOR U24231 ( .A(n24479), .B(n24483), .Z(n24481) );
  XNOR U24232 ( .A(n24465), .B(n24462), .Z(n24472) );
  AND U24233 ( .A(n24484), .B(n24485), .Z(n24462) );
  XOR U24234 ( .A(n24486), .B(n24487), .Z(n24465) );
  AND U24235 ( .A(n24488), .B(n24489), .Z(n24487) );
  XOR U24236 ( .A(n24486), .B(n24490), .Z(n24488) );
  XNOR U24237 ( .A(n24424), .B(n24468), .Z(n24470) );
  XNOR U24238 ( .A(n24491), .B(n24492), .Z(n24424) );
  AND U24239 ( .A(n567), .B(n24430), .Z(n24492) );
  XOR U24240 ( .A(n24491), .B(n24428), .Z(n24430) );
  XOR U24241 ( .A(n24493), .B(n24494), .Z(n24468) );
  AND U24242 ( .A(n24495), .B(n24496), .Z(n24494) );
  XNOR U24243 ( .A(n24493), .B(n24484), .Z(n24496) );
  IV U24244 ( .A(n24438), .Z(n24484) );
  XNOR U24245 ( .A(n24497), .B(n24477), .Z(n24438) );
  XNOR U24246 ( .A(n24498), .B(n24483), .Z(n24477) );
  XOR U24247 ( .A(n24499), .B(n24500), .Z(n24483) );
  NOR U24248 ( .A(n24501), .B(n24502), .Z(n24500) );
  XNOR U24249 ( .A(n24499), .B(n24503), .Z(n24501) );
  XNOR U24250 ( .A(n24482), .B(n24474), .Z(n24498) );
  XOR U24251 ( .A(n24504), .B(n24505), .Z(n24474) );
  AND U24252 ( .A(n24506), .B(n24507), .Z(n24505) );
  XNOR U24253 ( .A(n24504), .B(n24508), .Z(n24506) );
  XNOR U24254 ( .A(n24509), .B(n24479), .Z(n24482) );
  XOR U24255 ( .A(n24510), .B(n24511), .Z(n24479) );
  AND U24256 ( .A(n24512), .B(n24513), .Z(n24511) );
  XOR U24257 ( .A(n24510), .B(n24514), .Z(n24512) );
  XNOR U24258 ( .A(n24515), .B(n24516), .Z(n24509) );
  NOR U24259 ( .A(n24517), .B(n24518), .Z(n24516) );
  XOR U24260 ( .A(n24515), .B(n24519), .Z(n24517) );
  XNOR U24261 ( .A(n24478), .B(n24485), .Z(n24497) );
  NOR U24262 ( .A(n24446), .B(n24520), .Z(n24485) );
  XOR U24263 ( .A(n24490), .B(n24489), .Z(n24478) );
  XNOR U24264 ( .A(n24521), .B(n24486), .Z(n24489) );
  XOR U24265 ( .A(n24522), .B(n24523), .Z(n24486) );
  AND U24266 ( .A(n24524), .B(n24525), .Z(n24523) );
  XOR U24267 ( .A(n24522), .B(n24526), .Z(n24524) );
  XNOR U24268 ( .A(n24527), .B(n24528), .Z(n24521) );
  NOR U24269 ( .A(n24529), .B(n24530), .Z(n24528) );
  XNOR U24270 ( .A(n24527), .B(n24531), .Z(n24529) );
  XOR U24271 ( .A(n24532), .B(n24533), .Z(n24490) );
  NOR U24272 ( .A(n24534), .B(n24535), .Z(n24533) );
  XNOR U24273 ( .A(n24532), .B(n24536), .Z(n24534) );
  XNOR U24274 ( .A(n24435), .B(n24493), .Z(n24495) );
  XNOR U24275 ( .A(n24537), .B(n24538), .Z(n24435) );
  AND U24276 ( .A(n567), .B(n24442), .Z(n24538) );
  XOR U24277 ( .A(n24537), .B(n24440), .Z(n24442) );
  AND U24278 ( .A(n24443), .B(n24446), .Z(n24493) );
  XOR U24279 ( .A(n24539), .B(n24520), .Z(n24446) );
  XNOR U24280 ( .A(p_input[2048]), .B(p_input[768]), .Z(n24520) );
  XOR U24281 ( .A(n24508), .B(n24507), .Z(n24539) );
  XNOR U24282 ( .A(n24540), .B(n24514), .Z(n24507) );
  XNOR U24283 ( .A(n24503), .B(n24502), .Z(n24514) );
  XOR U24284 ( .A(n24541), .B(n24499), .Z(n24502) );
  XNOR U24285 ( .A(n16904), .B(p_input[778]), .Z(n24499) );
  XNOR U24286 ( .A(p_input[2059]), .B(p_input[779]), .Z(n24541) );
  XOR U24287 ( .A(p_input[2060]), .B(p_input[780]), .Z(n24503) );
  XNOR U24288 ( .A(n24513), .B(n24504), .Z(n24540) );
  XNOR U24289 ( .A(n17068), .B(p_input[769]), .Z(n24504) );
  XOR U24290 ( .A(n24542), .B(n24519), .Z(n24513) );
  XNOR U24291 ( .A(p_input[2063]), .B(p_input[783]), .Z(n24519) );
  XOR U24292 ( .A(n24510), .B(n24518), .Z(n24542) );
  XOR U24293 ( .A(n24543), .B(n24515), .Z(n24518) );
  XOR U24294 ( .A(p_input[2061]), .B(p_input[781]), .Z(n24515) );
  XNOR U24295 ( .A(p_input[2062]), .B(p_input[782]), .Z(n24543) );
  XNOR U24296 ( .A(n16738), .B(p_input[777]), .Z(n24510) );
  XNOR U24297 ( .A(n24526), .B(n24525), .Z(n24508) );
  XNOR U24298 ( .A(n24544), .B(n24531), .Z(n24525) );
  XOR U24299 ( .A(p_input[2056]), .B(p_input[776]), .Z(n24531) );
  XOR U24300 ( .A(n24522), .B(n24530), .Z(n24544) );
  XOR U24301 ( .A(n24545), .B(n24527), .Z(n24530) );
  XOR U24302 ( .A(p_input[2054]), .B(p_input[774]), .Z(n24527) );
  XNOR U24303 ( .A(p_input[2055]), .B(p_input[775]), .Z(n24545) );
  XNOR U24304 ( .A(n16741), .B(p_input[770]), .Z(n24522) );
  XNOR U24305 ( .A(n24536), .B(n24535), .Z(n24526) );
  XOR U24306 ( .A(n24546), .B(n24532), .Z(n24535) );
  XOR U24307 ( .A(p_input[2051]), .B(p_input[771]), .Z(n24532) );
  XNOR U24308 ( .A(p_input[2052]), .B(p_input[772]), .Z(n24546) );
  XOR U24309 ( .A(p_input[2053]), .B(p_input[773]), .Z(n24536) );
  XNOR U24310 ( .A(n24547), .B(n24548), .Z(n24443) );
  AND U24311 ( .A(n567), .B(n24549), .Z(n24548) );
  XNOR U24312 ( .A(n24550), .B(n24551), .Z(n567) );
  AND U24313 ( .A(n24552), .B(n24553), .Z(n24551) );
  XOR U24314 ( .A(n24550), .B(n24453), .Z(n24553) );
  XNOR U24315 ( .A(n24550), .B(n24407), .Z(n24552) );
  XOR U24316 ( .A(n24554), .B(n24555), .Z(n24550) );
  AND U24317 ( .A(n24556), .B(n24557), .Z(n24555) );
  XOR U24318 ( .A(n24554), .B(n24417), .Z(n24556) );
  XOR U24319 ( .A(n24558), .B(n24559), .Z(n24396) );
  AND U24320 ( .A(n571), .B(n24549), .Z(n24559) );
  XNOR U24321 ( .A(n24547), .B(n24558), .Z(n24549) );
  XNOR U24322 ( .A(n24560), .B(n24561), .Z(n571) );
  AND U24323 ( .A(n24562), .B(n24563), .Z(n24561) );
  XNOR U24324 ( .A(n24564), .B(n24560), .Z(n24563) );
  IV U24325 ( .A(n24453), .Z(n24564) );
  XNOR U24326 ( .A(n24565), .B(n24566), .Z(n24453) );
  AND U24327 ( .A(n574), .B(n24567), .Z(n24566) );
  XNOR U24328 ( .A(n24565), .B(n24568), .Z(n24567) );
  XNOR U24329 ( .A(n24407), .B(n24560), .Z(n24562) );
  XOR U24330 ( .A(n24569), .B(n24570), .Z(n24407) );
  AND U24331 ( .A(n582), .B(n24571), .Z(n24570) );
  XOR U24332 ( .A(n24554), .B(n24572), .Z(n24560) );
  AND U24333 ( .A(n24573), .B(n24557), .Z(n24572) );
  XNOR U24334 ( .A(n24466), .B(n24554), .Z(n24557) );
  XNOR U24335 ( .A(n24574), .B(n24575), .Z(n24466) );
  AND U24336 ( .A(n574), .B(n24576), .Z(n24575) );
  XOR U24337 ( .A(n24577), .B(n24574), .Z(n24576) );
  XNOR U24338 ( .A(n24578), .B(n24554), .Z(n24573) );
  IV U24339 ( .A(n24417), .Z(n24578) );
  XOR U24340 ( .A(n24579), .B(n24580), .Z(n24417) );
  AND U24341 ( .A(n582), .B(n24581), .Z(n24580) );
  XOR U24342 ( .A(n24582), .B(n24583), .Z(n24554) );
  AND U24343 ( .A(n24584), .B(n24585), .Z(n24583) );
  XNOR U24344 ( .A(n24491), .B(n24582), .Z(n24585) );
  XNOR U24345 ( .A(n24586), .B(n24587), .Z(n24491) );
  AND U24346 ( .A(n574), .B(n24588), .Z(n24587) );
  XNOR U24347 ( .A(n24589), .B(n24586), .Z(n24588) );
  XOR U24348 ( .A(n24582), .B(n24428), .Z(n24584) );
  XOR U24349 ( .A(n24590), .B(n24591), .Z(n24428) );
  AND U24350 ( .A(n582), .B(n24592), .Z(n24591) );
  XOR U24351 ( .A(n24593), .B(n24594), .Z(n24582) );
  AND U24352 ( .A(n24595), .B(n24596), .Z(n24594) );
  XNOR U24353 ( .A(n24593), .B(n24537), .Z(n24596) );
  XNOR U24354 ( .A(n24597), .B(n24598), .Z(n24537) );
  AND U24355 ( .A(n574), .B(n24599), .Z(n24598) );
  XOR U24356 ( .A(n24600), .B(n24597), .Z(n24599) );
  XNOR U24357 ( .A(n24601), .B(n24593), .Z(n24595) );
  IV U24358 ( .A(n24440), .Z(n24601) );
  XOR U24359 ( .A(n24602), .B(n24603), .Z(n24440) );
  AND U24360 ( .A(n582), .B(n24604), .Z(n24603) );
  AND U24361 ( .A(n24558), .B(n24547), .Z(n24593) );
  XNOR U24362 ( .A(n24605), .B(n24606), .Z(n24547) );
  AND U24363 ( .A(n574), .B(n24607), .Z(n24606) );
  XNOR U24364 ( .A(n24608), .B(n24605), .Z(n24607) );
  XNOR U24365 ( .A(n24609), .B(n24610), .Z(n574) );
  AND U24366 ( .A(n24611), .B(n24612), .Z(n24610) );
  XOR U24367 ( .A(n24568), .B(n24609), .Z(n24612) );
  AND U24368 ( .A(n24613), .B(n24614), .Z(n24568) );
  XOR U24369 ( .A(n24609), .B(n24565), .Z(n24611) );
  XNOR U24370 ( .A(n24615), .B(n24616), .Z(n24565) );
  AND U24371 ( .A(n578), .B(n24571), .Z(n24616) );
  XOR U24372 ( .A(n24569), .B(n24615), .Z(n24571) );
  XOR U24373 ( .A(n24617), .B(n24618), .Z(n24609) );
  AND U24374 ( .A(n24619), .B(n24620), .Z(n24618) );
  XNOR U24375 ( .A(n24617), .B(n24613), .Z(n24620) );
  IV U24376 ( .A(n24577), .Z(n24613) );
  XOR U24377 ( .A(n24621), .B(n24622), .Z(n24577) );
  XOR U24378 ( .A(n24623), .B(n24614), .Z(n24622) );
  AND U24379 ( .A(n24589), .B(n24624), .Z(n24614) );
  AND U24380 ( .A(n24625), .B(n24626), .Z(n24623) );
  XOR U24381 ( .A(n24627), .B(n24621), .Z(n24625) );
  XNOR U24382 ( .A(n24574), .B(n24617), .Z(n24619) );
  XNOR U24383 ( .A(n24628), .B(n24629), .Z(n24574) );
  AND U24384 ( .A(n578), .B(n24581), .Z(n24629) );
  XOR U24385 ( .A(n24628), .B(n24579), .Z(n24581) );
  XOR U24386 ( .A(n24630), .B(n24631), .Z(n24617) );
  AND U24387 ( .A(n24632), .B(n24633), .Z(n24631) );
  XNOR U24388 ( .A(n24630), .B(n24589), .Z(n24633) );
  XOR U24389 ( .A(n24634), .B(n24626), .Z(n24589) );
  XNOR U24390 ( .A(n24635), .B(n24621), .Z(n24626) );
  XOR U24391 ( .A(n24636), .B(n24637), .Z(n24621) );
  AND U24392 ( .A(n24638), .B(n24639), .Z(n24637) );
  XOR U24393 ( .A(n24640), .B(n24636), .Z(n24638) );
  XNOR U24394 ( .A(n24641), .B(n24642), .Z(n24635) );
  AND U24395 ( .A(n24643), .B(n24644), .Z(n24642) );
  XOR U24396 ( .A(n24641), .B(n24645), .Z(n24643) );
  XNOR U24397 ( .A(n24627), .B(n24624), .Z(n24634) );
  AND U24398 ( .A(n24646), .B(n24647), .Z(n24624) );
  XOR U24399 ( .A(n24648), .B(n24649), .Z(n24627) );
  AND U24400 ( .A(n24650), .B(n24651), .Z(n24649) );
  XOR U24401 ( .A(n24648), .B(n24652), .Z(n24650) );
  XNOR U24402 ( .A(n24586), .B(n24630), .Z(n24632) );
  XNOR U24403 ( .A(n24653), .B(n24654), .Z(n24586) );
  AND U24404 ( .A(n578), .B(n24592), .Z(n24654) );
  XOR U24405 ( .A(n24653), .B(n24590), .Z(n24592) );
  XOR U24406 ( .A(n24655), .B(n24656), .Z(n24630) );
  AND U24407 ( .A(n24657), .B(n24658), .Z(n24656) );
  XNOR U24408 ( .A(n24655), .B(n24646), .Z(n24658) );
  IV U24409 ( .A(n24600), .Z(n24646) );
  XNOR U24410 ( .A(n24659), .B(n24639), .Z(n24600) );
  XNOR U24411 ( .A(n24660), .B(n24645), .Z(n24639) );
  XOR U24412 ( .A(n24661), .B(n24662), .Z(n24645) );
  NOR U24413 ( .A(n24663), .B(n24664), .Z(n24662) );
  XNOR U24414 ( .A(n24661), .B(n24665), .Z(n24663) );
  XNOR U24415 ( .A(n24644), .B(n24636), .Z(n24660) );
  XOR U24416 ( .A(n24666), .B(n24667), .Z(n24636) );
  AND U24417 ( .A(n24668), .B(n24669), .Z(n24667) );
  XNOR U24418 ( .A(n24666), .B(n24670), .Z(n24668) );
  XNOR U24419 ( .A(n24671), .B(n24641), .Z(n24644) );
  XOR U24420 ( .A(n24672), .B(n24673), .Z(n24641) );
  AND U24421 ( .A(n24674), .B(n24675), .Z(n24673) );
  XOR U24422 ( .A(n24672), .B(n24676), .Z(n24674) );
  XNOR U24423 ( .A(n24677), .B(n24678), .Z(n24671) );
  NOR U24424 ( .A(n24679), .B(n24680), .Z(n24678) );
  XOR U24425 ( .A(n24677), .B(n24681), .Z(n24679) );
  XNOR U24426 ( .A(n24640), .B(n24647), .Z(n24659) );
  NOR U24427 ( .A(n24608), .B(n24682), .Z(n24647) );
  XOR U24428 ( .A(n24652), .B(n24651), .Z(n24640) );
  XNOR U24429 ( .A(n24683), .B(n24648), .Z(n24651) );
  XOR U24430 ( .A(n24684), .B(n24685), .Z(n24648) );
  AND U24431 ( .A(n24686), .B(n24687), .Z(n24685) );
  XOR U24432 ( .A(n24684), .B(n24688), .Z(n24686) );
  XNOR U24433 ( .A(n24689), .B(n24690), .Z(n24683) );
  NOR U24434 ( .A(n24691), .B(n24692), .Z(n24690) );
  XNOR U24435 ( .A(n24689), .B(n24693), .Z(n24691) );
  XOR U24436 ( .A(n24694), .B(n24695), .Z(n24652) );
  NOR U24437 ( .A(n24696), .B(n24697), .Z(n24695) );
  XNOR U24438 ( .A(n24694), .B(n24698), .Z(n24696) );
  XNOR U24439 ( .A(n24597), .B(n24655), .Z(n24657) );
  XNOR U24440 ( .A(n24699), .B(n24700), .Z(n24597) );
  AND U24441 ( .A(n578), .B(n24604), .Z(n24700) );
  XOR U24442 ( .A(n24699), .B(n24602), .Z(n24604) );
  AND U24443 ( .A(n24605), .B(n24608), .Z(n24655) );
  XOR U24444 ( .A(n24701), .B(n24682), .Z(n24608) );
  XNOR U24445 ( .A(p_input[2048]), .B(p_input[784]), .Z(n24682) );
  XOR U24446 ( .A(n24670), .B(n24669), .Z(n24701) );
  XNOR U24447 ( .A(n24702), .B(n24676), .Z(n24669) );
  XNOR U24448 ( .A(n24665), .B(n24664), .Z(n24676) );
  XOR U24449 ( .A(n24703), .B(n24661), .Z(n24664) );
  XNOR U24450 ( .A(n16904), .B(p_input[794]), .Z(n24661) );
  XNOR U24451 ( .A(p_input[2059]), .B(p_input[795]), .Z(n24703) );
  XOR U24452 ( .A(p_input[2060]), .B(p_input[796]), .Z(n24665) );
  XNOR U24453 ( .A(n24675), .B(n24666), .Z(n24702) );
  XNOR U24454 ( .A(n17068), .B(p_input[785]), .Z(n24666) );
  XOR U24455 ( .A(n24704), .B(n24681), .Z(n24675) );
  XNOR U24456 ( .A(p_input[2063]), .B(p_input[799]), .Z(n24681) );
  XOR U24457 ( .A(n24672), .B(n24680), .Z(n24704) );
  XOR U24458 ( .A(n24705), .B(n24677), .Z(n24680) );
  XOR U24459 ( .A(p_input[2061]), .B(p_input[797]), .Z(n24677) );
  XNOR U24460 ( .A(p_input[2062]), .B(p_input[798]), .Z(n24705) );
  XNOR U24461 ( .A(n16738), .B(p_input[793]), .Z(n24672) );
  XNOR U24462 ( .A(n24688), .B(n24687), .Z(n24670) );
  XNOR U24463 ( .A(n24706), .B(n24693), .Z(n24687) );
  XOR U24464 ( .A(p_input[2056]), .B(p_input[792]), .Z(n24693) );
  XOR U24465 ( .A(n24684), .B(n24692), .Z(n24706) );
  XOR U24466 ( .A(n24707), .B(n24689), .Z(n24692) );
  XOR U24467 ( .A(p_input[2054]), .B(p_input[790]), .Z(n24689) );
  XNOR U24468 ( .A(p_input[2055]), .B(p_input[791]), .Z(n24707) );
  XNOR U24469 ( .A(n16741), .B(p_input[786]), .Z(n24684) );
  XNOR U24470 ( .A(n24698), .B(n24697), .Z(n24688) );
  XOR U24471 ( .A(n24708), .B(n24694), .Z(n24697) );
  XOR U24472 ( .A(p_input[2051]), .B(p_input[787]), .Z(n24694) );
  XNOR U24473 ( .A(p_input[2052]), .B(p_input[788]), .Z(n24708) );
  XOR U24474 ( .A(p_input[2053]), .B(p_input[789]), .Z(n24698) );
  XNOR U24475 ( .A(n24709), .B(n24710), .Z(n24605) );
  AND U24476 ( .A(n578), .B(n24711), .Z(n24710) );
  XNOR U24477 ( .A(n24712), .B(n24713), .Z(n578) );
  AND U24478 ( .A(n24714), .B(n24715), .Z(n24713) );
  XOR U24479 ( .A(n24712), .B(n24615), .Z(n24715) );
  XNOR U24480 ( .A(n24712), .B(n24569), .Z(n24714) );
  XOR U24481 ( .A(n24716), .B(n24717), .Z(n24712) );
  AND U24482 ( .A(n24718), .B(n24719), .Z(n24717) );
  XOR U24483 ( .A(n24716), .B(n24579), .Z(n24718) );
  XOR U24484 ( .A(n24720), .B(n24721), .Z(n24558) );
  AND U24485 ( .A(n582), .B(n24711), .Z(n24721) );
  XNOR U24486 ( .A(n24709), .B(n24720), .Z(n24711) );
  XNOR U24487 ( .A(n24722), .B(n24723), .Z(n582) );
  AND U24488 ( .A(n24724), .B(n24725), .Z(n24723) );
  XNOR U24489 ( .A(n24726), .B(n24722), .Z(n24725) );
  IV U24490 ( .A(n24615), .Z(n24726) );
  XNOR U24491 ( .A(n24727), .B(n24728), .Z(n24615) );
  AND U24492 ( .A(n585), .B(n24729), .Z(n24728) );
  XNOR U24493 ( .A(n24727), .B(n24730), .Z(n24729) );
  XNOR U24494 ( .A(n24569), .B(n24722), .Z(n24724) );
  XOR U24495 ( .A(n24731), .B(n24732), .Z(n24569) );
  AND U24496 ( .A(n593), .B(n24733), .Z(n24732) );
  XOR U24497 ( .A(n24716), .B(n24734), .Z(n24722) );
  AND U24498 ( .A(n24735), .B(n24719), .Z(n24734) );
  XNOR U24499 ( .A(n24628), .B(n24716), .Z(n24719) );
  XNOR U24500 ( .A(n24736), .B(n24737), .Z(n24628) );
  AND U24501 ( .A(n585), .B(n24738), .Z(n24737) );
  XOR U24502 ( .A(n24739), .B(n24736), .Z(n24738) );
  XNOR U24503 ( .A(n24740), .B(n24716), .Z(n24735) );
  IV U24504 ( .A(n24579), .Z(n24740) );
  XOR U24505 ( .A(n24741), .B(n24742), .Z(n24579) );
  AND U24506 ( .A(n593), .B(n24743), .Z(n24742) );
  XOR U24507 ( .A(n24744), .B(n24745), .Z(n24716) );
  AND U24508 ( .A(n24746), .B(n24747), .Z(n24745) );
  XNOR U24509 ( .A(n24653), .B(n24744), .Z(n24747) );
  XNOR U24510 ( .A(n24748), .B(n24749), .Z(n24653) );
  AND U24511 ( .A(n585), .B(n24750), .Z(n24749) );
  XNOR U24512 ( .A(n24751), .B(n24748), .Z(n24750) );
  XOR U24513 ( .A(n24744), .B(n24590), .Z(n24746) );
  XOR U24514 ( .A(n24752), .B(n24753), .Z(n24590) );
  AND U24515 ( .A(n593), .B(n24754), .Z(n24753) );
  XOR U24516 ( .A(n24755), .B(n24756), .Z(n24744) );
  AND U24517 ( .A(n24757), .B(n24758), .Z(n24756) );
  XNOR U24518 ( .A(n24755), .B(n24699), .Z(n24758) );
  XNOR U24519 ( .A(n24759), .B(n24760), .Z(n24699) );
  AND U24520 ( .A(n585), .B(n24761), .Z(n24760) );
  XOR U24521 ( .A(n24762), .B(n24759), .Z(n24761) );
  XNOR U24522 ( .A(n24763), .B(n24755), .Z(n24757) );
  IV U24523 ( .A(n24602), .Z(n24763) );
  XOR U24524 ( .A(n24764), .B(n24765), .Z(n24602) );
  AND U24525 ( .A(n593), .B(n24766), .Z(n24765) );
  AND U24526 ( .A(n24720), .B(n24709), .Z(n24755) );
  XNOR U24527 ( .A(n24767), .B(n24768), .Z(n24709) );
  AND U24528 ( .A(n585), .B(n24769), .Z(n24768) );
  XNOR U24529 ( .A(n24770), .B(n24767), .Z(n24769) );
  XNOR U24530 ( .A(n24771), .B(n24772), .Z(n585) );
  AND U24531 ( .A(n24773), .B(n24774), .Z(n24772) );
  XOR U24532 ( .A(n24730), .B(n24771), .Z(n24774) );
  AND U24533 ( .A(n24775), .B(n24776), .Z(n24730) );
  XOR U24534 ( .A(n24771), .B(n24727), .Z(n24773) );
  XNOR U24535 ( .A(n24777), .B(n24778), .Z(n24727) );
  AND U24536 ( .A(n589), .B(n24733), .Z(n24778) );
  XOR U24537 ( .A(n24731), .B(n24777), .Z(n24733) );
  XOR U24538 ( .A(n24779), .B(n24780), .Z(n24771) );
  AND U24539 ( .A(n24781), .B(n24782), .Z(n24780) );
  XNOR U24540 ( .A(n24779), .B(n24775), .Z(n24782) );
  IV U24541 ( .A(n24739), .Z(n24775) );
  XOR U24542 ( .A(n24783), .B(n24784), .Z(n24739) );
  XOR U24543 ( .A(n24785), .B(n24776), .Z(n24784) );
  AND U24544 ( .A(n24751), .B(n24786), .Z(n24776) );
  AND U24545 ( .A(n24787), .B(n24788), .Z(n24785) );
  XOR U24546 ( .A(n24789), .B(n24783), .Z(n24787) );
  XNOR U24547 ( .A(n24736), .B(n24779), .Z(n24781) );
  XNOR U24548 ( .A(n24790), .B(n24791), .Z(n24736) );
  AND U24549 ( .A(n589), .B(n24743), .Z(n24791) );
  XOR U24550 ( .A(n24790), .B(n24741), .Z(n24743) );
  XOR U24551 ( .A(n24792), .B(n24793), .Z(n24779) );
  AND U24552 ( .A(n24794), .B(n24795), .Z(n24793) );
  XNOR U24553 ( .A(n24792), .B(n24751), .Z(n24795) );
  XOR U24554 ( .A(n24796), .B(n24788), .Z(n24751) );
  XNOR U24555 ( .A(n24797), .B(n24783), .Z(n24788) );
  XOR U24556 ( .A(n24798), .B(n24799), .Z(n24783) );
  AND U24557 ( .A(n24800), .B(n24801), .Z(n24799) );
  XOR U24558 ( .A(n24802), .B(n24798), .Z(n24800) );
  XNOR U24559 ( .A(n24803), .B(n24804), .Z(n24797) );
  AND U24560 ( .A(n24805), .B(n24806), .Z(n24804) );
  XOR U24561 ( .A(n24803), .B(n24807), .Z(n24805) );
  XNOR U24562 ( .A(n24789), .B(n24786), .Z(n24796) );
  AND U24563 ( .A(n24808), .B(n24809), .Z(n24786) );
  XOR U24564 ( .A(n24810), .B(n24811), .Z(n24789) );
  AND U24565 ( .A(n24812), .B(n24813), .Z(n24811) );
  XOR U24566 ( .A(n24810), .B(n24814), .Z(n24812) );
  XNOR U24567 ( .A(n24748), .B(n24792), .Z(n24794) );
  XNOR U24568 ( .A(n24815), .B(n24816), .Z(n24748) );
  AND U24569 ( .A(n589), .B(n24754), .Z(n24816) );
  XOR U24570 ( .A(n24815), .B(n24752), .Z(n24754) );
  XOR U24571 ( .A(n24817), .B(n24818), .Z(n24792) );
  AND U24572 ( .A(n24819), .B(n24820), .Z(n24818) );
  XNOR U24573 ( .A(n24817), .B(n24808), .Z(n24820) );
  IV U24574 ( .A(n24762), .Z(n24808) );
  XNOR U24575 ( .A(n24821), .B(n24801), .Z(n24762) );
  XNOR U24576 ( .A(n24822), .B(n24807), .Z(n24801) );
  XOR U24577 ( .A(n24823), .B(n24824), .Z(n24807) );
  NOR U24578 ( .A(n24825), .B(n24826), .Z(n24824) );
  XNOR U24579 ( .A(n24823), .B(n24827), .Z(n24825) );
  XNOR U24580 ( .A(n24806), .B(n24798), .Z(n24822) );
  XOR U24581 ( .A(n24828), .B(n24829), .Z(n24798) );
  AND U24582 ( .A(n24830), .B(n24831), .Z(n24829) );
  XNOR U24583 ( .A(n24828), .B(n24832), .Z(n24830) );
  XNOR U24584 ( .A(n24833), .B(n24803), .Z(n24806) );
  XOR U24585 ( .A(n24834), .B(n24835), .Z(n24803) );
  AND U24586 ( .A(n24836), .B(n24837), .Z(n24835) );
  XOR U24587 ( .A(n24834), .B(n24838), .Z(n24836) );
  XNOR U24588 ( .A(n24839), .B(n24840), .Z(n24833) );
  NOR U24589 ( .A(n24841), .B(n24842), .Z(n24840) );
  XOR U24590 ( .A(n24839), .B(n24843), .Z(n24841) );
  XNOR U24591 ( .A(n24802), .B(n24809), .Z(n24821) );
  NOR U24592 ( .A(n24770), .B(n24844), .Z(n24809) );
  XOR U24593 ( .A(n24814), .B(n24813), .Z(n24802) );
  XNOR U24594 ( .A(n24845), .B(n24810), .Z(n24813) );
  XOR U24595 ( .A(n24846), .B(n24847), .Z(n24810) );
  AND U24596 ( .A(n24848), .B(n24849), .Z(n24847) );
  XOR U24597 ( .A(n24846), .B(n24850), .Z(n24848) );
  XNOR U24598 ( .A(n24851), .B(n24852), .Z(n24845) );
  NOR U24599 ( .A(n24853), .B(n24854), .Z(n24852) );
  XNOR U24600 ( .A(n24851), .B(n24855), .Z(n24853) );
  XOR U24601 ( .A(n24856), .B(n24857), .Z(n24814) );
  NOR U24602 ( .A(n24858), .B(n24859), .Z(n24857) );
  XNOR U24603 ( .A(n24856), .B(n24860), .Z(n24858) );
  XNOR U24604 ( .A(n24759), .B(n24817), .Z(n24819) );
  XNOR U24605 ( .A(n24861), .B(n24862), .Z(n24759) );
  AND U24606 ( .A(n589), .B(n24766), .Z(n24862) );
  XOR U24607 ( .A(n24861), .B(n24764), .Z(n24766) );
  AND U24608 ( .A(n24767), .B(n24770), .Z(n24817) );
  XOR U24609 ( .A(n24863), .B(n24844), .Z(n24770) );
  XNOR U24610 ( .A(p_input[2048]), .B(p_input[800]), .Z(n24844) );
  XOR U24611 ( .A(n24832), .B(n24831), .Z(n24863) );
  XNOR U24612 ( .A(n24864), .B(n24838), .Z(n24831) );
  XNOR U24613 ( .A(n24827), .B(n24826), .Z(n24838) );
  XOR U24614 ( .A(n24865), .B(n24823), .Z(n24826) );
  XNOR U24615 ( .A(n16904), .B(p_input[810]), .Z(n24823) );
  XNOR U24616 ( .A(p_input[2059]), .B(p_input[811]), .Z(n24865) );
  XOR U24617 ( .A(p_input[2060]), .B(p_input[812]), .Z(n24827) );
  XNOR U24618 ( .A(n24837), .B(n24828), .Z(n24864) );
  XNOR U24619 ( .A(n17068), .B(p_input[801]), .Z(n24828) );
  XOR U24620 ( .A(n24866), .B(n24843), .Z(n24837) );
  XNOR U24621 ( .A(p_input[2063]), .B(p_input[815]), .Z(n24843) );
  XOR U24622 ( .A(n24834), .B(n24842), .Z(n24866) );
  XOR U24623 ( .A(n24867), .B(n24839), .Z(n24842) );
  XOR U24624 ( .A(p_input[2061]), .B(p_input[813]), .Z(n24839) );
  XNOR U24625 ( .A(p_input[2062]), .B(p_input[814]), .Z(n24867) );
  XNOR U24626 ( .A(n16738), .B(p_input[809]), .Z(n24834) );
  XNOR U24627 ( .A(n24850), .B(n24849), .Z(n24832) );
  XNOR U24628 ( .A(n24868), .B(n24855), .Z(n24849) );
  XOR U24629 ( .A(p_input[2056]), .B(p_input[808]), .Z(n24855) );
  XOR U24630 ( .A(n24846), .B(n24854), .Z(n24868) );
  XOR U24631 ( .A(n24869), .B(n24851), .Z(n24854) );
  XOR U24632 ( .A(p_input[2054]), .B(p_input[806]), .Z(n24851) );
  XNOR U24633 ( .A(p_input[2055]), .B(p_input[807]), .Z(n24869) );
  XNOR U24634 ( .A(n16741), .B(p_input[802]), .Z(n24846) );
  XNOR U24635 ( .A(n24860), .B(n24859), .Z(n24850) );
  XOR U24636 ( .A(n24870), .B(n24856), .Z(n24859) );
  XOR U24637 ( .A(p_input[2051]), .B(p_input[803]), .Z(n24856) );
  XNOR U24638 ( .A(p_input[2052]), .B(p_input[804]), .Z(n24870) );
  XOR U24639 ( .A(p_input[2053]), .B(p_input[805]), .Z(n24860) );
  XNOR U24640 ( .A(n24871), .B(n24872), .Z(n24767) );
  AND U24641 ( .A(n589), .B(n24873), .Z(n24872) );
  XNOR U24642 ( .A(n24874), .B(n24875), .Z(n589) );
  AND U24643 ( .A(n24876), .B(n24877), .Z(n24875) );
  XOR U24644 ( .A(n24874), .B(n24777), .Z(n24877) );
  XNOR U24645 ( .A(n24874), .B(n24731), .Z(n24876) );
  XOR U24646 ( .A(n24878), .B(n24879), .Z(n24874) );
  AND U24647 ( .A(n24880), .B(n24881), .Z(n24879) );
  XOR U24648 ( .A(n24878), .B(n24741), .Z(n24880) );
  XOR U24649 ( .A(n24882), .B(n24883), .Z(n24720) );
  AND U24650 ( .A(n593), .B(n24873), .Z(n24883) );
  XNOR U24651 ( .A(n24871), .B(n24882), .Z(n24873) );
  XNOR U24652 ( .A(n24884), .B(n24885), .Z(n593) );
  AND U24653 ( .A(n24886), .B(n24887), .Z(n24885) );
  XNOR U24654 ( .A(n24888), .B(n24884), .Z(n24887) );
  IV U24655 ( .A(n24777), .Z(n24888) );
  XNOR U24656 ( .A(n24889), .B(n24890), .Z(n24777) );
  AND U24657 ( .A(n596), .B(n24891), .Z(n24890) );
  XNOR U24658 ( .A(n24889), .B(n24892), .Z(n24891) );
  XNOR U24659 ( .A(n24731), .B(n24884), .Z(n24886) );
  XOR U24660 ( .A(n24893), .B(n24894), .Z(n24731) );
  AND U24661 ( .A(n604), .B(n24895), .Z(n24894) );
  XOR U24662 ( .A(n24878), .B(n24896), .Z(n24884) );
  AND U24663 ( .A(n24897), .B(n24881), .Z(n24896) );
  XNOR U24664 ( .A(n24790), .B(n24878), .Z(n24881) );
  XNOR U24665 ( .A(n24898), .B(n24899), .Z(n24790) );
  AND U24666 ( .A(n596), .B(n24900), .Z(n24899) );
  XOR U24667 ( .A(n24901), .B(n24898), .Z(n24900) );
  XNOR U24668 ( .A(n24902), .B(n24878), .Z(n24897) );
  IV U24669 ( .A(n24741), .Z(n24902) );
  XOR U24670 ( .A(n24903), .B(n24904), .Z(n24741) );
  AND U24671 ( .A(n604), .B(n24905), .Z(n24904) );
  XOR U24672 ( .A(n24906), .B(n24907), .Z(n24878) );
  AND U24673 ( .A(n24908), .B(n24909), .Z(n24907) );
  XNOR U24674 ( .A(n24815), .B(n24906), .Z(n24909) );
  XNOR U24675 ( .A(n24910), .B(n24911), .Z(n24815) );
  AND U24676 ( .A(n596), .B(n24912), .Z(n24911) );
  XNOR U24677 ( .A(n24913), .B(n24910), .Z(n24912) );
  XOR U24678 ( .A(n24906), .B(n24752), .Z(n24908) );
  XOR U24679 ( .A(n24914), .B(n24915), .Z(n24752) );
  AND U24680 ( .A(n604), .B(n24916), .Z(n24915) );
  XOR U24681 ( .A(n24917), .B(n24918), .Z(n24906) );
  AND U24682 ( .A(n24919), .B(n24920), .Z(n24918) );
  XNOR U24683 ( .A(n24917), .B(n24861), .Z(n24920) );
  XNOR U24684 ( .A(n24921), .B(n24922), .Z(n24861) );
  AND U24685 ( .A(n596), .B(n24923), .Z(n24922) );
  XOR U24686 ( .A(n24924), .B(n24921), .Z(n24923) );
  XNOR U24687 ( .A(n24925), .B(n24917), .Z(n24919) );
  IV U24688 ( .A(n24764), .Z(n24925) );
  XOR U24689 ( .A(n24926), .B(n24927), .Z(n24764) );
  AND U24690 ( .A(n604), .B(n24928), .Z(n24927) );
  AND U24691 ( .A(n24882), .B(n24871), .Z(n24917) );
  XNOR U24692 ( .A(n24929), .B(n24930), .Z(n24871) );
  AND U24693 ( .A(n596), .B(n24931), .Z(n24930) );
  XNOR U24694 ( .A(n24932), .B(n24929), .Z(n24931) );
  XNOR U24695 ( .A(n24933), .B(n24934), .Z(n596) );
  AND U24696 ( .A(n24935), .B(n24936), .Z(n24934) );
  XOR U24697 ( .A(n24892), .B(n24933), .Z(n24936) );
  AND U24698 ( .A(n24937), .B(n24938), .Z(n24892) );
  XOR U24699 ( .A(n24933), .B(n24889), .Z(n24935) );
  XNOR U24700 ( .A(n24939), .B(n24940), .Z(n24889) );
  AND U24701 ( .A(n600), .B(n24895), .Z(n24940) );
  XOR U24702 ( .A(n24893), .B(n24939), .Z(n24895) );
  XOR U24703 ( .A(n24941), .B(n24942), .Z(n24933) );
  AND U24704 ( .A(n24943), .B(n24944), .Z(n24942) );
  XNOR U24705 ( .A(n24941), .B(n24937), .Z(n24944) );
  IV U24706 ( .A(n24901), .Z(n24937) );
  XOR U24707 ( .A(n24945), .B(n24946), .Z(n24901) );
  XOR U24708 ( .A(n24947), .B(n24938), .Z(n24946) );
  AND U24709 ( .A(n24913), .B(n24948), .Z(n24938) );
  AND U24710 ( .A(n24949), .B(n24950), .Z(n24947) );
  XOR U24711 ( .A(n24951), .B(n24945), .Z(n24949) );
  XNOR U24712 ( .A(n24898), .B(n24941), .Z(n24943) );
  XNOR U24713 ( .A(n24952), .B(n24953), .Z(n24898) );
  AND U24714 ( .A(n600), .B(n24905), .Z(n24953) );
  XOR U24715 ( .A(n24952), .B(n24903), .Z(n24905) );
  XOR U24716 ( .A(n24954), .B(n24955), .Z(n24941) );
  AND U24717 ( .A(n24956), .B(n24957), .Z(n24955) );
  XNOR U24718 ( .A(n24954), .B(n24913), .Z(n24957) );
  XOR U24719 ( .A(n24958), .B(n24950), .Z(n24913) );
  XNOR U24720 ( .A(n24959), .B(n24945), .Z(n24950) );
  XOR U24721 ( .A(n24960), .B(n24961), .Z(n24945) );
  AND U24722 ( .A(n24962), .B(n24963), .Z(n24961) );
  XOR U24723 ( .A(n24964), .B(n24960), .Z(n24962) );
  XNOR U24724 ( .A(n24965), .B(n24966), .Z(n24959) );
  AND U24725 ( .A(n24967), .B(n24968), .Z(n24966) );
  XOR U24726 ( .A(n24965), .B(n24969), .Z(n24967) );
  XNOR U24727 ( .A(n24951), .B(n24948), .Z(n24958) );
  AND U24728 ( .A(n24970), .B(n24971), .Z(n24948) );
  XOR U24729 ( .A(n24972), .B(n24973), .Z(n24951) );
  AND U24730 ( .A(n24974), .B(n24975), .Z(n24973) );
  XOR U24731 ( .A(n24972), .B(n24976), .Z(n24974) );
  XNOR U24732 ( .A(n24910), .B(n24954), .Z(n24956) );
  XNOR U24733 ( .A(n24977), .B(n24978), .Z(n24910) );
  AND U24734 ( .A(n600), .B(n24916), .Z(n24978) );
  XOR U24735 ( .A(n24977), .B(n24914), .Z(n24916) );
  XOR U24736 ( .A(n24979), .B(n24980), .Z(n24954) );
  AND U24737 ( .A(n24981), .B(n24982), .Z(n24980) );
  XNOR U24738 ( .A(n24979), .B(n24970), .Z(n24982) );
  IV U24739 ( .A(n24924), .Z(n24970) );
  XNOR U24740 ( .A(n24983), .B(n24963), .Z(n24924) );
  XNOR U24741 ( .A(n24984), .B(n24969), .Z(n24963) );
  XOR U24742 ( .A(n24985), .B(n24986), .Z(n24969) );
  NOR U24743 ( .A(n24987), .B(n24988), .Z(n24986) );
  XNOR U24744 ( .A(n24985), .B(n24989), .Z(n24987) );
  XNOR U24745 ( .A(n24968), .B(n24960), .Z(n24984) );
  XOR U24746 ( .A(n24990), .B(n24991), .Z(n24960) );
  AND U24747 ( .A(n24992), .B(n24993), .Z(n24991) );
  XNOR U24748 ( .A(n24990), .B(n24994), .Z(n24992) );
  XNOR U24749 ( .A(n24995), .B(n24965), .Z(n24968) );
  XOR U24750 ( .A(n24996), .B(n24997), .Z(n24965) );
  AND U24751 ( .A(n24998), .B(n24999), .Z(n24997) );
  XOR U24752 ( .A(n24996), .B(n25000), .Z(n24998) );
  XNOR U24753 ( .A(n25001), .B(n25002), .Z(n24995) );
  NOR U24754 ( .A(n25003), .B(n25004), .Z(n25002) );
  XOR U24755 ( .A(n25001), .B(n25005), .Z(n25003) );
  XNOR U24756 ( .A(n24964), .B(n24971), .Z(n24983) );
  NOR U24757 ( .A(n24932), .B(n25006), .Z(n24971) );
  XOR U24758 ( .A(n24976), .B(n24975), .Z(n24964) );
  XNOR U24759 ( .A(n25007), .B(n24972), .Z(n24975) );
  XOR U24760 ( .A(n25008), .B(n25009), .Z(n24972) );
  AND U24761 ( .A(n25010), .B(n25011), .Z(n25009) );
  XOR U24762 ( .A(n25008), .B(n25012), .Z(n25010) );
  XNOR U24763 ( .A(n25013), .B(n25014), .Z(n25007) );
  NOR U24764 ( .A(n25015), .B(n25016), .Z(n25014) );
  XNOR U24765 ( .A(n25013), .B(n25017), .Z(n25015) );
  XOR U24766 ( .A(n25018), .B(n25019), .Z(n24976) );
  NOR U24767 ( .A(n25020), .B(n25021), .Z(n25019) );
  XNOR U24768 ( .A(n25018), .B(n25022), .Z(n25020) );
  XNOR U24769 ( .A(n24921), .B(n24979), .Z(n24981) );
  XNOR U24770 ( .A(n25023), .B(n25024), .Z(n24921) );
  AND U24771 ( .A(n600), .B(n24928), .Z(n25024) );
  XOR U24772 ( .A(n25023), .B(n24926), .Z(n24928) );
  AND U24773 ( .A(n24929), .B(n24932), .Z(n24979) );
  XOR U24774 ( .A(n25025), .B(n25006), .Z(n24932) );
  XNOR U24775 ( .A(p_input[2048]), .B(p_input[816]), .Z(n25006) );
  XOR U24776 ( .A(n24994), .B(n24993), .Z(n25025) );
  XNOR U24777 ( .A(n25026), .B(n25000), .Z(n24993) );
  XNOR U24778 ( .A(n24989), .B(n24988), .Z(n25000) );
  XOR U24779 ( .A(n25027), .B(n24985), .Z(n24988) );
  XNOR U24780 ( .A(n16904), .B(p_input[826]), .Z(n24985) );
  XNOR U24781 ( .A(p_input[2059]), .B(p_input[827]), .Z(n25027) );
  XOR U24782 ( .A(p_input[2060]), .B(p_input[828]), .Z(n24989) );
  XNOR U24783 ( .A(n24999), .B(n24990), .Z(n25026) );
  XNOR U24784 ( .A(n17068), .B(p_input[817]), .Z(n24990) );
  XOR U24785 ( .A(n25028), .B(n25005), .Z(n24999) );
  XNOR U24786 ( .A(p_input[2063]), .B(p_input[831]), .Z(n25005) );
  XOR U24787 ( .A(n24996), .B(n25004), .Z(n25028) );
  XOR U24788 ( .A(n25029), .B(n25001), .Z(n25004) );
  XOR U24789 ( .A(p_input[2061]), .B(p_input[829]), .Z(n25001) );
  XNOR U24790 ( .A(p_input[2062]), .B(p_input[830]), .Z(n25029) );
  XNOR U24791 ( .A(n16738), .B(p_input[825]), .Z(n24996) );
  XNOR U24792 ( .A(n25012), .B(n25011), .Z(n24994) );
  XNOR U24793 ( .A(n25030), .B(n25017), .Z(n25011) );
  XOR U24794 ( .A(p_input[2056]), .B(p_input[824]), .Z(n25017) );
  XOR U24795 ( .A(n25008), .B(n25016), .Z(n25030) );
  XOR U24796 ( .A(n25031), .B(n25013), .Z(n25016) );
  XOR U24797 ( .A(p_input[2054]), .B(p_input[822]), .Z(n25013) );
  XNOR U24798 ( .A(p_input[2055]), .B(p_input[823]), .Z(n25031) );
  XNOR U24799 ( .A(n16741), .B(p_input[818]), .Z(n25008) );
  XNOR U24800 ( .A(n25022), .B(n25021), .Z(n25012) );
  XOR U24801 ( .A(n25032), .B(n25018), .Z(n25021) );
  XOR U24802 ( .A(p_input[2051]), .B(p_input[819]), .Z(n25018) );
  XNOR U24803 ( .A(p_input[2052]), .B(p_input[820]), .Z(n25032) );
  XOR U24804 ( .A(p_input[2053]), .B(p_input[821]), .Z(n25022) );
  XNOR U24805 ( .A(n25033), .B(n25034), .Z(n24929) );
  AND U24806 ( .A(n600), .B(n25035), .Z(n25034) );
  XNOR U24807 ( .A(n25036), .B(n25037), .Z(n600) );
  AND U24808 ( .A(n25038), .B(n25039), .Z(n25037) );
  XOR U24809 ( .A(n25036), .B(n24939), .Z(n25039) );
  XNOR U24810 ( .A(n25036), .B(n24893), .Z(n25038) );
  XOR U24811 ( .A(n25040), .B(n25041), .Z(n25036) );
  AND U24812 ( .A(n25042), .B(n25043), .Z(n25041) );
  XOR U24813 ( .A(n25040), .B(n24903), .Z(n25042) );
  XOR U24814 ( .A(n25044), .B(n25045), .Z(n24882) );
  AND U24815 ( .A(n604), .B(n25035), .Z(n25045) );
  XNOR U24816 ( .A(n25033), .B(n25044), .Z(n25035) );
  XNOR U24817 ( .A(n25046), .B(n25047), .Z(n604) );
  AND U24818 ( .A(n25048), .B(n25049), .Z(n25047) );
  XNOR U24819 ( .A(n25050), .B(n25046), .Z(n25049) );
  IV U24820 ( .A(n24939), .Z(n25050) );
  XNOR U24821 ( .A(n25051), .B(n25052), .Z(n24939) );
  AND U24822 ( .A(n607), .B(n25053), .Z(n25052) );
  XNOR U24823 ( .A(n25051), .B(n25054), .Z(n25053) );
  XNOR U24824 ( .A(n24893), .B(n25046), .Z(n25048) );
  XOR U24825 ( .A(n25055), .B(n25056), .Z(n24893) );
  AND U24826 ( .A(n615), .B(n25057), .Z(n25056) );
  XOR U24827 ( .A(n25040), .B(n25058), .Z(n25046) );
  AND U24828 ( .A(n25059), .B(n25043), .Z(n25058) );
  XNOR U24829 ( .A(n24952), .B(n25040), .Z(n25043) );
  XNOR U24830 ( .A(n25060), .B(n25061), .Z(n24952) );
  AND U24831 ( .A(n607), .B(n25062), .Z(n25061) );
  XOR U24832 ( .A(n25063), .B(n25060), .Z(n25062) );
  XNOR U24833 ( .A(n25064), .B(n25040), .Z(n25059) );
  IV U24834 ( .A(n24903), .Z(n25064) );
  XOR U24835 ( .A(n25065), .B(n25066), .Z(n24903) );
  AND U24836 ( .A(n615), .B(n25067), .Z(n25066) );
  XOR U24837 ( .A(n25068), .B(n25069), .Z(n25040) );
  AND U24838 ( .A(n25070), .B(n25071), .Z(n25069) );
  XNOR U24839 ( .A(n24977), .B(n25068), .Z(n25071) );
  XNOR U24840 ( .A(n25072), .B(n25073), .Z(n24977) );
  AND U24841 ( .A(n607), .B(n25074), .Z(n25073) );
  XNOR U24842 ( .A(n25075), .B(n25072), .Z(n25074) );
  XOR U24843 ( .A(n25068), .B(n24914), .Z(n25070) );
  XOR U24844 ( .A(n25076), .B(n25077), .Z(n24914) );
  AND U24845 ( .A(n615), .B(n25078), .Z(n25077) );
  XOR U24846 ( .A(n25079), .B(n25080), .Z(n25068) );
  AND U24847 ( .A(n25081), .B(n25082), .Z(n25080) );
  XNOR U24848 ( .A(n25079), .B(n25023), .Z(n25082) );
  XNOR U24849 ( .A(n25083), .B(n25084), .Z(n25023) );
  AND U24850 ( .A(n607), .B(n25085), .Z(n25084) );
  XOR U24851 ( .A(n25086), .B(n25083), .Z(n25085) );
  XNOR U24852 ( .A(n25087), .B(n25079), .Z(n25081) );
  IV U24853 ( .A(n24926), .Z(n25087) );
  XOR U24854 ( .A(n25088), .B(n25089), .Z(n24926) );
  AND U24855 ( .A(n615), .B(n25090), .Z(n25089) );
  AND U24856 ( .A(n25044), .B(n25033), .Z(n25079) );
  XNOR U24857 ( .A(n25091), .B(n25092), .Z(n25033) );
  AND U24858 ( .A(n607), .B(n25093), .Z(n25092) );
  XNOR U24859 ( .A(n25094), .B(n25091), .Z(n25093) );
  XNOR U24860 ( .A(n25095), .B(n25096), .Z(n607) );
  AND U24861 ( .A(n25097), .B(n25098), .Z(n25096) );
  XOR U24862 ( .A(n25054), .B(n25095), .Z(n25098) );
  AND U24863 ( .A(n25099), .B(n25100), .Z(n25054) );
  XOR U24864 ( .A(n25095), .B(n25051), .Z(n25097) );
  XNOR U24865 ( .A(n25101), .B(n25102), .Z(n25051) );
  AND U24866 ( .A(n611), .B(n25057), .Z(n25102) );
  XOR U24867 ( .A(n25055), .B(n25101), .Z(n25057) );
  XOR U24868 ( .A(n25103), .B(n25104), .Z(n25095) );
  AND U24869 ( .A(n25105), .B(n25106), .Z(n25104) );
  XNOR U24870 ( .A(n25103), .B(n25099), .Z(n25106) );
  IV U24871 ( .A(n25063), .Z(n25099) );
  XOR U24872 ( .A(n25107), .B(n25108), .Z(n25063) );
  XOR U24873 ( .A(n25109), .B(n25100), .Z(n25108) );
  AND U24874 ( .A(n25075), .B(n25110), .Z(n25100) );
  AND U24875 ( .A(n25111), .B(n25112), .Z(n25109) );
  XOR U24876 ( .A(n25113), .B(n25107), .Z(n25111) );
  XNOR U24877 ( .A(n25060), .B(n25103), .Z(n25105) );
  XNOR U24878 ( .A(n25114), .B(n25115), .Z(n25060) );
  AND U24879 ( .A(n611), .B(n25067), .Z(n25115) );
  XOR U24880 ( .A(n25114), .B(n25065), .Z(n25067) );
  XOR U24881 ( .A(n25116), .B(n25117), .Z(n25103) );
  AND U24882 ( .A(n25118), .B(n25119), .Z(n25117) );
  XNOR U24883 ( .A(n25116), .B(n25075), .Z(n25119) );
  XOR U24884 ( .A(n25120), .B(n25112), .Z(n25075) );
  XNOR U24885 ( .A(n25121), .B(n25107), .Z(n25112) );
  XOR U24886 ( .A(n25122), .B(n25123), .Z(n25107) );
  AND U24887 ( .A(n25124), .B(n25125), .Z(n25123) );
  XOR U24888 ( .A(n25126), .B(n25122), .Z(n25124) );
  XNOR U24889 ( .A(n25127), .B(n25128), .Z(n25121) );
  AND U24890 ( .A(n25129), .B(n25130), .Z(n25128) );
  XOR U24891 ( .A(n25127), .B(n25131), .Z(n25129) );
  XNOR U24892 ( .A(n25113), .B(n25110), .Z(n25120) );
  AND U24893 ( .A(n25132), .B(n25133), .Z(n25110) );
  XOR U24894 ( .A(n25134), .B(n25135), .Z(n25113) );
  AND U24895 ( .A(n25136), .B(n25137), .Z(n25135) );
  XOR U24896 ( .A(n25134), .B(n25138), .Z(n25136) );
  XNOR U24897 ( .A(n25072), .B(n25116), .Z(n25118) );
  XNOR U24898 ( .A(n25139), .B(n25140), .Z(n25072) );
  AND U24899 ( .A(n611), .B(n25078), .Z(n25140) );
  XOR U24900 ( .A(n25139), .B(n25076), .Z(n25078) );
  XOR U24901 ( .A(n25141), .B(n25142), .Z(n25116) );
  AND U24902 ( .A(n25143), .B(n25144), .Z(n25142) );
  XNOR U24903 ( .A(n25141), .B(n25132), .Z(n25144) );
  IV U24904 ( .A(n25086), .Z(n25132) );
  XNOR U24905 ( .A(n25145), .B(n25125), .Z(n25086) );
  XNOR U24906 ( .A(n25146), .B(n25131), .Z(n25125) );
  XOR U24907 ( .A(n25147), .B(n25148), .Z(n25131) );
  NOR U24908 ( .A(n25149), .B(n25150), .Z(n25148) );
  XNOR U24909 ( .A(n25147), .B(n25151), .Z(n25149) );
  XNOR U24910 ( .A(n25130), .B(n25122), .Z(n25146) );
  XOR U24911 ( .A(n25152), .B(n25153), .Z(n25122) );
  AND U24912 ( .A(n25154), .B(n25155), .Z(n25153) );
  XNOR U24913 ( .A(n25152), .B(n25156), .Z(n25154) );
  XNOR U24914 ( .A(n25157), .B(n25127), .Z(n25130) );
  XOR U24915 ( .A(n25158), .B(n25159), .Z(n25127) );
  AND U24916 ( .A(n25160), .B(n25161), .Z(n25159) );
  XOR U24917 ( .A(n25158), .B(n25162), .Z(n25160) );
  XNOR U24918 ( .A(n25163), .B(n25164), .Z(n25157) );
  NOR U24919 ( .A(n25165), .B(n25166), .Z(n25164) );
  XOR U24920 ( .A(n25163), .B(n25167), .Z(n25165) );
  XNOR U24921 ( .A(n25126), .B(n25133), .Z(n25145) );
  NOR U24922 ( .A(n25094), .B(n25168), .Z(n25133) );
  XOR U24923 ( .A(n25138), .B(n25137), .Z(n25126) );
  XNOR U24924 ( .A(n25169), .B(n25134), .Z(n25137) );
  XOR U24925 ( .A(n25170), .B(n25171), .Z(n25134) );
  AND U24926 ( .A(n25172), .B(n25173), .Z(n25171) );
  XOR U24927 ( .A(n25170), .B(n25174), .Z(n25172) );
  XNOR U24928 ( .A(n25175), .B(n25176), .Z(n25169) );
  NOR U24929 ( .A(n25177), .B(n25178), .Z(n25176) );
  XNOR U24930 ( .A(n25175), .B(n25179), .Z(n25177) );
  XOR U24931 ( .A(n25180), .B(n25181), .Z(n25138) );
  NOR U24932 ( .A(n25182), .B(n25183), .Z(n25181) );
  XNOR U24933 ( .A(n25180), .B(n25184), .Z(n25182) );
  XNOR U24934 ( .A(n25083), .B(n25141), .Z(n25143) );
  XNOR U24935 ( .A(n25185), .B(n25186), .Z(n25083) );
  AND U24936 ( .A(n611), .B(n25090), .Z(n25186) );
  XOR U24937 ( .A(n25185), .B(n25088), .Z(n25090) );
  AND U24938 ( .A(n25091), .B(n25094), .Z(n25141) );
  XOR U24939 ( .A(n25187), .B(n25168), .Z(n25094) );
  XNOR U24940 ( .A(p_input[2048]), .B(p_input[832]), .Z(n25168) );
  XOR U24941 ( .A(n25156), .B(n25155), .Z(n25187) );
  XNOR U24942 ( .A(n25188), .B(n25162), .Z(n25155) );
  XNOR U24943 ( .A(n25151), .B(n25150), .Z(n25162) );
  XOR U24944 ( .A(n25189), .B(n25147), .Z(n25150) );
  XNOR U24945 ( .A(n16904), .B(p_input[842]), .Z(n25147) );
  XNOR U24946 ( .A(p_input[2059]), .B(p_input[843]), .Z(n25189) );
  XOR U24947 ( .A(p_input[2060]), .B(p_input[844]), .Z(n25151) );
  XNOR U24948 ( .A(n25161), .B(n25152), .Z(n25188) );
  XNOR U24949 ( .A(n17068), .B(p_input[833]), .Z(n25152) );
  XOR U24950 ( .A(n25190), .B(n25167), .Z(n25161) );
  XNOR U24951 ( .A(p_input[2063]), .B(p_input[847]), .Z(n25167) );
  XOR U24952 ( .A(n25158), .B(n25166), .Z(n25190) );
  XOR U24953 ( .A(n25191), .B(n25163), .Z(n25166) );
  XOR U24954 ( .A(p_input[2061]), .B(p_input[845]), .Z(n25163) );
  XNOR U24955 ( .A(p_input[2062]), .B(p_input[846]), .Z(n25191) );
  XNOR U24956 ( .A(n16738), .B(p_input[841]), .Z(n25158) );
  XNOR U24957 ( .A(n25174), .B(n25173), .Z(n25156) );
  XNOR U24958 ( .A(n25192), .B(n25179), .Z(n25173) );
  XOR U24959 ( .A(p_input[2056]), .B(p_input[840]), .Z(n25179) );
  XOR U24960 ( .A(n25170), .B(n25178), .Z(n25192) );
  XOR U24961 ( .A(n25193), .B(n25175), .Z(n25178) );
  XOR U24962 ( .A(p_input[2054]), .B(p_input[838]), .Z(n25175) );
  XNOR U24963 ( .A(p_input[2055]), .B(p_input[839]), .Z(n25193) );
  XNOR U24964 ( .A(n16741), .B(p_input[834]), .Z(n25170) );
  XNOR U24965 ( .A(n25184), .B(n25183), .Z(n25174) );
  XOR U24966 ( .A(n25194), .B(n25180), .Z(n25183) );
  XOR U24967 ( .A(p_input[2051]), .B(p_input[835]), .Z(n25180) );
  XNOR U24968 ( .A(p_input[2052]), .B(p_input[836]), .Z(n25194) );
  XOR U24969 ( .A(p_input[2053]), .B(p_input[837]), .Z(n25184) );
  XNOR U24970 ( .A(n25195), .B(n25196), .Z(n25091) );
  AND U24971 ( .A(n611), .B(n25197), .Z(n25196) );
  XNOR U24972 ( .A(n25198), .B(n25199), .Z(n611) );
  AND U24973 ( .A(n25200), .B(n25201), .Z(n25199) );
  XOR U24974 ( .A(n25198), .B(n25101), .Z(n25201) );
  XNOR U24975 ( .A(n25198), .B(n25055), .Z(n25200) );
  XOR U24976 ( .A(n25202), .B(n25203), .Z(n25198) );
  AND U24977 ( .A(n25204), .B(n25205), .Z(n25203) );
  XOR U24978 ( .A(n25202), .B(n25065), .Z(n25204) );
  XOR U24979 ( .A(n25206), .B(n25207), .Z(n25044) );
  AND U24980 ( .A(n615), .B(n25197), .Z(n25207) );
  XNOR U24981 ( .A(n25195), .B(n25206), .Z(n25197) );
  XNOR U24982 ( .A(n25208), .B(n25209), .Z(n615) );
  AND U24983 ( .A(n25210), .B(n25211), .Z(n25209) );
  XNOR U24984 ( .A(n25212), .B(n25208), .Z(n25211) );
  IV U24985 ( .A(n25101), .Z(n25212) );
  XNOR U24986 ( .A(n25213), .B(n25214), .Z(n25101) );
  AND U24987 ( .A(n618), .B(n25215), .Z(n25214) );
  XNOR U24988 ( .A(n25213), .B(n25216), .Z(n25215) );
  XNOR U24989 ( .A(n25055), .B(n25208), .Z(n25210) );
  XOR U24990 ( .A(n25217), .B(n25218), .Z(n25055) );
  AND U24991 ( .A(n626), .B(n25219), .Z(n25218) );
  XOR U24992 ( .A(n25202), .B(n25220), .Z(n25208) );
  AND U24993 ( .A(n25221), .B(n25205), .Z(n25220) );
  XNOR U24994 ( .A(n25114), .B(n25202), .Z(n25205) );
  XNOR U24995 ( .A(n25222), .B(n25223), .Z(n25114) );
  AND U24996 ( .A(n618), .B(n25224), .Z(n25223) );
  XOR U24997 ( .A(n25225), .B(n25222), .Z(n25224) );
  XNOR U24998 ( .A(n25226), .B(n25202), .Z(n25221) );
  IV U24999 ( .A(n25065), .Z(n25226) );
  XOR U25000 ( .A(n25227), .B(n25228), .Z(n25065) );
  AND U25001 ( .A(n626), .B(n25229), .Z(n25228) );
  XOR U25002 ( .A(n25230), .B(n25231), .Z(n25202) );
  AND U25003 ( .A(n25232), .B(n25233), .Z(n25231) );
  XNOR U25004 ( .A(n25139), .B(n25230), .Z(n25233) );
  XNOR U25005 ( .A(n25234), .B(n25235), .Z(n25139) );
  AND U25006 ( .A(n618), .B(n25236), .Z(n25235) );
  XNOR U25007 ( .A(n25237), .B(n25234), .Z(n25236) );
  XOR U25008 ( .A(n25230), .B(n25076), .Z(n25232) );
  XOR U25009 ( .A(n25238), .B(n25239), .Z(n25076) );
  AND U25010 ( .A(n626), .B(n25240), .Z(n25239) );
  XOR U25011 ( .A(n25241), .B(n25242), .Z(n25230) );
  AND U25012 ( .A(n25243), .B(n25244), .Z(n25242) );
  XNOR U25013 ( .A(n25241), .B(n25185), .Z(n25244) );
  XNOR U25014 ( .A(n25245), .B(n25246), .Z(n25185) );
  AND U25015 ( .A(n618), .B(n25247), .Z(n25246) );
  XOR U25016 ( .A(n25248), .B(n25245), .Z(n25247) );
  XNOR U25017 ( .A(n25249), .B(n25241), .Z(n25243) );
  IV U25018 ( .A(n25088), .Z(n25249) );
  XOR U25019 ( .A(n25250), .B(n25251), .Z(n25088) );
  AND U25020 ( .A(n626), .B(n25252), .Z(n25251) );
  AND U25021 ( .A(n25206), .B(n25195), .Z(n25241) );
  XNOR U25022 ( .A(n25253), .B(n25254), .Z(n25195) );
  AND U25023 ( .A(n618), .B(n25255), .Z(n25254) );
  XNOR U25024 ( .A(n25256), .B(n25253), .Z(n25255) );
  XNOR U25025 ( .A(n25257), .B(n25258), .Z(n618) );
  AND U25026 ( .A(n25259), .B(n25260), .Z(n25258) );
  XOR U25027 ( .A(n25216), .B(n25257), .Z(n25260) );
  AND U25028 ( .A(n25261), .B(n25262), .Z(n25216) );
  XOR U25029 ( .A(n25257), .B(n25213), .Z(n25259) );
  XNOR U25030 ( .A(n25263), .B(n25264), .Z(n25213) );
  AND U25031 ( .A(n622), .B(n25219), .Z(n25264) );
  XOR U25032 ( .A(n25217), .B(n25263), .Z(n25219) );
  XOR U25033 ( .A(n25265), .B(n25266), .Z(n25257) );
  AND U25034 ( .A(n25267), .B(n25268), .Z(n25266) );
  XNOR U25035 ( .A(n25265), .B(n25261), .Z(n25268) );
  IV U25036 ( .A(n25225), .Z(n25261) );
  XOR U25037 ( .A(n25269), .B(n25270), .Z(n25225) );
  XOR U25038 ( .A(n25271), .B(n25262), .Z(n25270) );
  AND U25039 ( .A(n25237), .B(n25272), .Z(n25262) );
  AND U25040 ( .A(n25273), .B(n25274), .Z(n25271) );
  XOR U25041 ( .A(n25275), .B(n25269), .Z(n25273) );
  XNOR U25042 ( .A(n25222), .B(n25265), .Z(n25267) );
  XNOR U25043 ( .A(n25276), .B(n25277), .Z(n25222) );
  AND U25044 ( .A(n622), .B(n25229), .Z(n25277) );
  XOR U25045 ( .A(n25276), .B(n25227), .Z(n25229) );
  XOR U25046 ( .A(n25278), .B(n25279), .Z(n25265) );
  AND U25047 ( .A(n25280), .B(n25281), .Z(n25279) );
  XNOR U25048 ( .A(n25278), .B(n25237), .Z(n25281) );
  XOR U25049 ( .A(n25282), .B(n25274), .Z(n25237) );
  XNOR U25050 ( .A(n25283), .B(n25269), .Z(n25274) );
  XOR U25051 ( .A(n25284), .B(n25285), .Z(n25269) );
  AND U25052 ( .A(n25286), .B(n25287), .Z(n25285) );
  XOR U25053 ( .A(n25288), .B(n25284), .Z(n25286) );
  XNOR U25054 ( .A(n25289), .B(n25290), .Z(n25283) );
  AND U25055 ( .A(n25291), .B(n25292), .Z(n25290) );
  XOR U25056 ( .A(n25289), .B(n25293), .Z(n25291) );
  XNOR U25057 ( .A(n25275), .B(n25272), .Z(n25282) );
  AND U25058 ( .A(n25294), .B(n25295), .Z(n25272) );
  XOR U25059 ( .A(n25296), .B(n25297), .Z(n25275) );
  AND U25060 ( .A(n25298), .B(n25299), .Z(n25297) );
  XOR U25061 ( .A(n25296), .B(n25300), .Z(n25298) );
  XNOR U25062 ( .A(n25234), .B(n25278), .Z(n25280) );
  XNOR U25063 ( .A(n25301), .B(n25302), .Z(n25234) );
  AND U25064 ( .A(n622), .B(n25240), .Z(n25302) );
  XOR U25065 ( .A(n25301), .B(n25238), .Z(n25240) );
  XOR U25066 ( .A(n25303), .B(n25304), .Z(n25278) );
  AND U25067 ( .A(n25305), .B(n25306), .Z(n25304) );
  XNOR U25068 ( .A(n25303), .B(n25294), .Z(n25306) );
  IV U25069 ( .A(n25248), .Z(n25294) );
  XNOR U25070 ( .A(n25307), .B(n25287), .Z(n25248) );
  XNOR U25071 ( .A(n25308), .B(n25293), .Z(n25287) );
  XOR U25072 ( .A(n25309), .B(n25310), .Z(n25293) );
  NOR U25073 ( .A(n25311), .B(n25312), .Z(n25310) );
  XNOR U25074 ( .A(n25309), .B(n25313), .Z(n25311) );
  XNOR U25075 ( .A(n25292), .B(n25284), .Z(n25308) );
  XOR U25076 ( .A(n25314), .B(n25315), .Z(n25284) );
  AND U25077 ( .A(n25316), .B(n25317), .Z(n25315) );
  XNOR U25078 ( .A(n25314), .B(n25318), .Z(n25316) );
  XNOR U25079 ( .A(n25319), .B(n25289), .Z(n25292) );
  XOR U25080 ( .A(n25320), .B(n25321), .Z(n25289) );
  AND U25081 ( .A(n25322), .B(n25323), .Z(n25321) );
  XOR U25082 ( .A(n25320), .B(n25324), .Z(n25322) );
  XNOR U25083 ( .A(n25325), .B(n25326), .Z(n25319) );
  NOR U25084 ( .A(n25327), .B(n25328), .Z(n25326) );
  XOR U25085 ( .A(n25325), .B(n25329), .Z(n25327) );
  XNOR U25086 ( .A(n25288), .B(n25295), .Z(n25307) );
  NOR U25087 ( .A(n25256), .B(n25330), .Z(n25295) );
  XOR U25088 ( .A(n25300), .B(n25299), .Z(n25288) );
  XNOR U25089 ( .A(n25331), .B(n25296), .Z(n25299) );
  XOR U25090 ( .A(n25332), .B(n25333), .Z(n25296) );
  AND U25091 ( .A(n25334), .B(n25335), .Z(n25333) );
  XOR U25092 ( .A(n25332), .B(n25336), .Z(n25334) );
  XNOR U25093 ( .A(n25337), .B(n25338), .Z(n25331) );
  NOR U25094 ( .A(n25339), .B(n25340), .Z(n25338) );
  XNOR U25095 ( .A(n25337), .B(n25341), .Z(n25339) );
  XOR U25096 ( .A(n25342), .B(n25343), .Z(n25300) );
  NOR U25097 ( .A(n25344), .B(n25345), .Z(n25343) );
  XNOR U25098 ( .A(n25342), .B(n25346), .Z(n25344) );
  XNOR U25099 ( .A(n25245), .B(n25303), .Z(n25305) );
  XNOR U25100 ( .A(n25347), .B(n25348), .Z(n25245) );
  AND U25101 ( .A(n622), .B(n25252), .Z(n25348) );
  XOR U25102 ( .A(n25347), .B(n25250), .Z(n25252) );
  AND U25103 ( .A(n25253), .B(n25256), .Z(n25303) );
  XOR U25104 ( .A(n25349), .B(n25330), .Z(n25256) );
  XNOR U25105 ( .A(p_input[2048]), .B(p_input[848]), .Z(n25330) );
  XOR U25106 ( .A(n25318), .B(n25317), .Z(n25349) );
  XNOR U25107 ( .A(n25350), .B(n25324), .Z(n25317) );
  XNOR U25108 ( .A(n25313), .B(n25312), .Z(n25324) );
  XOR U25109 ( .A(n25351), .B(n25309), .Z(n25312) );
  XNOR U25110 ( .A(n16904), .B(p_input[858]), .Z(n25309) );
  XNOR U25111 ( .A(p_input[2059]), .B(p_input[859]), .Z(n25351) );
  XOR U25112 ( .A(p_input[2060]), .B(p_input[860]), .Z(n25313) );
  XNOR U25113 ( .A(n25323), .B(n25314), .Z(n25350) );
  XNOR U25114 ( .A(n17068), .B(p_input[849]), .Z(n25314) );
  XOR U25115 ( .A(n25352), .B(n25329), .Z(n25323) );
  XNOR U25116 ( .A(p_input[2063]), .B(p_input[863]), .Z(n25329) );
  XOR U25117 ( .A(n25320), .B(n25328), .Z(n25352) );
  XOR U25118 ( .A(n25353), .B(n25325), .Z(n25328) );
  XOR U25119 ( .A(p_input[2061]), .B(p_input[861]), .Z(n25325) );
  XNOR U25120 ( .A(p_input[2062]), .B(p_input[862]), .Z(n25353) );
  XNOR U25121 ( .A(n16738), .B(p_input[857]), .Z(n25320) );
  XNOR U25122 ( .A(n25336), .B(n25335), .Z(n25318) );
  XNOR U25123 ( .A(n25354), .B(n25341), .Z(n25335) );
  XOR U25124 ( .A(p_input[2056]), .B(p_input[856]), .Z(n25341) );
  XOR U25125 ( .A(n25332), .B(n25340), .Z(n25354) );
  XOR U25126 ( .A(n25355), .B(n25337), .Z(n25340) );
  XOR U25127 ( .A(p_input[2054]), .B(p_input[854]), .Z(n25337) );
  XNOR U25128 ( .A(p_input[2055]), .B(p_input[855]), .Z(n25355) );
  XNOR U25129 ( .A(n16741), .B(p_input[850]), .Z(n25332) );
  XNOR U25130 ( .A(n25346), .B(n25345), .Z(n25336) );
  XOR U25131 ( .A(n25356), .B(n25342), .Z(n25345) );
  XOR U25132 ( .A(p_input[2051]), .B(p_input[851]), .Z(n25342) );
  XNOR U25133 ( .A(p_input[2052]), .B(p_input[852]), .Z(n25356) );
  XOR U25134 ( .A(p_input[2053]), .B(p_input[853]), .Z(n25346) );
  XNOR U25135 ( .A(n25357), .B(n25358), .Z(n25253) );
  AND U25136 ( .A(n622), .B(n25359), .Z(n25358) );
  XNOR U25137 ( .A(n25360), .B(n25361), .Z(n622) );
  AND U25138 ( .A(n25362), .B(n25363), .Z(n25361) );
  XOR U25139 ( .A(n25360), .B(n25263), .Z(n25363) );
  XNOR U25140 ( .A(n25360), .B(n25217), .Z(n25362) );
  XOR U25141 ( .A(n25364), .B(n25365), .Z(n25360) );
  AND U25142 ( .A(n25366), .B(n25367), .Z(n25365) );
  XOR U25143 ( .A(n25364), .B(n25227), .Z(n25366) );
  XOR U25144 ( .A(n25368), .B(n25369), .Z(n25206) );
  AND U25145 ( .A(n626), .B(n25359), .Z(n25369) );
  XNOR U25146 ( .A(n25357), .B(n25368), .Z(n25359) );
  XNOR U25147 ( .A(n25370), .B(n25371), .Z(n626) );
  AND U25148 ( .A(n25372), .B(n25373), .Z(n25371) );
  XNOR U25149 ( .A(n25374), .B(n25370), .Z(n25373) );
  IV U25150 ( .A(n25263), .Z(n25374) );
  XNOR U25151 ( .A(n25375), .B(n25376), .Z(n25263) );
  AND U25152 ( .A(n629), .B(n25377), .Z(n25376) );
  XNOR U25153 ( .A(n25375), .B(n25378), .Z(n25377) );
  XNOR U25154 ( .A(n25217), .B(n25370), .Z(n25372) );
  XOR U25155 ( .A(n25379), .B(n25380), .Z(n25217) );
  AND U25156 ( .A(n637), .B(n25381), .Z(n25380) );
  XOR U25157 ( .A(n25364), .B(n25382), .Z(n25370) );
  AND U25158 ( .A(n25383), .B(n25367), .Z(n25382) );
  XNOR U25159 ( .A(n25276), .B(n25364), .Z(n25367) );
  XNOR U25160 ( .A(n25384), .B(n25385), .Z(n25276) );
  AND U25161 ( .A(n629), .B(n25386), .Z(n25385) );
  XOR U25162 ( .A(n25387), .B(n25384), .Z(n25386) );
  XNOR U25163 ( .A(n25388), .B(n25364), .Z(n25383) );
  IV U25164 ( .A(n25227), .Z(n25388) );
  XOR U25165 ( .A(n25389), .B(n25390), .Z(n25227) );
  AND U25166 ( .A(n637), .B(n25391), .Z(n25390) );
  XOR U25167 ( .A(n25392), .B(n25393), .Z(n25364) );
  AND U25168 ( .A(n25394), .B(n25395), .Z(n25393) );
  XNOR U25169 ( .A(n25301), .B(n25392), .Z(n25395) );
  XNOR U25170 ( .A(n25396), .B(n25397), .Z(n25301) );
  AND U25171 ( .A(n629), .B(n25398), .Z(n25397) );
  XNOR U25172 ( .A(n25399), .B(n25396), .Z(n25398) );
  XOR U25173 ( .A(n25392), .B(n25238), .Z(n25394) );
  XOR U25174 ( .A(n25400), .B(n25401), .Z(n25238) );
  AND U25175 ( .A(n637), .B(n25402), .Z(n25401) );
  XOR U25176 ( .A(n25403), .B(n25404), .Z(n25392) );
  AND U25177 ( .A(n25405), .B(n25406), .Z(n25404) );
  XNOR U25178 ( .A(n25403), .B(n25347), .Z(n25406) );
  XNOR U25179 ( .A(n25407), .B(n25408), .Z(n25347) );
  AND U25180 ( .A(n629), .B(n25409), .Z(n25408) );
  XOR U25181 ( .A(n25410), .B(n25407), .Z(n25409) );
  XNOR U25182 ( .A(n25411), .B(n25403), .Z(n25405) );
  IV U25183 ( .A(n25250), .Z(n25411) );
  XOR U25184 ( .A(n25412), .B(n25413), .Z(n25250) );
  AND U25185 ( .A(n637), .B(n25414), .Z(n25413) );
  AND U25186 ( .A(n25368), .B(n25357), .Z(n25403) );
  XNOR U25187 ( .A(n25415), .B(n25416), .Z(n25357) );
  AND U25188 ( .A(n629), .B(n25417), .Z(n25416) );
  XNOR U25189 ( .A(n25418), .B(n25415), .Z(n25417) );
  XNOR U25190 ( .A(n25419), .B(n25420), .Z(n629) );
  AND U25191 ( .A(n25421), .B(n25422), .Z(n25420) );
  XOR U25192 ( .A(n25378), .B(n25419), .Z(n25422) );
  AND U25193 ( .A(n25423), .B(n25424), .Z(n25378) );
  XOR U25194 ( .A(n25419), .B(n25375), .Z(n25421) );
  XNOR U25195 ( .A(n25425), .B(n25426), .Z(n25375) );
  AND U25196 ( .A(n633), .B(n25381), .Z(n25426) );
  XOR U25197 ( .A(n25379), .B(n25425), .Z(n25381) );
  XOR U25198 ( .A(n25427), .B(n25428), .Z(n25419) );
  AND U25199 ( .A(n25429), .B(n25430), .Z(n25428) );
  XNOR U25200 ( .A(n25427), .B(n25423), .Z(n25430) );
  IV U25201 ( .A(n25387), .Z(n25423) );
  XOR U25202 ( .A(n25431), .B(n25432), .Z(n25387) );
  XOR U25203 ( .A(n25433), .B(n25424), .Z(n25432) );
  AND U25204 ( .A(n25399), .B(n25434), .Z(n25424) );
  AND U25205 ( .A(n25435), .B(n25436), .Z(n25433) );
  XOR U25206 ( .A(n25437), .B(n25431), .Z(n25435) );
  XNOR U25207 ( .A(n25384), .B(n25427), .Z(n25429) );
  XNOR U25208 ( .A(n25438), .B(n25439), .Z(n25384) );
  AND U25209 ( .A(n633), .B(n25391), .Z(n25439) );
  XOR U25210 ( .A(n25438), .B(n25389), .Z(n25391) );
  XOR U25211 ( .A(n25440), .B(n25441), .Z(n25427) );
  AND U25212 ( .A(n25442), .B(n25443), .Z(n25441) );
  XNOR U25213 ( .A(n25440), .B(n25399), .Z(n25443) );
  XOR U25214 ( .A(n25444), .B(n25436), .Z(n25399) );
  XNOR U25215 ( .A(n25445), .B(n25431), .Z(n25436) );
  XOR U25216 ( .A(n25446), .B(n25447), .Z(n25431) );
  AND U25217 ( .A(n25448), .B(n25449), .Z(n25447) );
  XOR U25218 ( .A(n25450), .B(n25446), .Z(n25448) );
  XNOR U25219 ( .A(n25451), .B(n25452), .Z(n25445) );
  AND U25220 ( .A(n25453), .B(n25454), .Z(n25452) );
  XOR U25221 ( .A(n25451), .B(n25455), .Z(n25453) );
  XNOR U25222 ( .A(n25437), .B(n25434), .Z(n25444) );
  AND U25223 ( .A(n25456), .B(n25457), .Z(n25434) );
  XOR U25224 ( .A(n25458), .B(n25459), .Z(n25437) );
  AND U25225 ( .A(n25460), .B(n25461), .Z(n25459) );
  XOR U25226 ( .A(n25458), .B(n25462), .Z(n25460) );
  XNOR U25227 ( .A(n25396), .B(n25440), .Z(n25442) );
  XNOR U25228 ( .A(n25463), .B(n25464), .Z(n25396) );
  AND U25229 ( .A(n633), .B(n25402), .Z(n25464) );
  XOR U25230 ( .A(n25463), .B(n25400), .Z(n25402) );
  XOR U25231 ( .A(n25465), .B(n25466), .Z(n25440) );
  AND U25232 ( .A(n25467), .B(n25468), .Z(n25466) );
  XNOR U25233 ( .A(n25465), .B(n25456), .Z(n25468) );
  IV U25234 ( .A(n25410), .Z(n25456) );
  XNOR U25235 ( .A(n25469), .B(n25449), .Z(n25410) );
  XNOR U25236 ( .A(n25470), .B(n25455), .Z(n25449) );
  XOR U25237 ( .A(n25471), .B(n25472), .Z(n25455) );
  NOR U25238 ( .A(n25473), .B(n25474), .Z(n25472) );
  XNOR U25239 ( .A(n25471), .B(n25475), .Z(n25473) );
  XNOR U25240 ( .A(n25454), .B(n25446), .Z(n25470) );
  XOR U25241 ( .A(n25476), .B(n25477), .Z(n25446) );
  AND U25242 ( .A(n25478), .B(n25479), .Z(n25477) );
  XNOR U25243 ( .A(n25476), .B(n25480), .Z(n25478) );
  XNOR U25244 ( .A(n25481), .B(n25451), .Z(n25454) );
  XOR U25245 ( .A(n25482), .B(n25483), .Z(n25451) );
  AND U25246 ( .A(n25484), .B(n25485), .Z(n25483) );
  XOR U25247 ( .A(n25482), .B(n25486), .Z(n25484) );
  XNOR U25248 ( .A(n25487), .B(n25488), .Z(n25481) );
  NOR U25249 ( .A(n25489), .B(n25490), .Z(n25488) );
  XOR U25250 ( .A(n25487), .B(n25491), .Z(n25489) );
  XNOR U25251 ( .A(n25450), .B(n25457), .Z(n25469) );
  NOR U25252 ( .A(n25418), .B(n25492), .Z(n25457) );
  XOR U25253 ( .A(n25462), .B(n25461), .Z(n25450) );
  XNOR U25254 ( .A(n25493), .B(n25458), .Z(n25461) );
  XOR U25255 ( .A(n25494), .B(n25495), .Z(n25458) );
  AND U25256 ( .A(n25496), .B(n25497), .Z(n25495) );
  XOR U25257 ( .A(n25494), .B(n25498), .Z(n25496) );
  XNOR U25258 ( .A(n25499), .B(n25500), .Z(n25493) );
  NOR U25259 ( .A(n25501), .B(n25502), .Z(n25500) );
  XNOR U25260 ( .A(n25499), .B(n25503), .Z(n25501) );
  XOR U25261 ( .A(n25504), .B(n25505), .Z(n25462) );
  NOR U25262 ( .A(n25506), .B(n25507), .Z(n25505) );
  XNOR U25263 ( .A(n25504), .B(n25508), .Z(n25506) );
  XNOR U25264 ( .A(n25407), .B(n25465), .Z(n25467) );
  XNOR U25265 ( .A(n25509), .B(n25510), .Z(n25407) );
  AND U25266 ( .A(n633), .B(n25414), .Z(n25510) );
  XOR U25267 ( .A(n25509), .B(n25412), .Z(n25414) );
  AND U25268 ( .A(n25415), .B(n25418), .Z(n25465) );
  XOR U25269 ( .A(n25511), .B(n25492), .Z(n25418) );
  XNOR U25270 ( .A(p_input[2048]), .B(p_input[864]), .Z(n25492) );
  XOR U25271 ( .A(n25480), .B(n25479), .Z(n25511) );
  XNOR U25272 ( .A(n25512), .B(n25486), .Z(n25479) );
  XNOR U25273 ( .A(n25475), .B(n25474), .Z(n25486) );
  XOR U25274 ( .A(n25513), .B(n25471), .Z(n25474) );
  XNOR U25275 ( .A(n16904), .B(p_input[874]), .Z(n25471) );
  XNOR U25276 ( .A(p_input[2059]), .B(p_input[875]), .Z(n25513) );
  XOR U25277 ( .A(p_input[2060]), .B(p_input[876]), .Z(n25475) );
  XNOR U25278 ( .A(n25485), .B(n25476), .Z(n25512) );
  XNOR U25279 ( .A(n17068), .B(p_input[865]), .Z(n25476) );
  XOR U25280 ( .A(n25514), .B(n25491), .Z(n25485) );
  XNOR U25281 ( .A(p_input[2063]), .B(p_input[879]), .Z(n25491) );
  XOR U25282 ( .A(n25482), .B(n25490), .Z(n25514) );
  XOR U25283 ( .A(n25515), .B(n25487), .Z(n25490) );
  XOR U25284 ( .A(p_input[2061]), .B(p_input[877]), .Z(n25487) );
  XNOR U25285 ( .A(p_input[2062]), .B(p_input[878]), .Z(n25515) );
  XNOR U25286 ( .A(n16738), .B(p_input[873]), .Z(n25482) );
  XNOR U25287 ( .A(n25498), .B(n25497), .Z(n25480) );
  XNOR U25288 ( .A(n25516), .B(n25503), .Z(n25497) );
  XOR U25289 ( .A(p_input[2056]), .B(p_input[872]), .Z(n25503) );
  XOR U25290 ( .A(n25494), .B(n25502), .Z(n25516) );
  XOR U25291 ( .A(n25517), .B(n25499), .Z(n25502) );
  XOR U25292 ( .A(p_input[2054]), .B(p_input[870]), .Z(n25499) );
  XNOR U25293 ( .A(p_input[2055]), .B(p_input[871]), .Z(n25517) );
  XNOR U25294 ( .A(n16741), .B(p_input[866]), .Z(n25494) );
  XNOR U25295 ( .A(n25508), .B(n25507), .Z(n25498) );
  XOR U25296 ( .A(n25518), .B(n25504), .Z(n25507) );
  XOR U25297 ( .A(p_input[2051]), .B(p_input[867]), .Z(n25504) );
  XNOR U25298 ( .A(p_input[2052]), .B(p_input[868]), .Z(n25518) );
  XOR U25299 ( .A(p_input[2053]), .B(p_input[869]), .Z(n25508) );
  XNOR U25300 ( .A(n25519), .B(n25520), .Z(n25415) );
  AND U25301 ( .A(n633), .B(n25521), .Z(n25520) );
  XNOR U25302 ( .A(n25522), .B(n25523), .Z(n633) );
  AND U25303 ( .A(n25524), .B(n25525), .Z(n25523) );
  XOR U25304 ( .A(n25522), .B(n25425), .Z(n25525) );
  XNOR U25305 ( .A(n25522), .B(n25379), .Z(n25524) );
  XOR U25306 ( .A(n25526), .B(n25527), .Z(n25522) );
  AND U25307 ( .A(n25528), .B(n25529), .Z(n25527) );
  XOR U25308 ( .A(n25526), .B(n25389), .Z(n25528) );
  XOR U25309 ( .A(n25530), .B(n25531), .Z(n25368) );
  AND U25310 ( .A(n637), .B(n25521), .Z(n25531) );
  XNOR U25311 ( .A(n25519), .B(n25530), .Z(n25521) );
  XNOR U25312 ( .A(n25532), .B(n25533), .Z(n637) );
  AND U25313 ( .A(n25534), .B(n25535), .Z(n25533) );
  XNOR U25314 ( .A(n25536), .B(n25532), .Z(n25535) );
  IV U25315 ( .A(n25425), .Z(n25536) );
  XNOR U25316 ( .A(n25537), .B(n25538), .Z(n25425) );
  AND U25317 ( .A(n640), .B(n25539), .Z(n25538) );
  XNOR U25318 ( .A(n25537), .B(n25540), .Z(n25539) );
  XNOR U25319 ( .A(n25379), .B(n25532), .Z(n25534) );
  XOR U25320 ( .A(n25541), .B(n25542), .Z(n25379) );
  AND U25321 ( .A(n648), .B(n25543), .Z(n25542) );
  XOR U25322 ( .A(n25526), .B(n25544), .Z(n25532) );
  AND U25323 ( .A(n25545), .B(n25529), .Z(n25544) );
  XNOR U25324 ( .A(n25438), .B(n25526), .Z(n25529) );
  XNOR U25325 ( .A(n25546), .B(n25547), .Z(n25438) );
  AND U25326 ( .A(n640), .B(n25548), .Z(n25547) );
  XOR U25327 ( .A(n25549), .B(n25546), .Z(n25548) );
  XNOR U25328 ( .A(n25550), .B(n25526), .Z(n25545) );
  IV U25329 ( .A(n25389), .Z(n25550) );
  XOR U25330 ( .A(n25551), .B(n25552), .Z(n25389) );
  AND U25331 ( .A(n648), .B(n25553), .Z(n25552) );
  XOR U25332 ( .A(n25554), .B(n25555), .Z(n25526) );
  AND U25333 ( .A(n25556), .B(n25557), .Z(n25555) );
  XNOR U25334 ( .A(n25463), .B(n25554), .Z(n25557) );
  XNOR U25335 ( .A(n25558), .B(n25559), .Z(n25463) );
  AND U25336 ( .A(n640), .B(n25560), .Z(n25559) );
  XNOR U25337 ( .A(n25561), .B(n25558), .Z(n25560) );
  XOR U25338 ( .A(n25554), .B(n25400), .Z(n25556) );
  XOR U25339 ( .A(n25562), .B(n25563), .Z(n25400) );
  AND U25340 ( .A(n648), .B(n25564), .Z(n25563) );
  XOR U25341 ( .A(n25565), .B(n25566), .Z(n25554) );
  AND U25342 ( .A(n25567), .B(n25568), .Z(n25566) );
  XNOR U25343 ( .A(n25565), .B(n25509), .Z(n25568) );
  XNOR U25344 ( .A(n25569), .B(n25570), .Z(n25509) );
  AND U25345 ( .A(n640), .B(n25571), .Z(n25570) );
  XOR U25346 ( .A(n25572), .B(n25569), .Z(n25571) );
  XNOR U25347 ( .A(n25573), .B(n25565), .Z(n25567) );
  IV U25348 ( .A(n25412), .Z(n25573) );
  XOR U25349 ( .A(n25574), .B(n25575), .Z(n25412) );
  AND U25350 ( .A(n648), .B(n25576), .Z(n25575) );
  AND U25351 ( .A(n25530), .B(n25519), .Z(n25565) );
  XNOR U25352 ( .A(n25577), .B(n25578), .Z(n25519) );
  AND U25353 ( .A(n640), .B(n25579), .Z(n25578) );
  XNOR U25354 ( .A(n25580), .B(n25577), .Z(n25579) );
  XNOR U25355 ( .A(n25581), .B(n25582), .Z(n640) );
  AND U25356 ( .A(n25583), .B(n25584), .Z(n25582) );
  XOR U25357 ( .A(n25540), .B(n25581), .Z(n25584) );
  AND U25358 ( .A(n25585), .B(n25586), .Z(n25540) );
  XOR U25359 ( .A(n25581), .B(n25537), .Z(n25583) );
  XNOR U25360 ( .A(n25587), .B(n25588), .Z(n25537) );
  AND U25361 ( .A(n644), .B(n25543), .Z(n25588) );
  XOR U25362 ( .A(n25541), .B(n25587), .Z(n25543) );
  XOR U25363 ( .A(n25589), .B(n25590), .Z(n25581) );
  AND U25364 ( .A(n25591), .B(n25592), .Z(n25590) );
  XNOR U25365 ( .A(n25589), .B(n25585), .Z(n25592) );
  IV U25366 ( .A(n25549), .Z(n25585) );
  XOR U25367 ( .A(n25593), .B(n25594), .Z(n25549) );
  XOR U25368 ( .A(n25595), .B(n25586), .Z(n25594) );
  AND U25369 ( .A(n25561), .B(n25596), .Z(n25586) );
  AND U25370 ( .A(n25597), .B(n25598), .Z(n25595) );
  XOR U25371 ( .A(n25599), .B(n25593), .Z(n25597) );
  XNOR U25372 ( .A(n25546), .B(n25589), .Z(n25591) );
  XNOR U25373 ( .A(n25600), .B(n25601), .Z(n25546) );
  AND U25374 ( .A(n644), .B(n25553), .Z(n25601) );
  XOR U25375 ( .A(n25600), .B(n25551), .Z(n25553) );
  XOR U25376 ( .A(n25602), .B(n25603), .Z(n25589) );
  AND U25377 ( .A(n25604), .B(n25605), .Z(n25603) );
  XNOR U25378 ( .A(n25602), .B(n25561), .Z(n25605) );
  XOR U25379 ( .A(n25606), .B(n25598), .Z(n25561) );
  XNOR U25380 ( .A(n25607), .B(n25593), .Z(n25598) );
  XOR U25381 ( .A(n25608), .B(n25609), .Z(n25593) );
  AND U25382 ( .A(n25610), .B(n25611), .Z(n25609) );
  XOR U25383 ( .A(n25612), .B(n25608), .Z(n25610) );
  XNOR U25384 ( .A(n25613), .B(n25614), .Z(n25607) );
  AND U25385 ( .A(n25615), .B(n25616), .Z(n25614) );
  XOR U25386 ( .A(n25613), .B(n25617), .Z(n25615) );
  XNOR U25387 ( .A(n25599), .B(n25596), .Z(n25606) );
  AND U25388 ( .A(n25618), .B(n25619), .Z(n25596) );
  XOR U25389 ( .A(n25620), .B(n25621), .Z(n25599) );
  AND U25390 ( .A(n25622), .B(n25623), .Z(n25621) );
  XOR U25391 ( .A(n25620), .B(n25624), .Z(n25622) );
  XNOR U25392 ( .A(n25558), .B(n25602), .Z(n25604) );
  XNOR U25393 ( .A(n25625), .B(n25626), .Z(n25558) );
  AND U25394 ( .A(n644), .B(n25564), .Z(n25626) );
  XOR U25395 ( .A(n25625), .B(n25562), .Z(n25564) );
  XOR U25396 ( .A(n25627), .B(n25628), .Z(n25602) );
  AND U25397 ( .A(n25629), .B(n25630), .Z(n25628) );
  XNOR U25398 ( .A(n25627), .B(n25618), .Z(n25630) );
  IV U25399 ( .A(n25572), .Z(n25618) );
  XNOR U25400 ( .A(n25631), .B(n25611), .Z(n25572) );
  XNOR U25401 ( .A(n25632), .B(n25617), .Z(n25611) );
  XOR U25402 ( .A(n25633), .B(n25634), .Z(n25617) );
  NOR U25403 ( .A(n25635), .B(n25636), .Z(n25634) );
  XNOR U25404 ( .A(n25633), .B(n25637), .Z(n25635) );
  XNOR U25405 ( .A(n25616), .B(n25608), .Z(n25632) );
  XOR U25406 ( .A(n25638), .B(n25639), .Z(n25608) );
  AND U25407 ( .A(n25640), .B(n25641), .Z(n25639) );
  XNOR U25408 ( .A(n25638), .B(n25642), .Z(n25640) );
  XNOR U25409 ( .A(n25643), .B(n25613), .Z(n25616) );
  XOR U25410 ( .A(n25644), .B(n25645), .Z(n25613) );
  AND U25411 ( .A(n25646), .B(n25647), .Z(n25645) );
  XOR U25412 ( .A(n25644), .B(n25648), .Z(n25646) );
  XNOR U25413 ( .A(n25649), .B(n25650), .Z(n25643) );
  NOR U25414 ( .A(n25651), .B(n25652), .Z(n25650) );
  XOR U25415 ( .A(n25649), .B(n25653), .Z(n25651) );
  XNOR U25416 ( .A(n25612), .B(n25619), .Z(n25631) );
  NOR U25417 ( .A(n25580), .B(n25654), .Z(n25619) );
  XOR U25418 ( .A(n25624), .B(n25623), .Z(n25612) );
  XNOR U25419 ( .A(n25655), .B(n25620), .Z(n25623) );
  XOR U25420 ( .A(n25656), .B(n25657), .Z(n25620) );
  AND U25421 ( .A(n25658), .B(n25659), .Z(n25657) );
  XOR U25422 ( .A(n25656), .B(n25660), .Z(n25658) );
  XNOR U25423 ( .A(n25661), .B(n25662), .Z(n25655) );
  NOR U25424 ( .A(n25663), .B(n25664), .Z(n25662) );
  XNOR U25425 ( .A(n25661), .B(n25665), .Z(n25663) );
  XOR U25426 ( .A(n25666), .B(n25667), .Z(n25624) );
  NOR U25427 ( .A(n25668), .B(n25669), .Z(n25667) );
  XNOR U25428 ( .A(n25666), .B(n25670), .Z(n25668) );
  XNOR U25429 ( .A(n25569), .B(n25627), .Z(n25629) );
  XNOR U25430 ( .A(n25671), .B(n25672), .Z(n25569) );
  AND U25431 ( .A(n644), .B(n25576), .Z(n25672) );
  XOR U25432 ( .A(n25671), .B(n25574), .Z(n25576) );
  AND U25433 ( .A(n25577), .B(n25580), .Z(n25627) );
  XOR U25434 ( .A(n25673), .B(n25654), .Z(n25580) );
  XNOR U25435 ( .A(p_input[2048]), .B(p_input[880]), .Z(n25654) );
  XOR U25436 ( .A(n25642), .B(n25641), .Z(n25673) );
  XNOR U25437 ( .A(n25674), .B(n25648), .Z(n25641) );
  XNOR U25438 ( .A(n25637), .B(n25636), .Z(n25648) );
  XOR U25439 ( .A(n25675), .B(n25633), .Z(n25636) );
  XNOR U25440 ( .A(n16904), .B(p_input[890]), .Z(n25633) );
  XNOR U25441 ( .A(p_input[2059]), .B(p_input[891]), .Z(n25675) );
  XOR U25442 ( .A(p_input[2060]), .B(p_input[892]), .Z(n25637) );
  XNOR U25443 ( .A(n25647), .B(n25638), .Z(n25674) );
  XNOR U25444 ( .A(n17068), .B(p_input[881]), .Z(n25638) );
  XOR U25445 ( .A(n25676), .B(n25653), .Z(n25647) );
  XNOR U25446 ( .A(p_input[2063]), .B(p_input[895]), .Z(n25653) );
  XOR U25447 ( .A(n25644), .B(n25652), .Z(n25676) );
  XOR U25448 ( .A(n25677), .B(n25649), .Z(n25652) );
  XOR U25449 ( .A(p_input[2061]), .B(p_input[893]), .Z(n25649) );
  XNOR U25450 ( .A(p_input[2062]), .B(p_input[894]), .Z(n25677) );
  XNOR U25451 ( .A(n16738), .B(p_input[889]), .Z(n25644) );
  XNOR U25452 ( .A(n25660), .B(n25659), .Z(n25642) );
  XNOR U25453 ( .A(n25678), .B(n25665), .Z(n25659) );
  XOR U25454 ( .A(p_input[2056]), .B(p_input[888]), .Z(n25665) );
  XOR U25455 ( .A(n25656), .B(n25664), .Z(n25678) );
  XOR U25456 ( .A(n25679), .B(n25661), .Z(n25664) );
  XOR U25457 ( .A(p_input[2054]), .B(p_input[886]), .Z(n25661) );
  XNOR U25458 ( .A(p_input[2055]), .B(p_input[887]), .Z(n25679) );
  XNOR U25459 ( .A(n16741), .B(p_input[882]), .Z(n25656) );
  XNOR U25460 ( .A(n25670), .B(n25669), .Z(n25660) );
  XOR U25461 ( .A(n25680), .B(n25666), .Z(n25669) );
  XOR U25462 ( .A(p_input[2051]), .B(p_input[883]), .Z(n25666) );
  XNOR U25463 ( .A(p_input[2052]), .B(p_input[884]), .Z(n25680) );
  XOR U25464 ( .A(p_input[2053]), .B(p_input[885]), .Z(n25670) );
  XNOR U25465 ( .A(n25681), .B(n25682), .Z(n25577) );
  AND U25466 ( .A(n644), .B(n25683), .Z(n25682) );
  XNOR U25467 ( .A(n25684), .B(n25685), .Z(n644) );
  AND U25468 ( .A(n25686), .B(n25687), .Z(n25685) );
  XOR U25469 ( .A(n25684), .B(n25587), .Z(n25687) );
  XNOR U25470 ( .A(n25684), .B(n25541), .Z(n25686) );
  XOR U25471 ( .A(n25688), .B(n25689), .Z(n25684) );
  AND U25472 ( .A(n25690), .B(n25691), .Z(n25689) );
  XOR U25473 ( .A(n25688), .B(n25551), .Z(n25690) );
  XOR U25474 ( .A(n25692), .B(n25693), .Z(n25530) );
  AND U25475 ( .A(n648), .B(n25683), .Z(n25693) );
  XNOR U25476 ( .A(n25681), .B(n25692), .Z(n25683) );
  XNOR U25477 ( .A(n25694), .B(n25695), .Z(n648) );
  AND U25478 ( .A(n25696), .B(n25697), .Z(n25695) );
  XNOR U25479 ( .A(n25698), .B(n25694), .Z(n25697) );
  IV U25480 ( .A(n25587), .Z(n25698) );
  XNOR U25481 ( .A(n25699), .B(n25700), .Z(n25587) );
  AND U25482 ( .A(n651), .B(n25701), .Z(n25700) );
  XNOR U25483 ( .A(n25699), .B(n25702), .Z(n25701) );
  XNOR U25484 ( .A(n25541), .B(n25694), .Z(n25696) );
  XOR U25485 ( .A(n25703), .B(n25704), .Z(n25541) );
  AND U25486 ( .A(n659), .B(n25705), .Z(n25704) );
  XOR U25487 ( .A(n25688), .B(n25706), .Z(n25694) );
  AND U25488 ( .A(n25707), .B(n25691), .Z(n25706) );
  XNOR U25489 ( .A(n25600), .B(n25688), .Z(n25691) );
  XNOR U25490 ( .A(n25708), .B(n25709), .Z(n25600) );
  AND U25491 ( .A(n651), .B(n25710), .Z(n25709) );
  XOR U25492 ( .A(n25711), .B(n25708), .Z(n25710) );
  XNOR U25493 ( .A(n25712), .B(n25688), .Z(n25707) );
  IV U25494 ( .A(n25551), .Z(n25712) );
  XOR U25495 ( .A(n25713), .B(n25714), .Z(n25551) );
  AND U25496 ( .A(n659), .B(n25715), .Z(n25714) );
  XOR U25497 ( .A(n25716), .B(n25717), .Z(n25688) );
  AND U25498 ( .A(n25718), .B(n25719), .Z(n25717) );
  XNOR U25499 ( .A(n25625), .B(n25716), .Z(n25719) );
  XNOR U25500 ( .A(n25720), .B(n25721), .Z(n25625) );
  AND U25501 ( .A(n651), .B(n25722), .Z(n25721) );
  XNOR U25502 ( .A(n25723), .B(n25720), .Z(n25722) );
  XOR U25503 ( .A(n25716), .B(n25562), .Z(n25718) );
  XOR U25504 ( .A(n25724), .B(n25725), .Z(n25562) );
  AND U25505 ( .A(n659), .B(n25726), .Z(n25725) );
  XOR U25506 ( .A(n25727), .B(n25728), .Z(n25716) );
  AND U25507 ( .A(n25729), .B(n25730), .Z(n25728) );
  XNOR U25508 ( .A(n25727), .B(n25671), .Z(n25730) );
  XNOR U25509 ( .A(n25731), .B(n25732), .Z(n25671) );
  AND U25510 ( .A(n651), .B(n25733), .Z(n25732) );
  XOR U25511 ( .A(n25734), .B(n25731), .Z(n25733) );
  XNOR U25512 ( .A(n25735), .B(n25727), .Z(n25729) );
  IV U25513 ( .A(n25574), .Z(n25735) );
  XOR U25514 ( .A(n25736), .B(n25737), .Z(n25574) );
  AND U25515 ( .A(n659), .B(n25738), .Z(n25737) );
  AND U25516 ( .A(n25692), .B(n25681), .Z(n25727) );
  XNOR U25517 ( .A(n25739), .B(n25740), .Z(n25681) );
  AND U25518 ( .A(n651), .B(n25741), .Z(n25740) );
  XNOR U25519 ( .A(n25742), .B(n25739), .Z(n25741) );
  XNOR U25520 ( .A(n25743), .B(n25744), .Z(n651) );
  AND U25521 ( .A(n25745), .B(n25746), .Z(n25744) );
  XOR U25522 ( .A(n25702), .B(n25743), .Z(n25746) );
  AND U25523 ( .A(n25747), .B(n25748), .Z(n25702) );
  XOR U25524 ( .A(n25743), .B(n25699), .Z(n25745) );
  XNOR U25525 ( .A(n25749), .B(n25750), .Z(n25699) );
  AND U25526 ( .A(n655), .B(n25705), .Z(n25750) );
  XOR U25527 ( .A(n25703), .B(n25749), .Z(n25705) );
  XOR U25528 ( .A(n25751), .B(n25752), .Z(n25743) );
  AND U25529 ( .A(n25753), .B(n25754), .Z(n25752) );
  XNOR U25530 ( .A(n25751), .B(n25747), .Z(n25754) );
  IV U25531 ( .A(n25711), .Z(n25747) );
  XOR U25532 ( .A(n25755), .B(n25756), .Z(n25711) );
  XOR U25533 ( .A(n25757), .B(n25748), .Z(n25756) );
  AND U25534 ( .A(n25723), .B(n25758), .Z(n25748) );
  AND U25535 ( .A(n25759), .B(n25760), .Z(n25757) );
  XOR U25536 ( .A(n25761), .B(n25755), .Z(n25759) );
  XNOR U25537 ( .A(n25708), .B(n25751), .Z(n25753) );
  XNOR U25538 ( .A(n25762), .B(n25763), .Z(n25708) );
  AND U25539 ( .A(n655), .B(n25715), .Z(n25763) );
  XOR U25540 ( .A(n25762), .B(n25713), .Z(n25715) );
  XOR U25541 ( .A(n25764), .B(n25765), .Z(n25751) );
  AND U25542 ( .A(n25766), .B(n25767), .Z(n25765) );
  XNOR U25543 ( .A(n25764), .B(n25723), .Z(n25767) );
  XOR U25544 ( .A(n25768), .B(n25760), .Z(n25723) );
  XNOR U25545 ( .A(n25769), .B(n25755), .Z(n25760) );
  XOR U25546 ( .A(n25770), .B(n25771), .Z(n25755) );
  AND U25547 ( .A(n25772), .B(n25773), .Z(n25771) );
  XOR U25548 ( .A(n25774), .B(n25770), .Z(n25772) );
  XNOR U25549 ( .A(n25775), .B(n25776), .Z(n25769) );
  AND U25550 ( .A(n25777), .B(n25778), .Z(n25776) );
  XOR U25551 ( .A(n25775), .B(n25779), .Z(n25777) );
  XNOR U25552 ( .A(n25761), .B(n25758), .Z(n25768) );
  AND U25553 ( .A(n25780), .B(n25781), .Z(n25758) );
  XOR U25554 ( .A(n25782), .B(n25783), .Z(n25761) );
  AND U25555 ( .A(n25784), .B(n25785), .Z(n25783) );
  XOR U25556 ( .A(n25782), .B(n25786), .Z(n25784) );
  XNOR U25557 ( .A(n25720), .B(n25764), .Z(n25766) );
  XNOR U25558 ( .A(n25787), .B(n25788), .Z(n25720) );
  AND U25559 ( .A(n655), .B(n25726), .Z(n25788) );
  XOR U25560 ( .A(n25787), .B(n25724), .Z(n25726) );
  XOR U25561 ( .A(n25789), .B(n25790), .Z(n25764) );
  AND U25562 ( .A(n25791), .B(n25792), .Z(n25790) );
  XNOR U25563 ( .A(n25789), .B(n25780), .Z(n25792) );
  IV U25564 ( .A(n25734), .Z(n25780) );
  XNOR U25565 ( .A(n25793), .B(n25773), .Z(n25734) );
  XNOR U25566 ( .A(n25794), .B(n25779), .Z(n25773) );
  XOR U25567 ( .A(n25795), .B(n25796), .Z(n25779) );
  NOR U25568 ( .A(n25797), .B(n25798), .Z(n25796) );
  XNOR U25569 ( .A(n25795), .B(n25799), .Z(n25797) );
  XNOR U25570 ( .A(n25778), .B(n25770), .Z(n25794) );
  XOR U25571 ( .A(n25800), .B(n25801), .Z(n25770) );
  AND U25572 ( .A(n25802), .B(n25803), .Z(n25801) );
  XNOR U25573 ( .A(n25800), .B(n25804), .Z(n25802) );
  XNOR U25574 ( .A(n25805), .B(n25775), .Z(n25778) );
  XOR U25575 ( .A(n25806), .B(n25807), .Z(n25775) );
  AND U25576 ( .A(n25808), .B(n25809), .Z(n25807) );
  XOR U25577 ( .A(n25806), .B(n25810), .Z(n25808) );
  XNOR U25578 ( .A(n25811), .B(n25812), .Z(n25805) );
  NOR U25579 ( .A(n25813), .B(n25814), .Z(n25812) );
  XOR U25580 ( .A(n25811), .B(n25815), .Z(n25813) );
  XNOR U25581 ( .A(n25774), .B(n25781), .Z(n25793) );
  NOR U25582 ( .A(n25742), .B(n25816), .Z(n25781) );
  XOR U25583 ( .A(n25786), .B(n25785), .Z(n25774) );
  XNOR U25584 ( .A(n25817), .B(n25782), .Z(n25785) );
  XOR U25585 ( .A(n25818), .B(n25819), .Z(n25782) );
  AND U25586 ( .A(n25820), .B(n25821), .Z(n25819) );
  XOR U25587 ( .A(n25818), .B(n25822), .Z(n25820) );
  XNOR U25588 ( .A(n25823), .B(n25824), .Z(n25817) );
  NOR U25589 ( .A(n25825), .B(n25826), .Z(n25824) );
  XNOR U25590 ( .A(n25823), .B(n25827), .Z(n25825) );
  XOR U25591 ( .A(n25828), .B(n25829), .Z(n25786) );
  NOR U25592 ( .A(n25830), .B(n25831), .Z(n25829) );
  XNOR U25593 ( .A(n25828), .B(n25832), .Z(n25830) );
  XNOR U25594 ( .A(n25731), .B(n25789), .Z(n25791) );
  XNOR U25595 ( .A(n25833), .B(n25834), .Z(n25731) );
  AND U25596 ( .A(n655), .B(n25738), .Z(n25834) );
  XOR U25597 ( .A(n25833), .B(n25736), .Z(n25738) );
  AND U25598 ( .A(n25739), .B(n25742), .Z(n25789) );
  XOR U25599 ( .A(n25835), .B(n25816), .Z(n25742) );
  XNOR U25600 ( .A(p_input[2048]), .B(p_input[896]), .Z(n25816) );
  XOR U25601 ( .A(n25804), .B(n25803), .Z(n25835) );
  XNOR U25602 ( .A(n25836), .B(n25810), .Z(n25803) );
  XNOR U25603 ( .A(n25799), .B(n25798), .Z(n25810) );
  XOR U25604 ( .A(n25837), .B(n25795), .Z(n25798) );
  XNOR U25605 ( .A(n16904), .B(p_input[906]), .Z(n25795) );
  XNOR U25606 ( .A(p_input[2059]), .B(p_input[907]), .Z(n25837) );
  XOR U25607 ( .A(p_input[2060]), .B(p_input[908]), .Z(n25799) );
  XNOR U25608 ( .A(n25809), .B(n25800), .Z(n25836) );
  XNOR U25609 ( .A(n17068), .B(p_input[897]), .Z(n25800) );
  XOR U25610 ( .A(n25838), .B(n25815), .Z(n25809) );
  XNOR U25611 ( .A(p_input[2063]), .B(p_input[911]), .Z(n25815) );
  XOR U25612 ( .A(n25806), .B(n25814), .Z(n25838) );
  XOR U25613 ( .A(n25839), .B(n25811), .Z(n25814) );
  XOR U25614 ( .A(p_input[2061]), .B(p_input[909]), .Z(n25811) );
  XNOR U25615 ( .A(p_input[2062]), .B(p_input[910]), .Z(n25839) );
  XNOR U25616 ( .A(n16738), .B(p_input[905]), .Z(n25806) );
  XNOR U25617 ( .A(n25822), .B(n25821), .Z(n25804) );
  XNOR U25618 ( .A(n25840), .B(n25827), .Z(n25821) );
  XOR U25619 ( .A(p_input[2056]), .B(p_input[904]), .Z(n25827) );
  XOR U25620 ( .A(n25818), .B(n25826), .Z(n25840) );
  XOR U25621 ( .A(n25841), .B(n25823), .Z(n25826) );
  XOR U25622 ( .A(p_input[2054]), .B(p_input[902]), .Z(n25823) );
  XNOR U25623 ( .A(p_input[2055]), .B(p_input[903]), .Z(n25841) );
  XNOR U25624 ( .A(n16741), .B(p_input[898]), .Z(n25818) );
  XNOR U25625 ( .A(n25832), .B(n25831), .Z(n25822) );
  XOR U25626 ( .A(n25842), .B(n25828), .Z(n25831) );
  XOR U25627 ( .A(p_input[2051]), .B(p_input[899]), .Z(n25828) );
  XNOR U25628 ( .A(p_input[2052]), .B(p_input[900]), .Z(n25842) );
  XOR U25629 ( .A(p_input[2053]), .B(p_input[901]), .Z(n25832) );
  XNOR U25630 ( .A(n25843), .B(n25844), .Z(n25739) );
  AND U25631 ( .A(n655), .B(n25845), .Z(n25844) );
  XNOR U25632 ( .A(n25846), .B(n25847), .Z(n655) );
  AND U25633 ( .A(n25848), .B(n25849), .Z(n25847) );
  XOR U25634 ( .A(n25846), .B(n25749), .Z(n25849) );
  XNOR U25635 ( .A(n25846), .B(n25703), .Z(n25848) );
  XOR U25636 ( .A(n25850), .B(n25851), .Z(n25846) );
  AND U25637 ( .A(n25852), .B(n25853), .Z(n25851) );
  XOR U25638 ( .A(n25850), .B(n25713), .Z(n25852) );
  XOR U25639 ( .A(n25854), .B(n25855), .Z(n25692) );
  AND U25640 ( .A(n659), .B(n25845), .Z(n25855) );
  XNOR U25641 ( .A(n25843), .B(n25854), .Z(n25845) );
  XNOR U25642 ( .A(n25856), .B(n25857), .Z(n659) );
  AND U25643 ( .A(n25858), .B(n25859), .Z(n25857) );
  XNOR U25644 ( .A(n25860), .B(n25856), .Z(n25859) );
  IV U25645 ( .A(n25749), .Z(n25860) );
  XNOR U25646 ( .A(n25861), .B(n25862), .Z(n25749) );
  AND U25647 ( .A(n662), .B(n25863), .Z(n25862) );
  XNOR U25648 ( .A(n25861), .B(n25864), .Z(n25863) );
  XNOR U25649 ( .A(n25703), .B(n25856), .Z(n25858) );
  XOR U25650 ( .A(n25865), .B(n25866), .Z(n25703) );
  AND U25651 ( .A(n670), .B(n25867), .Z(n25866) );
  XOR U25652 ( .A(n25850), .B(n25868), .Z(n25856) );
  AND U25653 ( .A(n25869), .B(n25853), .Z(n25868) );
  XNOR U25654 ( .A(n25762), .B(n25850), .Z(n25853) );
  XNOR U25655 ( .A(n25870), .B(n25871), .Z(n25762) );
  AND U25656 ( .A(n662), .B(n25872), .Z(n25871) );
  XOR U25657 ( .A(n25873), .B(n25870), .Z(n25872) );
  XNOR U25658 ( .A(n25874), .B(n25850), .Z(n25869) );
  IV U25659 ( .A(n25713), .Z(n25874) );
  XOR U25660 ( .A(n25875), .B(n25876), .Z(n25713) );
  AND U25661 ( .A(n670), .B(n25877), .Z(n25876) );
  XOR U25662 ( .A(n25878), .B(n25879), .Z(n25850) );
  AND U25663 ( .A(n25880), .B(n25881), .Z(n25879) );
  XNOR U25664 ( .A(n25787), .B(n25878), .Z(n25881) );
  XNOR U25665 ( .A(n25882), .B(n25883), .Z(n25787) );
  AND U25666 ( .A(n662), .B(n25884), .Z(n25883) );
  XNOR U25667 ( .A(n25885), .B(n25882), .Z(n25884) );
  XOR U25668 ( .A(n25878), .B(n25724), .Z(n25880) );
  XOR U25669 ( .A(n25886), .B(n25887), .Z(n25724) );
  AND U25670 ( .A(n670), .B(n25888), .Z(n25887) );
  XOR U25671 ( .A(n25889), .B(n25890), .Z(n25878) );
  AND U25672 ( .A(n25891), .B(n25892), .Z(n25890) );
  XNOR U25673 ( .A(n25889), .B(n25833), .Z(n25892) );
  XNOR U25674 ( .A(n25893), .B(n25894), .Z(n25833) );
  AND U25675 ( .A(n662), .B(n25895), .Z(n25894) );
  XOR U25676 ( .A(n25896), .B(n25893), .Z(n25895) );
  XNOR U25677 ( .A(n25897), .B(n25889), .Z(n25891) );
  IV U25678 ( .A(n25736), .Z(n25897) );
  XOR U25679 ( .A(n25898), .B(n25899), .Z(n25736) );
  AND U25680 ( .A(n670), .B(n25900), .Z(n25899) );
  AND U25681 ( .A(n25854), .B(n25843), .Z(n25889) );
  XNOR U25682 ( .A(n25901), .B(n25902), .Z(n25843) );
  AND U25683 ( .A(n662), .B(n25903), .Z(n25902) );
  XNOR U25684 ( .A(n25904), .B(n25901), .Z(n25903) );
  XNOR U25685 ( .A(n25905), .B(n25906), .Z(n662) );
  AND U25686 ( .A(n25907), .B(n25908), .Z(n25906) );
  XOR U25687 ( .A(n25864), .B(n25905), .Z(n25908) );
  AND U25688 ( .A(n25909), .B(n25910), .Z(n25864) );
  XOR U25689 ( .A(n25905), .B(n25861), .Z(n25907) );
  XNOR U25690 ( .A(n25911), .B(n25912), .Z(n25861) );
  AND U25691 ( .A(n666), .B(n25867), .Z(n25912) );
  XOR U25692 ( .A(n25865), .B(n25911), .Z(n25867) );
  XOR U25693 ( .A(n25913), .B(n25914), .Z(n25905) );
  AND U25694 ( .A(n25915), .B(n25916), .Z(n25914) );
  XNOR U25695 ( .A(n25913), .B(n25909), .Z(n25916) );
  IV U25696 ( .A(n25873), .Z(n25909) );
  XOR U25697 ( .A(n25917), .B(n25918), .Z(n25873) );
  XOR U25698 ( .A(n25919), .B(n25910), .Z(n25918) );
  AND U25699 ( .A(n25885), .B(n25920), .Z(n25910) );
  AND U25700 ( .A(n25921), .B(n25922), .Z(n25919) );
  XOR U25701 ( .A(n25923), .B(n25917), .Z(n25921) );
  XNOR U25702 ( .A(n25870), .B(n25913), .Z(n25915) );
  XNOR U25703 ( .A(n25924), .B(n25925), .Z(n25870) );
  AND U25704 ( .A(n666), .B(n25877), .Z(n25925) );
  XOR U25705 ( .A(n25924), .B(n25875), .Z(n25877) );
  XOR U25706 ( .A(n25926), .B(n25927), .Z(n25913) );
  AND U25707 ( .A(n25928), .B(n25929), .Z(n25927) );
  XNOR U25708 ( .A(n25926), .B(n25885), .Z(n25929) );
  XOR U25709 ( .A(n25930), .B(n25922), .Z(n25885) );
  XNOR U25710 ( .A(n25931), .B(n25917), .Z(n25922) );
  XOR U25711 ( .A(n25932), .B(n25933), .Z(n25917) );
  AND U25712 ( .A(n25934), .B(n25935), .Z(n25933) );
  XOR U25713 ( .A(n25936), .B(n25932), .Z(n25934) );
  XNOR U25714 ( .A(n25937), .B(n25938), .Z(n25931) );
  AND U25715 ( .A(n25939), .B(n25940), .Z(n25938) );
  XOR U25716 ( .A(n25937), .B(n25941), .Z(n25939) );
  XNOR U25717 ( .A(n25923), .B(n25920), .Z(n25930) );
  AND U25718 ( .A(n25942), .B(n25943), .Z(n25920) );
  XOR U25719 ( .A(n25944), .B(n25945), .Z(n25923) );
  AND U25720 ( .A(n25946), .B(n25947), .Z(n25945) );
  XOR U25721 ( .A(n25944), .B(n25948), .Z(n25946) );
  XNOR U25722 ( .A(n25882), .B(n25926), .Z(n25928) );
  XNOR U25723 ( .A(n25949), .B(n25950), .Z(n25882) );
  AND U25724 ( .A(n666), .B(n25888), .Z(n25950) );
  XOR U25725 ( .A(n25949), .B(n25886), .Z(n25888) );
  XOR U25726 ( .A(n25951), .B(n25952), .Z(n25926) );
  AND U25727 ( .A(n25953), .B(n25954), .Z(n25952) );
  XNOR U25728 ( .A(n25951), .B(n25942), .Z(n25954) );
  IV U25729 ( .A(n25896), .Z(n25942) );
  XNOR U25730 ( .A(n25955), .B(n25935), .Z(n25896) );
  XNOR U25731 ( .A(n25956), .B(n25941), .Z(n25935) );
  XOR U25732 ( .A(n25957), .B(n25958), .Z(n25941) );
  NOR U25733 ( .A(n25959), .B(n25960), .Z(n25958) );
  XNOR U25734 ( .A(n25957), .B(n25961), .Z(n25959) );
  XNOR U25735 ( .A(n25940), .B(n25932), .Z(n25956) );
  XOR U25736 ( .A(n25962), .B(n25963), .Z(n25932) );
  AND U25737 ( .A(n25964), .B(n25965), .Z(n25963) );
  XNOR U25738 ( .A(n25962), .B(n25966), .Z(n25964) );
  XNOR U25739 ( .A(n25967), .B(n25937), .Z(n25940) );
  XOR U25740 ( .A(n25968), .B(n25969), .Z(n25937) );
  AND U25741 ( .A(n25970), .B(n25971), .Z(n25969) );
  XOR U25742 ( .A(n25968), .B(n25972), .Z(n25970) );
  XNOR U25743 ( .A(n25973), .B(n25974), .Z(n25967) );
  NOR U25744 ( .A(n25975), .B(n25976), .Z(n25974) );
  XOR U25745 ( .A(n25973), .B(n25977), .Z(n25975) );
  XNOR U25746 ( .A(n25936), .B(n25943), .Z(n25955) );
  NOR U25747 ( .A(n25904), .B(n25978), .Z(n25943) );
  XOR U25748 ( .A(n25948), .B(n25947), .Z(n25936) );
  XNOR U25749 ( .A(n25979), .B(n25944), .Z(n25947) );
  XOR U25750 ( .A(n25980), .B(n25981), .Z(n25944) );
  AND U25751 ( .A(n25982), .B(n25983), .Z(n25981) );
  XOR U25752 ( .A(n25980), .B(n25984), .Z(n25982) );
  XNOR U25753 ( .A(n25985), .B(n25986), .Z(n25979) );
  NOR U25754 ( .A(n25987), .B(n25988), .Z(n25986) );
  XNOR U25755 ( .A(n25985), .B(n25989), .Z(n25987) );
  XOR U25756 ( .A(n25990), .B(n25991), .Z(n25948) );
  NOR U25757 ( .A(n25992), .B(n25993), .Z(n25991) );
  XNOR U25758 ( .A(n25990), .B(n25994), .Z(n25992) );
  XNOR U25759 ( .A(n25893), .B(n25951), .Z(n25953) );
  XNOR U25760 ( .A(n25995), .B(n25996), .Z(n25893) );
  AND U25761 ( .A(n666), .B(n25900), .Z(n25996) );
  XOR U25762 ( .A(n25995), .B(n25898), .Z(n25900) );
  AND U25763 ( .A(n25901), .B(n25904), .Z(n25951) );
  XOR U25764 ( .A(n25997), .B(n25978), .Z(n25904) );
  XNOR U25765 ( .A(p_input[2048]), .B(p_input[912]), .Z(n25978) );
  XOR U25766 ( .A(n25966), .B(n25965), .Z(n25997) );
  XNOR U25767 ( .A(n25998), .B(n25972), .Z(n25965) );
  XNOR U25768 ( .A(n25961), .B(n25960), .Z(n25972) );
  XOR U25769 ( .A(n25999), .B(n25957), .Z(n25960) );
  XNOR U25770 ( .A(n16904), .B(p_input[922]), .Z(n25957) );
  XNOR U25771 ( .A(p_input[2059]), .B(p_input[923]), .Z(n25999) );
  XOR U25772 ( .A(p_input[2060]), .B(p_input[924]), .Z(n25961) );
  XNOR U25773 ( .A(n25971), .B(n25962), .Z(n25998) );
  XNOR U25774 ( .A(n17068), .B(p_input[913]), .Z(n25962) );
  XOR U25775 ( .A(n26000), .B(n25977), .Z(n25971) );
  XNOR U25776 ( .A(p_input[2063]), .B(p_input[927]), .Z(n25977) );
  XOR U25777 ( .A(n25968), .B(n25976), .Z(n26000) );
  XOR U25778 ( .A(n26001), .B(n25973), .Z(n25976) );
  XOR U25779 ( .A(p_input[2061]), .B(p_input[925]), .Z(n25973) );
  XNOR U25780 ( .A(p_input[2062]), .B(p_input[926]), .Z(n26001) );
  XNOR U25781 ( .A(n16738), .B(p_input[921]), .Z(n25968) );
  XNOR U25782 ( .A(n25984), .B(n25983), .Z(n25966) );
  XNOR U25783 ( .A(n26002), .B(n25989), .Z(n25983) );
  XOR U25784 ( .A(p_input[2056]), .B(p_input[920]), .Z(n25989) );
  XOR U25785 ( .A(n25980), .B(n25988), .Z(n26002) );
  XOR U25786 ( .A(n26003), .B(n25985), .Z(n25988) );
  XOR U25787 ( .A(p_input[2054]), .B(p_input[918]), .Z(n25985) );
  XNOR U25788 ( .A(p_input[2055]), .B(p_input[919]), .Z(n26003) );
  XNOR U25789 ( .A(n16741), .B(p_input[914]), .Z(n25980) );
  XNOR U25790 ( .A(n25994), .B(n25993), .Z(n25984) );
  XOR U25791 ( .A(n26004), .B(n25990), .Z(n25993) );
  XOR U25792 ( .A(p_input[2051]), .B(p_input[915]), .Z(n25990) );
  XNOR U25793 ( .A(p_input[2052]), .B(p_input[916]), .Z(n26004) );
  XOR U25794 ( .A(p_input[2053]), .B(p_input[917]), .Z(n25994) );
  XNOR U25795 ( .A(n26005), .B(n26006), .Z(n25901) );
  AND U25796 ( .A(n666), .B(n26007), .Z(n26006) );
  XNOR U25797 ( .A(n26008), .B(n26009), .Z(n666) );
  AND U25798 ( .A(n26010), .B(n26011), .Z(n26009) );
  XOR U25799 ( .A(n26008), .B(n25911), .Z(n26011) );
  XNOR U25800 ( .A(n26008), .B(n25865), .Z(n26010) );
  XOR U25801 ( .A(n26012), .B(n26013), .Z(n26008) );
  AND U25802 ( .A(n26014), .B(n26015), .Z(n26013) );
  XOR U25803 ( .A(n26012), .B(n25875), .Z(n26014) );
  XOR U25804 ( .A(n26016), .B(n26017), .Z(n25854) );
  AND U25805 ( .A(n670), .B(n26007), .Z(n26017) );
  XNOR U25806 ( .A(n26005), .B(n26016), .Z(n26007) );
  XNOR U25807 ( .A(n26018), .B(n26019), .Z(n670) );
  AND U25808 ( .A(n26020), .B(n26021), .Z(n26019) );
  XNOR U25809 ( .A(n26022), .B(n26018), .Z(n26021) );
  IV U25810 ( .A(n25911), .Z(n26022) );
  XNOR U25811 ( .A(n26023), .B(n26024), .Z(n25911) );
  AND U25812 ( .A(n673), .B(n26025), .Z(n26024) );
  XNOR U25813 ( .A(n26023), .B(n26026), .Z(n26025) );
  XNOR U25814 ( .A(n25865), .B(n26018), .Z(n26020) );
  XOR U25815 ( .A(n26027), .B(n26028), .Z(n25865) );
  AND U25816 ( .A(n681), .B(n26029), .Z(n26028) );
  XOR U25817 ( .A(n26012), .B(n26030), .Z(n26018) );
  AND U25818 ( .A(n26031), .B(n26015), .Z(n26030) );
  XNOR U25819 ( .A(n25924), .B(n26012), .Z(n26015) );
  XNOR U25820 ( .A(n26032), .B(n26033), .Z(n25924) );
  AND U25821 ( .A(n673), .B(n26034), .Z(n26033) );
  XOR U25822 ( .A(n26035), .B(n26032), .Z(n26034) );
  XNOR U25823 ( .A(n26036), .B(n26012), .Z(n26031) );
  IV U25824 ( .A(n25875), .Z(n26036) );
  XOR U25825 ( .A(n26037), .B(n26038), .Z(n25875) );
  AND U25826 ( .A(n681), .B(n26039), .Z(n26038) );
  XOR U25827 ( .A(n26040), .B(n26041), .Z(n26012) );
  AND U25828 ( .A(n26042), .B(n26043), .Z(n26041) );
  XNOR U25829 ( .A(n25949), .B(n26040), .Z(n26043) );
  XNOR U25830 ( .A(n26044), .B(n26045), .Z(n25949) );
  AND U25831 ( .A(n673), .B(n26046), .Z(n26045) );
  XNOR U25832 ( .A(n26047), .B(n26044), .Z(n26046) );
  XOR U25833 ( .A(n26040), .B(n25886), .Z(n26042) );
  XOR U25834 ( .A(n26048), .B(n26049), .Z(n25886) );
  AND U25835 ( .A(n681), .B(n26050), .Z(n26049) );
  XOR U25836 ( .A(n26051), .B(n26052), .Z(n26040) );
  AND U25837 ( .A(n26053), .B(n26054), .Z(n26052) );
  XNOR U25838 ( .A(n26051), .B(n25995), .Z(n26054) );
  XNOR U25839 ( .A(n26055), .B(n26056), .Z(n25995) );
  AND U25840 ( .A(n673), .B(n26057), .Z(n26056) );
  XOR U25841 ( .A(n26058), .B(n26055), .Z(n26057) );
  XNOR U25842 ( .A(n26059), .B(n26051), .Z(n26053) );
  IV U25843 ( .A(n25898), .Z(n26059) );
  XOR U25844 ( .A(n26060), .B(n26061), .Z(n25898) );
  AND U25845 ( .A(n681), .B(n26062), .Z(n26061) );
  AND U25846 ( .A(n26016), .B(n26005), .Z(n26051) );
  XNOR U25847 ( .A(n26063), .B(n26064), .Z(n26005) );
  AND U25848 ( .A(n673), .B(n26065), .Z(n26064) );
  XNOR U25849 ( .A(n26066), .B(n26063), .Z(n26065) );
  XNOR U25850 ( .A(n26067), .B(n26068), .Z(n673) );
  AND U25851 ( .A(n26069), .B(n26070), .Z(n26068) );
  XOR U25852 ( .A(n26026), .B(n26067), .Z(n26070) );
  AND U25853 ( .A(n26071), .B(n26072), .Z(n26026) );
  XOR U25854 ( .A(n26067), .B(n26023), .Z(n26069) );
  XNOR U25855 ( .A(n26073), .B(n26074), .Z(n26023) );
  AND U25856 ( .A(n677), .B(n26029), .Z(n26074) );
  XOR U25857 ( .A(n26027), .B(n26073), .Z(n26029) );
  XOR U25858 ( .A(n26075), .B(n26076), .Z(n26067) );
  AND U25859 ( .A(n26077), .B(n26078), .Z(n26076) );
  XNOR U25860 ( .A(n26075), .B(n26071), .Z(n26078) );
  IV U25861 ( .A(n26035), .Z(n26071) );
  XOR U25862 ( .A(n26079), .B(n26080), .Z(n26035) );
  XOR U25863 ( .A(n26081), .B(n26072), .Z(n26080) );
  AND U25864 ( .A(n26047), .B(n26082), .Z(n26072) );
  AND U25865 ( .A(n26083), .B(n26084), .Z(n26081) );
  XOR U25866 ( .A(n26085), .B(n26079), .Z(n26083) );
  XNOR U25867 ( .A(n26032), .B(n26075), .Z(n26077) );
  XNOR U25868 ( .A(n26086), .B(n26087), .Z(n26032) );
  AND U25869 ( .A(n677), .B(n26039), .Z(n26087) );
  XOR U25870 ( .A(n26086), .B(n26037), .Z(n26039) );
  XOR U25871 ( .A(n26088), .B(n26089), .Z(n26075) );
  AND U25872 ( .A(n26090), .B(n26091), .Z(n26089) );
  XNOR U25873 ( .A(n26088), .B(n26047), .Z(n26091) );
  XOR U25874 ( .A(n26092), .B(n26084), .Z(n26047) );
  XNOR U25875 ( .A(n26093), .B(n26079), .Z(n26084) );
  XOR U25876 ( .A(n26094), .B(n26095), .Z(n26079) );
  AND U25877 ( .A(n26096), .B(n26097), .Z(n26095) );
  XOR U25878 ( .A(n26098), .B(n26094), .Z(n26096) );
  XNOR U25879 ( .A(n26099), .B(n26100), .Z(n26093) );
  AND U25880 ( .A(n26101), .B(n26102), .Z(n26100) );
  XOR U25881 ( .A(n26099), .B(n26103), .Z(n26101) );
  XNOR U25882 ( .A(n26085), .B(n26082), .Z(n26092) );
  AND U25883 ( .A(n26104), .B(n26105), .Z(n26082) );
  XOR U25884 ( .A(n26106), .B(n26107), .Z(n26085) );
  AND U25885 ( .A(n26108), .B(n26109), .Z(n26107) );
  XOR U25886 ( .A(n26106), .B(n26110), .Z(n26108) );
  XNOR U25887 ( .A(n26044), .B(n26088), .Z(n26090) );
  XNOR U25888 ( .A(n26111), .B(n26112), .Z(n26044) );
  AND U25889 ( .A(n677), .B(n26050), .Z(n26112) );
  XOR U25890 ( .A(n26111), .B(n26048), .Z(n26050) );
  XOR U25891 ( .A(n26113), .B(n26114), .Z(n26088) );
  AND U25892 ( .A(n26115), .B(n26116), .Z(n26114) );
  XNOR U25893 ( .A(n26113), .B(n26104), .Z(n26116) );
  IV U25894 ( .A(n26058), .Z(n26104) );
  XNOR U25895 ( .A(n26117), .B(n26097), .Z(n26058) );
  XNOR U25896 ( .A(n26118), .B(n26103), .Z(n26097) );
  XOR U25897 ( .A(n26119), .B(n26120), .Z(n26103) );
  NOR U25898 ( .A(n26121), .B(n26122), .Z(n26120) );
  XNOR U25899 ( .A(n26119), .B(n26123), .Z(n26121) );
  XNOR U25900 ( .A(n26102), .B(n26094), .Z(n26118) );
  XOR U25901 ( .A(n26124), .B(n26125), .Z(n26094) );
  AND U25902 ( .A(n26126), .B(n26127), .Z(n26125) );
  XNOR U25903 ( .A(n26124), .B(n26128), .Z(n26126) );
  XNOR U25904 ( .A(n26129), .B(n26099), .Z(n26102) );
  XOR U25905 ( .A(n26130), .B(n26131), .Z(n26099) );
  AND U25906 ( .A(n26132), .B(n26133), .Z(n26131) );
  XOR U25907 ( .A(n26130), .B(n26134), .Z(n26132) );
  XNOR U25908 ( .A(n26135), .B(n26136), .Z(n26129) );
  NOR U25909 ( .A(n26137), .B(n26138), .Z(n26136) );
  XOR U25910 ( .A(n26135), .B(n26139), .Z(n26137) );
  XNOR U25911 ( .A(n26098), .B(n26105), .Z(n26117) );
  NOR U25912 ( .A(n26066), .B(n26140), .Z(n26105) );
  XOR U25913 ( .A(n26110), .B(n26109), .Z(n26098) );
  XNOR U25914 ( .A(n26141), .B(n26106), .Z(n26109) );
  XOR U25915 ( .A(n26142), .B(n26143), .Z(n26106) );
  AND U25916 ( .A(n26144), .B(n26145), .Z(n26143) );
  XOR U25917 ( .A(n26142), .B(n26146), .Z(n26144) );
  XNOR U25918 ( .A(n26147), .B(n26148), .Z(n26141) );
  NOR U25919 ( .A(n26149), .B(n26150), .Z(n26148) );
  XNOR U25920 ( .A(n26147), .B(n26151), .Z(n26149) );
  XOR U25921 ( .A(n26152), .B(n26153), .Z(n26110) );
  NOR U25922 ( .A(n26154), .B(n26155), .Z(n26153) );
  XNOR U25923 ( .A(n26152), .B(n26156), .Z(n26154) );
  XNOR U25924 ( .A(n26055), .B(n26113), .Z(n26115) );
  XNOR U25925 ( .A(n26157), .B(n26158), .Z(n26055) );
  AND U25926 ( .A(n677), .B(n26062), .Z(n26158) );
  XOR U25927 ( .A(n26157), .B(n26060), .Z(n26062) );
  AND U25928 ( .A(n26063), .B(n26066), .Z(n26113) );
  XOR U25929 ( .A(n26159), .B(n26140), .Z(n26066) );
  XNOR U25930 ( .A(p_input[2048]), .B(p_input[928]), .Z(n26140) );
  XOR U25931 ( .A(n26128), .B(n26127), .Z(n26159) );
  XNOR U25932 ( .A(n26160), .B(n26134), .Z(n26127) );
  XNOR U25933 ( .A(n26123), .B(n26122), .Z(n26134) );
  XOR U25934 ( .A(n26161), .B(n26119), .Z(n26122) );
  XNOR U25935 ( .A(n16904), .B(p_input[938]), .Z(n26119) );
  XNOR U25936 ( .A(p_input[2059]), .B(p_input[939]), .Z(n26161) );
  XOR U25937 ( .A(p_input[2060]), .B(p_input[940]), .Z(n26123) );
  XNOR U25938 ( .A(n26133), .B(n26124), .Z(n26160) );
  XNOR U25939 ( .A(n17068), .B(p_input[929]), .Z(n26124) );
  XOR U25940 ( .A(n26162), .B(n26139), .Z(n26133) );
  XNOR U25941 ( .A(p_input[2063]), .B(p_input[943]), .Z(n26139) );
  XOR U25942 ( .A(n26130), .B(n26138), .Z(n26162) );
  XOR U25943 ( .A(n26163), .B(n26135), .Z(n26138) );
  XOR U25944 ( .A(p_input[2061]), .B(p_input[941]), .Z(n26135) );
  XNOR U25945 ( .A(p_input[2062]), .B(p_input[942]), .Z(n26163) );
  XNOR U25946 ( .A(n16738), .B(p_input[937]), .Z(n26130) );
  XNOR U25947 ( .A(n26146), .B(n26145), .Z(n26128) );
  XNOR U25948 ( .A(n26164), .B(n26151), .Z(n26145) );
  XOR U25949 ( .A(p_input[2056]), .B(p_input[936]), .Z(n26151) );
  XOR U25950 ( .A(n26142), .B(n26150), .Z(n26164) );
  XOR U25951 ( .A(n26165), .B(n26147), .Z(n26150) );
  XOR U25952 ( .A(p_input[2054]), .B(p_input[934]), .Z(n26147) );
  XNOR U25953 ( .A(p_input[2055]), .B(p_input[935]), .Z(n26165) );
  XNOR U25954 ( .A(n16741), .B(p_input[930]), .Z(n26142) );
  XNOR U25955 ( .A(n26156), .B(n26155), .Z(n26146) );
  XOR U25956 ( .A(n26166), .B(n26152), .Z(n26155) );
  XOR U25957 ( .A(p_input[2051]), .B(p_input[931]), .Z(n26152) );
  XNOR U25958 ( .A(p_input[2052]), .B(p_input[932]), .Z(n26166) );
  XOR U25959 ( .A(p_input[2053]), .B(p_input[933]), .Z(n26156) );
  XNOR U25960 ( .A(n26167), .B(n26168), .Z(n26063) );
  AND U25961 ( .A(n677), .B(n26169), .Z(n26168) );
  XNOR U25962 ( .A(n26170), .B(n26171), .Z(n677) );
  AND U25963 ( .A(n26172), .B(n26173), .Z(n26171) );
  XOR U25964 ( .A(n26170), .B(n26073), .Z(n26173) );
  XNOR U25965 ( .A(n26170), .B(n26027), .Z(n26172) );
  XOR U25966 ( .A(n26174), .B(n26175), .Z(n26170) );
  AND U25967 ( .A(n26176), .B(n26177), .Z(n26175) );
  XOR U25968 ( .A(n26174), .B(n26037), .Z(n26176) );
  XOR U25969 ( .A(n26178), .B(n26179), .Z(n26016) );
  AND U25970 ( .A(n681), .B(n26169), .Z(n26179) );
  XNOR U25971 ( .A(n26167), .B(n26178), .Z(n26169) );
  XNOR U25972 ( .A(n26180), .B(n26181), .Z(n681) );
  AND U25973 ( .A(n26182), .B(n26183), .Z(n26181) );
  XNOR U25974 ( .A(n26184), .B(n26180), .Z(n26183) );
  IV U25975 ( .A(n26073), .Z(n26184) );
  XNOR U25976 ( .A(n26185), .B(n26186), .Z(n26073) );
  AND U25977 ( .A(n684), .B(n26187), .Z(n26186) );
  XNOR U25978 ( .A(n26185), .B(n26188), .Z(n26187) );
  XNOR U25979 ( .A(n26027), .B(n26180), .Z(n26182) );
  XOR U25980 ( .A(n26189), .B(n26190), .Z(n26027) );
  AND U25981 ( .A(n692), .B(n26191), .Z(n26190) );
  XOR U25982 ( .A(n26174), .B(n26192), .Z(n26180) );
  AND U25983 ( .A(n26193), .B(n26177), .Z(n26192) );
  XNOR U25984 ( .A(n26086), .B(n26174), .Z(n26177) );
  XNOR U25985 ( .A(n26194), .B(n26195), .Z(n26086) );
  AND U25986 ( .A(n684), .B(n26196), .Z(n26195) );
  XOR U25987 ( .A(n26197), .B(n26194), .Z(n26196) );
  XNOR U25988 ( .A(n26198), .B(n26174), .Z(n26193) );
  IV U25989 ( .A(n26037), .Z(n26198) );
  XOR U25990 ( .A(n26199), .B(n26200), .Z(n26037) );
  AND U25991 ( .A(n692), .B(n26201), .Z(n26200) );
  XOR U25992 ( .A(n26202), .B(n26203), .Z(n26174) );
  AND U25993 ( .A(n26204), .B(n26205), .Z(n26203) );
  XNOR U25994 ( .A(n26111), .B(n26202), .Z(n26205) );
  XNOR U25995 ( .A(n26206), .B(n26207), .Z(n26111) );
  AND U25996 ( .A(n684), .B(n26208), .Z(n26207) );
  XNOR U25997 ( .A(n26209), .B(n26206), .Z(n26208) );
  XOR U25998 ( .A(n26202), .B(n26048), .Z(n26204) );
  XOR U25999 ( .A(n26210), .B(n26211), .Z(n26048) );
  AND U26000 ( .A(n692), .B(n26212), .Z(n26211) );
  XOR U26001 ( .A(n26213), .B(n26214), .Z(n26202) );
  AND U26002 ( .A(n26215), .B(n26216), .Z(n26214) );
  XNOR U26003 ( .A(n26213), .B(n26157), .Z(n26216) );
  XNOR U26004 ( .A(n26217), .B(n26218), .Z(n26157) );
  AND U26005 ( .A(n684), .B(n26219), .Z(n26218) );
  XOR U26006 ( .A(n26220), .B(n26217), .Z(n26219) );
  XNOR U26007 ( .A(n26221), .B(n26213), .Z(n26215) );
  IV U26008 ( .A(n26060), .Z(n26221) );
  XOR U26009 ( .A(n26222), .B(n26223), .Z(n26060) );
  AND U26010 ( .A(n692), .B(n26224), .Z(n26223) );
  AND U26011 ( .A(n26178), .B(n26167), .Z(n26213) );
  XNOR U26012 ( .A(n26225), .B(n26226), .Z(n26167) );
  AND U26013 ( .A(n684), .B(n26227), .Z(n26226) );
  XNOR U26014 ( .A(n26228), .B(n26225), .Z(n26227) );
  XNOR U26015 ( .A(n26229), .B(n26230), .Z(n684) );
  AND U26016 ( .A(n26231), .B(n26232), .Z(n26230) );
  XOR U26017 ( .A(n26188), .B(n26229), .Z(n26232) );
  AND U26018 ( .A(n26233), .B(n26234), .Z(n26188) );
  XOR U26019 ( .A(n26229), .B(n26185), .Z(n26231) );
  XNOR U26020 ( .A(n26235), .B(n26236), .Z(n26185) );
  AND U26021 ( .A(n688), .B(n26191), .Z(n26236) );
  XOR U26022 ( .A(n26189), .B(n26235), .Z(n26191) );
  XOR U26023 ( .A(n26237), .B(n26238), .Z(n26229) );
  AND U26024 ( .A(n26239), .B(n26240), .Z(n26238) );
  XNOR U26025 ( .A(n26237), .B(n26233), .Z(n26240) );
  IV U26026 ( .A(n26197), .Z(n26233) );
  XOR U26027 ( .A(n26241), .B(n26242), .Z(n26197) );
  XOR U26028 ( .A(n26243), .B(n26234), .Z(n26242) );
  AND U26029 ( .A(n26209), .B(n26244), .Z(n26234) );
  AND U26030 ( .A(n26245), .B(n26246), .Z(n26243) );
  XOR U26031 ( .A(n26247), .B(n26241), .Z(n26245) );
  XNOR U26032 ( .A(n26194), .B(n26237), .Z(n26239) );
  XNOR U26033 ( .A(n26248), .B(n26249), .Z(n26194) );
  AND U26034 ( .A(n688), .B(n26201), .Z(n26249) );
  XOR U26035 ( .A(n26248), .B(n26199), .Z(n26201) );
  XOR U26036 ( .A(n26250), .B(n26251), .Z(n26237) );
  AND U26037 ( .A(n26252), .B(n26253), .Z(n26251) );
  XNOR U26038 ( .A(n26250), .B(n26209), .Z(n26253) );
  XOR U26039 ( .A(n26254), .B(n26246), .Z(n26209) );
  XNOR U26040 ( .A(n26255), .B(n26241), .Z(n26246) );
  XOR U26041 ( .A(n26256), .B(n26257), .Z(n26241) );
  AND U26042 ( .A(n26258), .B(n26259), .Z(n26257) );
  XOR U26043 ( .A(n26260), .B(n26256), .Z(n26258) );
  XNOR U26044 ( .A(n26261), .B(n26262), .Z(n26255) );
  AND U26045 ( .A(n26263), .B(n26264), .Z(n26262) );
  XOR U26046 ( .A(n26261), .B(n26265), .Z(n26263) );
  XNOR U26047 ( .A(n26247), .B(n26244), .Z(n26254) );
  AND U26048 ( .A(n26266), .B(n26267), .Z(n26244) );
  XOR U26049 ( .A(n26268), .B(n26269), .Z(n26247) );
  AND U26050 ( .A(n26270), .B(n26271), .Z(n26269) );
  XOR U26051 ( .A(n26268), .B(n26272), .Z(n26270) );
  XNOR U26052 ( .A(n26206), .B(n26250), .Z(n26252) );
  XNOR U26053 ( .A(n26273), .B(n26274), .Z(n26206) );
  AND U26054 ( .A(n688), .B(n26212), .Z(n26274) );
  XOR U26055 ( .A(n26273), .B(n26210), .Z(n26212) );
  XOR U26056 ( .A(n26275), .B(n26276), .Z(n26250) );
  AND U26057 ( .A(n26277), .B(n26278), .Z(n26276) );
  XNOR U26058 ( .A(n26275), .B(n26266), .Z(n26278) );
  IV U26059 ( .A(n26220), .Z(n26266) );
  XNOR U26060 ( .A(n26279), .B(n26259), .Z(n26220) );
  XNOR U26061 ( .A(n26280), .B(n26265), .Z(n26259) );
  XOR U26062 ( .A(n26281), .B(n26282), .Z(n26265) );
  NOR U26063 ( .A(n26283), .B(n26284), .Z(n26282) );
  XNOR U26064 ( .A(n26281), .B(n26285), .Z(n26283) );
  XNOR U26065 ( .A(n26264), .B(n26256), .Z(n26280) );
  XOR U26066 ( .A(n26286), .B(n26287), .Z(n26256) );
  AND U26067 ( .A(n26288), .B(n26289), .Z(n26287) );
  XNOR U26068 ( .A(n26286), .B(n26290), .Z(n26288) );
  XNOR U26069 ( .A(n26291), .B(n26261), .Z(n26264) );
  XOR U26070 ( .A(n26292), .B(n26293), .Z(n26261) );
  AND U26071 ( .A(n26294), .B(n26295), .Z(n26293) );
  XOR U26072 ( .A(n26292), .B(n26296), .Z(n26294) );
  XNOR U26073 ( .A(n26297), .B(n26298), .Z(n26291) );
  NOR U26074 ( .A(n26299), .B(n26300), .Z(n26298) );
  XOR U26075 ( .A(n26297), .B(n26301), .Z(n26299) );
  XNOR U26076 ( .A(n26260), .B(n26267), .Z(n26279) );
  NOR U26077 ( .A(n26228), .B(n26302), .Z(n26267) );
  XOR U26078 ( .A(n26272), .B(n26271), .Z(n26260) );
  XNOR U26079 ( .A(n26303), .B(n26268), .Z(n26271) );
  XOR U26080 ( .A(n26304), .B(n26305), .Z(n26268) );
  AND U26081 ( .A(n26306), .B(n26307), .Z(n26305) );
  XOR U26082 ( .A(n26304), .B(n26308), .Z(n26306) );
  XNOR U26083 ( .A(n26309), .B(n26310), .Z(n26303) );
  NOR U26084 ( .A(n26311), .B(n26312), .Z(n26310) );
  XNOR U26085 ( .A(n26309), .B(n26313), .Z(n26311) );
  XOR U26086 ( .A(n26314), .B(n26315), .Z(n26272) );
  NOR U26087 ( .A(n26316), .B(n26317), .Z(n26315) );
  XNOR U26088 ( .A(n26314), .B(n26318), .Z(n26316) );
  XNOR U26089 ( .A(n26217), .B(n26275), .Z(n26277) );
  XNOR U26090 ( .A(n26319), .B(n26320), .Z(n26217) );
  AND U26091 ( .A(n688), .B(n26224), .Z(n26320) );
  XOR U26092 ( .A(n26319), .B(n26222), .Z(n26224) );
  AND U26093 ( .A(n26225), .B(n26228), .Z(n26275) );
  XOR U26094 ( .A(n26321), .B(n26302), .Z(n26228) );
  XNOR U26095 ( .A(p_input[2048]), .B(p_input[944]), .Z(n26302) );
  XOR U26096 ( .A(n26290), .B(n26289), .Z(n26321) );
  XNOR U26097 ( .A(n26322), .B(n26296), .Z(n26289) );
  XNOR U26098 ( .A(n26285), .B(n26284), .Z(n26296) );
  XOR U26099 ( .A(n26323), .B(n26281), .Z(n26284) );
  XNOR U26100 ( .A(n16904), .B(p_input[954]), .Z(n26281) );
  XNOR U26101 ( .A(p_input[2059]), .B(p_input[955]), .Z(n26323) );
  XOR U26102 ( .A(p_input[2060]), .B(p_input[956]), .Z(n26285) );
  XNOR U26103 ( .A(n26295), .B(n26286), .Z(n26322) );
  XNOR U26104 ( .A(n17068), .B(p_input[945]), .Z(n26286) );
  XOR U26105 ( .A(n26324), .B(n26301), .Z(n26295) );
  XNOR U26106 ( .A(p_input[2063]), .B(p_input[959]), .Z(n26301) );
  XOR U26107 ( .A(n26292), .B(n26300), .Z(n26324) );
  XOR U26108 ( .A(n26325), .B(n26297), .Z(n26300) );
  XOR U26109 ( .A(p_input[2061]), .B(p_input[957]), .Z(n26297) );
  XNOR U26110 ( .A(p_input[2062]), .B(p_input[958]), .Z(n26325) );
  XNOR U26111 ( .A(n16738), .B(p_input[953]), .Z(n26292) );
  XNOR U26112 ( .A(n26308), .B(n26307), .Z(n26290) );
  XNOR U26113 ( .A(n26326), .B(n26313), .Z(n26307) );
  XOR U26114 ( .A(p_input[2056]), .B(p_input[952]), .Z(n26313) );
  XOR U26115 ( .A(n26304), .B(n26312), .Z(n26326) );
  XOR U26116 ( .A(n26327), .B(n26309), .Z(n26312) );
  XOR U26117 ( .A(p_input[2054]), .B(p_input[950]), .Z(n26309) );
  XNOR U26118 ( .A(p_input[2055]), .B(p_input[951]), .Z(n26327) );
  XNOR U26119 ( .A(n16741), .B(p_input[946]), .Z(n26304) );
  XNOR U26120 ( .A(n26318), .B(n26317), .Z(n26308) );
  XOR U26121 ( .A(n26328), .B(n26314), .Z(n26317) );
  XOR U26122 ( .A(p_input[2051]), .B(p_input[947]), .Z(n26314) );
  XNOR U26123 ( .A(p_input[2052]), .B(p_input[948]), .Z(n26328) );
  XOR U26124 ( .A(p_input[2053]), .B(p_input[949]), .Z(n26318) );
  XNOR U26125 ( .A(n26329), .B(n26330), .Z(n26225) );
  AND U26126 ( .A(n688), .B(n26331), .Z(n26330) );
  XNOR U26127 ( .A(n26332), .B(n26333), .Z(n688) );
  AND U26128 ( .A(n26334), .B(n26335), .Z(n26333) );
  XOR U26129 ( .A(n26332), .B(n26235), .Z(n26335) );
  XNOR U26130 ( .A(n26332), .B(n26189), .Z(n26334) );
  XOR U26131 ( .A(n26336), .B(n26337), .Z(n26332) );
  AND U26132 ( .A(n26338), .B(n26339), .Z(n26337) );
  XOR U26133 ( .A(n26336), .B(n26199), .Z(n26338) );
  XOR U26134 ( .A(n26340), .B(n26341), .Z(n26178) );
  AND U26135 ( .A(n692), .B(n26331), .Z(n26341) );
  XNOR U26136 ( .A(n26329), .B(n26340), .Z(n26331) );
  XNOR U26137 ( .A(n26342), .B(n26343), .Z(n692) );
  AND U26138 ( .A(n26344), .B(n26345), .Z(n26343) );
  XNOR U26139 ( .A(n26346), .B(n26342), .Z(n26345) );
  IV U26140 ( .A(n26235), .Z(n26346) );
  XNOR U26141 ( .A(n26347), .B(n26348), .Z(n26235) );
  AND U26142 ( .A(n695), .B(n26349), .Z(n26348) );
  XNOR U26143 ( .A(n26347), .B(n26350), .Z(n26349) );
  XNOR U26144 ( .A(n26189), .B(n26342), .Z(n26344) );
  XOR U26145 ( .A(n26351), .B(n26352), .Z(n26189) );
  AND U26146 ( .A(n703), .B(n26353), .Z(n26352) );
  XOR U26147 ( .A(n26336), .B(n26354), .Z(n26342) );
  AND U26148 ( .A(n26355), .B(n26339), .Z(n26354) );
  XNOR U26149 ( .A(n26248), .B(n26336), .Z(n26339) );
  XNOR U26150 ( .A(n26356), .B(n26357), .Z(n26248) );
  AND U26151 ( .A(n695), .B(n26358), .Z(n26357) );
  XOR U26152 ( .A(n26359), .B(n26356), .Z(n26358) );
  XNOR U26153 ( .A(n26360), .B(n26336), .Z(n26355) );
  IV U26154 ( .A(n26199), .Z(n26360) );
  XOR U26155 ( .A(n26361), .B(n26362), .Z(n26199) );
  AND U26156 ( .A(n703), .B(n26363), .Z(n26362) );
  XOR U26157 ( .A(n26364), .B(n26365), .Z(n26336) );
  AND U26158 ( .A(n26366), .B(n26367), .Z(n26365) );
  XNOR U26159 ( .A(n26273), .B(n26364), .Z(n26367) );
  XNOR U26160 ( .A(n26368), .B(n26369), .Z(n26273) );
  AND U26161 ( .A(n695), .B(n26370), .Z(n26369) );
  XNOR U26162 ( .A(n26371), .B(n26368), .Z(n26370) );
  XOR U26163 ( .A(n26364), .B(n26210), .Z(n26366) );
  XOR U26164 ( .A(n26372), .B(n26373), .Z(n26210) );
  AND U26165 ( .A(n703), .B(n26374), .Z(n26373) );
  XOR U26166 ( .A(n26375), .B(n26376), .Z(n26364) );
  AND U26167 ( .A(n26377), .B(n26378), .Z(n26376) );
  XNOR U26168 ( .A(n26375), .B(n26319), .Z(n26378) );
  XNOR U26169 ( .A(n26379), .B(n26380), .Z(n26319) );
  AND U26170 ( .A(n695), .B(n26381), .Z(n26380) );
  XOR U26171 ( .A(n26382), .B(n26379), .Z(n26381) );
  XNOR U26172 ( .A(n26383), .B(n26375), .Z(n26377) );
  IV U26173 ( .A(n26222), .Z(n26383) );
  XOR U26174 ( .A(n26384), .B(n26385), .Z(n26222) );
  AND U26175 ( .A(n703), .B(n26386), .Z(n26385) );
  AND U26176 ( .A(n26340), .B(n26329), .Z(n26375) );
  XNOR U26177 ( .A(n26387), .B(n26388), .Z(n26329) );
  AND U26178 ( .A(n695), .B(n26389), .Z(n26388) );
  XNOR U26179 ( .A(n26390), .B(n26387), .Z(n26389) );
  XNOR U26180 ( .A(n26391), .B(n26392), .Z(n695) );
  AND U26181 ( .A(n26393), .B(n26394), .Z(n26392) );
  XOR U26182 ( .A(n26350), .B(n26391), .Z(n26394) );
  AND U26183 ( .A(n26395), .B(n26396), .Z(n26350) );
  XOR U26184 ( .A(n26391), .B(n26347), .Z(n26393) );
  XNOR U26185 ( .A(n26397), .B(n26398), .Z(n26347) );
  AND U26186 ( .A(n699), .B(n26353), .Z(n26398) );
  XOR U26187 ( .A(n26351), .B(n26397), .Z(n26353) );
  XOR U26188 ( .A(n26399), .B(n26400), .Z(n26391) );
  AND U26189 ( .A(n26401), .B(n26402), .Z(n26400) );
  XNOR U26190 ( .A(n26399), .B(n26395), .Z(n26402) );
  IV U26191 ( .A(n26359), .Z(n26395) );
  XOR U26192 ( .A(n26403), .B(n26404), .Z(n26359) );
  XOR U26193 ( .A(n26405), .B(n26396), .Z(n26404) );
  AND U26194 ( .A(n26371), .B(n26406), .Z(n26396) );
  AND U26195 ( .A(n26407), .B(n26408), .Z(n26405) );
  XOR U26196 ( .A(n26409), .B(n26403), .Z(n26407) );
  XNOR U26197 ( .A(n26356), .B(n26399), .Z(n26401) );
  XNOR U26198 ( .A(n26410), .B(n26411), .Z(n26356) );
  AND U26199 ( .A(n699), .B(n26363), .Z(n26411) );
  XOR U26200 ( .A(n26410), .B(n26361), .Z(n26363) );
  XOR U26201 ( .A(n26412), .B(n26413), .Z(n26399) );
  AND U26202 ( .A(n26414), .B(n26415), .Z(n26413) );
  XNOR U26203 ( .A(n26412), .B(n26371), .Z(n26415) );
  XOR U26204 ( .A(n26416), .B(n26408), .Z(n26371) );
  XNOR U26205 ( .A(n26417), .B(n26403), .Z(n26408) );
  XOR U26206 ( .A(n26418), .B(n26419), .Z(n26403) );
  AND U26207 ( .A(n26420), .B(n26421), .Z(n26419) );
  XOR U26208 ( .A(n26422), .B(n26418), .Z(n26420) );
  XNOR U26209 ( .A(n26423), .B(n26424), .Z(n26417) );
  AND U26210 ( .A(n26425), .B(n26426), .Z(n26424) );
  XOR U26211 ( .A(n26423), .B(n26427), .Z(n26425) );
  XNOR U26212 ( .A(n26409), .B(n26406), .Z(n26416) );
  AND U26213 ( .A(n26428), .B(n26429), .Z(n26406) );
  XOR U26214 ( .A(n26430), .B(n26431), .Z(n26409) );
  AND U26215 ( .A(n26432), .B(n26433), .Z(n26431) );
  XOR U26216 ( .A(n26430), .B(n26434), .Z(n26432) );
  XNOR U26217 ( .A(n26368), .B(n26412), .Z(n26414) );
  XNOR U26218 ( .A(n26435), .B(n26436), .Z(n26368) );
  AND U26219 ( .A(n699), .B(n26374), .Z(n26436) );
  XOR U26220 ( .A(n26435), .B(n26372), .Z(n26374) );
  XOR U26221 ( .A(n26437), .B(n26438), .Z(n26412) );
  AND U26222 ( .A(n26439), .B(n26440), .Z(n26438) );
  XNOR U26223 ( .A(n26437), .B(n26428), .Z(n26440) );
  IV U26224 ( .A(n26382), .Z(n26428) );
  XNOR U26225 ( .A(n26441), .B(n26421), .Z(n26382) );
  XNOR U26226 ( .A(n26442), .B(n26427), .Z(n26421) );
  XOR U26227 ( .A(n26443), .B(n26444), .Z(n26427) );
  NOR U26228 ( .A(n26445), .B(n26446), .Z(n26444) );
  XNOR U26229 ( .A(n26443), .B(n26447), .Z(n26445) );
  XNOR U26230 ( .A(n26426), .B(n26418), .Z(n26442) );
  XOR U26231 ( .A(n26448), .B(n26449), .Z(n26418) );
  AND U26232 ( .A(n26450), .B(n26451), .Z(n26449) );
  XNOR U26233 ( .A(n26448), .B(n26452), .Z(n26450) );
  XNOR U26234 ( .A(n26453), .B(n26423), .Z(n26426) );
  XOR U26235 ( .A(n26454), .B(n26455), .Z(n26423) );
  AND U26236 ( .A(n26456), .B(n26457), .Z(n26455) );
  XOR U26237 ( .A(n26454), .B(n26458), .Z(n26456) );
  XNOR U26238 ( .A(n26459), .B(n26460), .Z(n26453) );
  NOR U26239 ( .A(n26461), .B(n26462), .Z(n26460) );
  XOR U26240 ( .A(n26459), .B(n26463), .Z(n26461) );
  XNOR U26241 ( .A(n26422), .B(n26429), .Z(n26441) );
  NOR U26242 ( .A(n26390), .B(n26464), .Z(n26429) );
  XOR U26243 ( .A(n26434), .B(n26433), .Z(n26422) );
  XNOR U26244 ( .A(n26465), .B(n26430), .Z(n26433) );
  XOR U26245 ( .A(n26466), .B(n26467), .Z(n26430) );
  AND U26246 ( .A(n26468), .B(n26469), .Z(n26467) );
  XOR U26247 ( .A(n26466), .B(n26470), .Z(n26468) );
  XNOR U26248 ( .A(n26471), .B(n26472), .Z(n26465) );
  NOR U26249 ( .A(n26473), .B(n26474), .Z(n26472) );
  XNOR U26250 ( .A(n26471), .B(n26475), .Z(n26473) );
  XOR U26251 ( .A(n26476), .B(n26477), .Z(n26434) );
  NOR U26252 ( .A(n26478), .B(n26479), .Z(n26477) );
  XNOR U26253 ( .A(n26476), .B(n26480), .Z(n26478) );
  XNOR U26254 ( .A(n26379), .B(n26437), .Z(n26439) );
  XNOR U26255 ( .A(n26481), .B(n26482), .Z(n26379) );
  AND U26256 ( .A(n699), .B(n26386), .Z(n26482) );
  XOR U26257 ( .A(n26481), .B(n26384), .Z(n26386) );
  AND U26258 ( .A(n26387), .B(n26390), .Z(n26437) );
  XOR U26259 ( .A(n26483), .B(n26464), .Z(n26390) );
  XNOR U26260 ( .A(p_input[2048]), .B(p_input[960]), .Z(n26464) );
  XOR U26261 ( .A(n26452), .B(n26451), .Z(n26483) );
  XNOR U26262 ( .A(n26484), .B(n26458), .Z(n26451) );
  XNOR U26263 ( .A(n26447), .B(n26446), .Z(n26458) );
  XOR U26264 ( .A(n26485), .B(n26443), .Z(n26446) );
  XNOR U26265 ( .A(n16904), .B(p_input[970]), .Z(n26443) );
  XNOR U26266 ( .A(p_input[2059]), .B(p_input[971]), .Z(n26485) );
  XOR U26267 ( .A(p_input[2060]), .B(p_input[972]), .Z(n26447) );
  XNOR U26268 ( .A(n26457), .B(n26448), .Z(n26484) );
  XNOR U26269 ( .A(n17068), .B(p_input[961]), .Z(n26448) );
  XOR U26270 ( .A(n26486), .B(n26463), .Z(n26457) );
  XNOR U26271 ( .A(p_input[2063]), .B(p_input[975]), .Z(n26463) );
  XOR U26272 ( .A(n26454), .B(n26462), .Z(n26486) );
  XOR U26273 ( .A(n26487), .B(n26459), .Z(n26462) );
  XOR U26274 ( .A(p_input[2061]), .B(p_input[973]), .Z(n26459) );
  XNOR U26275 ( .A(p_input[2062]), .B(p_input[974]), .Z(n26487) );
  XNOR U26276 ( .A(n16738), .B(p_input[969]), .Z(n26454) );
  XNOR U26277 ( .A(n26470), .B(n26469), .Z(n26452) );
  XNOR U26278 ( .A(n26488), .B(n26475), .Z(n26469) );
  XOR U26279 ( .A(p_input[2056]), .B(p_input[968]), .Z(n26475) );
  XOR U26280 ( .A(n26466), .B(n26474), .Z(n26488) );
  XOR U26281 ( .A(n26489), .B(n26471), .Z(n26474) );
  XOR U26282 ( .A(p_input[2054]), .B(p_input[966]), .Z(n26471) );
  XNOR U26283 ( .A(p_input[2055]), .B(p_input[967]), .Z(n26489) );
  XNOR U26284 ( .A(n16741), .B(p_input[962]), .Z(n26466) );
  XNOR U26285 ( .A(n26480), .B(n26479), .Z(n26470) );
  XOR U26286 ( .A(n26490), .B(n26476), .Z(n26479) );
  XOR U26287 ( .A(p_input[2051]), .B(p_input[963]), .Z(n26476) );
  XNOR U26288 ( .A(p_input[2052]), .B(p_input[964]), .Z(n26490) );
  XOR U26289 ( .A(p_input[2053]), .B(p_input[965]), .Z(n26480) );
  XNOR U26290 ( .A(n26491), .B(n26492), .Z(n26387) );
  AND U26291 ( .A(n699), .B(n26493), .Z(n26492) );
  XNOR U26292 ( .A(n26494), .B(n26495), .Z(n699) );
  AND U26293 ( .A(n26496), .B(n26497), .Z(n26495) );
  XOR U26294 ( .A(n26494), .B(n26397), .Z(n26497) );
  XNOR U26295 ( .A(n26494), .B(n26351), .Z(n26496) );
  XOR U26296 ( .A(n26498), .B(n26499), .Z(n26494) );
  AND U26297 ( .A(n26500), .B(n26501), .Z(n26499) );
  XOR U26298 ( .A(n26498), .B(n26361), .Z(n26500) );
  XOR U26299 ( .A(n26502), .B(n26503), .Z(n26340) );
  AND U26300 ( .A(n703), .B(n26493), .Z(n26503) );
  XNOR U26301 ( .A(n26491), .B(n26502), .Z(n26493) );
  XNOR U26302 ( .A(n26504), .B(n26505), .Z(n703) );
  AND U26303 ( .A(n26506), .B(n26507), .Z(n26505) );
  XNOR U26304 ( .A(n26508), .B(n26504), .Z(n26507) );
  IV U26305 ( .A(n26397), .Z(n26508) );
  XNOR U26306 ( .A(n26509), .B(n26510), .Z(n26397) );
  AND U26307 ( .A(n706), .B(n26511), .Z(n26510) );
  XNOR U26308 ( .A(n26509), .B(n26512), .Z(n26511) );
  XNOR U26309 ( .A(n26351), .B(n26504), .Z(n26506) );
  XOR U26310 ( .A(n26513), .B(n26514), .Z(n26351) );
  AND U26311 ( .A(n714), .B(n26515), .Z(n26514) );
  XOR U26312 ( .A(n26498), .B(n26516), .Z(n26504) );
  AND U26313 ( .A(n26517), .B(n26501), .Z(n26516) );
  XNOR U26314 ( .A(n26410), .B(n26498), .Z(n26501) );
  XNOR U26315 ( .A(n26518), .B(n26519), .Z(n26410) );
  AND U26316 ( .A(n706), .B(n26520), .Z(n26519) );
  XOR U26317 ( .A(n26521), .B(n26518), .Z(n26520) );
  XNOR U26318 ( .A(n26522), .B(n26498), .Z(n26517) );
  IV U26319 ( .A(n26361), .Z(n26522) );
  XOR U26320 ( .A(n26523), .B(n26524), .Z(n26361) );
  AND U26321 ( .A(n714), .B(n26525), .Z(n26524) );
  XOR U26322 ( .A(n26526), .B(n26527), .Z(n26498) );
  AND U26323 ( .A(n26528), .B(n26529), .Z(n26527) );
  XNOR U26324 ( .A(n26435), .B(n26526), .Z(n26529) );
  XNOR U26325 ( .A(n26530), .B(n26531), .Z(n26435) );
  AND U26326 ( .A(n706), .B(n26532), .Z(n26531) );
  XNOR U26327 ( .A(n26533), .B(n26530), .Z(n26532) );
  XOR U26328 ( .A(n26526), .B(n26372), .Z(n26528) );
  XOR U26329 ( .A(n26534), .B(n26535), .Z(n26372) );
  AND U26330 ( .A(n714), .B(n26536), .Z(n26535) );
  XOR U26331 ( .A(n26537), .B(n26538), .Z(n26526) );
  AND U26332 ( .A(n26539), .B(n26540), .Z(n26538) );
  XNOR U26333 ( .A(n26537), .B(n26481), .Z(n26540) );
  XNOR U26334 ( .A(n26541), .B(n26542), .Z(n26481) );
  AND U26335 ( .A(n706), .B(n26543), .Z(n26542) );
  XOR U26336 ( .A(n26544), .B(n26541), .Z(n26543) );
  XNOR U26337 ( .A(n26545), .B(n26537), .Z(n26539) );
  IV U26338 ( .A(n26384), .Z(n26545) );
  XOR U26339 ( .A(n26546), .B(n26547), .Z(n26384) );
  AND U26340 ( .A(n714), .B(n26548), .Z(n26547) );
  AND U26341 ( .A(n26502), .B(n26491), .Z(n26537) );
  XNOR U26342 ( .A(n26549), .B(n26550), .Z(n26491) );
  AND U26343 ( .A(n706), .B(n26551), .Z(n26550) );
  XNOR U26344 ( .A(n26552), .B(n26549), .Z(n26551) );
  XNOR U26345 ( .A(n26553), .B(n26554), .Z(n706) );
  AND U26346 ( .A(n26555), .B(n26556), .Z(n26554) );
  XOR U26347 ( .A(n26512), .B(n26553), .Z(n26556) );
  AND U26348 ( .A(n26557), .B(n26558), .Z(n26512) );
  XOR U26349 ( .A(n26553), .B(n26509), .Z(n26555) );
  XNOR U26350 ( .A(n26559), .B(n26560), .Z(n26509) );
  AND U26351 ( .A(n710), .B(n26515), .Z(n26560) );
  XOR U26352 ( .A(n26513), .B(n26559), .Z(n26515) );
  XOR U26353 ( .A(n26561), .B(n26562), .Z(n26553) );
  AND U26354 ( .A(n26563), .B(n26564), .Z(n26562) );
  XNOR U26355 ( .A(n26561), .B(n26557), .Z(n26564) );
  IV U26356 ( .A(n26521), .Z(n26557) );
  XOR U26357 ( .A(n26565), .B(n26566), .Z(n26521) );
  XOR U26358 ( .A(n26567), .B(n26558), .Z(n26566) );
  AND U26359 ( .A(n26533), .B(n26568), .Z(n26558) );
  AND U26360 ( .A(n26569), .B(n26570), .Z(n26567) );
  XOR U26361 ( .A(n26571), .B(n26565), .Z(n26569) );
  XNOR U26362 ( .A(n26518), .B(n26561), .Z(n26563) );
  XNOR U26363 ( .A(n26572), .B(n26573), .Z(n26518) );
  AND U26364 ( .A(n710), .B(n26525), .Z(n26573) );
  XOR U26365 ( .A(n26572), .B(n26523), .Z(n26525) );
  XOR U26366 ( .A(n26574), .B(n26575), .Z(n26561) );
  AND U26367 ( .A(n26576), .B(n26577), .Z(n26575) );
  XNOR U26368 ( .A(n26574), .B(n26533), .Z(n26577) );
  XOR U26369 ( .A(n26578), .B(n26570), .Z(n26533) );
  XNOR U26370 ( .A(n26579), .B(n26565), .Z(n26570) );
  XOR U26371 ( .A(n26580), .B(n26581), .Z(n26565) );
  AND U26372 ( .A(n26582), .B(n26583), .Z(n26581) );
  XOR U26373 ( .A(n26584), .B(n26580), .Z(n26582) );
  XNOR U26374 ( .A(n26585), .B(n26586), .Z(n26579) );
  AND U26375 ( .A(n26587), .B(n26588), .Z(n26586) );
  XOR U26376 ( .A(n26585), .B(n26589), .Z(n26587) );
  XNOR U26377 ( .A(n26571), .B(n26568), .Z(n26578) );
  AND U26378 ( .A(n26590), .B(n26591), .Z(n26568) );
  XOR U26379 ( .A(n26592), .B(n26593), .Z(n26571) );
  AND U26380 ( .A(n26594), .B(n26595), .Z(n26593) );
  XOR U26381 ( .A(n26592), .B(n26596), .Z(n26594) );
  XNOR U26382 ( .A(n26530), .B(n26574), .Z(n26576) );
  XNOR U26383 ( .A(n26597), .B(n26598), .Z(n26530) );
  AND U26384 ( .A(n710), .B(n26536), .Z(n26598) );
  XOR U26385 ( .A(n26597), .B(n26534), .Z(n26536) );
  XOR U26386 ( .A(n26599), .B(n26600), .Z(n26574) );
  AND U26387 ( .A(n26601), .B(n26602), .Z(n26600) );
  XNOR U26388 ( .A(n26599), .B(n26590), .Z(n26602) );
  IV U26389 ( .A(n26544), .Z(n26590) );
  XNOR U26390 ( .A(n26603), .B(n26583), .Z(n26544) );
  XNOR U26391 ( .A(n26604), .B(n26589), .Z(n26583) );
  XOR U26392 ( .A(n26605), .B(n26606), .Z(n26589) );
  NOR U26393 ( .A(n26607), .B(n26608), .Z(n26606) );
  XNOR U26394 ( .A(n26605), .B(n26609), .Z(n26607) );
  XNOR U26395 ( .A(n26588), .B(n26580), .Z(n26604) );
  XOR U26396 ( .A(n26610), .B(n26611), .Z(n26580) );
  AND U26397 ( .A(n26612), .B(n26613), .Z(n26611) );
  XNOR U26398 ( .A(n26610), .B(n26614), .Z(n26612) );
  XNOR U26399 ( .A(n26615), .B(n26585), .Z(n26588) );
  XOR U26400 ( .A(n26616), .B(n26617), .Z(n26585) );
  AND U26401 ( .A(n26618), .B(n26619), .Z(n26617) );
  XOR U26402 ( .A(n26616), .B(n26620), .Z(n26618) );
  XNOR U26403 ( .A(n26621), .B(n26622), .Z(n26615) );
  NOR U26404 ( .A(n26623), .B(n26624), .Z(n26622) );
  XOR U26405 ( .A(n26621), .B(n26625), .Z(n26623) );
  XNOR U26406 ( .A(n26584), .B(n26591), .Z(n26603) );
  NOR U26407 ( .A(n26552), .B(n26626), .Z(n26591) );
  XOR U26408 ( .A(n26596), .B(n26595), .Z(n26584) );
  XNOR U26409 ( .A(n26627), .B(n26592), .Z(n26595) );
  XOR U26410 ( .A(n26628), .B(n26629), .Z(n26592) );
  AND U26411 ( .A(n26630), .B(n26631), .Z(n26629) );
  XOR U26412 ( .A(n26628), .B(n26632), .Z(n26630) );
  XNOR U26413 ( .A(n26633), .B(n26634), .Z(n26627) );
  NOR U26414 ( .A(n26635), .B(n26636), .Z(n26634) );
  XNOR U26415 ( .A(n26633), .B(n26637), .Z(n26635) );
  XOR U26416 ( .A(n26638), .B(n26639), .Z(n26596) );
  NOR U26417 ( .A(n26640), .B(n26641), .Z(n26639) );
  XNOR U26418 ( .A(n26638), .B(n26642), .Z(n26640) );
  XNOR U26419 ( .A(n26541), .B(n26599), .Z(n26601) );
  XNOR U26420 ( .A(n26643), .B(n26644), .Z(n26541) );
  AND U26421 ( .A(n710), .B(n26548), .Z(n26644) );
  XOR U26422 ( .A(n26643), .B(n26546), .Z(n26548) );
  AND U26423 ( .A(n26549), .B(n26552), .Z(n26599) );
  XOR U26424 ( .A(n26645), .B(n26626), .Z(n26552) );
  XNOR U26425 ( .A(p_input[2048]), .B(p_input[976]), .Z(n26626) );
  XOR U26426 ( .A(n26614), .B(n26613), .Z(n26645) );
  XNOR U26427 ( .A(n26646), .B(n26620), .Z(n26613) );
  XNOR U26428 ( .A(n26609), .B(n26608), .Z(n26620) );
  XOR U26429 ( .A(n26647), .B(n26605), .Z(n26608) );
  XNOR U26430 ( .A(n16904), .B(p_input[986]), .Z(n26605) );
  XNOR U26431 ( .A(p_input[2059]), .B(p_input[987]), .Z(n26647) );
  XOR U26432 ( .A(p_input[2060]), .B(p_input[988]), .Z(n26609) );
  XNOR U26433 ( .A(n26619), .B(n26610), .Z(n26646) );
  XNOR U26434 ( .A(n17068), .B(p_input[977]), .Z(n26610) );
  XOR U26435 ( .A(n26648), .B(n26625), .Z(n26619) );
  XNOR U26436 ( .A(p_input[2063]), .B(p_input[991]), .Z(n26625) );
  XOR U26437 ( .A(n26616), .B(n26624), .Z(n26648) );
  XOR U26438 ( .A(n26649), .B(n26621), .Z(n26624) );
  XOR U26439 ( .A(p_input[2061]), .B(p_input[989]), .Z(n26621) );
  XNOR U26440 ( .A(p_input[2062]), .B(p_input[990]), .Z(n26649) );
  XNOR U26441 ( .A(n16738), .B(p_input[985]), .Z(n26616) );
  IV U26442 ( .A(p_input[2057]), .Z(n16738) );
  XNOR U26443 ( .A(n26632), .B(n26631), .Z(n26614) );
  XNOR U26444 ( .A(n26650), .B(n26637), .Z(n26631) );
  XOR U26445 ( .A(p_input[2056]), .B(p_input[984]), .Z(n26637) );
  XOR U26446 ( .A(n26628), .B(n26636), .Z(n26650) );
  XOR U26447 ( .A(n26651), .B(n26633), .Z(n26636) );
  XOR U26448 ( .A(p_input[2054]), .B(p_input[982]), .Z(n26633) );
  XNOR U26449 ( .A(p_input[2055]), .B(p_input[983]), .Z(n26651) );
  XNOR U26450 ( .A(n16741), .B(p_input[978]), .Z(n26628) );
  XNOR U26451 ( .A(n26642), .B(n26641), .Z(n26632) );
  XOR U26452 ( .A(n26652), .B(n26638), .Z(n26641) );
  XOR U26453 ( .A(p_input[2051]), .B(p_input[979]), .Z(n26638) );
  XNOR U26454 ( .A(p_input[2052]), .B(p_input[980]), .Z(n26652) );
  XOR U26455 ( .A(p_input[2053]), .B(p_input[981]), .Z(n26642) );
  XNOR U26456 ( .A(n26653), .B(n26654), .Z(n26549) );
  AND U26457 ( .A(n710), .B(n26655), .Z(n26654) );
  XNOR U26458 ( .A(n26656), .B(n26657), .Z(n710) );
  AND U26459 ( .A(n26658), .B(n26659), .Z(n26657) );
  XOR U26460 ( .A(n26656), .B(n26559), .Z(n26659) );
  XNOR U26461 ( .A(n26656), .B(n26513), .Z(n26658) );
  XOR U26462 ( .A(n26660), .B(n26661), .Z(n26656) );
  AND U26463 ( .A(n26662), .B(n26663), .Z(n26661) );
  XOR U26464 ( .A(n26660), .B(n26523), .Z(n26662) );
  XOR U26465 ( .A(n26664), .B(n26665), .Z(n26502) );
  AND U26466 ( .A(n714), .B(n26655), .Z(n26665) );
  XNOR U26467 ( .A(n26653), .B(n26664), .Z(n26655) );
  XNOR U26468 ( .A(n26666), .B(n26667), .Z(n714) );
  AND U26469 ( .A(n26668), .B(n26669), .Z(n26667) );
  XNOR U26470 ( .A(n26670), .B(n26666), .Z(n26669) );
  IV U26471 ( .A(n26559), .Z(n26670) );
  XNOR U26472 ( .A(n26671), .B(n26672), .Z(n26559) );
  AND U26473 ( .A(n717), .B(n26673), .Z(n26672) );
  XNOR U26474 ( .A(n26671), .B(n26674), .Z(n26673) );
  XNOR U26475 ( .A(n26513), .B(n26666), .Z(n26668) );
  XOR U26476 ( .A(n26675), .B(n26676), .Z(n26513) );
  AND U26477 ( .A(n725), .B(n26677), .Z(n26676) );
  XOR U26478 ( .A(n26660), .B(n26678), .Z(n26666) );
  AND U26479 ( .A(n26679), .B(n26663), .Z(n26678) );
  XNOR U26480 ( .A(n26572), .B(n26660), .Z(n26663) );
  XNOR U26481 ( .A(n26680), .B(n26681), .Z(n26572) );
  AND U26482 ( .A(n717), .B(n26682), .Z(n26681) );
  XOR U26483 ( .A(n26683), .B(n26680), .Z(n26682) );
  XNOR U26484 ( .A(n26684), .B(n26660), .Z(n26679) );
  IV U26485 ( .A(n26523), .Z(n26684) );
  XOR U26486 ( .A(n26685), .B(n26686), .Z(n26523) );
  AND U26487 ( .A(n725), .B(n26687), .Z(n26686) );
  XOR U26488 ( .A(n26688), .B(n26689), .Z(n26660) );
  AND U26489 ( .A(n26690), .B(n26691), .Z(n26689) );
  XNOR U26490 ( .A(n26597), .B(n26688), .Z(n26691) );
  XNOR U26491 ( .A(n26692), .B(n26693), .Z(n26597) );
  AND U26492 ( .A(n717), .B(n26694), .Z(n26693) );
  XNOR U26493 ( .A(n26695), .B(n26692), .Z(n26694) );
  XOR U26494 ( .A(n26688), .B(n26534), .Z(n26690) );
  XOR U26495 ( .A(n26696), .B(n26697), .Z(n26534) );
  AND U26496 ( .A(n725), .B(n26698), .Z(n26697) );
  XOR U26497 ( .A(n26699), .B(n26700), .Z(n26688) );
  AND U26498 ( .A(n26701), .B(n26702), .Z(n26700) );
  XNOR U26499 ( .A(n26699), .B(n26643), .Z(n26702) );
  XNOR U26500 ( .A(n26703), .B(n26704), .Z(n26643) );
  AND U26501 ( .A(n717), .B(n26705), .Z(n26704) );
  XOR U26502 ( .A(n26706), .B(n26703), .Z(n26705) );
  XNOR U26503 ( .A(n26707), .B(n26699), .Z(n26701) );
  IV U26504 ( .A(n26546), .Z(n26707) );
  XOR U26505 ( .A(n26708), .B(n26709), .Z(n26546) );
  AND U26506 ( .A(n725), .B(n26710), .Z(n26709) );
  AND U26507 ( .A(n26664), .B(n26653), .Z(n26699) );
  XNOR U26508 ( .A(n26711), .B(n26712), .Z(n26653) );
  AND U26509 ( .A(n717), .B(n26713), .Z(n26712) );
  XNOR U26510 ( .A(n26714), .B(n26711), .Z(n26713) );
  XNOR U26511 ( .A(n26715), .B(n26716), .Z(n717) );
  AND U26512 ( .A(n26717), .B(n26718), .Z(n26716) );
  XOR U26513 ( .A(n26674), .B(n26715), .Z(n26718) );
  AND U26514 ( .A(n26719), .B(n26720), .Z(n26674) );
  XOR U26515 ( .A(n26715), .B(n26671), .Z(n26717) );
  XNOR U26516 ( .A(n26721), .B(n26722), .Z(n26671) );
  AND U26517 ( .A(n721), .B(n26677), .Z(n26722) );
  XOR U26518 ( .A(n26675), .B(n26721), .Z(n26677) );
  XOR U26519 ( .A(n26723), .B(n26724), .Z(n26715) );
  AND U26520 ( .A(n26725), .B(n26726), .Z(n26724) );
  XNOR U26521 ( .A(n26723), .B(n26719), .Z(n26726) );
  IV U26522 ( .A(n26683), .Z(n26719) );
  XOR U26523 ( .A(n26727), .B(n26728), .Z(n26683) );
  XOR U26524 ( .A(n26729), .B(n26720), .Z(n26728) );
  AND U26525 ( .A(n26695), .B(n26730), .Z(n26720) );
  AND U26526 ( .A(n26731), .B(n26732), .Z(n26729) );
  XOR U26527 ( .A(n26733), .B(n26727), .Z(n26731) );
  XNOR U26528 ( .A(n26680), .B(n26723), .Z(n26725) );
  XNOR U26529 ( .A(n26734), .B(n26735), .Z(n26680) );
  AND U26530 ( .A(n721), .B(n26687), .Z(n26735) );
  XOR U26531 ( .A(n26734), .B(n26685), .Z(n26687) );
  XOR U26532 ( .A(n26736), .B(n26737), .Z(n26723) );
  AND U26533 ( .A(n26738), .B(n26739), .Z(n26737) );
  XNOR U26534 ( .A(n26736), .B(n26695), .Z(n26739) );
  XOR U26535 ( .A(n26740), .B(n26732), .Z(n26695) );
  XNOR U26536 ( .A(n26741), .B(n26727), .Z(n26732) );
  XOR U26537 ( .A(n26742), .B(n26743), .Z(n26727) );
  AND U26538 ( .A(n26744), .B(n26745), .Z(n26743) );
  XOR U26539 ( .A(n26746), .B(n26742), .Z(n26744) );
  XNOR U26540 ( .A(n26747), .B(n26748), .Z(n26741) );
  AND U26541 ( .A(n26749), .B(n26750), .Z(n26748) );
  XOR U26542 ( .A(n26747), .B(n26751), .Z(n26749) );
  XNOR U26543 ( .A(n26733), .B(n26730), .Z(n26740) );
  AND U26544 ( .A(n26752), .B(n26753), .Z(n26730) );
  XOR U26545 ( .A(n26754), .B(n26755), .Z(n26733) );
  AND U26546 ( .A(n26756), .B(n26757), .Z(n26755) );
  XOR U26547 ( .A(n26754), .B(n26758), .Z(n26756) );
  XNOR U26548 ( .A(n26692), .B(n26736), .Z(n26738) );
  XNOR U26549 ( .A(n26759), .B(n26760), .Z(n26692) );
  AND U26550 ( .A(n721), .B(n26698), .Z(n26760) );
  XOR U26551 ( .A(n26759), .B(n26696), .Z(n26698) );
  XOR U26552 ( .A(n26761), .B(n26762), .Z(n26736) );
  AND U26553 ( .A(n26763), .B(n26764), .Z(n26762) );
  XNOR U26554 ( .A(n26761), .B(n26752), .Z(n26764) );
  IV U26555 ( .A(n26706), .Z(n26752) );
  XNOR U26556 ( .A(n26765), .B(n26745), .Z(n26706) );
  XNOR U26557 ( .A(n26766), .B(n26751), .Z(n26745) );
  XNOR U26558 ( .A(n26767), .B(n26768), .Z(n26751) );
  NOR U26559 ( .A(n26769), .B(n26770), .Z(n26768) );
  XOR U26560 ( .A(n26767), .B(n26771), .Z(n26769) );
  XNOR U26561 ( .A(n26750), .B(n26742), .Z(n26766) );
  XOR U26562 ( .A(n26772), .B(n26773), .Z(n26742) );
  AND U26563 ( .A(n26774), .B(n26775), .Z(n26773) );
  XOR U26564 ( .A(n26772), .B(n26776), .Z(n26774) );
  XNOR U26565 ( .A(n26777), .B(n26747), .Z(n26750) );
  XOR U26566 ( .A(n26778), .B(n26779), .Z(n26747) );
  AND U26567 ( .A(n26780), .B(n26781), .Z(n26779) );
  XNOR U26568 ( .A(n26782), .B(n26783), .Z(n26780) );
  IV U26569 ( .A(n26778), .Z(n26782) );
  XNOR U26570 ( .A(n26784), .B(n26785), .Z(n26777) );
  NOR U26571 ( .A(n26786), .B(n26787), .Z(n26785) );
  XNOR U26572 ( .A(n26784), .B(n26788), .Z(n26786) );
  XNOR U26573 ( .A(n26746), .B(n26753), .Z(n26765) );
  NOR U26574 ( .A(n26714), .B(n26789), .Z(n26753) );
  XOR U26575 ( .A(n26758), .B(n26757), .Z(n26746) );
  XNOR U26576 ( .A(n26790), .B(n26754), .Z(n26757) );
  XOR U26577 ( .A(n26791), .B(n26792), .Z(n26754) );
  AND U26578 ( .A(n26793), .B(n26794), .Z(n26792) );
  XOR U26579 ( .A(n26791), .B(n26795), .Z(n26793) );
  XNOR U26580 ( .A(n26796), .B(n26797), .Z(n26790) );
  NOR U26581 ( .A(n26798), .B(n26799), .Z(n26797) );
  XNOR U26582 ( .A(n26796), .B(n26800), .Z(n26798) );
  XOR U26583 ( .A(n26801), .B(n26802), .Z(n26758) );
  NOR U26584 ( .A(n26803), .B(n26804), .Z(n26802) );
  XNOR U26585 ( .A(n26801), .B(n26805), .Z(n26803) );
  XNOR U26586 ( .A(n26703), .B(n26761), .Z(n26763) );
  XNOR U26587 ( .A(n26806), .B(n26807), .Z(n26703) );
  AND U26588 ( .A(n721), .B(n26710), .Z(n26807) );
  XOR U26589 ( .A(n26806), .B(n26708), .Z(n26710) );
  AND U26590 ( .A(n26711), .B(n26714), .Z(n26761) );
  XOR U26591 ( .A(n26808), .B(n26789), .Z(n26714) );
  XNOR U26592 ( .A(p_input[2048]), .B(p_input[992]), .Z(n26789) );
  XNOR U26593 ( .A(n26776), .B(n26775), .Z(n26808) );
  XNOR U26594 ( .A(n26809), .B(n26783), .Z(n26775) );
  XNOR U26595 ( .A(n26771), .B(n26770), .Z(n26783) );
  XNOR U26596 ( .A(n26810), .B(n26767), .Z(n26770) );
  XNOR U26597 ( .A(p_input[1002]), .B(p_input[2058]), .Z(n26767) );
  XOR U26598 ( .A(p_input[1003]), .B(n16732), .Z(n26810) );
  XOR U26599 ( .A(p_input[1004]), .B(p_input[2060]), .Z(n26771) );
  XNOR U26600 ( .A(n26781), .B(n26772), .Z(n26809) );
  XNOR U26601 ( .A(n17068), .B(p_input[993]), .Z(n26772) );
  IV U26602 ( .A(p_input[2049]), .Z(n17068) );
  XNOR U26603 ( .A(n26811), .B(n26788), .Z(n26781) );
  XNOR U26604 ( .A(p_input[1007]), .B(n16735), .Z(n26788) );
  XOR U26605 ( .A(n26778), .B(n26787), .Z(n26811) );
  XOR U26606 ( .A(n26812), .B(n26784), .Z(n26787) );
  XOR U26607 ( .A(p_input[1005]), .B(p_input[2061]), .Z(n26784) );
  XOR U26608 ( .A(p_input[1006]), .B(n16737), .Z(n26812) );
  XOR U26609 ( .A(p_input[1001]), .B(p_input[2057]), .Z(n26778) );
  XOR U26610 ( .A(n26795), .B(n26794), .Z(n26776) );
  XNOR U26611 ( .A(n26813), .B(n26800), .Z(n26794) );
  XOR U26612 ( .A(p_input[1000]), .B(p_input[2056]), .Z(n26800) );
  XOR U26613 ( .A(n26791), .B(n26799), .Z(n26813) );
  XOR U26614 ( .A(n26814), .B(n26796), .Z(n26799) );
  XOR U26615 ( .A(p_input[2054]), .B(p_input[998]), .Z(n26796) );
  XNOR U26616 ( .A(p_input[2055]), .B(p_input[999]), .Z(n26814) );
  XNOR U26617 ( .A(n16741), .B(p_input[994]), .Z(n26791) );
  IV U26618 ( .A(p_input[2050]), .Z(n16741) );
  XNOR U26619 ( .A(n26805), .B(n26804), .Z(n26795) );
  XOR U26620 ( .A(n26815), .B(n26801), .Z(n26804) );
  XOR U26621 ( .A(p_input[2051]), .B(p_input[995]), .Z(n26801) );
  XNOR U26622 ( .A(p_input[2052]), .B(p_input[996]), .Z(n26815) );
  XOR U26623 ( .A(p_input[2053]), .B(p_input[997]), .Z(n26805) );
  XNOR U26624 ( .A(n26816), .B(n26817), .Z(n26711) );
  AND U26625 ( .A(n721), .B(n26818), .Z(n26817) );
  XNOR U26626 ( .A(n26819), .B(n26820), .Z(n721) );
  AND U26627 ( .A(n26821), .B(n26822), .Z(n26820) );
  XOR U26628 ( .A(n26819), .B(n26721), .Z(n26822) );
  XNOR U26629 ( .A(n26819), .B(n26675), .Z(n26821) );
  XOR U26630 ( .A(n26823), .B(n26824), .Z(n26819) );
  AND U26631 ( .A(n26825), .B(n26826), .Z(n26824) );
  XOR U26632 ( .A(n26823), .B(n26685), .Z(n26825) );
  XOR U26633 ( .A(n26827), .B(n26828), .Z(n26664) );
  AND U26634 ( .A(n725), .B(n26818), .Z(n26828) );
  XNOR U26635 ( .A(n26816), .B(n26827), .Z(n26818) );
  XNOR U26636 ( .A(n26829), .B(n26830), .Z(n725) );
  AND U26637 ( .A(n26831), .B(n26832), .Z(n26830) );
  XNOR U26638 ( .A(n26833), .B(n26829), .Z(n26832) );
  IV U26639 ( .A(n26721), .Z(n26833) );
  XNOR U26640 ( .A(n26834), .B(n26835), .Z(n26721) );
  AND U26641 ( .A(n728), .B(n26836), .Z(n26835) );
  XNOR U26642 ( .A(n26834), .B(n26837), .Z(n26836) );
  XNOR U26643 ( .A(n26675), .B(n26829), .Z(n26831) );
  XOR U26644 ( .A(n26838), .B(n26839), .Z(n26675) );
  AND U26645 ( .A(n736), .B(n26840), .Z(n26839) );
  XOR U26646 ( .A(n26823), .B(n26841), .Z(n26829) );
  AND U26647 ( .A(n26842), .B(n26826), .Z(n26841) );
  XNOR U26648 ( .A(n26734), .B(n26823), .Z(n26826) );
  XNOR U26649 ( .A(n26843), .B(n26844), .Z(n26734) );
  AND U26650 ( .A(n728), .B(n26845), .Z(n26844) );
  XOR U26651 ( .A(n26846), .B(n26843), .Z(n26845) );
  XNOR U26652 ( .A(n26847), .B(n26823), .Z(n26842) );
  IV U26653 ( .A(n26685), .Z(n26847) );
  XOR U26654 ( .A(n26848), .B(n26849), .Z(n26685) );
  AND U26655 ( .A(n736), .B(n26850), .Z(n26849) );
  XOR U26656 ( .A(n26851), .B(n26852), .Z(n26823) );
  AND U26657 ( .A(n26853), .B(n26854), .Z(n26852) );
  XNOR U26658 ( .A(n26759), .B(n26851), .Z(n26854) );
  XNOR U26659 ( .A(n26855), .B(n26856), .Z(n26759) );
  AND U26660 ( .A(n728), .B(n26857), .Z(n26856) );
  XNOR U26661 ( .A(n26858), .B(n26855), .Z(n26857) );
  XOR U26662 ( .A(n26851), .B(n26696), .Z(n26853) );
  XOR U26663 ( .A(n26859), .B(n26860), .Z(n26696) );
  AND U26664 ( .A(n736), .B(n26861), .Z(n26860) );
  XOR U26665 ( .A(n26862), .B(n26863), .Z(n26851) );
  AND U26666 ( .A(n26864), .B(n26865), .Z(n26863) );
  XNOR U26667 ( .A(n26862), .B(n26806), .Z(n26865) );
  XNOR U26668 ( .A(n26866), .B(n26867), .Z(n26806) );
  AND U26669 ( .A(n728), .B(n26868), .Z(n26867) );
  XOR U26670 ( .A(n26869), .B(n26866), .Z(n26868) );
  XNOR U26671 ( .A(n26870), .B(n26862), .Z(n26864) );
  IV U26672 ( .A(n26708), .Z(n26870) );
  XOR U26673 ( .A(n26871), .B(n26872), .Z(n26708) );
  AND U26674 ( .A(n736), .B(n26873), .Z(n26872) );
  AND U26675 ( .A(n26827), .B(n26816), .Z(n26862) );
  XNOR U26676 ( .A(n26874), .B(n26875), .Z(n26816) );
  AND U26677 ( .A(n728), .B(n26876), .Z(n26875) );
  XNOR U26678 ( .A(n26877), .B(n26874), .Z(n26876) );
  XNOR U26679 ( .A(n26878), .B(n26879), .Z(n728) );
  AND U26680 ( .A(n26880), .B(n26881), .Z(n26879) );
  XOR U26681 ( .A(n26837), .B(n26878), .Z(n26881) );
  AND U26682 ( .A(n26882), .B(n26883), .Z(n26837) );
  XOR U26683 ( .A(n26878), .B(n26834), .Z(n26880) );
  XNOR U26684 ( .A(n26884), .B(n26885), .Z(n26834) );
  AND U26685 ( .A(n732), .B(n26840), .Z(n26885) );
  XOR U26686 ( .A(n26838), .B(n26884), .Z(n26840) );
  XOR U26687 ( .A(n26886), .B(n26887), .Z(n26878) );
  AND U26688 ( .A(n26888), .B(n26889), .Z(n26887) );
  XNOR U26689 ( .A(n26886), .B(n26882), .Z(n26889) );
  IV U26690 ( .A(n26846), .Z(n26882) );
  XOR U26691 ( .A(n26890), .B(n26891), .Z(n26846) );
  XOR U26692 ( .A(n26892), .B(n26883), .Z(n26891) );
  AND U26693 ( .A(n26858), .B(n26893), .Z(n26883) );
  AND U26694 ( .A(n26894), .B(n26895), .Z(n26892) );
  XOR U26695 ( .A(n26896), .B(n26890), .Z(n26894) );
  XNOR U26696 ( .A(n26843), .B(n26886), .Z(n26888) );
  XNOR U26697 ( .A(n26897), .B(n26898), .Z(n26843) );
  AND U26698 ( .A(n732), .B(n26850), .Z(n26898) );
  XOR U26699 ( .A(n26897), .B(n26848), .Z(n26850) );
  XOR U26700 ( .A(n26899), .B(n26900), .Z(n26886) );
  AND U26701 ( .A(n26901), .B(n26902), .Z(n26900) );
  XNOR U26702 ( .A(n26899), .B(n26858), .Z(n26902) );
  XOR U26703 ( .A(n26903), .B(n26895), .Z(n26858) );
  XNOR U26704 ( .A(n26904), .B(n26890), .Z(n26895) );
  XOR U26705 ( .A(n26905), .B(n26906), .Z(n26890) );
  AND U26706 ( .A(n26907), .B(n26908), .Z(n26906) );
  XOR U26707 ( .A(n26909), .B(n26905), .Z(n26907) );
  XNOR U26708 ( .A(n26910), .B(n26911), .Z(n26904) );
  AND U26709 ( .A(n26912), .B(n26913), .Z(n26911) );
  XOR U26710 ( .A(n26910), .B(n26914), .Z(n26912) );
  XNOR U26711 ( .A(n26896), .B(n26893), .Z(n26903) );
  AND U26712 ( .A(n26915), .B(n26916), .Z(n26893) );
  XOR U26713 ( .A(n26917), .B(n26918), .Z(n26896) );
  AND U26714 ( .A(n26919), .B(n26920), .Z(n26918) );
  XOR U26715 ( .A(n26917), .B(n26921), .Z(n26919) );
  XNOR U26716 ( .A(n26855), .B(n26899), .Z(n26901) );
  XNOR U26717 ( .A(n26922), .B(n26923), .Z(n26855) );
  AND U26718 ( .A(n732), .B(n26861), .Z(n26923) );
  XOR U26719 ( .A(n26922), .B(n26859), .Z(n26861) );
  XOR U26720 ( .A(n26924), .B(n26925), .Z(n26899) );
  AND U26721 ( .A(n26926), .B(n26927), .Z(n26925) );
  XNOR U26722 ( .A(n26924), .B(n26915), .Z(n26927) );
  IV U26723 ( .A(n26869), .Z(n26915) );
  XNOR U26724 ( .A(n26928), .B(n26908), .Z(n26869) );
  XNOR U26725 ( .A(n26929), .B(n26914), .Z(n26908) );
  XNOR U26726 ( .A(n26930), .B(n26931), .Z(n26914) );
  NOR U26727 ( .A(n26932), .B(n26933), .Z(n26931) );
  XOR U26728 ( .A(n26930), .B(n26934), .Z(n26932) );
  XNOR U26729 ( .A(n26913), .B(n26905), .Z(n26929) );
  XOR U26730 ( .A(n26935), .B(n26936), .Z(n26905) );
  AND U26731 ( .A(n26937), .B(n26938), .Z(n26936) );
  XOR U26732 ( .A(n26935), .B(n26939), .Z(n26937) );
  XNOR U26733 ( .A(n26940), .B(n26910), .Z(n26913) );
  XOR U26734 ( .A(n26941), .B(n26942), .Z(n26910) );
  AND U26735 ( .A(n26943), .B(n26944), .Z(n26942) );
  XNOR U26736 ( .A(n26945), .B(n26946), .Z(n26943) );
  IV U26737 ( .A(n26941), .Z(n26945) );
  XNOR U26738 ( .A(n26947), .B(n26948), .Z(n26940) );
  NOR U26739 ( .A(n26949), .B(n26950), .Z(n26948) );
  XNOR U26740 ( .A(n26947), .B(n26951), .Z(n26949) );
  XNOR U26741 ( .A(n26909), .B(n26916), .Z(n26928) );
  NOR U26742 ( .A(n26877), .B(n26952), .Z(n26916) );
  XOR U26743 ( .A(n26921), .B(n26920), .Z(n26909) );
  XNOR U26744 ( .A(n26953), .B(n26917), .Z(n26920) );
  XOR U26745 ( .A(n26954), .B(n26955), .Z(n26917) );
  AND U26746 ( .A(n26956), .B(n26957), .Z(n26955) );
  XNOR U26747 ( .A(n26958), .B(n26959), .Z(n26956) );
  IV U26748 ( .A(n26954), .Z(n26958) );
  XNOR U26749 ( .A(n26960), .B(n26961), .Z(n26953) );
  NOR U26750 ( .A(n26962), .B(n26963), .Z(n26961) );
  XNOR U26751 ( .A(n26960), .B(n26964), .Z(n26962) );
  XOR U26752 ( .A(n26965), .B(n26966), .Z(n26921) );
  NOR U26753 ( .A(n26967), .B(n26968), .Z(n26966) );
  XNOR U26754 ( .A(n26965), .B(n26969), .Z(n26967) );
  XNOR U26755 ( .A(n26866), .B(n26924), .Z(n26926) );
  XNOR U26756 ( .A(n26970), .B(n26971), .Z(n26866) );
  AND U26757 ( .A(n732), .B(n26873), .Z(n26971) );
  XOR U26758 ( .A(n26970), .B(n26871), .Z(n26873) );
  AND U26759 ( .A(n26874), .B(n26877), .Z(n26924) );
  XOR U26760 ( .A(n26972), .B(n26952), .Z(n26877) );
  XNOR U26761 ( .A(p_input[1008]), .B(p_input[2048]), .Z(n26952) );
  XNOR U26762 ( .A(n26939), .B(n26938), .Z(n26972) );
  XNOR U26763 ( .A(n26973), .B(n26946), .Z(n26938) );
  XNOR U26764 ( .A(n26934), .B(n26933), .Z(n26946) );
  XNOR U26765 ( .A(n26974), .B(n26930), .Z(n26933) );
  XNOR U26766 ( .A(p_input[1018]), .B(p_input[2058]), .Z(n26930) );
  XOR U26767 ( .A(p_input[1019]), .B(n16732), .Z(n26974) );
  XOR U26768 ( .A(p_input[1020]), .B(p_input[2060]), .Z(n26934) );
  XOR U26769 ( .A(n26944), .B(n26975), .Z(n26973) );
  IV U26770 ( .A(n26935), .Z(n26975) );
  XOR U26771 ( .A(p_input[1009]), .B(p_input[2049]), .Z(n26935) );
  XNOR U26772 ( .A(n26976), .B(n26951), .Z(n26944) );
  XNOR U26773 ( .A(p_input[1023]), .B(n16735), .Z(n26951) );
  XOR U26774 ( .A(n26941), .B(n26950), .Z(n26976) );
  XOR U26775 ( .A(n26977), .B(n26947), .Z(n26950) );
  XOR U26776 ( .A(p_input[1021]), .B(p_input[2061]), .Z(n26947) );
  XOR U26777 ( .A(p_input[1022]), .B(n16737), .Z(n26977) );
  XOR U26778 ( .A(p_input[1017]), .B(p_input[2057]), .Z(n26941) );
  XOR U26779 ( .A(n26959), .B(n26957), .Z(n26939) );
  XNOR U26780 ( .A(n26978), .B(n26964), .Z(n26957) );
  XOR U26781 ( .A(p_input[1016]), .B(p_input[2056]), .Z(n26964) );
  XOR U26782 ( .A(n26954), .B(n26963), .Z(n26978) );
  XOR U26783 ( .A(n26979), .B(n26960), .Z(n26963) );
  XOR U26784 ( .A(p_input[1014]), .B(p_input[2054]), .Z(n26960) );
  XOR U26785 ( .A(p_input[1015]), .B(n17722), .Z(n26979) );
  XOR U26786 ( .A(p_input[1010]), .B(p_input[2050]), .Z(n26954) );
  XNOR U26787 ( .A(n26969), .B(n26968), .Z(n26959) );
  XOR U26788 ( .A(n26980), .B(n26965), .Z(n26968) );
  XOR U26789 ( .A(p_input[1011]), .B(p_input[2051]), .Z(n26965) );
  XOR U26790 ( .A(p_input[1012]), .B(n17724), .Z(n26980) );
  XOR U26791 ( .A(p_input[1013]), .B(p_input[2053]), .Z(n26969) );
  XNOR U26792 ( .A(n26981), .B(n26982), .Z(n26874) );
  AND U26793 ( .A(n732), .B(n26983), .Z(n26982) );
  XNOR U26794 ( .A(n26984), .B(n26985), .Z(n732) );
  AND U26795 ( .A(n26986), .B(n26987), .Z(n26985) );
  XOR U26796 ( .A(n26984), .B(n26884), .Z(n26987) );
  XNOR U26797 ( .A(n26984), .B(n26838), .Z(n26986) );
  XOR U26798 ( .A(n26988), .B(n26989), .Z(n26984) );
  AND U26799 ( .A(n26990), .B(n26991), .Z(n26989) );
  XOR U26800 ( .A(n26988), .B(n26848), .Z(n26990) );
  XOR U26801 ( .A(n26992), .B(n26993), .Z(n26827) );
  AND U26802 ( .A(n736), .B(n26983), .Z(n26993) );
  XNOR U26803 ( .A(n26981), .B(n26992), .Z(n26983) );
  XNOR U26804 ( .A(n26994), .B(n26995), .Z(n736) );
  AND U26805 ( .A(n26996), .B(n26997), .Z(n26995) );
  XNOR U26806 ( .A(n26998), .B(n26994), .Z(n26997) );
  IV U26807 ( .A(n26884), .Z(n26998) );
  XNOR U26808 ( .A(n26999), .B(n27000), .Z(n26884) );
  AND U26809 ( .A(n739), .B(n27001), .Z(n27000) );
  XNOR U26810 ( .A(n26999), .B(n27002), .Z(n27001) );
  XNOR U26811 ( .A(n26838), .B(n26994), .Z(n26996) );
  XOR U26812 ( .A(n27003), .B(n27004), .Z(n26838) );
  AND U26813 ( .A(n747), .B(n27005), .Z(n27004) );
  XOR U26814 ( .A(n26988), .B(n27006), .Z(n26994) );
  AND U26815 ( .A(n27007), .B(n26991), .Z(n27006) );
  XNOR U26816 ( .A(n26897), .B(n26988), .Z(n26991) );
  XNOR U26817 ( .A(n27008), .B(n27009), .Z(n26897) );
  AND U26818 ( .A(n739), .B(n27010), .Z(n27009) );
  XOR U26819 ( .A(n27011), .B(n27008), .Z(n27010) );
  XNOR U26820 ( .A(n27012), .B(n26988), .Z(n27007) );
  IV U26821 ( .A(n26848), .Z(n27012) );
  XOR U26822 ( .A(n27013), .B(n27014), .Z(n26848) );
  AND U26823 ( .A(n747), .B(n27015), .Z(n27014) );
  XOR U26824 ( .A(n27016), .B(n27017), .Z(n26988) );
  AND U26825 ( .A(n27018), .B(n27019), .Z(n27017) );
  XNOR U26826 ( .A(n26922), .B(n27016), .Z(n27019) );
  XNOR U26827 ( .A(n27020), .B(n27021), .Z(n26922) );
  AND U26828 ( .A(n739), .B(n27022), .Z(n27021) );
  XNOR U26829 ( .A(n27023), .B(n27020), .Z(n27022) );
  XOR U26830 ( .A(n27016), .B(n26859), .Z(n27018) );
  XOR U26831 ( .A(n27024), .B(n27025), .Z(n26859) );
  AND U26832 ( .A(n747), .B(n27026), .Z(n27025) );
  XOR U26833 ( .A(n27027), .B(n27028), .Z(n27016) );
  AND U26834 ( .A(n27029), .B(n27030), .Z(n27028) );
  XNOR U26835 ( .A(n27027), .B(n26970), .Z(n27030) );
  XNOR U26836 ( .A(n27031), .B(n27032), .Z(n26970) );
  AND U26837 ( .A(n739), .B(n27033), .Z(n27032) );
  XOR U26838 ( .A(n27034), .B(n27031), .Z(n27033) );
  XNOR U26839 ( .A(n27035), .B(n27027), .Z(n27029) );
  IV U26840 ( .A(n26871), .Z(n27035) );
  XOR U26841 ( .A(n27036), .B(n27037), .Z(n26871) );
  AND U26842 ( .A(n747), .B(n27038), .Z(n27037) );
  AND U26843 ( .A(n26992), .B(n26981), .Z(n27027) );
  XNOR U26844 ( .A(n27039), .B(n27040), .Z(n26981) );
  AND U26845 ( .A(n739), .B(n27041), .Z(n27040) );
  XNOR U26846 ( .A(n27042), .B(n27039), .Z(n27041) );
  XNOR U26847 ( .A(n27043), .B(n27044), .Z(n739) );
  AND U26848 ( .A(n27045), .B(n27046), .Z(n27044) );
  XOR U26849 ( .A(n27002), .B(n27043), .Z(n27046) );
  AND U26850 ( .A(n27047), .B(n27048), .Z(n27002) );
  XOR U26851 ( .A(n27043), .B(n26999), .Z(n27045) );
  XNOR U26852 ( .A(n27049), .B(n27050), .Z(n26999) );
  AND U26853 ( .A(n743), .B(n27005), .Z(n27050) );
  XOR U26854 ( .A(n27003), .B(n27049), .Z(n27005) );
  XOR U26855 ( .A(n27051), .B(n27052), .Z(n27043) );
  AND U26856 ( .A(n27053), .B(n27054), .Z(n27052) );
  XNOR U26857 ( .A(n27051), .B(n27047), .Z(n27054) );
  IV U26858 ( .A(n27011), .Z(n27047) );
  XOR U26859 ( .A(n27055), .B(n27056), .Z(n27011) );
  XOR U26860 ( .A(n27057), .B(n27048), .Z(n27056) );
  AND U26861 ( .A(n27023), .B(n27058), .Z(n27048) );
  AND U26862 ( .A(n27059), .B(n27060), .Z(n27057) );
  XOR U26863 ( .A(n27061), .B(n27055), .Z(n27059) );
  XNOR U26864 ( .A(n27008), .B(n27051), .Z(n27053) );
  XNOR U26865 ( .A(n27062), .B(n27063), .Z(n27008) );
  AND U26866 ( .A(n743), .B(n27015), .Z(n27063) );
  XOR U26867 ( .A(n27062), .B(n27013), .Z(n27015) );
  XOR U26868 ( .A(n27064), .B(n27065), .Z(n27051) );
  AND U26869 ( .A(n27066), .B(n27067), .Z(n27065) );
  XNOR U26870 ( .A(n27064), .B(n27023), .Z(n27067) );
  XOR U26871 ( .A(n27068), .B(n27060), .Z(n27023) );
  XNOR U26872 ( .A(n27069), .B(n27055), .Z(n27060) );
  XOR U26873 ( .A(n27070), .B(n27071), .Z(n27055) );
  AND U26874 ( .A(n27072), .B(n27073), .Z(n27071) );
  XOR U26875 ( .A(n27074), .B(n27070), .Z(n27072) );
  XNOR U26876 ( .A(n27075), .B(n27076), .Z(n27069) );
  AND U26877 ( .A(n27077), .B(n27078), .Z(n27076) );
  XOR U26878 ( .A(n27075), .B(n27079), .Z(n27077) );
  XNOR U26879 ( .A(n27061), .B(n27058), .Z(n27068) );
  AND U26880 ( .A(n27080), .B(n27081), .Z(n27058) );
  XOR U26881 ( .A(n27082), .B(n27083), .Z(n27061) );
  AND U26882 ( .A(n27084), .B(n27085), .Z(n27083) );
  XOR U26883 ( .A(n27082), .B(n27086), .Z(n27084) );
  XNOR U26884 ( .A(n27020), .B(n27064), .Z(n27066) );
  XNOR U26885 ( .A(n27087), .B(n27088), .Z(n27020) );
  AND U26886 ( .A(n743), .B(n27026), .Z(n27088) );
  XOR U26887 ( .A(n27087), .B(n27024), .Z(n27026) );
  XOR U26888 ( .A(n27089), .B(n27090), .Z(n27064) );
  AND U26889 ( .A(n27091), .B(n27092), .Z(n27090) );
  XNOR U26890 ( .A(n27089), .B(n27080), .Z(n27092) );
  IV U26891 ( .A(n27034), .Z(n27080) );
  XNOR U26892 ( .A(n27093), .B(n27073), .Z(n27034) );
  XNOR U26893 ( .A(n27094), .B(n27079), .Z(n27073) );
  XNOR U26894 ( .A(n27095), .B(n27096), .Z(n27079) );
  NOR U26895 ( .A(n27097), .B(n27098), .Z(n27096) );
  XOR U26896 ( .A(n27095), .B(n27099), .Z(n27097) );
  XNOR U26897 ( .A(n27078), .B(n27070), .Z(n27094) );
  XOR U26898 ( .A(n27100), .B(n27101), .Z(n27070) );
  AND U26899 ( .A(n27102), .B(n27103), .Z(n27101) );
  XOR U26900 ( .A(n27100), .B(n27104), .Z(n27102) );
  XNOR U26901 ( .A(n27105), .B(n27075), .Z(n27078) );
  XOR U26902 ( .A(n27106), .B(n27107), .Z(n27075) );
  AND U26903 ( .A(n27108), .B(n27109), .Z(n27107) );
  XNOR U26904 ( .A(n27110), .B(n27111), .Z(n27108) );
  IV U26905 ( .A(n27106), .Z(n27110) );
  XNOR U26906 ( .A(n27112), .B(n27113), .Z(n27105) );
  NOR U26907 ( .A(n27114), .B(n27115), .Z(n27113) );
  XNOR U26908 ( .A(n27112), .B(n27116), .Z(n27114) );
  XNOR U26909 ( .A(n27074), .B(n27081), .Z(n27093) );
  NOR U26910 ( .A(n27042), .B(n27117), .Z(n27081) );
  XOR U26911 ( .A(n27086), .B(n27085), .Z(n27074) );
  XNOR U26912 ( .A(n27118), .B(n27082), .Z(n27085) );
  XOR U26913 ( .A(n27119), .B(n27120), .Z(n27082) );
  AND U26914 ( .A(n27121), .B(n27122), .Z(n27120) );
  XNOR U26915 ( .A(n27123), .B(n27124), .Z(n27121) );
  IV U26916 ( .A(n27119), .Z(n27123) );
  XNOR U26917 ( .A(n27125), .B(n27126), .Z(n27118) );
  NOR U26918 ( .A(n27127), .B(n27128), .Z(n27126) );
  XNOR U26919 ( .A(n27125), .B(n27129), .Z(n27127) );
  XOR U26920 ( .A(n27130), .B(n27131), .Z(n27086) );
  NOR U26921 ( .A(n27132), .B(n27133), .Z(n27131) );
  XNOR U26922 ( .A(n27130), .B(n27134), .Z(n27132) );
  XNOR U26923 ( .A(n27031), .B(n27089), .Z(n27091) );
  XNOR U26924 ( .A(n27135), .B(n27136), .Z(n27031) );
  AND U26925 ( .A(n743), .B(n27038), .Z(n27136) );
  XOR U26926 ( .A(n27135), .B(n27036), .Z(n27038) );
  AND U26927 ( .A(n27039), .B(n27042), .Z(n27089) );
  XOR U26928 ( .A(n27137), .B(n27117), .Z(n27042) );
  XNOR U26929 ( .A(p_input[1024]), .B(p_input[2048]), .Z(n27117) );
  XNOR U26930 ( .A(n27104), .B(n27103), .Z(n27137) );
  XNOR U26931 ( .A(n27138), .B(n27111), .Z(n27103) );
  XNOR U26932 ( .A(n27099), .B(n27098), .Z(n27111) );
  XNOR U26933 ( .A(n27139), .B(n27095), .Z(n27098) );
  XNOR U26934 ( .A(p_input[1034]), .B(p_input[2058]), .Z(n27095) );
  XOR U26935 ( .A(p_input[1035]), .B(n16732), .Z(n27139) );
  XOR U26936 ( .A(p_input[1036]), .B(p_input[2060]), .Z(n27099) );
  XOR U26937 ( .A(n27109), .B(n27140), .Z(n27138) );
  IV U26938 ( .A(n27100), .Z(n27140) );
  XOR U26939 ( .A(p_input[1025]), .B(p_input[2049]), .Z(n27100) );
  XNOR U26940 ( .A(n27141), .B(n27116), .Z(n27109) );
  XNOR U26941 ( .A(p_input[1039]), .B(n16735), .Z(n27116) );
  XOR U26942 ( .A(n27106), .B(n27115), .Z(n27141) );
  XOR U26943 ( .A(n27142), .B(n27112), .Z(n27115) );
  XOR U26944 ( .A(p_input[1037]), .B(p_input[2061]), .Z(n27112) );
  XOR U26945 ( .A(p_input[1038]), .B(n16737), .Z(n27142) );
  XOR U26946 ( .A(p_input[1033]), .B(p_input[2057]), .Z(n27106) );
  XOR U26947 ( .A(n27124), .B(n27122), .Z(n27104) );
  XNOR U26948 ( .A(n27143), .B(n27129), .Z(n27122) );
  XOR U26949 ( .A(p_input[1032]), .B(p_input[2056]), .Z(n27129) );
  XOR U26950 ( .A(n27119), .B(n27128), .Z(n27143) );
  XOR U26951 ( .A(n27144), .B(n27125), .Z(n27128) );
  XOR U26952 ( .A(p_input[1030]), .B(p_input[2054]), .Z(n27125) );
  XOR U26953 ( .A(p_input[1031]), .B(n17722), .Z(n27144) );
  XOR U26954 ( .A(p_input[1026]), .B(p_input[2050]), .Z(n27119) );
  XNOR U26955 ( .A(n27134), .B(n27133), .Z(n27124) );
  XOR U26956 ( .A(n27145), .B(n27130), .Z(n27133) );
  XOR U26957 ( .A(p_input[1027]), .B(p_input[2051]), .Z(n27130) );
  XOR U26958 ( .A(p_input[1028]), .B(n17724), .Z(n27145) );
  XOR U26959 ( .A(p_input[1029]), .B(p_input[2053]), .Z(n27134) );
  XNOR U26960 ( .A(n27146), .B(n27147), .Z(n27039) );
  AND U26961 ( .A(n743), .B(n27148), .Z(n27147) );
  XNOR U26962 ( .A(n27149), .B(n27150), .Z(n743) );
  AND U26963 ( .A(n27151), .B(n27152), .Z(n27150) );
  XOR U26964 ( .A(n27149), .B(n27049), .Z(n27152) );
  XNOR U26965 ( .A(n27149), .B(n27003), .Z(n27151) );
  XOR U26966 ( .A(n27153), .B(n27154), .Z(n27149) );
  AND U26967 ( .A(n27155), .B(n27156), .Z(n27154) );
  XOR U26968 ( .A(n27153), .B(n27013), .Z(n27155) );
  XOR U26969 ( .A(n27157), .B(n27158), .Z(n26992) );
  AND U26970 ( .A(n747), .B(n27148), .Z(n27158) );
  XNOR U26971 ( .A(n27146), .B(n27157), .Z(n27148) );
  XNOR U26972 ( .A(n27159), .B(n27160), .Z(n747) );
  AND U26973 ( .A(n27161), .B(n27162), .Z(n27160) );
  XNOR U26974 ( .A(n27163), .B(n27159), .Z(n27162) );
  IV U26975 ( .A(n27049), .Z(n27163) );
  XNOR U26976 ( .A(n27164), .B(n27165), .Z(n27049) );
  AND U26977 ( .A(n750), .B(n27166), .Z(n27165) );
  XNOR U26978 ( .A(n27164), .B(n27167), .Z(n27166) );
  XNOR U26979 ( .A(n27003), .B(n27159), .Z(n27161) );
  XOR U26980 ( .A(n27168), .B(n27169), .Z(n27003) );
  AND U26981 ( .A(n758), .B(n27170), .Z(n27169) );
  XOR U26982 ( .A(n27153), .B(n27171), .Z(n27159) );
  AND U26983 ( .A(n27172), .B(n27156), .Z(n27171) );
  XNOR U26984 ( .A(n27062), .B(n27153), .Z(n27156) );
  XNOR U26985 ( .A(n27173), .B(n27174), .Z(n27062) );
  AND U26986 ( .A(n750), .B(n27175), .Z(n27174) );
  XOR U26987 ( .A(n27176), .B(n27173), .Z(n27175) );
  XNOR U26988 ( .A(n27177), .B(n27153), .Z(n27172) );
  IV U26989 ( .A(n27013), .Z(n27177) );
  XOR U26990 ( .A(n27178), .B(n27179), .Z(n27013) );
  AND U26991 ( .A(n758), .B(n27180), .Z(n27179) );
  XOR U26992 ( .A(n27181), .B(n27182), .Z(n27153) );
  AND U26993 ( .A(n27183), .B(n27184), .Z(n27182) );
  XNOR U26994 ( .A(n27087), .B(n27181), .Z(n27184) );
  XNOR U26995 ( .A(n27185), .B(n27186), .Z(n27087) );
  AND U26996 ( .A(n750), .B(n27187), .Z(n27186) );
  XNOR U26997 ( .A(n27188), .B(n27185), .Z(n27187) );
  XOR U26998 ( .A(n27181), .B(n27024), .Z(n27183) );
  XOR U26999 ( .A(n27189), .B(n27190), .Z(n27024) );
  AND U27000 ( .A(n758), .B(n27191), .Z(n27190) );
  XOR U27001 ( .A(n27192), .B(n27193), .Z(n27181) );
  AND U27002 ( .A(n27194), .B(n27195), .Z(n27193) );
  XNOR U27003 ( .A(n27192), .B(n27135), .Z(n27195) );
  XNOR U27004 ( .A(n27196), .B(n27197), .Z(n27135) );
  AND U27005 ( .A(n750), .B(n27198), .Z(n27197) );
  XOR U27006 ( .A(n27199), .B(n27196), .Z(n27198) );
  XNOR U27007 ( .A(n27200), .B(n27192), .Z(n27194) );
  IV U27008 ( .A(n27036), .Z(n27200) );
  XOR U27009 ( .A(n27201), .B(n27202), .Z(n27036) );
  AND U27010 ( .A(n758), .B(n27203), .Z(n27202) );
  AND U27011 ( .A(n27157), .B(n27146), .Z(n27192) );
  XNOR U27012 ( .A(n27204), .B(n27205), .Z(n27146) );
  AND U27013 ( .A(n750), .B(n27206), .Z(n27205) );
  XNOR U27014 ( .A(n27207), .B(n27204), .Z(n27206) );
  XNOR U27015 ( .A(n27208), .B(n27209), .Z(n750) );
  AND U27016 ( .A(n27210), .B(n27211), .Z(n27209) );
  XOR U27017 ( .A(n27167), .B(n27208), .Z(n27211) );
  AND U27018 ( .A(n27212), .B(n27213), .Z(n27167) );
  XOR U27019 ( .A(n27208), .B(n27164), .Z(n27210) );
  XNOR U27020 ( .A(n27214), .B(n27215), .Z(n27164) );
  AND U27021 ( .A(n754), .B(n27170), .Z(n27215) );
  XOR U27022 ( .A(n27168), .B(n27214), .Z(n27170) );
  XOR U27023 ( .A(n27216), .B(n27217), .Z(n27208) );
  AND U27024 ( .A(n27218), .B(n27219), .Z(n27217) );
  XNOR U27025 ( .A(n27216), .B(n27212), .Z(n27219) );
  IV U27026 ( .A(n27176), .Z(n27212) );
  XOR U27027 ( .A(n27220), .B(n27221), .Z(n27176) );
  XOR U27028 ( .A(n27222), .B(n27213), .Z(n27221) );
  AND U27029 ( .A(n27188), .B(n27223), .Z(n27213) );
  AND U27030 ( .A(n27224), .B(n27225), .Z(n27222) );
  XOR U27031 ( .A(n27226), .B(n27220), .Z(n27224) );
  XNOR U27032 ( .A(n27173), .B(n27216), .Z(n27218) );
  XNOR U27033 ( .A(n27227), .B(n27228), .Z(n27173) );
  AND U27034 ( .A(n754), .B(n27180), .Z(n27228) );
  XOR U27035 ( .A(n27227), .B(n27178), .Z(n27180) );
  XOR U27036 ( .A(n27229), .B(n27230), .Z(n27216) );
  AND U27037 ( .A(n27231), .B(n27232), .Z(n27230) );
  XNOR U27038 ( .A(n27229), .B(n27188), .Z(n27232) );
  XOR U27039 ( .A(n27233), .B(n27225), .Z(n27188) );
  XNOR U27040 ( .A(n27234), .B(n27220), .Z(n27225) );
  XOR U27041 ( .A(n27235), .B(n27236), .Z(n27220) );
  AND U27042 ( .A(n27237), .B(n27238), .Z(n27236) );
  XOR U27043 ( .A(n27239), .B(n27235), .Z(n27237) );
  XNOR U27044 ( .A(n27240), .B(n27241), .Z(n27234) );
  AND U27045 ( .A(n27242), .B(n27243), .Z(n27241) );
  XOR U27046 ( .A(n27240), .B(n27244), .Z(n27242) );
  XNOR U27047 ( .A(n27226), .B(n27223), .Z(n27233) );
  AND U27048 ( .A(n27245), .B(n27246), .Z(n27223) );
  XOR U27049 ( .A(n27247), .B(n27248), .Z(n27226) );
  AND U27050 ( .A(n27249), .B(n27250), .Z(n27248) );
  XOR U27051 ( .A(n27247), .B(n27251), .Z(n27249) );
  XNOR U27052 ( .A(n27185), .B(n27229), .Z(n27231) );
  XNOR U27053 ( .A(n27252), .B(n27253), .Z(n27185) );
  AND U27054 ( .A(n754), .B(n27191), .Z(n27253) );
  XOR U27055 ( .A(n27252), .B(n27189), .Z(n27191) );
  XOR U27056 ( .A(n27254), .B(n27255), .Z(n27229) );
  AND U27057 ( .A(n27256), .B(n27257), .Z(n27255) );
  XNOR U27058 ( .A(n27254), .B(n27245), .Z(n27257) );
  IV U27059 ( .A(n27199), .Z(n27245) );
  XNOR U27060 ( .A(n27258), .B(n27238), .Z(n27199) );
  XNOR U27061 ( .A(n27259), .B(n27244), .Z(n27238) );
  XNOR U27062 ( .A(n27260), .B(n27261), .Z(n27244) );
  NOR U27063 ( .A(n27262), .B(n27263), .Z(n27261) );
  XOR U27064 ( .A(n27260), .B(n27264), .Z(n27262) );
  XNOR U27065 ( .A(n27243), .B(n27235), .Z(n27259) );
  XOR U27066 ( .A(n27265), .B(n27266), .Z(n27235) );
  AND U27067 ( .A(n27267), .B(n27268), .Z(n27266) );
  XOR U27068 ( .A(n27265), .B(n27269), .Z(n27267) );
  XNOR U27069 ( .A(n27270), .B(n27240), .Z(n27243) );
  XOR U27070 ( .A(n27271), .B(n27272), .Z(n27240) );
  AND U27071 ( .A(n27273), .B(n27274), .Z(n27272) );
  XNOR U27072 ( .A(n27275), .B(n27276), .Z(n27273) );
  IV U27073 ( .A(n27271), .Z(n27275) );
  XNOR U27074 ( .A(n27277), .B(n27278), .Z(n27270) );
  NOR U27075 ( .A(n27279), .B(n27280), .Z(n27278) );
  XNOR U27076 ( .A(n27277), .B(n27281), .Z(n27279) );
  XNOR U27077 ( .A(n27239), .B(n27246), .Z(n27258) );
  NOR U27078 ( .A(n27207), .B(n27282), .Z(n27246) );
  XOR U27079 ( .A(n27251), .B(n27250), .Z(n27239) );
  XNOR U27080 ( .A(n27283), .B(n27247), .Z(n27250) );
  XOR U27081 ( .A(n27284), .B(n27285), .Z(n27247) );
  AND U27082 ( .A(n27286), .B(n27287), .Z(n27285) );
  XNOR U27083 ( .A(n27288), .B(n27289), .Z(n27286) );
  IV U27084 ( .A(n27284), .Z(n27288) );
  XNOR U27085 ( .A(n27290), .B(n27291), .Z(n27283) );
  NOR U27086 ( .A(n27292), .B(n27293), .Z(n27291) );
  XNOR U27087 ( .A(n27290), .B(n27294), .Z(n27292) );
  XOR U27088 ( .A(n27295), .B(n27296), .Z(n27251) );
  NOR U27089 ( .A(n27297), .B(n27298), .Z(n27296) );
  XNOR U27090 ( .A(n27295), .B(n27299), .Z(n27297) );
  XNOR U27091 ( .A(n27196), .B(n27254), .Z(n27256) );
  XNOR U27092 ( .A(n27300), .B(n27301), .Z(n27196) );
  AND U27093 ( .A(n754), .B(n27203), .Z(n27301) );
  XOR U27094 ( .A(n27300), .B(n27201), .Z(n27203) );
  AND U27095 ( .A(n27204), .B(n27207), .Z(n27254) );
  XOR U27096 ( .A(n27302), .B(n27282), .Z(n27207) );
  XNOR U27097 ( .A(p_input[1040]), .B(p_input[2048]), .Z(n27282) );
  XNOR U27098 ( .A(n27269), .B(n27268), .Z(n27302) );
  XNOR U27099 ( .A(n27303), .B(n27276), .Z(n27268) );
  XNOR U27100 ( .A(n27264), .B(n27263), .Z(n27276) );
  XNOR U27101 ( .A(n27304), .B(n27260), .Z(n27263) );
  XNOR U27102 ( .A(p_input[1050]), .B(p_input[2058]), .Z(n27260) );
  XOR U27103 ( .A(p_input[1051]), .B(n16732), .Z(n27304) );
  XOR U27104 ( .A(p_input[1052]), .B(p_input[2060]), .Z(n27264) );
  XOR U27105 ( .A(n27274), .B(n27305), .Z(n27303) );
  IV U27106 ( .A(n27265), .Z(n27305) );
  XOR U27107 ( .A(p_input[1041]), .B(p_input[2049]), .Z(n27265) );
  XNOR U27108 ( .A(n27306), .B(n27281), .Z(n27274) );
  XNOR U27109 ( .A(p_input[1055]), .B(n16735), .Z(n27281) );
  XOR U27110 ( .A(n27271), .B(n27280), .Z(n27306) );
  XOR U27111 ( .A(n27307), .B(n27277), .Z(n27280) );
  XOR U27112 ( .A(p_input[1053]), .B(p_input[2061]), .Z(n27277) );
  XOR U27113 ( .A(p_input[1054]), .B(n16737), .Z(n27307) );
  XOR U27114 ( .A(p_input[1049]), .B(p_input[2057]), .Z(n27271) );
  XOR U27115 ( .A(n27289), .B(n27287), .Z(n27269) );
  XNOR U27116 ( .A(n27308), .B(n27294), .Z(n27287) );
  XOR U27117 ( .A(p_input[1048]), .B(p_input[2056]), .Z(n27294) );
  XOR U27118 ( .A(n27284), .B(n27293), .Z(n27308) );
  XOR U27119 ( .A(n27309), .B(n27290), .Z(n27293) );
  XOR U27120 ( .A(p_input[1046]), .B(p_input[2054]), .Z(n27290) );
  XOR U27121 ( .A(p_input[1047]), .B(n17722), .Z(n27309) );
  XOR U27122 ( .A(p_input[1042]), .B(p_input[2050]), .Z(n27284) );
  XNOR U27123 ( .A(n27299), .B(n27298), .Z(n27289) );
  XOR U27124 ( .A(n27310), .B(n27295), .Z(n27298) );
  XOR U27125 ( .A(p_input[1043]), .B(p_input[2051]), .Z(n27295) );
  XOR U27126 ( .A(p_input[1044]), .B(n17724), .Z(n27310) );
  XOR U27127 ( .A(p_input[1045]), .B(p_input[2053]), .Z(n27299) );
  XNOR U27128 ( .A(n27311), .B(n27312), .Z(n27204) );
  AND U27129 ( .A(n754), .B(n27313), .Z(n27312) );
  XNOR U27130 ( .A(n27314), .B(n27315), .Z(n754) );
  AND U27131 ( .A(n27316), .B(n27317), .Z(n27315) );
  XOR U27132 ( .A(n27314), .B(n27214), .Z(n27317) );
  XNOR U27133 ( .A(n27314), .B(n27168), .Z(n27316) );
  XOR U27134 ( .A(n27318), .B(n27319), .Z(n27314) );
  AND U27135 ( .A(n27320), .B(n27321), .Z(n27319) );
  XOR U27136 ( .A(n27318), .B(n27178), .Z(n27320) );
  XOR U27137 ( .A(n27322), .B(n27323), .Z(n27157) );
  AND U27138 ( .A(n758), .B(n27313), .Z(n27323) );
  XNOR U27139 ( .A(n27311), .B(n27322), .Z(n27313) );
  XNOR U27140 ( .A(n27324), .B(n27325), .Z(n758) );
  AND U27141 ( .A(n27326), .B(n27327), .Z(n27325) );
  XNOR U27142 ( .A(n27328), .B(n27324), .Z(n27327) );
  IV U27143 ( .A(n27214), .Z(n27328) );
  XNOR U27144 ( .A(n27329), .B(n27330), .Z(n27214) );
  AND U27145 ( .A(n761), .B(n27331), .Z(n27330) );
  XNOR U27146 ( .A(n27329), .B(n27332), .Z(n27331) );
  XNOR U27147 ( .A(n27168), .B(n27324), .Z(n27326) );
  XOR U27148 ( .A(n27333), .B(n27334), .Z(n27168) );
  AND U27149 ( .A(n769), .B(n27335), .Z(n27334) );
  XOR U27150 ( .A(n27318), .B(n27336), .Z(n27324) );
  AND U27151 ( .A(n27337), .B(n27321), .Z(n27336) );
  XNOR U27152 ( .A(n27227), .B(n27318), .Z(n27321) );
  XNOR U27153 ( .A(n27338), .B(n27339), .Z(n27227) );
  AND U27154 ( .A(n761), .B(n27340), .Z(n27339) );
  XOR U27155 ( .A(n27341), .B(n27338), .Z(n27340) );
  XNOR U27156 ( .A(n27342), .B(n27318), .Z(n27337) );
  IV U27157 ( .A(n27178), .Z(n27342) );
  XOR U27158 ( .A(n27343), .B(n27344), .Z(n27178) );
  AND U27159 ( .A(n769), .B(n27345), .Z(n27344) );
  XOR U27160 ( .A(n27346), .B(n27347), .Z(n27318) );
  AND U27161 ( .A(n27348), .B(n27349), .Z(n27347) );
  XNOR U27162 ( .A(n27252), .B(n27346), .Z(n27349) );
  XNOR U27163 ( .A(n27350), .B(n27351), .Z(n27252) );
  AND U27164 ( .A(n761), .B(n27352), .Z(n27351) );
  XNOR U27165 ( .A(n27353), .B(n27350), .Z(n27352) );
  XOR U27166 ( .A(n27346), .B(n27189), .Z(n27348) );
  XOR U27167 ( .A(n27354), .B(n27355), .Z(n27189) );
  AND U27168 ( .A(n769), .B(n27356), .Z(n27355) );
  XOR U27169 ( .A(n27357), .B(n27358), .Z(n27346) );
  AND U27170 ( .A(n27359), .B(n27360), .Z(n27358) );
  XNOR U27171 ( .A(n27357), .B(n27300), .Z(n27360) );
  XNOR U27172 ( .A(n27361), .B(n27362), .Z(n27300) );
  AND U27173 ( .A(n761), .B(n27363), .Z(n27362) );
  XOR U27174 ( .A(n27364), .B(n27361), .Z(n27363) );
  XNOR U27175 ( .A(n27365), .B(n27357), .Z(n27359) );
  IV U27176 ( .A(n27201), .Z(n27365) );
  XOR U27177 ( .A(n27366), .B(n27367), .Z(n27201) );
  AND U27178 ( .A(n769), .B(n27368), .Z(n27367) );
  AND U27179 ( .A(n27322), .B(n27311), .Z(n27357) );
  XNOR U27180 ( .A(n27369), .B(n27370), .Z(n27311) );
  AND U27181 ( .A(n761), .B(n27371), .Z(n27370) );
  XNOR U27182 ( .A(n27372), .B(n27369), .Z(n27371) );
  XNOR U27183 ( .A(n27373), .B(n27374), .Z(n761) );
  AND U27184 ( .A(n27375), .B(n27376), .Z(n27374) );
  XOR U27185 ( .A(n27332), .B(n27373), .Z(n27376) );
  AND U27186 ( .A(n27377), .B(n27378), .Z(n27332) );
  XOR U27187 ( .A(n27373), .B(n27329), .Z(n27375) );
  XNOR U27188 ( .A(n27379), .B(n27380), .Z(n27329) );
  AND U27189 ( .A(n765), .B(n27335), .Z(n27380) );
  XOR U27190 ( .A(n27333), .B(n27379), .Z(n27335) );
  XOR U27191 ( .A(n27381), .B(n27382), .Z(n27373) );
  AND U27192 ( .A(n27383), .B(n27384), .Z(n27382) );
  XNOR U27193 ( .A(n27381), .B(n27377), .Z(n27384) );
  IV U27194 ( .A(n27341), .Z(n27377) );
  XOR U27195 ( .A(n27385), .B(n27386), .Z(n27341) );
  XOR U27196 ( .A(n27387), .B(n27378), .Z(n27386) );
  AND U27197 ( .A(n27353), .B(n27388), .Z(n27378) );
  AND U27198 ( .A(n27389), .B(n27390), .Z(n27387) );
  XOR U27199 ( .A(n27391), .B(n27385), .Z(n27389) );
  XNOR U27200 ( .A(n27338), .B(n27381), .Z(n27383) );
  XNOR U27201 ( .A(n27392), .B(n27393), .Z(n27338) );
  AND U27202 ( .A(n765), .B(n27345), .Z(n27393) );
  XOR U27203 ( .A(n27392), .B(n27343), .Z(n27345) );
  XOR U27204 ( .A(n27394), .B(n27395), .Z(n27381) );
  AND U27205 ( .A(n27396), .B(n27397), .Z(n27395) );
  XNOR U27206 ( .A(n27394), .B(n27353), .Z(n27397) );
  XOR U27207 ( .A(n27398), .B(n27390), .Z(n27353) );
  XNOR U27208 ( .A(n27399), .B(n27385), .Z(n27390) );
  XOR U27209 ( .A(n27400), .B(n27401), .Z(n27385) );
  AND U27210 ( .A(n27402), .B(n27403), .Z(n27401) );
  XOR U27211 ( .A(n27404), .B(n27400), .Z(n27402) );
  XNOR U27212 ( .A(n27405), .B(n27406), .Z(n27399) );
  AND U27213 ( .A(n27407), .B(n27408), .Z(n27406) );
  XOR U27214 ( .A(n27405), .B(n27409), .Z(n27407) );
  XNOR U27215 ( .A(n27391), .B(n27388), .Z(n27398) );
  AND U27216 ( .A(n27410), .B(n27411), .Z(n27388) );
  XOR U27217 ( .A(n27412), .B(n27413), .Z(n27391) );
  AND U27218 ( .A(n27414), .B(n27415), .Z(n27413) );
  XOR U27219 ( .A(n27412), .B(n27416), .Z(n27414) );
  XNOR U27220 ( .A(n27350), .B(n27394), .Z(n27396) );
  XNOR U27221 ( .A(n27417), .B(n27418), .Z(n27350) );
  AND U27222 ( .A(n765), .B(n27356), .Z(n27418) );
  XOR U27223 ( .A(n27417), .B(n27354), .Z(n27356) );
  XOR U27224 ( .A(n27419), .B(n27420), .Z(n27394) );
  AND U27225 ( .A(n27421), .B(n27422), .Z(n27420) );
  XNOR U27226 ( .A(n27419), .B(n27410), .Z(n27422) );
  IV U27227 ( .A(n27364), .Z(n27410) );
  XNOR U27228 ( .A(n27423), .B(n27403), .Z(n27364) );
  XNOR U27229 ( .A(n27424), .B(n27409), .Z(n27403) );
  XNOR U27230 ( .A(n27425), .B(n27426), .Z(n27409) );
  NOR U27231 ( .A(n27427), .B(n27428), .Z(n27426) );
  XOR U27232 ( .A(n27425), .B(n27429), .Z(n27427) );
  XNOR U27233 ( .A(n27408), .B(n27400), .Z(n27424) );
  XOR U27234 ( .A(n27430), .B(n27431), .Z(n27400) );
  AND U27235 ( .A(n27432), .B(n27433), .Z(n27431) );
  XOR U27236 ( .A(n27430), .B(n27434), .Z(n27432) );
  XNOR U27237 ( .A(n27435), .B(n27405), .Z(n27408) );
  XOR U27238 ( .A(n27436), .B(n27437), .Z(n27405) );
  AND U27239 ( .A(n27438), .B(n27439), .Z(n27437) );
  XNOR U27240 ( .A(n27440), .B(n27441), .Z(n27438) );
  IV U27241 ( .A(n27436), .Z(n27440) );
  XNOR U27242 ( .A(n27442), .B(n27443), .Z(n27435) );
  NOR U27243 ( .A(n27444), .B(n27445), .Z(n27443) );
  XNOR U27244 ( .A(n27442), .B(n27446), .Z(n27444) );
  XNOR U27245 ( .A(n27404), .B(n27411), .Z(n27423) );
  NOR U27246 ( .A(n27372), .B(n27447), .Z(n27411) );
  XOR U27247 ( .A(n27416), .B(n27415), .Z(n27404) );
  XNOR U27248 ( .A(n27448), .B(n27412), .Z(n27415) );
  XOR U27249 ( .A(n27449), .B(n27450), .Z(n27412) );
  AND U27250 ( .A(n27451), .B(n27452), .Z(n27450) );
  XNOR U27251 ( .A(n27453), .B(n27454), .Z(n27451) );
  IV U27252 ( .A(n27449), .Z(n27453) );
  XNOR U27253 ( .A(n27455), .B(n27456), .Z(n27448) );
  NOR U27254 ( .A(n27457), .B(n27458), .Z(n27456) );
  XNOR U27255 ( .A(n27455), .B(n27459), .Z(n27457) );
  XOR U27256 ( .A(n27460), .B(n27461), .Z(n27416) );
  NOR U27257 ( .A(n27462), .B(n27463), .Z(n27461) );
  XNOR U27258 ( .A(n27460), .B(n27464), .Z(n27462) );
  XNOR U27259 ( .A(n27361), .B(n27419), .Z(n27421) );
  XNOR U27260 ( .A(n27465), .B(n27466), .Z(n27361) );
  AND U27261 ( .A(n765), .B(n27368), .Z(n27466) );
  XOR U27262 ( .A(n27465), .B(n27366), .Z(n27368) );
  AND U27263 ( .A(n27369), .B(n27372), .Z(n27419) );
  XOR U27264 ( .A(n27467), .B(n27447), .Z(n27372) );
  XNOR U27265 ( .A(p_input[1056]), .B(p_input[2048]), .Z(n27447) );
  XNOR U27266 ( .A(n27434), .B(n27433), .Z(n27467) );
  XNOR U27267 ( .A(n27468), .B(n27441), .Z(n27433) );
  XNOR U27268 ( .A(n27429), .B(n27428), .Z(n27441) );
  XNOR U27269 ( .A(n27469), .B(n27425), .Z(n27428) );
  XNOR U27270 ( .A(p_input[1066]), .B(p_input[2058]), .Z(n27425) );
  XOR U27271 ( .A(p_input[1067]), .B(n16732), .Z(n27469) );
  XOR U27272 ( .A(p_input[1068]), .B(p_input[2060]), .Z(n27429) );
  XOR U27273 ( .A(n27439), .B(n27470), .Z(n27468) );
  IV U27274 ( .A(n27430), .Z(n27470) );
  XOR U27275 ( .A(p_input[1057]), .B(p_input[2049]), .Z(n27430) );
  XNOR U27276 ( .A(n27471), .B(n27446), .Z(n27439) );
  XNOR U27277 ( .A(p_input[1071]), .B(n16735), .Z(n27446) );
  XOR U27278 ( .A(n27436), .B(n27445), .Z(n27471) );
  XOR U27279 ( .A(n27472), .B(n27442), .Z(n27445) );
  XOR U27280 ( .A(p_input[1069]), .B(p_input[2061]), .Z(n27442) );
  XOR U27281 ( .A(p_input[1070]), .B(n16737), .Z(n27472) );
  XOR U27282 ( .A(p_input[1065]), .B(p_input[2057]), .Z(n27436) );
  XOR U27283 ( .A(n27454), .B(n27452), .Z(n27434) );
  XNOR U27284 ( .A(n27473), .B(n27459), .Z(n27452) );
  XOR U27285 ( .A(p_input[1064]), .B(p_input[2056]), .Z(n27459) );
  XOR U27286 ( .A(n27449), .B(n27458), .Z(n27473) );
  XOR U27287 ( .A(n27474), .B(n27455), .Z(n27458) );
  XOR U27288 ( .A(p_input[1062]), .B(p_input[2054]), .Z(n27455) );
  XOR U27289 ( .A(p_input[1063]), .B(n17722), .Z(n27474) );
  XOR U27290 ( .A(p_input[1058]), .B(p_input[2050]), .Z(n27449) );
  XNOR U27291 ( .A(n27464), .B(n27463), .Z(n27454) );
  XOR U27292 ( .A(n27475), .B(n27460), .Z(n27463) );
  XOR U27293 ( .A(p_input[1059]), .B(p_input[2051]), .Z(n27460) );
  XOR U27294 ( .A(p_input[1060]), .B(n17724), .Z(n27475) );
  XOR U27295 ( .A(p_input[1061]), .B(p_input[2053]), .Z(n27464) );
  XNOR U27296 ( .A(n27476), .B(n27477), .Z(n27369) );
  AND U27297 ( .A(n765), .B(n27478), .Z(n27477) );
  XNOR U27298 ( .A(n27479), .B(n27480), .Z(n765) );
  AND U27299 ( .A(n27481), .B(n27482), .Z(n27480) );
  XOR U27300 ( .A(n27479), .B(n27379), .Z(n27482) );
  XNOR U27301 ( .A(n27479), .B(n27333), .Z(n27481) );
  XOR U27302 ( .A(n27483), .B(n27484), .Z(n27479) );
  AND U27303 ( .A(n27485), .B(n27486), .Z(n27484) );
  XOR U27304 ( .A(n27483), .B(n27343), .Z(n27485) );
  XOR U27305 ( .A(n27487), .B(n27488), .Z(n27322) );
  AND U27306 ( .A(n769), .B(n27478), .Z(n27488) );
  XNOR U27307 ( .A(n27476), .B(n27487), .Z(n27478) );
  XNOR U27308 ( .A(n27489), .B(n27490), .Z(n769) );
  AND U27309 ( .A(n27491), .B(n27492), .Z(n27490) );
  XNOR U27310 ( .A(n27493), .B(n27489), .Z(n27492) );
  IV U27311 ( .A(n27379), .Z(n27493) );
  XNOR U27312 ( .A(n27494), .B(n27495), .Z(n27379) );
  AND U27313 ( .A(n772), .B(n27496), .Z(n27495) );
  XNOR U27314 ( .A(n27494), .B(n27497), .Z(n27496) );
  XNOR U27315 ( .A(n27333), .B(n27489), .Z(n27491) );
  XOR U27316 ( .A(n27498), .B(n27499), .Z(n27333) );
  AND U27317 ( .A(n780), .B(n27500), .Z(n27499) );
  XOR U27318 ( .A(n27483), .B(n27501), .Z(n27489) );
  AND U27319 ( .A(n27502), .B(n27486), .Z(n27501) );
  XNOR U27320 ( .A(n27392), .B(n27483), .Z(n27486) );
  XNOR U27321 ( .A(n27503), .B(n27504), .Z(n27392) );
  AND U27322 ( .A(n772), .B(n27505), .Z(n27504) );
  XOR U27323 ( .A(n27506), .B(n27503), .Z(n27505) );
  XNOR U27324 ( .A(n27507), .B(n27483), .Z(n27502) );
  IV U27325 ( .A(n27343), .Z(n27507) );
  XOR U27326 ( .A(n27508), .B(n27509), .Z(n27343) );
  AND U27327 ( .A(n780), .B(n27510), .Z(n27509) );
  XOR U27328 ( .A(n27511), .B(n27512), .Z(n27483) );
  AND U27329 ( .A(n27513), .B(n27514), .Z(n27512) );
  XNOR U27330 ( .A(n27417), .B(n27511), .Z(n27514) );
  XNOR U27331 ( .A(n27515), .B(n27516), .Z(n27417) );
  AND U27332 ( .A(n772), .B(n27517), .Z(n27516) );
  XNOR U27333 ( .A(n27518), .B(n27515), .Z(n27517) );
  XOR U27334 ( .A(n27511), .B(n27354), .Z(n27513) );
  XOR U27335 ( .A(n27519), .B(n27520), .Z(n27354) );
  AND U27336 ( .A(n780), .B(n27521), .Z(n27520) );
  XOR U27337 ( .A(n27522), .B(n27523), .Z(n27511) );
  AND U27338 ( .A(n27524), .B(n27525), .Z(n27523) );
  XNOR U27339 ( .A(n27522), .B(n27465), .Z(n27525) );
  XNOR U27340 ( .A(n27526), .B(n27527), .Z(n27465) );
  AND U27341 ( .A(n772), .B(n27528), .Z(n27527) );
  XOR U27342 ( .A(n27529), .B(n27526), .Z(n27528) );
  XNOR U27343 ( .A(n27530), .B(n27522), .Z(n27524) );
  IV U27344 ( .A(n27366), .Z(n27530) );
  XOR U27345 ( .A(n27531), .B(n27532), .Z(n27366) );
  AND U27346 ( .A(n780), .B(n27533), .Z(n27532) );
  AND U27347 ( .A(n27487), .B(n27476), .Z(n27522) );
  XNOR U27348 ( .A(n27534), .B(n27535), .Z(n27476) );
  AND U27349 ( .A(n772), .B(n27536), .Z(n27535) );
  XNOR U27350 ( .A(n27537), .B(n27534), .Z(n27536) );
  XNOR U27351 ( .A(n27538), .B(n27539), .Z(n772) );
  AND U27352 ( .A(n27540), .B(n27541), .Z(n27539) );
  XOR U27353 ( .A(n27497), .B(n27538), .Z(n27541) );
  AND U27354 ( .A(n27542), .B(n27543), .Z(n27497) );
  XOR U27355 ( .A(n27538), .B(n27494), .Z(n27540) );
  XNOR U27356 ( .A(n27544), .B(n27545), .Z(n27494) );
  AND U27357 ( .A(n776), .B(n27500), .Z(n27545) );
  XOR U27358 ( .A(n27498), .B(n27544), .Z(n27500) );
  XOR U27359 ( .A(n27546), .B(n27547), .Z(n27538) );
  AND U27360 ( .A(n27548), .B(n27549), .Z(n27547) );
  XNOR U27361 ( .A(n27546), .B(n27542), .Z(n27549) );
  IV U27362 ( .A(n27506), .Z(n27542) );
  XOR U27363 ( .A(n27550), .B(n27551), .Z(n27506) );
  XOR U27364 ( .A(n27552), .B(n27543), .Z(n27551) );
  AND U27365 ( .A(n27518), .B(n27553), .Z(n27543) );
  AND U27366 ( .A(n27554), .B(n27555), .Z(n27552) );
  XOR U27367 ( .A(n27556), .B(n27550), .Z(n27554) );
  XNOR U27368 ( .A(n27503), .B(n27546), .Z(n27548) );
  XNOR U27369 ( .A(n27557), .B(n27558), .Z(n27503) );
  AND U27370 ( .A(n776), .B(n27510), .Z(n27558) );
  XOR U27371 ( .A(n27557), .B(n27508), .Z(n27510) );
  XOR U27372 ( .A(n27559), .B(n27560), .Z(n27546) );
  AND U27373 ( .A(n27561), .B(n27562), .Z(n27560) );
  XNOR U27374 ( .A(n27559), .B(n27518), .Z(n27562) );
  XOR U27375 ( .A(n27563), .B(n27555), .Z(n27518) );
  XNOR U27376 ( .A(n27564), .B(n27550), .Z(n27555) );
  XOR U27377 ( .A(n27565), .B(n27566), .Z(n27550) );
  AND U27378 ( .A(n27567), .B(n27568), .Z(n27566) );
  XOR U27379 ( .A(n27569), .B(n27565), .Z(n27567) );
  XNOR U27380 ( .A(n27570), .B(n27571), .Z(n27564) );
  AND U27381 ( .A(n27572), .B(n27573), .Z(n27571) );
  XOR U27382 ( .A(n27570), .B(n27574), .Z(n27572) );
  XNOR U27383 ( .A(n27556), .B(n27553), .Z(n27563) );
  AND U27384 ( .A(n27575), .B(n27576), .Z(n27553) );
  XOR U27385 ( .A(n27577), .B(n27578), .Z(n27556) );
  AND U27386 ( .A(n27579), .B(n27580), .Z(n27578) );
  XOR U27387 ( .A(n27577), .B(n27581), .Z(n27579) );
  XNOR U27388 ( .A(n27515), .B(n27559), .Z(n27561) );
  XNOR U27389 ( .A(n27582), .B(n27583), .Z(n27515) );
  AND U27390 ( .A(n776), .B(n27521), .Z(n27583) );
  XOR U27391 ( .A(n27582), .B(n27519), .Z(n27521) );
  XOR U27392 ( .A(n27584), .B(n27585), .Z(n27559) );
  AND U27393 ( .A(n27586), .B(n27587), .Z(n27585) );
  XNOR U27394 ( .A(n27584), .B(n27575), .Z(n27587) );
  IV U27395 ( .A(n27529), .Z(n27575) );
  XNOR U27396 ( .A(n27588), .B(n27568), .Z(n27529) );
  XNOR U27397 ( .A(n27589), .B(n27574), .Z(n27568) );
  XNOR U27398 ( .A(n27590), .B(n27591), .Z(n27574) );
  NOR U27399 ( .A(n27592), .B(n27593), .Z(n27591) );
  XOR U27400 ( .A(n27590), .B(n27594), .Z(n27592) );
  XNOR U27401 ( .A(n27573), .B(n27565), .Z(n27589) );
  XOR U27402 ( .A(n27595), .B(n27596), .Z(n27565) );
  AND U27403 ( .A(n27597), .B(n27598), .Z(n27596) );
  XOR U27404 ( .A(n27595), .B(n27599), .Z(n27597) );
  XNOR U27405 ( .A(n27600), .B(n27570), .Z(n27573) );
  XOR U27406 ( .A(n27601), .B(n27602), .Z(n27570) );
  AND U27407 ( .A(n27603), .B(n27604), .Z(n27602) );
  XNOR U27408 ( .A(n27605), .B(n27606), .Z(n27603) );
  IV U27409 ( .A(n27601), .Z(n27605) );
  XNOR U27410 ( .A(n27607), .B(n27608), .Z(n27600) );
  NOR U27411 ( .A(n27609), .B(n27610), .Z(n27608) );
  XNOR U27412 ( .A(n27607), .B(n27611), .Z(n27609) );
  XNOR U27413 ( .A(n27569), .B(n27576), .Z(n27588) );
  NOR U27414 ( .A(n27537), .B(n27612), .Z(n27576) );
  XOR U27415 ( .A(n27581), .B(n27580), .Z(n27569) );
  XNOR U27416 ( .A(n27613), .B(n27577), .Z(n27580) );
  XOR U27417 ( .A(n27614), .B(n27615), .Z(n27577) );
  AND U27418 ( .A(n27616), .B(n27617), .Z(n27615) );
  XNOR U27419 ( .A(n27618), .B(n27619), .Z(n27616) );
  IV U27420 ( .A(n27614), .Z(n27618) );
  XNOR U27421 ( .A(n27620), .B(n27621), .Z(n27613) );
  NOR U27422 ( .A(n27622), .B(n27623), .Z(n27621) );
  XNOR U27423 ( .A(n27620), .B(n27624), .Z(n27622) );
  XOR U27424 ( .A(n27625), .B(n27626), .Z(n27581) );
  NOR U27425 ( .A(n27627), .B(n27628), .Z(n27626) );
  XNOR U27426 ( .A(n27625), .B(n27629), .Z(n27627) );
  XNOR U27427 ( .A(n27526), .B(n27584), .Z(n27586) );
  XNOR U27428 ( .A(n27630), .B(n27631), .Z(n27526) );
  AND U27429 ( .A(n776), .B(n27533), .Z(n27631) );
  XOR U27430 ( .A(n27630), .B(n27531), .Z(n27533) );
  AND U27431 ( .A(n27534), .B(n27537), .Z(n27584) );
  XOR U27432 ( .A(n27632), .B(n27612), .Z(n27537) );
  XNOR U27433 ( .A(p_input[1072]), .B(p_input[2048]), .Z(n27612) );
  XNOR U27434 ( .A(n27599), .B(n27598), .Z(n27632) );
  XNOR U27435 ( .A(n27633), .B(n27606), .Z(n27598) );
  XNOR U27436 ( .A(n27594), .B(n27593), .Z(n27606) );
  XNOR U27437 ( .A(n27634), .B(n27590), .Z(n27593) );
  XNOR U27438 ( .A(p_input[1082]), .B(p_input[2058]), .Z(n27590) );
  XOR U27439 ( .A(p_input[1083]), .B(n16732), .Z(n27634) );
  XOR U27440 ( .A(p_input[1084]), .B(p_input[2060]), .Z(n27594) );
  XOR U27441 ( .A(n27604), .B(n27635), .Z(n27633) );
  IV U27442 ( .A(n27595), .Z(n27635) );
  XOR U27443 ( .A(p_input[1073]), .B(p_input[2049]), .Z(n27595) );
  XNOR U27444 ( .A(n27636), .B(n27611), .Z(n27604) );
  XNOR U27445 ( .A(p_input[1087]), .B(n16735), .Z(n27611) );
  XOR U27446 ( .A(n27601), .B(n27610), .Z(n27636) );
  XOR U27447 ( .A(n27637), .B(n27607), .Z(n27610) );
  XOR U27448 ( .A(p_input[1085]), .B(p_input[2061]), .Z(n27607) );
  XOR U27449 ( .A(p_input[1086]), .B(n16737), .Z(n27637) );
  XOR U27450 ( .A(p_input[1081]), .B(p_input[2057]), .Z(n27601) );
  XOR U27451 ( .A(n27619), .B(n27617), .Z(n27599) );
  XNOR U27452 ( .A(n27638), .B(n27624), .Z(n27617) );
  XOR U27453 ( .A(p_input[1080]), .B(p_input[2056]), .Z(n27624) );
  XOR U27454 ( .A(n27614), .B(n27623), .Z(n27638) );
  XOR U27455 ( .A(n27639), .B(n27620), .Z(n27623) );
  XOR U27456 ( .A(p_input[1078]), .B(p_input[2054]), .Z(n27620) );
  XOR U27457 ( .A(p_input[1079]), .B(n17722), .Z(n27639) );
  XOR U27458 ( .A(p_input[1074]), .B(p_input[2050]), .Z(n27614) );
  XNOR U27459 ( .A(n27629), .B(n27628), .Z(n27619) );
  XOR U27460 ( .A(n27640), .B(n27625), .Z(n27628) );
  XOR U27461 ( .A(p_input[1075]), .B(p_input[2051]), .Z(n27625) );
  XOR U27462 ( .A(p_input[1076]), .B(n17724), .Z(n27640) );
  XOR U27463 ( .A(p_input[1077]), .B(p_input[2053]), .Z(n27629) );
  XNOR U27464 ( .A(n27641), .B(n27642), .Z(n27534) );
  AND U27465 ( .A(n776), .B(n27643), .Z(n27642) );
  XNOR U27466 ( .A(n27644), .B(n27645), .Z(n776) );
  AND U27467 ( .A(n27646), .B(n27647), .Z(n27645) );
  XOR U27468 ( .A(n27644), .B(n27544), .Z(n27647) );
  XNOR U27469 ( .A(n27644), .B(n27498), .Z(n27646) );
  XOR U27470 ( .A(n27648), .B(n27649), .Z(n27644) );
  AND U27471 ( .A(n27650), .B(n27651), .Z(n27649) );
  XOR U27472 ( .A(n27648), .B(n27508), .Z(n27650) );
  XOR U27473 ( .A(n27652), .B(n27653), .Z(n27487) );
  AND U27474 ( .A(n780), .B(n27643), .Z(n27653) );
  XNOR U27475 ( .A(n27641), .B(n27652), .Z(n27643) );
  XNOR U27476 ( .A(n27654), .B(n27655), .Z(n780) );
  AND U27477 ( .A(n27656), .B(n27657), .Z(n27655) );
  XNOR U27478 ( .A(n27658), .B(n27654), .Z(n27657) );
  IV U27479 ( .A(n27544), .Z(n27658) );
  XNOR U27480 ( .A(n27659), .B(n27660), .Z(n27544) );
  AND U27481 ( .A(n783), .B(n27661), .Z(n27660) );
  XNOR U27482 ( .A(n27659), .B(n27662), .Z(n27661) );
  XNOR U27483 ( .A(n27498), .B(n27654), .Z(n27656) );
  XOR U27484 ( .A(n27663), .B(n27664), .Z(n27498) );
  AND U27485 ( .A(n791), .B(n27665), .Z(n27664) );
  XOR U27486 ( .A(n27648), .B(n27666), .Z(n27654) );
  AND U27487 ( .A(n27667), .B(n27651), .Z(n27666) );
  XNOR U27488 ( .A(n27557), .B(n27648), .Z(n27651) );
  XNOR U27489 ( .A(n27668), .B(n27669), .Z(n27557) );
  AND U27490 ( .A(n783), .B(n27670), .Z(n27669) );
  XOR U27491 ( .A(n27671), .B(n27668), .Z(n27670) );
  XNOR U27492 ( .A(n27672), .B(n27648), .Z(n27667) );
  IV U27493 ( .A(n27508), .Z(n27672) );
  XOR U27494 ( .A(n27673), .B(n27674), .Z(n27508) );
  AND U27495 ( .A(n791), .B(n27675), .Z(n27674) );
  XOR U27496 ( .A(n27676), .B(n27677), .Z(n27648) );
  AND U27497 ( .A(n27678), .B(n27679), .Z(n27677) );
  XNOR U27498 ( .A(n27582), .B(n27676), .Z(n27679) );
  XNOR U27499 ( .A(n27680), .B(n27681), .Z(n27582) );
  AND U27500 ( .A(n783), .B(n27682), .Z(n27681) );
  XNOR U27501 ( .A(n27683), .B(n27680), .Z(n27682) );
  XOR U27502 ( .A(n27676), .B(n27519), .Z(n27678) );
  XOR U27503 ( .A(n27684), .B(n27685), .Z(n27519) );
  AND U27504 ( .A(n791), .B(n27686), .Z(n27685) );
  XOR U27505 ( .A(n27687), .B(n27688), .Z(n27676) );
  AND U27506 ( .A(n27689), .B(n27690), .Z(n27688) );
  XNOR U27507 ( .A(n27687), .B(n27630), .Z(n27690) );
  XNOR U27508 ( .A(n27691), .B(n27692), .Z(n27630) );
  AND U27509 ( .A(n783), .B(n27693), .Z(n27692) );
  XOR U27510 ( .A(n27694), .B(n27691), .Z(n27693) );
  XNOR U27511 ( .A(n27695), .B(n27687), .Z(n27689) );
  IV U27512 ( .A(n27531), .Z(n27695) );
  XOR U27513 ( .A(n27696), .B(n27697), .Z(n27531) );
  AND U27514 ( .A(n791), .B(n27698), .Z(n27697) );
  AND U27515 ( .A(n27652), .B(n27641), .Z(n27687) );
  XNOR U27516 ( .A(n27699), .B(n27700), .Z(n27641) );
  AND U27517 ( .A(n783), .B(n27701), .Z(n27700) );
  XNOR U27518 ( .A(n27702), .B(n27699), .Z(n27701) );
  XNOR U27519 ( .A(n27703), .B(n27704), .Z(n783) );
  AND U27520 ( .A(n27705), .B(n27706), .Z(n27704) );
  XOR U27521 ( .A(n27662), .B(n27703), .Z(n27706) );
  AND U27522 ( .A(n27707), .B(n27708), .Z(n27662) );
  XOR U27523 ( .A(n27703), .B(n27659), .Z(n27705) );
  XNOR U27524 ( .A(n27709), .B(n27710), .Z(n27659) );
  AND U27525 ( .A(n787), .B(n27665), .Z(n27710) );
  XOR U27526 ( .A(n27663), .B(n27709), .Z(n27665) );
  XOR U27527 ( .A(n27711), .B(n27712), .Z(n27703) );
  AND U27528 ( .A(n27713), .B(n27714), .Z(n27712) );
  XNOR U27529 ( .A(n27711), .B(n27707), .Z(n27714) );
  IV U27530 ( .A(n27671), .Z(n27707) );
  XOR U27531 ( .A(n27715), .B(n27716), .Z(n27671) );
  XOR U27532 ( .A(n27717), .B(n27708), .Z(n27716) );
  AND U27533 ( .A(n27683), .B(n27718), .Z(n27708) );
  AND U27534 ( .A(n27719), .B(n27720), .Z(n27717) );
  XOR U27535 ( .A(n27721), .B(n27715), .Z(n27719) );
  XNOR U27536 ( .A(n27668), .B(n27711), .Z(n27713) );
  XNOR U27537 ( .A(n27722), .B(n27723), .Z(n27668) );
  AND U27538 ( .A(n787), .B(n27675), .Z(n27723) );
  XOR U27539 ( .A(n27722), .B(n27673), .Z(n27675) );
  XOR U27540 ( .A(n27724), .B(n27725), .Z(n27711) );
  AND U27541 ( .A(n27726), .B(n27727), .Z(n27725) );
  XNOR U27542 ( .A(n27724), .B(n27683), .Z(n27727) );
  XOR U27543 ( .A(n27728), .B(n27720), .Z(n27683) );
  XNOR U27544 ( .A(n27729), .B(n27715), .Z(n27720) );
  XOR U27545 ( .A(n27730), .B(n27731), .Z(n27715) );
  AND U27546 ( .A(n27732), .B(n27733), .Z(n27731) );
  XOR U27547 ( .A(n27734), .B(n27730), .Z(n27732) );
  XNOR U27548 ( .A(n27735), .B(n27736), .Z(n27729) );
  AND U27549 ( .A(n27737), .B(n27738), .Z(n27736) );
  XOR U27550 ( .A(n27735), .B(n27739), .Z(n27737) );
  XNOR U27551 ( .A(n27721), .B(n27718), .Z(n27728) );
  AND U27552 ( .A(n27740), .B(n27741), .Z(n27718) );
  XOR U27553 ( .A(n27742), .B(n27743), .Z(n27721) );
  AND U27554 ( .A(n27744), .B(n27745), .Z(n27743) );
  XOR U27555 ( .A(n27742), .B(n27746), .Z(n27744) );
  XNOR U27556 ( .A(n27680), .B(n27724), .Z(n27726) );
  XNOR U27557 ( .A(n27747), .B(n27748), .Z(n27680) );
  AND U27558 ( .A(n787), .B(n27686), .Z(n27748) );
  XOR U27559 ( .A(n27747), .B(n27684), .Z(n27686) );
  XOR U27560 ( .A(n27749), .B(n27750), .Z(n27724) );
  AND U27561 ( .A(n27751), .B(n27752), .Z(n27750) );
  XNOR U27562 ( .A(n27749), .B(n27740), .Z(n27752) );
  IV U27563 ( .A(n27694), .Z(n27740) );
  XNOR U27564 ( .A(n27753), .B(n27733), .Z(n27694) );
  XNOR U27565 ( .A(n27754), .B(n27739), .Z(n27733) );
  XNOR U27566 ( .A(n27755), .B(n27756), .Z(n27739) );
  NOR U27567 ( .A(n27757), .B(n27758), .Z(n27756) );
  XOR U27568 ( .A(n27755), .B(n27759), .Z(n27757) );
  XNOR U27569 ( .A(n27738), .B(n27730), .Z(n27754) );
  XOR U27570 ( .A(n27760), .B(n27761), .Z(n27730) );
  AND U27571 ( .A(n27762), .B(n27763), .Z(n27761) );
  XOR U27572 ( .A(n27760), .B(n27764), .Z(n27762) );
  XNOR U27573 ( .A(n27765), .B(n27735), .Z(n27738) );
  XOR U27574 ( .A(n27766), .B(n27767), .Z(n27735) );
  AND U27575 ( .A(n27768), .B(n27769), .Z(n27767) );
  XNOR U27576 ( .A(n27770), .B(n27771), .Z(n27768) );
  IV U27577 ( .A(n27766), .Z(n27770) );
  XNOR U27578 ( .A(n27772), .B(n27773), .Z(n27765) );
  NOR U27579 ( .A(n27774), .B(n27775), .Z(n27773) );
  XNOR U27580 ( .A(n27772), .B(n27776), .Z(n27774) );
  XNOR U27581 ( .A(n27734), .B(n27741), .Z(n27753) );
  NOR U27582 ( .A(n27702), .B(n27777), .Z(n27741) );
  XOR U27583 ( .A(n27746), .B(n27745), .Z(n27734) );
  XNOR U27584 ( .A(n27778), .B(n27742), .Z(n27745) );
  XOR U27585 ( .A(n27779), .B(n27780), .Z(n27742) );
  AND U27586 ( .A(n27781), .B(n27782), .Z(n27780) );
  XNOR U27587 ( .A(n27783), .B(n27784), .Z(n27781) );
  IV U27588 ( .A(n27779), .Z(n27783) );
  XNOR U27589 ( .A(n27785), .B(n27786), .Z(n27778) );
  NOR U27590 ( .A(n27787), .B(n27788), .Z(n27786) );
  XNOR U27591 ( .A(n27785), .B(n27789), .Z(n27787) );
  XOR U27592 ( .A(n27790), .B(n27791), .Z(n27746) );
  NOR U27593 ( .A(n27792), .B(n27793), .Z(n27791) );
  XNOR U27594 ( .A(n27790), .B(n27794), .Z(n27792) );
  XNOR U27595 ( .A(n27691), .B(n27749), .Z(n27751) );
  XNOR U27596 ( .A(n27795), .B(n27796), .Z(n27691) );
  AND U27597 ( .A(n787), .B(n27698), .Z(n27796) );
  XOR U27598 ( .A(n27795), .B(n27696), .Z(n27698) );
  AND U27599 ( .A(n27699), .B(n27702), .Z(n27749) );
  XOR U27600 ( .A(n27797), .B(n27777), .Z(n27702) );
  XNOR U27601 ( .A(p_input[1088]), .B(p_input[2048]), .Z(n27777) );
  XNOR U27602 ( .A(n27764), .B(n27763), .Z(n27797) );
  XNOR U27603 ( .A(n27798), .B(n27771), .Z(n27763) );
  XNOR U27604 ( .A(n27759), .B(n27758), .Z(n27771) );
  XNOR U27605 ( .A(n27799), .B(n27755), .Z(n27758) );
  XNOR U27606 ( .A(p_input[1098]), .B(p_input[2058]), .Z(n27755) );
  XOR U27607 ( .A(p_input[1099]), .B(n16732), .Z(n27799) );
  XOR U27608 ( .A(p_input[1100]), .B(p_input[2060]), .Z(n27759) );
  XOR U27609 ( .A(n27769), .B(n27800), .Z(n27798) );
  IV U27610 ( .A(n27760), .Z(n27800) );
  XOR U27611 ( .A(p_input[1089]), .B(p_input[2049]), .Z(n27760) );
  XNOR U27612 ( .A(n27801), .B(n27776), .Z(n27769) );
  XNOR U27613 ( .A(p_input[1103]), .B(n16735), .Z(n27776) );
  XOR U27614 ( .A(n27766), .B(n27775), .Z(n27801) );
  XOR U27615 ( .A(n27802), .B(n27772), .Z(n27775) );
  XOR U27616 ( .A(p_input[1101]), .B(p_input[2061]), .Z(n27772) );
  XOR U27617 ( .A(p_input[1102]), .B(n16737), .Z(n27802) );
  XOR U27618 ( .A(p_input[1097]), .B(p_input[2057]), .Z(n27766) );
  XOR U27619 ( .A(n27784), .B(n27782), .Z(n27764) );
  XNOR U27620 ( .A(n27803), .B(n27789), .Z(n27782) );
  XOR U27621 ( .A(p_input[1096]), .B(p_input[2056]), .Z(n27789) );
  XOR U27622 ( .A(n27779), .B(n27788), .Z(n27803) );
  XOR U27623 ( .A(n27804), .B(n27785), .Z(n27788) );
  XOR U27624 ( .A(p_input[1094]), .B(p_input[2054]), .Z(n27785) );
  XOR U27625 ( .A(p_input[1095]), .B(n17722), .Z(n27804) );
  XOR U27626 ( .A(p_input[1090]), .B(p_input[2050]), .Z(n27779) );
  XNOR U27627 ( .A(n27794), .B(n27793), .Z(n27784) );
  XOR U27628 ( .A(n27805), .B(n27790), .Z(n27793) );
  XOR U27629 ( .A(p_input[1091]), .B(p_input[2051]), .Z(n27790) );
  XOR U27630 ( .A(p_input[1092]), .B(n17724), .Z(n27805) );
  XOR U27631 ( .A(p_input[1093]), .B(p_input[2053]), .Z(n27794) );
  XNOR U27632 ( .A(n27806), .B(n27807), .Z(n27699) );
  AND U27633 ( .A(n787), .B(n27808), .Z(n27807) );
  XNOR U27634 ( .A(n27809), .B(n27810), .Z(n787) );
  AND U27635 ( .A(n27811), .B(n27812), .Z(n27810) );
  XOR U27636 ( .A(n27809), .B(n27709), .Z(n27812) );
  XNOR U27637 ( .A(n27809), .B(n27663), .Z(n27811) );
  XOR U27638 ( .A(n27813), .B(n27814), .Z(n27809) );
  AND U27639 ( .A(n27815), .B(n27816), .Z(n27814) );
  XOR U27640 ( .A(n27813), .B(n27673), .Z(n27815) );
  XOR U27641 ( .A(n27817), .B(n27818), .Z(n27652) );
  AND U27642 ( .A(n791), .B(n27808), .Z(n27818) );
  XNOR U27643 ( .A(n27806), .B(n27817), .Z(n27808) );
  XNOR U27644 ( .A(n27819), .B(n27820), .Z(n791) );
  AND U27645 ( .A(n27821), .B(n27822), .Z(n27820) );
  XNOR U27646 ( .A(n27823), .B(n27819), .Z(n27822) );
  IV U27647 ( .A(n27709), .Z(n27823) );
  XNOR U27648 ( .A(n27824), .B(n27825), .Z(n27709) );
  AND U27649 ( .A(n794), .B(n27826), .Z(n27825) );
  XNOR U27650 ( .A(n27824), .B(n27827), .Z(n27826) );
  XNOR U27651 ( .A(n27663), .B(n27819), .Z(n27821) );
  XOR U27652 ( .A(n27828), .B(n27829), .Z(n27663) );
  AND U27653 ( .A(n802), .B(n27830), .Z(n27829) );
  XOR U27654 ( .A(n27813), .B(n27831), .Z(n27819) );
  AND U27655 ( .A(n27832), .B(n27816), .Z(n27831) );
  XNOR U27656 ( .A(n27722), .B(n27813), .Z(n27816) );
  XNOR U27657 ( .A(n27833), .B(n27834), .Z(n27722) );
  AND U27658 ( .A(n794), .B(n27835), .Z(n27834) );
  XOR U27659 ( .A(n27836), .B(n27833), .Z(n27835) );
  XNOR U27660 ( .A(n27837), .B(n27813), .Z(n27832) );
  IV U27661 ( .A(n27673), .Z(n27837) );
  XOR U27662 ( .A(n27838), .B(n27839), .Z(n27673) );
  AND U27663 ( .A(n802), .B(n27840), .Z(n27839) );
  XOR U27664 ( .A(n27841), .B(n27842), .Z(n27813) );
  AND U27665 ( .A(n27843), .B(n27844), .Z(n27842) );
  XNOR U27666 ( .A(n27747), .B(n27841), .Z(n27844) );
  XNOR U27667 ( .A(n27845), .B(n27846), .Z(n27747) );
  AND U27668 ( .A(n794), .B(n27847), .Z(n27846) );
  XNOR U27669 ( .A(n27848), .B(n27845), .Z(n27847) );
  XOR U27670 ( .A(n27841), .B(n27684), .Z(n27843) );
  XOR U27671 ( .A(n27849), .B(n27850), .Z(n27684) );
  AND U27672 ( .A(n802), .B(n27851), .Z(n27850) );
  XOR U27673 ( .A(n27852), .B(n27853), .Z(n27841) );
  AND U27674 ( .A(n27854), .B(n27855), .Z(n27853) );
  XNOR U27675 ( .A(n27852), .B(n27795), .Z(n27855) );
  XNOR U27676 ( .A(n27856), .B(n27857), .Z(n27795) );
  AND U27677 ( .A(n794), .B(n27858), .Z(n27857) );
  XOR U27678 ( .A(n27859), .B(n27856), .Z(n27858) );
  XNOR U27679 ( .A(n27860), .B(n27852), .Z(n27854) );
  IV U27680 ( .A(n27696), .Z(n27860) );
  XOR U27681 ( .A(n27861), .B(n27862), .Z(n27696) );
  AND U27682 ( .A(n802), .B(n27863), .Z(n27862) );
  AND U27683 ( .A(n27817), .B(n27806), .Z(n27852) );
  XNOR U27684 ( .A(n27864), .B(n27865), .Z(n27806) );
  AND U27685 ( .A(n794), .B(n27866), .Z(n27865) );
  XNOR U27686 ( .A(n27867), .B(n27864), .Z(n27866) );
  XNOR U27687 ( .A(n27868), .B(n27869), .Z(n794) );
  AND U27688 ( .A(n27870), .B(n27871), .Z(n27869) );
  XOR U27689 ( .A(n27827), .B(n27868), .Z(n27871) );
  AND U27690 ( .A(n27872), .B(n27873), .Z(n27827) );
  XOR U27691 ( .A(n27868), .B(n27824), .Z(n27870) );
  XNOR U27692 ( .A(n27874), .B(n27875), .Z(n27824) );
  AND U27693 ( .A(n798), .B(n27830), .Z(n27875) );
  XOR U27694 ( .A(n27828), .B(n27874), .Z(n27830) );
  XOR U27695 ( .A(n27876), .B(n27877), .Z(n27868) );
  AND U27696 ( .A(n27878), .B(n27879), .Z(n27877) );
  XNOR U27697 ( .A(n27876), .B(n27872), .Z(n27879) );
  IV U27698 ( .A(n27836), .Z(n27872) );
  XOR U27699 ( .A(n27880), .B(n27881), .Z(n27836) );
  XOR U27700 ( .A(n27882), .B(n27873), .Z(n27881) );
  AND U27701 ( .A(n27848), .B(n27883), .Z(n27873) );
  AND U27702 ( .A(n27884), .B(n27885), .Z(n27882) );
  XOR U27703 ( .A(n27886), .B(n27880), .Z(n27884) );
  XNOR U27704 ( .A(n27833), .B(n27876), .Z(n27878) );
  XNOR U27705 ( .A(n27887), .B(n27888), .Z(n27833) );
  AND U27706 ( .A(n798), .B(n27840), .Z(n27888) );
  XOR U27707 ( .A(n27887), .B(n27838), .Z(n27840) );
  XOR U27708 ( .A(n27889), .B(n27890), .Z(n27876) );
  AND U27709 ( .A(n27891), .B(n27892), .Z(n27890) );
  XNOR U27710 ( .A(n27889), .B(n27848), .Z(n27892) );
  XOR U27711 ( .A(n27893), .B(n27885), .Z(n27848) );
  XNOR U27712 ( .A(n27894), .B(n27880), .Z(n27885) );
  XOR U27713 ( .A(n27895), .B(n27896), .Z(n27880) );
  AND U27714 ( .A(n27897), .B(n27898), .Z(n27896) );
  XOR U27715 ( .A(n27899), .B(n27895), .Z(n27897) );
  XNOR U27716 ( .A(n27900), .B(n27901), .Z(n27894) );
  AND U27717 ( .A(n27902), .B(n27903), .Z(n27901) );
  XOR U27718 ( .A(n27900), .B(n27904), .Z(n27902) );
  XNOR U27719 ( .A(n27886), .B(n27883), .Z(n27893) );
  AND U27720 ( .A(n27905), .B(n27906), .Z(n27883) );
  XOR U27721 ( .A(n27907), .B(n27908), .Z(n27886) );
  AND U27722 ( .A(n27909), .B(n27910), .Z(n27908) );
  XOR U27723 ( .A(n27907), .B(n27911), .Z(n27909) );
  XNOR U27724 ( .A(n27845), .B(n27889), .Z(n27891) );
  XNOR U27725 ( .A(n27912), .B(n27913), .Z(n27845) );
  AND U27726 ( .A(n798), .B(n27851), .Z(n27913) );
  XOR U27727 ( .A(n27912), .B(n27849), .Z(n27851) );
  XOR U27728 ( .A(n27914), .B(n27915), .Z(n27889) );
  AND U27729 ( .A(n27916), .B(n27917), .Z(n27915) );
  XNOR U27730 ( .A(n27914), .B(n27905), .Z(n27917) );
  IV U27731 ( .A(n27859), .Z(n27905) );
  XNOR U27732 ( .A(n27918), .B(n27898), .Z(n27859) );
  XNOR U27733 ( .A(n27919), .B(n27904), .Z(n27898) );
  XNOR U27734 ( .A(n27920), .B(n27921), .Z(n27904) );
  NOR U27735 ( .A(n27922), .B(n27923), .Z(n27921) );
  XOR U27736 ( .A(n27920), .B(n27924), .Z(n27922) );
  XNOR U27737 ( .A(n27903), .B(n27895), .Z(n27919) );
  XOR U27738 ( .A(n27925), .B(n27926), .Z(n27895) );
  AND U27739 ( .A(n27927), .B(n27928), .Z(n27926) );
  XOR U27740 ( .A(n27925), .B(n27929), .Z(n27927) );
  XNOR U27741 ( .A(n27930), .B(n27900), .Z(n27903) );
  XOR U27742 ( .A(n27931), .B(n27932), .Z(n27900) );
  AND U27743 ( .A(n27933), .B(n27934), .Z(n27932) );
  XNOR U27744 ( .A(n27935), .B(n27936), .Z(n27933) );
  IV U27745 ( .A(n27931), .Z(n27935) );
  XNOR U27746 ( .A(n27937), .B(n27938), .Z(n27930) );
  NOR U27747 ( .A(n27939), .B(n27940), .Z(n27938) );
  XNOR U27748 ( .A(n27937), .B(n27941), .Z(n27939) );
  XNOR U27749 ( .A(n27899), .B(n27906), .Z(n27918) );
  NOR U27750 ( .A(n27867), .B(n27942), .Z(n27906) );
  XOR U27751 ( .A(n27911), .B(n27910), .Z(n27899) );
  XNOR U27752 ( .A(n27943), .B(n27907), .Z(n27910) );
  XOR U27753 ( .A(n27944), .B(n27945), .Z(n27907) );
  AND U27754 ( .A(n27946), .B(n27947), .Z(n27945) );
  XNOR U27755 ( .A(n27948), .B(n27949), .Z(n27946) );
  IV U27756 ( .A(n27944), .Z(n27948) );
  XNOR U27757 ( .A(n27950), .B(n27951), .Z(n27943) );
  NOR U27758 ( .A(n27952), .B(n27953), .Z(n27951) );
  XNOR U27759 ( .A(n27950), .B(n27954), .Z(n27952) );
  XOR U27760 ( .A(n27955), .B(n27956), .Z(n27911) );
  NOR U27761 ( .A(n27957), .B(n27958), .Z(n27956) );
  XNOR U27762 ( .A(n27955), .B(n27959), .Z(n27957) );
  XNOR U27763 ( .A(n27856), .B(n27914), .Z(n27916) );
  XNOR U27764 ( .A(n27960), .B(n27961), .Z(n27856) );
  AND U27765 ( .A(n798), .B(n27863), .Z(n27961) );
  XOR U27766 ( .A(n27960), .B(n27861), .Z(n27863) );
  AND U27767 ( .A(n27864), .B(n27867), .Z(n27914) );
  XOR U27768 ( .A(n27962), .B(n27942), .Z(n27867) );
  XNOR U27769 ( .A(p_input[1104]), .B(p_input[2048]), .Z(n27942) );
  XNOR U27770 ( .A(n27929), .B(n27928), .Z(n27962) );
  XNOR U27771 ( .A(n27963), .B(n27936), .Z(n27928) );
  XNOR U27772 ( .A(n27924), .B(n27923), .Z(n27936) );
  XNOR U27773 ( .A(n27964), .B(n27920), .Z(n27923) );
  XNOR U27774 ( .A(p_input[1114]), .B(p_input[2058]), .Z(n27920) );
  XOR U27775 ( .A(p_input[1115]), .B(n16732), .Z(n27964) );
  XOR U27776 ( .A(p_input[1116]), .B(p_input[2060]), .Z(n27924) );
  XOR U27777 ( .A(n27934), .B(n27965), .Z(n27963) );
  IV U27778 ( .A(n27925), .Z(n27965) );
  XOR U27779 ( .A(p_input[1105]), .B(p_input[2049]), .Z(n27925) );
  XNOR U27780 ( .A(n27966), .B(n27941), .Z(n27934) );
  XNOR U27781 ( .A(p_input[1119]), .B(n16735), .Z(n27941) );
  XOR U27782 ( .A(n27931), .B(n27940), .Z(n27966) );
  XOR U27783 ( .A(n27967), .B(n27937), .Z(n27940) );
  XOR U27784 ( .A(p_input[1117]), .B(p_input[2061]), .Z(n27937) );
  XOR U27785 ( .A(p_input[1118]), .B(n16737), .Z(n27967) );
  XOR U27786 ( .A(p_input[1113]), .B(p_input[2057]), .Z(n27931) );
  XOR U27787 ( .A(n27949), .B(n27947), .Z(n27929) );
  XNOR U27788 ( .A(n27968), .B(n27954), .Z(n27947) );
  XOR U27789 ( .A(p_input[1112]), .B(p_input[2056]), .Z(n27954) );
  XOR U27790 ( .A(n27944), .B(n27953), .Z(n27968) );
  XOR U27791 ( .A(n27969), .B(n27950), .Z(n27953) );
  XOR U27792 ( .A(p_input[1110]), .B(p_input[2054]), .Z(n27950) );
  XOR U27793 ( .A(p_input[1111]), .B(n17722), .Z(n27969) );
  XOR U27794 ( .A(p_input[1106]), .B(p_input[2050]), .Z(n27944) );
  XNOR U27795 ( .A(n27959), .B(n27958), .Z(n27949) );
  XOR U27796 ( .A(n27970), .B(n27955), .Z(n27958) );
  XOR U27797 ( .A(p_input[1107]), .B(p_input[2051]), .Z(n27955) );
  XOR U27798 ( .A(p_input[1108]), .B(n17724), .Z(n27970) );
  XOR U27799 ( .A(p_input[1109]), .B(p_input[2053]), .Z(n27959) );
  XNOR U27800 ( .A(n27971), .B(n27972), .Z(n27864) );
  AND U27801 ( .A(n798), .B(n27973), .Z(n27972) );
  XNOR U27802 ( .A(n27974), .B(n27975), .Z(n798) );
  AND U27803 ( .A(n27976), .B(n27977), .Z(n27975) );
  XOR U27804 ( .A(n27974), .B(n27874), .Z(n27977) );
  XNOR U27805 ( .A(n27974), .B(n27828), .Z(n27976) );
  XOR U27806 ( .A(n27978), .B(n27979), .Z(n27974) );
  AND U27807 ( .A(n27980), .B(n27981), .Z(n27979) );
  XOR U27808 ( .A(n27978), .B(n27838), .Z(n27980) );
  XOR U27809 ( .A(n27982), .B(n27983), .Z(n27817) );
  AND U27810 ( .A(n802), .B(n27973), .Z(n27983) );
  XNOR U27811 ( .A(n27971), .B(n27982), .Z(n27973) );
  XNOR U27812 ( .A(n27984), .B(n27985), .Z(n802) );
  AND U27813 ( .A(n27986), .B(n27987), .Z(n27985) );
  XNOR U27814 ( .A(n27988), .B(n27984), .Z(n27987) );
  IV U27815 ( .A(n27874), .Z(n27988) );
  XNOR U27816 ( .A(n27989), .B(n27990), .Z(n27874) );
  AND U27817 ( .A(n805), .B(n27991), .Z(n27990) );
  XNOR U27818 ( .A(n27989), .B(n27992), .Z(n27991) );
  XNOR U27819 ( .A(n27828), .B(n27984), .Z(n27986) );
  XOR U27820 ( .A(n27993), .B(n27994), .Z(n27828) );
  AND U27821 ( .A(n813), .B(n27995), .Z(n27994) );
  XOR U27822 ( .A(n27978), .B(n27996), .Z(n27984) );
  AND U27823 ( .A(n27997), .B(n27981), .Z(n27996) );
  XNOR U27824 ( .A(n27887), .B(n27978), .Z(n27981) );
  XNOR U27825 ( .A(n27998), .B(n27999), .Z(n27887) );
  AND U27826 ( .A(n805), .B(n28000), .Z(n27999) );
  XOR U27827 ( .A(n28001), .B(n27998), .Z(n28000) );
  XNOR U27828 ( .A(n28002), .B(n27978), .Z(n27997) );
  IV U27829 ( .A(n27838), .Z(n28002) );
  XOR U27830 ( .A(n28003), .B(n28004), .Z(n27838) );
  AND U27831 ( .A(n813), .B(n28005), .Z(n28004) );
  XOR U27832 ( .A(n28006), .B(n28007), .Z(n27978) );
  AND U27833 ( .A(n28008), .B(n28009), .Z(n28007) );
  XNOR U27834 ( .A(n27912), .B(n28006), .Z(n28009) );
  XNOR U27835 ( .A(n28010), .B(n28011), .Z(n27912) );
  AND U27836 ( .A(n805), .B(n28012), .Z(n28011) );
  XNOR U27837 ( .A(n28013), .B(n28010), .Z(n28012) );
  XOR U27838 ( .A(n28006), .B(n27849), .Z(n28008) );
  XOR U27839 ( .A(n28014), .B(n28015), .Z(n27849) );
  AND U27840 ( .A(n813), .B(n28016), .Z(n28015) );
  XOR U27841 ( .A(n28017), .B(n28018), .Z(n28006) );
  AND U27842 ( .A(n28019), .B(n28020), .Z(n28018) );
  XNOR U27843 ( .A(n28017), .B(n27960), .Z(n28020) );
  XNOR U27844 ( .A(n28021), .B(n28022), .Z(n27960) );
  AND U27845 ( .A(n805), .B(n28023), .Z(n28022) );
  XOR U27846 ( .A(n28024), .B(n28021), .Z(n28023) );
  XNOR U27847 ( .A(n28025), .B(n28017), .Z(n28019) );
  IV U27848 ( .A(n27861), .Z(n28025) );
  XOR U27849 ( .A(n28026), .B(n28027), .Z(n27861) );
  AND U27850 ( .A(n813), .B(n28028), .Z(n28027) );
  AND U27851 ( .A(n27982), .B(n27971), .Z(n28017) );
  XNOR U27852 ( .A(n28029), .B(n28030), .Z(n27971) );
  AND U27853 ( .A(n805), .B(n28031), .Z(n28030) );
  XNOR U27854 ( .A(n28032), .B(n28029), .Z(n28031) );
  XNOR U27855 ( .A(n28033), .B(n28034), .Z(n805) );
  AND U27856 ( .A(n28035), .B(n28036), .Z(n28034) );
  XOR U27857 ( .A(n27992), .B(n28033), .Z(n28036) );
  AND U27858 ( .A(n28037), .B(n28038), .Z(n27992) );
  XOR U27859 ( .A(n28033), .B(n27989), .Z(n28035) );
  XNOR U27860 ( .A(n28039), .B(n28040), .Z(n27989) );
  AND U27861 ( .A(n809), .B(n27995), .Z(n28040) );
  XOR U27862 ( .A(n27993), .B(n28039), .Z(n27995) );
  XOR U27863 ( .A(n28041), .B(n28042), .Z(n28033) );
  AND U27864 ( .A(n28043), .B(n28044), .Z(n28042) );
  XNOR U27865 ( .A(n28041), .B(n28037), .Z(n28044) );
  IV U27866 ( .A(n28001), .Z(n28037) );
  XOR U27867 ( .A(n28045), .B(n28046), .Z(n28001) );
  XOR U27868 ( .A(n28047), .B(n28038), .Z(n28046) );
  AND U27869 ( .A(n28013), .B(n28048), .Z(n28038) );
  AND U27870 ( .A(n28049), .B(n28050), .Z(n28047) );
  XOR U27871 ( .A(n28051), .B(n28045), .Z(n28049) );
  XNOR U27872 ( .A(n27998), .B(n28041), .Z(n28043) );
  XNOR U27873 ( .A(n28052), .B(n28053), .Z(n27998) );
  AND U27874 ( .A(n809), .B(n28005), .Z(n28053) );
  XOR U27875 ( .A(n28052), .B(n28003), .Z(n28005) );
  XOR U27876 ( .A(n28054), .B(n28055), .Z(n28041) );
  AND U27877 ( .A(n28056), .B(n28057), .Z(n28055) );
  XNOR U27878 ( .A(n28054), .B(n28013), .Z(n28057) );
  XOR U27879 ( .A(n28058), .B(n28050), .Z(n28013) );
  XNOR U27880 ( .A(n28059), .B(n28045), .Z(n28050) );
  XOR U27881 ( .A(n28060), .B(n28061), .Z(n28045) );
  AND U27882 ( .A(n28062), .B(n28063), .Z(n28061) );
  XOR U27883 ( .A(n28064), .B(n28060), .Z(n28062) );
  XNOR U27884 ( .A(n28065), .B(n28066), .Z(n28059) );
  AND U27885 ( .A(n28067), .B(n28068), .Z(n28066) );
  XOR U27886 ( .A(n28065), .B(n28069), .Z(n28067) );
  XNOR U27887 ( .A(n28051), .B(n28048), .Z(n28058) );
  AND U27888 ( .A(n28070), .B(n28071), .Z(n28048) );
  XOR U27889 ( .A(n28072), .B(n28073), .Z(n28051) );
  AND U27890 ( .A(n28074), .B(n28075), .Z(n28073) );
  XOR U27891 ( .A(n28072), .B(n28076), .Z(n28074) );
  XNOR U27892 ( .A(n28010), .B(n28054), .Z(n28056) );
  XNOR U27893 ( .A(n28077), .B(n28078), .Z(n28010) );
  AND U27894 ( .A(n809), .B(n28016), .Z(n28078) );
  XOR U27895 ( .A(n28077), .B(n28014), .Z(n28016) );
  XOR U27896 ( .A(n28079), .B(n28080), .Z(n28054) );
  AND U27897 ( .A(n28081), .B(n28082), .Z(n28080) );
  XNOR U27898 ( .A(n28079), .B(n28070), .Z(n28082) );
  IV U27899 ( .A(n28024), .Z(n28070) );
  XNOR U27900 ( .A(n28083), .B(n28063), .Z(n28024) );
  XNOR U27901 ( .A(n28084), .B(n28069), .Z(n28063) );
  XNOR U27902 ( .A(n28085), .B(n28086), .Z(n28069) );
  NOR U27903 ( .A(n28087), .B(n28088), .Z(n28086) );
  XOR U27904 ( .A(n28085), .B(n28089), .Z(n28087) );
  XNOR U27905 ( .A(n28068), .B(n28060), .Z(n28084) );
  XOR U27906 ( .A(n28090), .B(n28091), .Z(n28060) );
  AND U27907 ( .A(n28092), .B(n28093), .Z(n28091) );
  XOR U27908 ( .A(n28090), .B(n28094), .Z(n28092) );
  XNOR U27909 ( .A(n28095), .B(n28065), .Z(n28068) );
  XOR U27910 ( .A(n28096), .B(n28097), .Z(n28065) );
  AND U27911 ( .A(n28098), .B(n28099), .Z(n28097) );
  XNOR U27912 ( .A(n28100), .B(n28101), .Z(n28098) );
  IV U27913 ( .A(n28096), .Z(n28100) );
  XNOR U27914 ( .A(n28102), .B(n28103), .Z(n28095) );
  NOR U27915 ( .A(n28104), .B(n28105), .Z(n28103) );
  XNOR U27916 ( .A(n28102), .B(n28106), .Z(n28104) );
  XNOR U27917 ( .A(n28064), .B(n28071), .Z(n28083) );
  NOR U27918 ( .A(n28032), .B(n28107), .Z(n28071) );
  XOR U27919 ( .A(n28076), .B(n28075), .Z(n28064) );
  XNOR U27920 ( .A(n28108), .B(n28072), .Z(n28075) );
  XOR U27921 ( .A(n28109), .B(n28110), .Z(n28072) );
  AND U27922 ( .A(n28111), .B(n28112), .Z(n28110) );
  XNOR U27923 ( .A(n28113), .B(n28114), .Z(n28111) );
  IV U27924 ( .A(n28109), .Z(n28113) );
  XNOR U27925 ( .A(n28115), .B(n28116), .Z(n28108) );
  NOR U27926 ( .A(n28117), .B(n28118), .Z(n28116) );
  XNOR U27927 ( .A(n28115), .B(n28119), .Z(n28117) );
  XOR U27928 ( .A(n28120), .B(n28121), .Z(n28076) );
  NOR U27929 ( .A(n28122), .B(n28123), .Z(n28121) );
  XNOR U27930 ( .A(n28120), .B(n28124), .Z(n28122) );
  XNOR U27931 ( .A(n28021), .B(n28079), .Z(n28081) );
  XNOR U27932 ( .A(n28125), .B(n28126), .Z(n28021) );
  AND U27933 ( .A(n809), .B(n28028), .Z(n28126) );
  XOR U27934 ( .A(n28125), .B(n28026), .Z(n28028) );
  AND U27935 ( .A(n28029), .B(n28032), .Z(n28079) );
  XOR U27936 ( .A(n28127), .B(n28107), .Z(n28032) );
  XNOR U27937 ( .A(p_input[1120]), .B(p_input[2048]), .Z(n28107) );
  XNOR U27938 ( .A(n28094), .B(n28093), .Z(n28127) );
  XNOR U27939 ( .A(n28128), .B(n28101), .Z(n28093) );
  XNOR U27940 ( .A(n28089), .B(n28088), .Z(n28101) );
  XNOR U27941 ( .A(n28129), .B(n28085), .Z(n28088) );
  XNOR U27942 ( .A(p_input[1130]), .B(p_input[2058]), .Z(n28085) );
  XOR U27943 ( .A(p_input[1131]), .B(n16732), .Z(n28129) );
  XOR U27944 ( .A(p_input[1132]), .B(p_input[2060]), .Z(n28089) );
  XOR U27945 ( .A(n28099), .B(n28130), .Z(n28128) );
  IV U27946 ( .A(n28090), .Z(n28130) );
  XOR U27947 ( .A(p_input[1121]), .B(p_input[2049]), .Z(n28090) );
  XNOR U27948 ( .A(n28131), .B(n28106), .Z(n28099) );
  XNOR U27949 ( .A(p_input[1135]), .B(n16735), .Z(n28106) );
  XOR U27950 ( .A(n28096), .B(n28105), .Z(n28131) );
  XOR U27951 ( .A(n28132), .B(n28102), .Z(n28105) );
  XOR U27952 ( .A(p_input[1133]), .B(p_input[2061]), .Z(n28102) );
  XOR U27953 ( .A(p_input[1134]), .B(n16737), .Z(n28132) );
  XOR U27954 ( .A(p_input[1129]), .B(p_input[2057]), .Z(n28096) );
  XOR U27955 ( .A(n28114), .B(n28112), .Z(n28094) );
  XNOR U27956 ( .A(n28133), .B(n28119), .Z(n28112) );
  XOR U27957 ( .A(p_input[1128]), .B(p_input[2056]), .Z(n28119) );
  XOR U27958 ( .A(n28109), .B(n28118), .Z(n28133) );
  XOR U27959 ( .A(n28134), .B(n28115), .Z(n28118) );
  XOR U27960 ( .A(p_input[1126]), .B(p_input[2054]), .Z(n28115) );
  XOR U27961 ( .A(p_input[1127]), .B(n17722), .Z(n28134) );
  XOR U27962 ( .A(p_input[1122]), .B(p_input[2050]), .Z(n28109) );
  XNOR U27963 ( .A(n28124), .B(n28123), .Z(n28114) );
  XOR U27964 ( .A(n28135), .B(n28120), .Z(n28123) );
  XOR U27965 ( .A(p_input[1123]), .B(p_input[2051]), .Z(n28120) );
  XOR U27966 ( .A(p_input[1124]), .B(n17724), .Z(n28135) );
  XOR U27967 ( .A(p_input[1125]), .B(p_input[2053]), .Z(n28124) );
  XNOR U27968 ( .A(n28136), .B(n28137), .Z(n28029) );
  AND U27969 ( .A(n809), .B(n28138), .Z(n28137) );
  XNOR U27970 ( .A(n28139), .B(n28140), .Z(n809) );
  AND U27971 ( .A(n28141), .B(n28142), .Z(n28140) );
  XOR U27972 ( .A(n28139), .B(n28039), .Z(n28142) );
  XNOR U27973 ( .A(n28139), .B(n27993), .Z(n28141) );
  XOR U27974 ( .A(n28143), .B(n28144), .Z(n28139) );
  AND U27975 ( .A(n28145), .B(n28146), .Z(n28144) );
  XOR U27976 ( .A(n28143), .B(n28003), .Z(n28145) );
  XOR U27977 ( .A(n28147), .B(n28148), .Z(n27982) );
  AND U27978 ( .A(n813), .B(n28138), .Z(n28148) );
  XNOR U27979 ( .A(n28136), .B(n28147), .Z(n28138) );
  XNOR U27980 ( .A(n28149), .B(n28150), .Z(n813) );
  AND U27981 ( .A(n28151), .B(n28152), .Z(n28150) );
  XNOR U27982 ( .A(n28153), .B(n28149), .Z(n28152) );
  IV U27983 ( .A(n28039), .Z(n28153) );
  XNOR U27984 ( .A(n28154), .B(n28155), .Z(n28039) );
  AND U27985 ( .A(n816), .B(n28156), .Z(n28155) );
  XNOR U27986 ( .A(n28154), .B(n28157), .Z(n28156) );
  XNOR U27987 ( .A(n27993), .B(n28149), .Z(n28151) );
  XOR U27988 ( .A(n28158), .B(n28159), .Z(n27993) );
  AND U27989 ( .A(n824), .B(n28160), .Z(n28159) );
  XOR U27990 ( .A(n28143), .B(n28161), .Z(n28149) );
  AND U27991 ( .A(n28162), .B(n28146), .Z(n28161) );
  XNOR U27992 ( .A(n28052), .B(n28143), .Z(n28146) );
  XNOR U27993 ( .A(n28163), .B(n28164), .Z(n28052) );
  AND U27994 ( .A(n816), .B(n28165), .Z(n28164) );
  XOR U27995 ( .A(n28166), .B(n28163), .Z(n28165) );
  XNOR U27996 ( .A(n28167), .B(n28143), .Z(n28162) );
  IV U27997 ( .A(n28003), .Z(n28167) );
  XOR U27998 ( .A(n28168), .B(n28169), .Z(n28003) );
  AND U27999 ( .A(n824), .B(n28170), .Z(n28169) );
  XOR U28000 ( .A(n28171), .B(n28172), .Z(n28143) );
  AND U28001 ( .A(n28173), .B(n28174), .Z(n28172) );
  XNOR U28002 ( .A(n28077), .B(n28171), .Z(n28174) );
  XNOR U28003 ( .A(n28175), .B(n28176), .Z(n28077) );
  AND U28004 ( .A(n816), .B(n28177), .Z(n28176) );
  XNOR U28005 ( .A(n28178), .B(n28175), .Z(n28177) );
  XOR U28006 ( .A(n28171), .B(n28014), .Z(n28173) );
  XOR U28007 ( .A(n28179), .B(n28180), .Z(n28014) );
  AND U28008 ( .A(n824), .B(n28181), .Z(n28180) );
  XOR U28009 ( .A(n28182), .B(n28183), .Z(n28171) );
  AND U28010 ( .A(n28184), .B(n28185), .Z(n28183) );
  XNOR U28011 ( .A(n28182), .B(n28125), .Z(n28185) );
  XNOR U28012 ( .A(n28186), .B(n28187), .Z(n28125) );
  AND U28013 ( .A(n816), .B(n28188), .Z(n28187) );
  XOR U28014 ( .A(n28189), .B(n28186), .Z(n28188) );
  XNOR U28015 ( .A(n28190), .B(n28182), .Z(n28184) );
  IV U28016 ( .A(n28026), .Z(n28190) );
  XOR U28017 ( .A(n28191), .B(n28192), .Z(n28026) );
  AND U28018 ( .A(n824), .B(n28193), .Z(n28192) );
  AND U28019 ( .A(n28147), .B(n28136), .Z(n28182) );
  XNOR U28020 ( .A(n28194), .B(n28195), .Z(n28136) );
  AND U28021 ( .A(n816), .B(n28196), .Z(n28195) );
  XNOR U28022 ( .A(n28197), .B(n28194), .Z(n28196) );
  XNOR U28023 ( .A(n28198), .B(n28199), .Z(n816) );
  AND U28024 ( .A(n28200), .B(n28201), .Z(n28199) );
  XOR U28025 ( .A(n28157), .B(n28198), .Z(n28201) );
  AND U28026 ( .A(n28202), .B(n28203), .Z(n28157) );
  XOR U28027 ( .A(n28198), .B(n28154), .Z(n28200) );
  XNOR U28028 ( .A(n28204), .B(n28205), .Z(n28154) );
  AND U28029 ( .A(n820), .B(n28160), .Z(n28205) );
  XOR U28030 ( .A(n28158), .B(n28204), .Z(n28160) );
  XOR U28031 ( .A(n28206), .B(n28207), .Z(n28198) );
  AND U28032 ( .A(n28208), .B(n28209), .Z(n28207) );
  XNOR U28033 ( .A(n28206), .B(n28202), .Z(n28209) );
  IV U28034 ( .A(n28166), .Z(n28202) );
  XOR U28035 ( .A(n28210), .B(n28211), .Z(n28166) );
  XOR U28036 ( .A(n28212), .B(n28203), .Z(n28211) );
  AND U28037 ( .A(n28178), .B(n28213), .Z(n28203) );
  AND U28038 ( .A(n28214), .B(n28215), .Z(n28212) );
  XOR U28039 ( .A(n28216), .B(n28210), .Z(n28214) );
  XNOR U28040 ( .A(n28163), .B(n28206), .Z(n28208) );
  XNOR U28041 ( .A(n28217), .B(n28218), .Z(n28163) );
  AND U28042 ( .A(n820), .B(n28170), .Z(n28218) );
  XOR U28043 ( .A(n28217), .B(n28168), .Z(n28170) );
  XOR U28044 ( .A(n28219), .B(n28220), .Z(n28206) );
  AND U28045 ( .A(n28221), .B(n28222), .Z(n28220) );
  XNOR U28046 ( .A(n28219), .B(n28178), .Z(n28222) );
  XOR U28047 ( .A(n28223), .B(n28215), .Z(n28178) );
  XNOR U28048 ( .A(n28224), .B(n28210), .Z(n28215) );
  XOR U28049 ( .A(n28225), .B(n28226), .Z(n28210) );
  AND U28050 ( .A(n28227), .B(n28228), .Z(n28226) );
  XOR U28051 ( .A(n28229), .B(n28225), .Z(n28227) );
  XNOR U28052 ( .A(n28230), .B(n28231), .Z(n28224) );
  AND U28053 ( .A(n28232), .B(n28233), .Z(n28231) );
  XOR U28054 ( .A(n28230), .B(n28234), .Z(n28232) );
  XNOR U28055 ( .A(n28216), .B(n28213), .Z(n28223) );
  AND U28056 ( .A(n28235), .B(n28236), .Z(n28213) );
  XOR U28057 ( .A(n28237), .B(n28238), .Z(n28216) );
  AND U28058 ( .A(n28239), .B(n28240), .Z(n28238) );
  XOR U28059 ( .A(n28237), .B(n28241), .Z(n28239) );
  XNOR U28060 ( .A(n28175), .B(n28219), .Z(n28221) );
  XNOR U28061 ( .A(n28242), .B(n28243), .Z(n28175) );
  AND U28062 ( .A(n820), .B(n28181), .Z(n28243) );
  XOR U28063 ( .A(n28242), .B(n28179), .Z(n28181) );
  XOR U28064 ( .A(n28244), .B(n28245), .Z(n28219) );
  AND U28065 ( .A(n28246), .B(n28247), .Z(n28245) );
  XNOR U28066 ( .A(n28244), .B(n28235), .Z(n28247) );
  IV U28067 ( .A(n28189), .Z(n28235) );
  XNOR U28068 ( .A(n28248), .B(n28228), .Z(n28189) );
  XNOR U28069 ( .A(n28249), .B(n28234), .Z(n28228) );
  XNOR U28070 ( .A(n28250), .B(n28251), .Z(n28234) );
  NOR U28071 ( .A(n28252), .B(n28253), .Z(n28251) );
  XOR U28072 ( .A(n28250), .B(n28254), .Z(n28252) );
  XNOR U28073 ( .A(n28233), .B(n28225), .Z(n28249) );
  XOR U28074 ( .A(n28255), .B(n28256), .Z(n28225) );
  AND U28075 ( .A(n28257), .B(n28258), .Z(n28256) );
  XOR U28076 ( .A(n28255), .B(n28259), .Z(n28257) );
  XNOR U28077 ( .A(n28260), .B(n28230), .Z(n28233) );
  XOR U28078 ( .A(n28261), .B(n28262), .Z(n28230) );
  AND U28079 ( .A(n28263), .B(n28264), .Z(n28262) );
  XNOR U28080 ( .A(n28265), .B(n28266), .Z(n28263) );
  IV U28081 ( .A(n28261), .Z(n28265) );
  XNOR U28082 ( .A(n28267), .B(n28268), .Z(n28260) );
  NOR U28083 ( .A(n28269), .B(n28270), .Z(n28268) );
  XNOR U28084 ( .A(n28267), .B(n28271), .Z(n28269) );
  XNOR U28085 ( .A(n28229), .B(n28236), .Z(n28248) );
  NOR U28086 ( .A(n28197), .B(n28272), .Z(n28236) );
  XOR U28087 ( .A(n28241), .B(n28240), .Z(n28229) );
  XNOR U28088 ( .A(n28273), .B(n28237), .Z(n28240) );
  XOR U28089 ( .A(n28274), .B(n28275), .Z(n28237) );
  AND U28090 ( .A(n28276), .B(n28277), .Z(n28275) );
  XNOR U28091 ( .A(n28278), .B(n28279), .Z(n28276) );
  IV U28092 ( .A(n28274), .Z(n28278) );
  XNOR U28093 ( .A(n28280), .B(n28281), .Z(n28273) );
  NOR U28094 ( .A(n28282), .B(n28283), .Z(n28281) );
  XNOR U28095 ( .A(n28280), .B(n28284), .Z(n28282) );
  XOR U28096 ( .A(n28285), .B(n28286), .Z(n28241) );
  NOR U28097 ( .A(n28287), .B(n28288), .Z(n28286) );
  XNOR U28098 ( .A(n28285), .B(n28289), .Z(n28287) );
  XNOR U28099 ( .A(n28186), .B(n28244), .Z(n28246) );
  XNOR U28100 ( .A(n28290), .B(n28291), .Z(n28186) );
  AND U28101 ( .A(n820), .B(n28193), .Z(n28291) );
  XOR U28102 ( .A(n28290), .B(n28191), .Z(n28193) );
  AND U28103 ( .A(n28194), .B(n28197), .Z(n28244) );
  XOR U28104 ( .A(n28292), .B(n28272), .Z(n28197) );
  XNOR U28105 ( .A(p_input[1136]), .B(p_input[2048]), .Z(n28272) );
  XNOR U28106 ( .A(n28259), .B(n28258), .Z(n28292) );
  XNOR U28107 ( .A(n28293), .B(n28266), .Z(n28258) );
  XNOR U28108 ( .A(n28254), .B(n28253), .Z(n28266) );
  XNOR U28109 ( .A(n28294), .B(n28250), .Z(n28253) );
  XNOR U28110 ( .A(p_input[1146]), .B(p_input[2058]), .Z(n28250) );
  XOR U28111 ( .A(p_input[1147]), .B(n16732), .Z(n28294) );
  XOR U28112 ( .A(p_input[1148]), .B(p_input[2060]), .Z(n28254) );
  XOR U28113 ( .A(n28264), .B(n28295), .Z(n28293) );
  IV U28114 ( .A(n28255), .Z(n28295) );
  XOR U28115 ( .A(p_input[1137]), .B(p_input[2049]), .Z(n28255) );
  XNOR U28116 ( .A(n28296), .B(n28271), .Z(n28264) );
  XNOR U28117 ( .A(p_input[1151]), .B(n16735), .Z(n28271) );
  XOR U28118 ( .A(n28261), .B(n28270), .Z(n28296) );
  XOR U28119 ( .A(n28297), .B(n28267), .Z(n28270) );
  XOR U28120 ( .A(p_input[1149]), .B(p_input[2061]), .Z(n28267) );
  XOR U28121 ( .A(p_input[1150]), .B(n16737), .Z(n28297) );
  XOR U28122 ( .A(p_input[1145]), .B(p_input[2057]), .Z(n28261) );
  XOR U28123 ( .A(n28279), .B(n28277), .Z(n28259) );
  XNOR U28124 ( .A(n28298), .B(n28284), .Z(n28277) );
  XOR U28125 ( .A(p_input[1144]), .B(p_input[2056]), .Z(n28284) );
  XOR U28126 ( .A(n28274), .B(n28283), .Z(n28298) );
  XOR U28127 ( .A(n28299), .B(n28280), .Z(n28283) );
  XOR U28128 ( .A(p_input[1142]), .B(p_input[2054]), .Z(n28280) );
  XOR U28129 ( .A(p_input[1143]), .B(n17722), .Z(n28299) );
  XOR U28130 ( .A(p_input[1138]), .B(p_input[2050]), .Z(n28274) );
  XNOR U28131 ( .A(n28289), .B(n28288), .Z(n28279) );
  XOR U28132 ( .A(n28300), .B(n28285), .Z(n28288) );
  XOR U28133 ( .A(p_input[1139]), .B(p_input[2051]), .Z(n28285) );
  XOR U28134 ( .A(p_input[1140]), .B(n17724), .Z(n28300) );
  XOR U28135 ( .A(p_input[1141]), .B(p_input[2053]), .Z(n28289) );
  XNOR U28136 ( .A(n28301), .B(n28302), .Z(n28194) );
  AND U28137 ( .A(n820), .B(n28303), .Z(n28302) );
  XNOR U28138 ( .A(n28304), .B(n28305), .Z(n820) );
  AND U28139 ( .A(n28306), .B(n28307), .Z(n28305) );
  XOR U28140 ( .A(n28304), .B(n28204), .Z(n28307) );
  XNOR U28141 ( .A(n28304), .B(n28158), .Z(n28306) );
  XOR U28142 ( .A(n28308), .B(n28309), .Z(n28304) );
  AND U28143 ( .A(n28310), .B(n28311), .Z(n28309) );
  XOR U28144 ( .A(n28308), .B(n28168), .Z(n28310) );
  XOR U28145 ( .A(n28312), .B(n28313), .Z(n28147) );
  AND U28146 ( .A(n824), .B(n28303), .Z(n28313) );
  XNOR U28147 ( .A(n28301), .B(n28312), .Z(n28303) );
  XNOR U28148 ( .A(n28314), .B(n28315), .Z(n824) );
  AND U28149 ( .A(n28316), .B(n28317), .Z(n28315) );
  XNOR U28150 ( .A(n28318), .B(n28314), .Z(n28317) );
  IV U28151 ( .A(n28204), .Z(n28318) );
  XNOR U28152 ( .A(n28319), .B(n28320), .Z(n28204) );
  AND U28153 ( .A(n827), .B(n28321), .Z(n28320) );
  XNOR U28154 ( .A(n28319), .B(n28322), .Z(n28321) );
  XNOR U28155 ( .A(n28158), .B(n28314), .Z(n28316) );
  XOR U28156 ( .A(n28323), .B(n28324), .Z(n28158) );
  AND U28157 ( .A(n835), .B(n28325), .Z(n28324) );
  XOR U28158 ( .A(n28308), .B(n28326), .Z(n28314) );
  AND U28159 ( .A(n28327), .B(n28311), .Z(n28326) );
  XNOR U28160 ( .A(n28217), .B(n28308), .Z(n28311) );
  XNOR U28161 ( .A(n28328), .B(n28329), .Z(n28217) );
  AND U28162 ( .A(n827), .B(n28330), .Z(n28329) );
  XOR U28163 ( .A(n28331), .B(n28328), .Z(n28330) );
  XNOR U28164 ( .A(n28332), .B(n28308), .Z(n28327) );
  IV U28165 ( .A(n28168), .Z(n28332) );
  XOR U28166 ( .A(n28333), .B(n28334), .Z(n28168) );
  AND U28167 ( .A(n835), .B(n28335), .Z(n28334) );
  XOR U28168 ( .A(n28336), .B(n28337), .Z(n28308) );
  AND U28169 ( .A(n28338), .B(n28339), .Z(n28337) );
  XNOR U28170 ( .A(n28242), .B(n28336), .Z(n28339) );
  XNOR U28171 ( .A(n28340), .B(n28341), .Z(n28242) );
  AND U28172 ( .A(n827), .B(n28342), .Z(n28341) );
  XNOR U28173 ( .A(n28343), .B(n28340), .Z(n28342) );
  XOR U28174 ( .A(n28336), .B(n28179), .Z(n28338) );
  XOR U28175 ( .A(n28344), .B(n28345), .Z(n28179) );
  AND U28176 ( .A(n835), .B(n28346), .Z(n28345) );
  XOR U28177 ( .A(n28347), .B(n28348), .Z(n28336) );
  AND U28178 ( .A(n28349), .B(n28350), .Z(n28348) );
  XNOR U28179 ( .A(n28347), .B(n28290), .Z(n28350) );
  XNOR U28180 ( .A(n28351), .B(n28352), .Z(n28290) );
  AND U28181 ( .A(n827), .B(n28353), .Z(n28352) );
  XOR U28182 ( .A(n28354), .B(n28351), .Z(n28353) );
  XNOR U28183 ( .A(n28355), .B(n28347), .Z(n28349) );
  IV U28184 ( .A(n28191), .Z(n28355) );
  XOR U28185 ( .A(n28356), .B(n28357), .Z(n28191) );
  AND U28186 ( .A(n835), .B(n28358), .Z(n28357) );
  AND U28187 ( .A(n28312), .B(n28301), .Z(n28347) );
  XNOR U28188 ( .A(n28359), .B(n28360), .Z(n28301) );
  AND U28189 ( .A(n827), .B(n28361), .Z(n28360) );
  XNOR U28190 ( .A(n28362), .B(n28359), .Z(n28361) );
  XNOR U28191 ( .A(n28363), .B(n28364), .Z(n827) );
  AND U28192 ( .A(n28365), .B(n28366), .Z(n28364) );
  XOR U28193 ( .A(n28322), .B(n28363), .Z(n28366) );
  AND U28194 ( .A(n28367), .B(n28368), .Z(n28322) );
  XOR U28195 ( .A(n28363), .B(n28319), .Z(n28365) );
  XNOR U28196 ( .A(n28369), .B(n28370), .Z(n28319) );
  AND U28197 ( .A(n831), .B(n28325), .Z(n28370) );
  XOR U28198 ( .A(n28323), .B(n28369), .Z(n28325) );
  XOR U28199 ( .A(n28371), .B(n28372), .Z(n28363) );
  AND U28200 ( .A(n28373), .B(n28374), .Z(n28372) );
  XNOR U28201 ( .A(n28371), .B(n28367), .Z(n28374) );
  IV U28202 ( .A(n28331), .Z(n28367) );
  XOR U28203 ( .A(n28375), .B(n28376), .Z(n28331) );
  XOR U28204 ( .A(n28377), .B(n28368), .Z(n28376) );
  AND U28205 ( .A(n28343), .B(n28378), .Z(n28368) );
  AND U28206 ( .A(n28379), .B(n28380), .Z(n28377) );
  XOR U28207 ( .A(n28381), .B(n28375), .Z(n28379) );
  XNOR U28208 ( .A(n28328), .B(n28371), .Z(n28373) );
  XNOR U28209 ( .A(n28382), .B(n28383), .Z(n28328) );
  AND U28210 ( .A(n831), .B(n28335), .Z(n28383) );
  XOR U28211 ( .A(n28382), .B(n28333), .Z(n28335) );
  XOR U28212 ( .A(n28384), .B(n28385), .Z(n28371) );
  AND U28213 ( .A(n28386), .B(n28387), .Z(n28385) );
  XNOR U28214 ( .A(n28384), .B(n28343), .Z(n28387) );
  XOR U28215 ( .A(n28388), .B(n28380), .Z(n28343) );
  XNOR U28216 ( .A(n28389), .B(n28375), .Z(n28380) );
  XOR U28217 ( .A(n28390), .B(n28391), .Z(n28375) );
  AND U28218 ( .A(n28392), .B(n28393), .Z(n28391) );
  XOR U28219 ( .A(n28394), .B(n28390), .Z(n28392) );
  XNOR U28220 ( .A(n28395), .B(n28396), .Z(n28389) );
  AND U28221 ( .A(n28397), .B(n28398), .Z(n28396) );
  XOR U28222 ( .A(n28395), .B(n28399), .Z(n28397) );
  XNOR U28223 ( .A(n28381), .B(n28378), .Z(n28388) );
  AND U28224 ( .A(n28400), .B(n28401), .Z(n28378) );
  XOR U28225 ( .A(n28402), .B(n28403), .Z(n28381) );
  AND U28226 ( .A(n28404), .B(n28405), .Z(n28403) );
  XOR U28227 ( .A(n28402), .B(n28406), .Z(n28404) );
  XNOR U28228 ( .A(n28340), .B(n28384), .Z(n28386) );
  XNOR U28229 ( .A(n28407), .B(n28408), .Z(n28340) );
  AND U28230 ( .A(n831), .B(n28346), .Z(n28408) );
  XOR U28231 ( .A(n28407), .B(n28344), .Z(n28346) );
  XOR U28232 ( .A(n28409), .B(n28410), .Z(n28384) );
  AND U28233 ( .A(n28411), .B(n28412), .Z(n28410) );
  XNOR U28234 ( .A(n28409), .B(n28400), .Z(n28412) );
  IV U28235 ( .A(n28354), .Z(n28400) );
  XNOR U28236 ( .A(n28413), .B(n28393), .Z(n28354) );
  XNOR U28237 ( .A(n28414), .B(n28399), .Z(n28393) );
  XNOR U28238 ( .A(n28415), .B(n28416), .Z(n28399) );
  NOR U28239 ( .A(n28417), .B(n28418), .Z(n28416) );
  XOR U28240 ( .A(n28415), .B(n28419), .Z(n28417) );
  XNOR U28241 ( .A(n28398), .B(n28390), .Z(n28414) );
  XOR U28242 ( .A(n28420), .B(n28421), .Z(n28390) );
  AND U28243 ( .A(n28422), .B(n28423), .Z(n28421) );
  XOR U28244 ( .A(n28420), .B(n28424), .Z(n28422) );
  XNOR U28245 ( .A(n28425), .B(n28395), .Z(n28398) );
  XOR U28246 ( .A(n28426), .B(n28427), .Z(n28395) );
  AND U28247 ( .A(n28428), .B(n28429), .Z(n28427) );
  XNOR U28248 ( .A(n28430), .B(n28431), .Z(n28428) );
  IV U28249 ( .A(n28426), .Z(n28430) );
  XNOR U28250 ( .A(n28432), .B(n28433), .Z(n28425) );
  NOR U28251 ( .A(n28434), .B(n28435), .Z(n28433) );
  XNOR U28252 ( .A(n28432), .B(n28436), .Z(n28434) );
  XNOR U28253 ( .A(n28394), .B(n28401), .Z(n28413) );
  NOR U28254 ( .A(n28362), .B(n28437), .Z(n28401) );
  XOR U28255 ( .A(n28406), .B(n28405), .Z(n28394) );
  XNOR U28256 ( .A(n28438), .B(n28402), .Z(n28405) );
  XOR U28257 ( .A(n28439), .B(n28440), .Z(n28402) );
  AND U28258 ( .A(n28441), .B(n28442), .Z(n28440) );
  XNOR U28259 ( .A(n28443), .B(n28444), .Z(n28441) );
  IV U28260 ( .A(n28439), .Z(n28443) );
  XNOR U28261 ( .A(n28445), .B(n28446), .Z(n28438) );
  NOR U28262 ( .A(n28447), .B(n28448), .Z(n28446) );
  XNOR U28263 ( .A(n28445), .B(n28449), .Z(n28447) );
  XOR U28264 ( .A(n28450), .B(n28451), .Z(n28406) );
  NOR U28265 ( .A(n28452), .B(n28453), .Z(n28451) );
  XNOR U28266 ( .A(n28450), .B(n28454), .Z(n28452) );
  XNOR U28267 ( .A(n28351), .B(n28409), .Z(n28411) );
  XNOR U28268 ( .A(n28455), .B(n28456), .Z(n28351) );
  AND U28269 ( .A(n831), .B(n28358), .Z(n28456) );
  XOR U28270 ( .A(n28455), .B(n28356), .Z(n28358) );
  AND U28271 ( .A(n28359), .B(n28362), .Z(n28409) );
  XOR U28272 ( .A(n28457), .B(n28437), .Z(n28362) );
  XNOR U28273 ( .A(p_input[1152]), .B(p_input[2048]), .Z(n28437) );
  XNOR U28274 ( .A(n28424), .B(n28423), .Z(n28457) );
  XNOR U28275 ( .A(n28458), .B(n28431), .Z(n28423) );
  XNOR U28276 ( .A(n28419), .B(n28418), .Z(n28431) );
  XNOR U28277 ( .A(n28459), .B(n28415), .Z(n28418) );
  XNOR U28278 ( .A(p_input[1162]), .B(p_input[2058]), .Z(n28415) );
  XOR U28279 ( .A(p_input[1163]), .B(n16732), .Z(n28459) );
  XOR U28280 ( .A(p_input[1164]), .B(p_input[2060]), .Z(n28419) );
  XOR U28281 ( .A(n28429), .B(n28460), .Z(n28458) );
  IV U28282 ( .A(n28420), .Z(n28460) );
  XOR U28283 ( .A(p_input[1153]), .B(p_input[2049]), .Z(n28420) );
  XNOR U28284 ( .A(n28461), .B(n28436), .Z(n28429) );
  XNOR U28285 ( .A(p_input[1167]), .B(n16735), .Z(n28436) );
  XOR U28286 ( .A(n28426), .B(n28435), .Z(n28461) );
  XOR U28287 ( .A(n28462), .B(n28432), .Z(n28435) );
  XOR U28288 ( .A(p_input[1165]), .B(p_input[2061]), .Z(n28432) );
  XOR U28289 ( .A(p_input[1166]), .B(n16737), .Z(n28462) );
  XOR U28290 ( .A(p_input[1161]), .B(p_input[2057]), .Z(n28426) );
  XOR U28291 ( .A(n28444), .B(n28442), .Z(n28424) );
  XNOR U28292 ( .A(n28463), .B(n28449), .Z(n28442) );
  XOR U28293 ( .A(p_input[1160]), .B(p_input[2056]), .Z(n28449) );
  XOR U28294 ( .A(n28439), .B(n28448), .Z(n28463) );
  XOR U28295 ( .A(n28464), .B(n28445), .Z(n28448) );
  XOR U28296 ( .A(p_input[1158]), .B(p_input[2054]), .Z(n28445) );
  XOR U28297 ( .A(p_input[1159]), .B(n17722), .Z(n28464) );
  XOR U28298 ( .A(p_input[1154]), .B(p_input[2050]), .Z(n28439) );
  XNOR U28299 ( .A(n28454), .B(n28453), .Z(n28444) );
  XOR U28300 ( .A(n28465), .B(n28450), .Z(n28453) );
  XOR U28301 ( .A(p_input[1155]), .B(p_input[2051]), .Z(n28450) );
  XOR U28302 ( .A(p_input[1156]), .B(n17724), .Z(n28465) );
  XOR U28303 ( .A(p_input[1157]), .B(p_input[2053]), .Z(n28454) );
  XNOR U28304 ( .A(n28466), .B(n28467), .Z(n28359) );
  AND U28305 ( .A(n831), .B(n28468), .Z(n28467) );
  XNOR U28306 ( .A(n28469), .B(n28470), .Z(n831) );
  AND U28307 ( .A(n28471), .B(n28472), .Z(n28470) );
  XOR U28308 ( .A(n28469), .B(n28369), .Z(n28472) );
  XNOR U28309 ( .A(n28469), .B(n28323), .Z(n28471) );
  XOR U28310 ( .A(n28473), .B(n28474), .Z(n28469) );
  AND U28311 ( .A(n28475), .B(n28476), .Z(n28474) );
  XOR U28312 ( .A(n28473), .B(n28333), .Z(n28475) );
  XOR U28313 ( .A(n28477), .B(n28478), .Z(n28312) );
  AND U28314 ( .A(n835), .B(n28468), .Z(n28478) );
  XNOR U28315 ( .A(n28466), .B(n28477), .Z(n28468) );
  XNOR U28316 ( .A(n28479), .B(n28480), .Z(n835) );
  AND U28317 ( .A(n28481), .B(n28482), .Z(n28480) );
  XNOR U28318 ( .A(n28483), .B(n28479), .Z(n28482) );
  IV U28319 ( .A(n28369), .Z(n28483) );
  XNOR U28320 ( .A(n28484), .B(n28485), .Z(n28369) );
  AND U28321 ( .A(n838), .B(n28486), .Z(n28485) );
  XNOR U28322 ( .A(n28484), .B(n28487), .Z(n28486) );
  XNOR U28323 ( .A(n28323), .B(n28479), .Z(n28481) );
  XOR U28324 ( .A(n28488), .B(n28489), .Z(n28323) );
  AND U28325 ( .A(n846), .B(n28490), .Z(n28489) );
  XOR U28326 ( .A(n28473), .B(n28491), .Z(n28479) );
  AND U28327 ( .A(n28492), .B(n28476), .Z(n28491) );
  XNOR U28328 ( .A(n28382), .B(n28473), .Z(n28476) );
  XNOR U28329 ( .A(n28493), .B(n28494), .Z(n28382) );
  AND U28330 ( .A(n838), .B(n28495), .Z(n28494) );
  XOR U28331 ( .A(n28496), .B(n28493), .Z(n28495) );
  XNOR U28332 ( .A(n28497), .B(n28473), .Z(n28492) );
  IV U28333 ( .A(n28333), .Z(n28497) );
  XOR U28334 ( .A(n28498), .B(n28499), .Z(n28333) );
  AND U28335 ( .A(n846), .B(n28500), .Z(n28499) );
  XOR U28336 ( .A(n28501), .B(n28502), .Z(n28473) );
  AND U28337 ( .A(n28503), .B(n28504), .Z(n28502) );
  XNOR U28338 ( .A(n28407), .B(n28501), .Z(n28504) );
  XNOR U28339 ( .A(n28505), .B(n28506), .Z(n28407) );
  AND U28340 ( .A(n838), .B(n28507), .Z(n28506) );
  XNOR U28341 ( .A(n28508), .B(n28505), .Z(n28507) );
  XOR U28342 ( .A(n28501), .B(n28344), .Z(n28503) );
  XOR U28343 ( .A(n28509), .B(n28510), .Z(n28344) );
  AND U28344 ( .A(n846), .B(n28511), .Z(n28510) );
  XOR U28345 ( .A(n28512), .B(n28513), .Z(n28501) );
  AND U28346 ( .A(n28514), .B(n28515), .Z(n28513) );
  XNOR U28347 ( .A(n28512), .B(n28455), .Z(n28515) );
  XNOR U28348 ( .A(n28516), .B(n28517), .Z(n28455) );
  AND U28349 ( .A(n838), .B(n28518), .Z(n28517) );
  XOR U28350 ( .A(n28519), .B(n28516), .Z(n28518) );
  XNOR U28351 ( .A(n28520), .B(n28512), .Z(n28514) );
  IV U28352 ( .A(n28356), .Z(n28520) );
  XOR U28353 ( .A(n28521), .B(n28522), .Z(n28356) );
  AND U28354 ( .A(n846), .B(n28523), .Z(n28522) );
  AND U28355 ( .A(n28477), .B(n28466), .Z(n28512) );
  XNOR U28356 ( .A(n28524), .B(n28525), .Z(n28466) );
  AND U28357 ( .A(n838), .B(n28526), .Z(n28525) );
  XNOR U28358 ( .A(n28527), .B(n28524), .Z(n28526) );
  XNOR U28359 ( .A(n28528), .B(n28529), .Z(n838) );
  AND U28360 ( .A(n28530), .B(n28531), .Z(n28529) );
  XOR U28361 ( .A(n28487), .B(n28528), .Z(n28531) );
  AND U28362 ( .A(n28532), .B(n28533), .Z(n28487) );
  XOR U28363 ( .A(n28528), .B(n28484), .Z(n28530) );
  XNOR U28364 ( .A(n28534), .B(n28535), .Z(n28484) );
  AND U28365 ( .A(n842), .B(n28490), .Z(n28535) );
  XOR U28366 ( .A(n28488), .B(n28534), .Z(n28490) );
  XOR U28367 ( .A(n28536), .B(n28537), .Z(n28528) );
  AND U28368 ( .A(n28538), .B(n28539), .Z(n28537) );
  XNOR U28369 ( .A(n28536), .B(n28532), .Z(n28539) );
  IV U28370 ( .A(n28496), .Z(n28532) );
  XOR U28371 ( .A(n28540), .B(n28541), .Z(n28496) );
  XOR U28372 ( .A(n28542), .B(n28533), .Z(n28541) );
  AND U28373 ( .A(n28508), .B(n28543), .Z(n28533) );
  AND U28374 ( .A(n28544), .B(n28545), .Z(n28542) );
  XOR U28375 ( .A(n28546), .B(n28540), .Z(n28544) );
  XNOR U28376 ( .A(n28493), .B(n28536), .Z(n28538) );
  XNOR U28377 ( .A(n28547), .B(n28548), .Z(n28493) );
  AND U28378 ( .A(n842), .B(n28500), .Z(n28548) );
  XOR U28379 ( .A(n28547), .B(n28498), .Z(n28500) );
  XOR U28380 ( .A(n28549), .B(n28550), .Z(n28536) );
  AND U28381 ( .A(n28551), .B(n28552), .Z(n28550) );
  XNOR U28382 ( .A(n28549), .B(n28508), .Z(n28552) );
  XOR U28383 ( .A(n28553), .B(n28545), .Z(n28508) );
  XNOR U28384 ( .A(n28554), .B(n28540), .Z(n28545) );
  XOR U28385 ( .A(n28555), .B(n28556), .Z(n28540) );
  AND U28386 ( .A(n28557), .B(n28558), .Z(n28556) );
  XOR U28387 ( .A(n28559), .B(n28555), .Z(n28557) );
  XNOR U28388 ( .A(n28560), .B(n28561), .Z(n28554) );
  AND U28389 ( .A(n28562), .B(n28563), .Z(n28561) );
  XOR U28390 ( .A(n28560), .B(n28564), .Z(n28562) );
  XNOR U28391 ( .A(n28546), .B(n28543), .Z(n28553) );
  AND U28392 ( .A(n28565), .B(n28566), .Z(n28543) );
  XOR U28393 ( .A(n28567), .B(n28568), .Z(n28546) );
  AND U28394 ( .A(n28569), .B(n28570), .Z(n28568) );
  XOR U28395 ( .A(n28567), .B(n28571), .Z(n28569) );
  XNOR U28396 ( .A(n28505), .B(n28549), .Z(n28551) );
  XNOR U28397 ( .A(n28572), .B(n28573), .Z(n28505) );
  AND U28398 ( .A(n842), .B(n28511), .Z(n28573) );
  XOR U28399 ( .A(n28572), .B(n28509), .Z(n28511) );
  XOR U28400 ( .A(n28574), .B(n28575), .Z(n28549) );
  AND U28401 ( .A(n28576), .B(n28577), .Z(n28575) );
  XNOR U28402 ( .A(n28574), .B(n28565), .Z(n28577) );
  IV U28403 ( .A(n28519), .Z(n28565) );
  XNOR U28404 ( .A(n28578), .B(n28558), .Z(n28519) );
  XNOR U28405 ( .A(n28579), .B(n28564), .Z(n28558) );
  XNOR U28406 ( .A(n28580), .B(n28581), .Z(n28564) );
  NOR U28407 ( .A(n28582), .B(n28583), .Z(n28581) );
  XOR U28408 ( .A(n28580), .B(n28584), .Z(n28582) );
  XNOR U28409 ( .A(n28563), .B(n28555), .Z(n28579) );
  XOR U28410 ( .A(n28585), .B(n28586), .Z(n28555) );
  AND U28411 ( .A(n28587), .B(n28588), .Z(n28586) );
  XOR U28412 ( .A(n28585), .B(n28589), .Z(n28587) );
  XNOR U28413 ( .A(n28590), .B(n28560), .Z(n28563) );
  XOR U28414 ( .A(n28591), .B(n28592), .Z(n28560) );
  AND U28415 ( .A(n28593), .B(n28594), .Z(n28592) );
  XNOR U28416 ( .A(n28595), .B(n28596), .Z(n28593) );
  IV U28417 ( .A(n28591), .Z(n28595) );
  XNOR U28418 ( .A(n28597), .B(n28598), .Z(n28590) );
  NOR U28419 ( .A(n28599), .B(n28600), .Z(n28598) );
  XNOR U28420 ( .A(n28597), .B(n28601), .Z(n28599) );
  XNOR U28421 ( .A(n28559), .B(n28566), .Z(n28578) );
  NOR U28422 ( .A(n28527), .B(n28602), .Z(n28566) );
  XOR U28423 ( .A(n28571), .B(n28570), .Z(n28559) );
  XNOR U28424 ( .A(n28603), .B(n28567), .Z(n28570) );
  XOR U28425 ( .A(n28604), .B(n28605), .Z(n28567) );
  AND U28426 ( .A(n28606), .B(n28607), .Z(n28605) );
  XNOR U28427 ( .A(n28608), .B(n28609), .Z(n28606) );
  IV U28428 ( .A(n28604), .Z(n28608) );
  XNOR U28429 ( .A(n28610), .B(n28611), .Z(n28603) );
  NOR U28430 ( .A(n28612), .B(n28613), .Z(n28611) );
  XNOR U28431 ( .A(n28610), .B(n28614), .Z(n28612) );
  XOR U28432 ( .A(n28615), .B(n28616), .Z(n28571) );
  NOR U28433 ( .A(n28617), .B(n28618), .Z(n28616) );
  XNOR U28434 ( .A(n28615), .B(n28619), .Z(n28617) );
  XNOR U28435 ( .A(n28516), .B(n28574), .Z(n28576) );
  XNOR U28436 ( .A(n28620), .B(n28621), .Z(n28516) );
  AND U28437 ( .A(n842), .B(n28523), .Z(n28621) );
  XOR U28438 ( .A(n28620), .B(n28521), .Z(n28523) );
  AND U28439 ( .A(n28524), .B(n28527), .Z(n28574) );
  XOR U28440 ( .A(n28622), .B(n28602), .Z(n28527) );
  XNOR U28441 ( .A(p_input[1168]), .B(p_input[2048]), .Z(n28602) );
  XNOR U28442 ( .A(n28589), .B(n28588), .Z(n28622) );
  XNOR U28443 ( .A(n28623), .B(n28596), .Z(n28588) );
  XNOR U28444 ( .A(n28584), .B(n28583), .Z(n28596) );
  XNOR U28445 ( .A(n28624), .B(n28580), .Z(n28583) );
  XNOR U28446 ( .A(p_input[1178]), .B(p_input[2058]), .Z(n28580) );
  XOR U28447 ( .A(p_input[1179]), .B(n16732), .Z(n28624) );
  XOR U28448 ( .A(p_input[1180]), .B(p_input[2060]), .Z(n28584) );
  XOR U28449 ( .A(n28594), .B(n28625), .Z(n28623) );
  IV U28450 ( .A(n28585), .Z(n28625) );
  XOR U28451 ( .A(p_input[1169]), .B(p_input[2049]), .Z(n28585) );
  XNOR U28452 ( .A(n28626), .B(n28601), .Z(n28594) );
  XNOR U28453 ( .A(p_input[1183]), .B(n16735), .Z(n28601) );
  XOR U28454 ( .A(n28591), .B(n28600), .Z(n28626) );
  XOR U28455 ( .A(n28627), .B(n28597), .Z(n28600) );
  XOR U28456 ( .A(p_input[1181]), .B(p_input[2061]), .Z(n28597) );
  XOR U28457 ( .A(p_input[1182]), .B(n16737), .Z(n28627) );
  XOR U28458 ( .A(p_input[1177]), .B(p_input[2057]), .Z(n28591) );
  XOR U28459 ( .A(n28609), .B(n28607), .Z(n28589) );
  XNOR U28460 ( .A(n28628), .B(n28614), .Z(n28607) );
  XOR U28461 ( .A(p_input[1176]), .B(p_input[2056]), .Z(n28614) );
  XOR U28462 ( .A(n28604), .B(n28613), .Z(n28628) );
  XOR U28463 ( .A(n28629), .B(n28610), .Z(n28613) );
  XOR U28464 ( .A(p_input[1174]), .B(p_input[2054]), .Z(n28610) );
  XOR U28465 ( .A(p_input[1175]), .B(n17722), .Z(n28629) );
  XOR U28466 ( .A(p_input[1170]), .B(p_input[2050]), .Z(n28604) );
  XNOR U28467 ( .A(n28619), .B(n28618), .Z(n28609) );
  XOR U28468 ( .A(n28630), .B(n28615), .Z(n28618) );
  XOR U28469 ( .A(p_input[1171]), .B(p_input[2051]), .Z(n28615) );
  XOR U28470 ( .A(p_input[1172]), .B(n17724), .Z(n28630) );
  XOR U28471 ( .A(p_input[1173]), .B(p_input[2053]), .Z(n28619) );
  XNOR U28472 ( .A(n28631), .B(n28632), .Z(n28524) );
  AND U28473 ( .A(n842), .B(n28633), .Z(n28632) );
  XNOR U28474 ( .A(n28634), .B(n28635), .Z(n842) );
  AND U28475 ( .A(n28636), .B(n28637), .Z(n28635) );
  XOR U28476 ( .A(n28634), .B(n28534), .Z(n28637) );
  XNOR U28477 ( .A(n28634), .B(n28488), .Z(n28636) );
  XOR U28478 ( .A(n28638), .B(n28639), .Z(n28634) );
  AND U28479 ( .A(n28640), .B(n28641), .Z(n28639) );
  XOR U28480 ( .A(n28638), .B(n28498), .Z(n28640) );
  XOR U28481 ( .A(n28642), .B(n28643), .Z(n28477) );
  AND U28482 ( .A(n846), .B(n28633), .Z(n28643) );
  XNOR U28483 ( .A(n28631), .B(n28642), .Z(n28633) );
  XNOR U28484 ( .A(n28644), .B(n28645), .Z(n846) );
  AND U28485 ( .A(n28646), .B(n28647), .Z(n28645) );
  XNOR U28486 ( .A(n28648), .B(n28644), .Z(n28647) );
  IV U28487 ( .A(n28534), .Z(n28648) );
  XNOR U28488 ( .A(n28649), .B(n28650), .Z(n28534) );
  AND U28489 ( .A(n849), .B(n28651), .Z(n28650) );
  XNOR U28490 ( .A(n28649), .B(n28652), .Z(n28651) );
  XNOR U28491 ( .A(n28488), .B(n28644), .Z(n28646) );
  XOR U28492 ( .A(n28653), .B(n28654), .Z(n28488) );
  AND U28493 ( .A(n857), .B(n28655), .Z(n28654) );
  XOR U28494 ( .A(n28638), .B(n28656), .Z(n28644) );
  AND U28495 ( .A(n28657), .B(n28641), .Z(n28656) );
  XNOR U28496 ( .A(n28547), .B(n28638), .Z(n28641) );
  XNOR U28497 ( .A(n28658), .B(n28659), .Z(n28547) );
  AND U28498 ( .A(n849), .B(n28660), .Z(n28659) );
  XOR U28499 ( .A(n28661), .B(n28658), .Z(n28660) );
  XNOR U28500 ( .A(n28662), .B(n28638), .Z(n28657) );
  IV U28501 ( .A(n28498), .Z(n28662) );
  XOR U28502 ( .A(n28663), .B(n28664), .Z(n28498) );
  AND U28503 ( .A(n857), .B(n28665), .Z(n28664) );
  XOR U28504 ( .A(n28666), .B(n28667), .Z(n28638) );
  AND U28505 ( .A(n28668), .B(n28669), .Z(n28667) );
  XNOR U28506 ( .A(n28572), .B(n28666), .Z(n28669) );
  XNOR U28507 ( .A(n28670), .B(n28671), .Z(n28572) );
  AND U28508 ( .A(n849), .B(n28672), .Z(n28671) );
  XNOR U28509 ( .A(n28673), .B(n28670), .Z(n28672) );
  XOR U28510 ( .A(n28666), .B(n28509), .Z(n28668) );
  XOR U28511 ( .A(n28674), .B(n28675), .Z(n28509) );
  AND U28512 ( .A(n857), .B(n28676), .Z(n28675) );
  XOR U28513 ( .A(n28677), .B(n28678), .Z(n28666) );
  AND U28514 ( .A(n28679), .B(n28680), .Z(n28678) );
  XNOR U28515 ( .A(n28677), .B(n28620), .Z(n28680) );
  XNOR U28516 ( .A(n28681), .B(n28682), .Z(n28620) );
  AND U28517 ( .A(n849), .B(n28683), .Z(n28682) );
  XOR U28518 ( .A(n28684), .B(n28681), .Z(n28683) );
  XNOR U28519 ( .A(n28685), .B(n28677), .Z(n28679) );
  IV U28520 ( .A(n28521), .Z(n28685) );
  XOR U28521 ( .A(n28686), .B(n28687), .Z(n28521) );
  AND U28522 ( .A(n857), .B(n28688), .Z(n28687) );
  AND U28523 ( .A(n28642), .B(n28631), .Z(n28677) );
  XNOR U28524 ( .A(n28689), .B(n28690), .Z(n28631) );
  AND U28525 ( .A(n849), .B(n28691), .Z(n28690) );
  XNOR U28526 ( .A(n28692), .B(n28689), .Z(n28691) );
  XNOR U28527 ( .A(n28693), .B(n28694), .Z(n849) );
  AND U28528 ( .A(n28695), .B(n28696), .Z(n28694) );
  XOR U28529 ( .A(n28652), .B(n28693), .Z(n28696) );
  AND U28530 ( .A(n28697), .B(n28698), .Z(n28652) );
  XOR U28531 ( .A(n28693), .B(n28649), .Z(n28695) );
  XNOR U28532 ( .A(n28699), .B(n28700), .Z(n28649) );
  AND U28533 ( .A(n853), .B(n28655), .Z(n28700) );
  XOR U28534 ( .A(n28653), .B(n28699), .Z(n28655) );
  XOR U28535 ( .A(n28701), .B(n28702), .Z(n28693) );
  AND U28536 ( .A(n28703), .B(n28704), .Z(n28702) );
  XNOR U28537 ( .A(n28701), .B(n28697), .Z(n28704) );
  IV U28538 ( .A(n28661), .Z(n28697) );
  XOR U28539 ( .A(n28705), .B(n28706), .Z(n28661) );
  XOR U28540 ( .A(n28707), .B(n28698), .Z(n28706) );
  AND U28541 ( .A(n28673), .B(n28708), .Z(n28698) );
  AND U28542 ( .A(n28709), .B(n28710), .Z(n28707) );
  XOR U28543 ( .A(n28711), .B(n28705), .Z(n28709) );
  XNOR U28544 ( .A(n28658), .B(n28701), .Z(n28703) );
  XNOR U28545 ( .A(n28712), .B(n28713), .Z(n28658) );
  AND U28546 ( .A(n853), .B(n28665), .Z(n28713) );
  XOR U28547 ( .A(n28712), .B(n28663), .Z(n28665) );
  XOR U28548 ( .A(n28714), .B(n28715), .Z(n28701) );
  AND U28549 ( .A(n28716), .B(n28717), .Z(n28715) );
  XNOR U28550 ( .A(n28714), .B(n28673), .Z(n28717) );
  XOR U28551 ( .A(n28718), .B(n28710), .Z(n28673) );
  XNOR U28552 ( .A(n28719), .B(n28705), .Z(n28710) );
  XOR U28553 ( .A(n28720), .B(n28721), .Z(n28705) );
  AND U28554 ( .A(n28722), .B(n28723), .Z(n28721) );
  XOR U28555 ( .A(n28724), .B(n28720), .Z(n28722) );
  XNOR U28556 ( .A(n28725), .B(n28726), .Z(n28719) );
  AND U28557 ( .A(n28727), .B(n28728), .Z(n28726) );
  XOR U28558 ( .A(n28725), .B(n28729), .Z(n28727) );
  XNOR U28559 ( .A(n28711), .B(n28708), .Z(n28718) );
  AND U28560 ( .A(n28730), .B(n28731), .Z(n28708) );
  XOR U28561 ( .A(n28732), .B(n28733), .Z(n28711) );
  AND U28562 ( .A(n28734), .B(n28735), .Z(n28733) );
  XOR U28563 ( .A(n28732), .B(n28736), .Z(n28734) );
  XNOR U28564 ( .A(n28670), .B(n28714), .Z(n28716) );
  XNOR U28565 ( .A(n28737), .B(n28738), .Z(n28670) );
  AND U28566 ( .A(n853), .B(n28676), .Z(n28738) );
  XOR U28567 ( .A(n28737), .B(n28674), .Z(n28676) );
  XOR U28568 ( .A(n28739), .B(n28740), .Z(n28714) );
  AND U28569 ( .A(n28741), .B(n28742), .Z(n28740) );
  XNOR U28570 ( .A(n28739), .B(n28730), .Z(n28742) );
  IV U28571 ( .A(n28684), .Z(n28730) );
  XNOR U28572 ( .A(n28743), .B(n28723), .Z(n28684) );
  XNOR U28573 ( .A(n28744), .B(n28729), .Z(n28723) );
  XNOR U28574 ( .A(n28745), .B(n28746), .Z(n28729) );
  NOR U28575 ( .A(n28747), .B(n28748), .Z(n28746) );
  XOR U28576 ( .A(n28745), .B(n28749), .Z(n28747) );
  XNOR U28577 ( .A(n28728), .B(n28720), .Z(n28744) );
  XOR U28578 ( .A(n28750), .B(n28751), .Z(n28720) );
  AND U28579 ( .A(n28752), .B(n28753), .Z(n28751) );
  XOR U28580 ( .A(n28750), .B(n28754), .Z(n28752) );
  XNOR U28581 ( .A(n28755), .B(n28725), .Z(n28728) );
  XOR U28582 ( .A(n28756), .B(n28757), .Z(n28725) );
  AND U28583 ( .A(n28758), .B(n28759), .Z(n28757) );
  XNOR U28584 ( .A(n28760), .B(n28761), .Z(n28758) );
  IV U28585 ( .A(n28756), .Z(n28760) );
  XNOR U28586 ( .A(n28762), .B(n28763), .Z(n28755) );
  NOR U28587 ( .A(n28764), .B(n28765), .Z(n28763) );
  XNOR U28588 ( .A(n28762), .B(n28766), .Z(n28764) );
  XNOR U28589 ( .A(n28724), .B(n28731), .Z(n28743) );
  NOR U28590 ( .A(n28692), .B(n28767), .Z(n28731) );
  XOR U28591 ( .A(n28736), .B(n28735), .Z(n28724) );
  XNOR U28592 ( .A(n28768), .B(n28732), .Z(n28735) );
  XOR U28593 ( .A(n28769), .B(n28770), .Z(n28732) );
  AND U28594 ( .A(n28771), .B(n28772), .Z(n28770) );
  XNOR U28595 ( .A(n28773), .B(n28774), .Z(n28771) );
  IV U28596 ( .A(n28769), .Z(n28773) );
  XNOR U28597 ( .A(n28775), .B(n28776), .Z(n28768) );
  NOR U28598 ( .A(n28777), .B(n28778), .Z(n28776) );
  XNOR U28599 ( .A(n28775), .B(n28779), .Z(n28777) );
  XOR U28600 ( .A(n28780), .B(n28781), .Z(n28736) );
  NOR U28601 ( .A(n28782), .B(n28783), .Z(n28781) );
  XNOR U28602 ( .A(n28780), .B(n28784), .Z(n28782) );
  XNOR U28603 ( .A(n28681), .B(n28739), .Z(n28741) );
  XNOR U28604 ( .A(n28785), .B(n28786), .Z(n28681) );
  AND U28605 ( .A(n853), .B(n28688), .Z(n28786) );
  XOR U28606 ( .A(n28785), .B(n28686), .Z(n28688) );
  AND U28607 ( .A(n28689), .B(n28692), .Z(n28739) );
  XOR U28608 ( .A(n28787), .B(n28767), .Z(n28692) );
  XNOR U28609 ( .A(p_input[1184]), .B(p_input[2048]), .Z(n28767) );
  XNOR U28610 ( .A(n28754), .B(n28753), .Z(n28787) );
  XNOR U28611 ( .A(n28788), .B(n28761), .Z(n28753) );
  XNOR U28612 ( .A(n28749), .B(n28748), .Z(n28761) );
  XNOR U28613 ( .A(n28789), .B(n28745), .Z(n28748) );
  XNOR U28614 ( .A(p_input[1194]), .B(p_input[2058]), .Z(n28745) );
  XOR U28615 ( .A(p_input[1195]), .B(n16732), .Z(n28789) );
  XOR U28616 ( .A(p_input[1196]), .B(p_input[2060]), .Z(n28749) );
  XOR U28617 ( .A(n28759), .B(n28790), .Z(n28788) );
  IV U28618 ( .A(n28750), .Z(n28790) );
  XOR U28619 ( .A(p_input[1185]), .B(p_input[2049]), .Z(n28750) );
  XNOR U28620 ( .A(n28791), .B(n28766), .Z(n28759) );
  XNOR U28621 ( .A(p_input[1199]), .B(n16735), .Z(n28766) );
  XOR U28622 ( .A(n28756), .B(n28765), .Z(n28791) );
  XOR U28623 ( .A(n28792), .B(n28762), .Z(n28765) );
  XOR U28624 ( .A(p_input[1197]), .B(p_input[2061]), .Z(n28762) );
  XOR U28625 ( .A(p_input[1198]), .B(n16737), .Z(n28792) );
  XOR U28626 ( .A(p_input[1193]), .B(p_input[2057]), .Z(n28756) );
  XOR U28627 ( .A(n28774), .B(n28772), .Z(n28754) );
  XNOR U28628 ( .A(n28793), .B(n28779), .Z(n28772) );
  XOR U28629 ( .A(p_input[1192]), .B(p_input[2056]), .Z(n28779) );
  XOR U28630 ( .A(n28769), .B(n28778), .Z(n28793) );
  XOR U28631 ( .A(n28794), .B(n28775), .Z(n28778) );
  XOR U28632 ( .A(p_input[1190]), .B(p_input[2054]), .Z(n28775) );
  XOR U28633 ( .A(p_input[1191]), .B(n17722), .Z(n28794) );
  XOR U28634 ( .A(p_input[1186]), .B(p_input[2050]), .Z(n28769) );
  XNOR U28635 ( .A(n28784), .B(n28783), .Z(n28774) );
  XOR U28636 ( .A(n28795), .B(n28780), .Z(n28783) );
  XOR U28637 ( .A(p_input[1187]), .B(p_input[2051]), .Z(n28780) );
  XOR U28638 ( .A(p_input[1188]), .B(n17724), .Z(n28795) );
  XOR U28639 ( .A(p_input[1189]), .B(p_input[2053]), .Z(n28784) );
  XNOR U28640 ( .A(n28796), .B(n28797), .Z(n28689) );
  AND U28641 ( .A(n853), .B(n28798), .Z(n28797) );
  XNOR U28642 ( .A(n28799), .B(n28800), .Z(n853) );
  AND U28643 ( .A(n28801), .B(n28802), .Z(n28800) );
  XOR U28644 ( .A(n28799), .B(n28699), .Z(n28802) );
  XNOR U28645 ( .A(n28799), .B(n28653), .Z(n28801) );
  XOR U28646 ( .A(n28803), .B(n28804), .Z(n28799) );
  AND U28647 ( .A(n28805), .B(n28806), .Z(n28804) );
  XOR U28648 ( .A(n28803), .B(n28663), .Z(n28805) );
  XOR U28649 ( .A(n28807), .B(n28808), .Z(n28642) );
  AND U28650 ( .A(n857), .B(n28798), .Z(n28808) );
  XNOR U28651 ( .A(n28796), .B(n28807), .Z(n28798) );
  XNOR U28652 ( .A(n28809), .B(n28810), .Z(n857) );
  AND U28653 ( .A(n28811), .B(n28812), .Z(n28810) );
  XNOR U28654 ( .A(n28813), .B(n28809), .Z(n28812) );
  IV U28655 ( .A(n28699), .Z(n28813) );
  XNOR U28656 ( .A(n28814), .B(n28815), .Z(n28699) );
  AND U28657 ( .A(n860), .B(n28816), .Z(n28815) );
  XNOR U28658 ( .A(n28814), .B(n28817), .Z(n28816) );
  XNOR U28659 ( .A(n28653), .B(n28809), .Z(n28811) );
  XOR U28660 ( .A(n28818), .B(n28819), .Z(n28653) );
  AND U28661 ( .A(n868), .B(n28820), .Z(n28819) );
  XOR U28662 ( .A(n28803), .B(n28821), .Z(n28809) );
  AND U28663 ( .A(n28822), .B(n28806), .Z(n28821) );
  XNOR U28664 ( .A(n28712), .B(n28803), .Z(n28806) );
  XNOR U28665 ( .A(n28823), .B(n28824), .Z(n28712) );
  AND U28666 ( .A(n860), .B(n28825), .Z(n28824) );
  XOR U28667 ( .A(n28826), .B(n28823), .Z(n28825) );
  XNOR U28668 ( .A(n28827), .B(n28803), .Z(n28822) );
  IV U28669 ( .A(n28663), .Z(n28827) );
  XOR U28670 ( .A(n28828), .B(n28829), .Z(n28663) );
  AND U28671 ( .A(n868), .B(n28830), .Z(n28829) );
  XOR U28672 ( .A(n28831), .B(n28832), .Z(n28803) );
  AND U28673 ( .A(n28833), .B(n28834), .Z(n28832) );
  XNOR U28674 ( .A(n28737), .B(n28831), .Z(n28834) );
  XNOR U28675 ( .A(n28835), .B(n28836), .Z(n28737) );
  AND U28676 ( .A(n860), .B(n28837), .Z(n28836) );
  XNOR U28677 ( .A(n28838), .B(n28835), .Z(n28837) );
  XOR U28678 ( .A(n28831), .B(n28674), .Z(n28833) );
  XOR U28679 ( .A(n28839), .B(n28840), .Z(n28674) );
  AND U28680 ( .A(n868), .B(n28841), .Z(n28840) );
  XOR U28681 ( .A(n28842), .B(n28843), .Z(n28831) );
  AND U28682 ( .A(n28844), .B(n28845), .Z(n28843) );
  XNOR U28683 ( .A(n28842), .B(n28785), .Z(n28845) );
  XNOR U28684 ( .A(n28846), .B(n28847), .Z(n28785) );
  AND U28685 ( .A(n860), .B(n28848), .Z(n28847) );
  XOR U28686 ( .A(n28849), .B(n28846), .Z(n28848) );
  XNOR U28687 ( .A(n28850), .B(n28842), .Z(n28844) );
  IV U28688 ( .A(n28686), .Z(n28850) );
  XOR U28689 ( .A(n28851), .B(n28852), .Z(n28686) );
  AND U28690 ( .A(n868), .B(n28853), .Z(n28852) );
  AND U28691 ( .A(n28807), .B(n28796), .Z(n28842) );
  XNOR U28692 ( .A(n28854), .B(n28855), .Z(n28796) );
  AND U28693 ( .A(n860), .B(n28856), .Z(n28855) );
  XNOR U28694 ( .A(n28857), .B(n28854), .Z(n28856) );
  XNOR U28695 ( .A(n28858), .B(n28859), .Z(n860) );
  AND U28696 ( .A(n28860), .B(n28861), .Z(n28859) );
  XOR U28697 ( .A(n28817), .B(n28858), .Z(n28861) );
  AND U28698 ( .A(n28862), .B(n28863), .Z(n28817) );
  XOR U28699 ( .A(n28858), .B(n28814), .Z(n28860) );
  XNOR U28700 ( .A(n28864), .B(n28865), .Z(n28814) );
  AND U28701 ( .A(n864), .B(n28820), .Z(n28865) );
  XOR U28702 ( .A(n28818), .B(n28864), .Z(n28820) );
  XOR U28703 ( .A(n28866), .B(n28867), .Z(n28858) );
  AND U28704 ( .A(n28868), .B(n28869), .Z(n28867) );
  XNOR U28705 ( .A(n28866), .B(n28862), .Z(n28869) );
  IV U28706 ( .A(n28826), .Z(n28862) );
  XOR U28707 ( .A(n28870), .B(n28871), .Z(n28826) );
  XOR U28708 ( .A(n28872), .B(n28863), .Z(n28871) );
  AND U28709 ( .A(n28838), .B(n28873), .Z(n28863) );
  AND U28710 ( .A(n28874), .B(n28875), .Z(n28872) );
  XOR U28711 ( .A(n28876), .B(n28870), .Z(n28874) );
  XNOR U28712 ( .A(n28823), .B(n28866), .Z(n28868) );
  XNOR U28713 ( .A(n28877), .B(n28878), .Z(n28823) );
  AND U28714 ( .A(n864), .B(n28830), .Z(n28878) );
  XOR U28715 ( .A(n28877), .B(n28828), .Z(n28830) );
  XOR U28716 ( .A(n28879), .B(n28880), .Z(n28866) );
  AND U28717 ( .A(n28881), .B(n28882), .Z(n28880) );
  XNOR U28718 ( .A(n28879), .B(n28838), .Z(n28882) );
  XOR U28719 ( .A(n28883), .B(n28875), .Z(n28838) );
  XNOR U28720 ( .A(n28884), .B(n28870), .Z(n28875) );
  XOR U28721 ( .A(n28885), .B(n28886), .Z(n28870) );
  AND U28722 ( .A(n28887), .B(n28888), .Z(n28886) );
  XOR U28723 ( .A(n28889), .B(n28885), .Z(n28887) );
  XNOR U28724 ( .A(n28890), .B(n28891), .Z(n28884) );
  AND U28725 ( .A(n28892), .B(n28893), .Z(n28891) );
  XOR U28726 ( .A(n28890), .B(n28894), .Z(n28892) );
  XNOR U28727 ( .A(n28876), .B(n28873), .Z(n28883) );
  AND U28728 ( .A(n28895), .B(n28896), .Z(n28873) );
  XOR U28729 ( .A(n28897), .B(n28898), .Z(n28876) );
  AND U28730 ( .A(n28899), .B(n28900), .Z(n28898) );
  XOR U28731 ( .A(n28897), .B(n28901), .Z(n28899) );
  XNOR U28732 ( .A(n28835), .B(n28879), .Z(n28881) );
  XNOR U28733 ( .A(n28902), .B(n28903), .Z(n28835) );
  AND U28734 ( .A(n864), .B(n28841), .Z(n28903) );
  XOR U28735 ( .A(n28902), .B(n28839), .Z(n28841) );
  XOR U28736 ( .A(n28904), .B(n28905), .Z(n28879) );
  AND U28737 ( .A(n28906), .B(n28907), .Z(n28905) );
  XNOR U28738 ( .A(n28904), .B(n28895), .Z(n28907) );
  IV U28739 ( .A(n28849), .Z(n28895) );
  XNOR U28740 ( .A(n28908), .B(n28888), .Z(n28849) );
  XNOR U28741 ( .A(n28909), .B(n28894), .Z(n28888) );
  XNOR U28742 ( .A(n28910), .B(n28911), .Z(n28894) );
  NOR U28743 ( .A(n28912), .B(n28913), .Z(n28911) );
  XOR U28744 ( .A(n28910), .B(n28914), .Z(n28912) );
  XNOR U28745 ( .A(n28893), .B(n28885), .Z(n28909) );
  XOR U28746 ( .A(n28915), .B(n28916), .Z(n28885) );
  AND U28747 ( .A(n28917), .B(n28918), .Z(n28916) );
  XOR U28748 ( .A(n28915), .B(n28919), .Z(n28917) );
  XNOR U28749 ( .A(n28920), .B(n28890), .Z(n28893) );
  XOR U28750 ( .A(n28921), .B(n28922), .Z(n28890) );
  AND U28751 ( .A(n28923), .B(n28924), .Z(n28922) );
  XNOR U28752 ( .A(n28925), .B(n28926), .Z(n28923) );
  IV U28753 ( .A(n28921), .Z(n28925) );
  XNOR U28754 ( .A(n28927), .B(n28928), .Z(n28920) );
  NOR U28755 ( .A(n28929), .B(n28930), .Z(n28928) );
  XNOR U28756 ( .A(n28927), .B(n28931), .Z(n28929) );
  XNOR U28757 ( .A(n28889), .B(n28896), .Z(n28908) );
  NOR U28758 ( .A(n28857), .B(n28932), .Z(n28896) );
  XOR U28759 ( .A(n28901), .B(n28900), .Z(n28889) );
  XNOR U28760 ( .A(n28933), .B(n28897), .Z(n28900) );
  XOR U28761 ( .A(n28934), .B(n28935), .Z(n28897) );
  AND U28762 ( .A(n28936), .B(n28937), .Z(n28935) );
  XNOR U28763 ( .A(n28938), .B(n28939), .Z(n28936) );
  IV U28764 ( .A(n28934), .Z(n28938) );
  XNOR U28765 ( .A(n28940), .B(n28941), .Z(n28933) );
  NOR U28766 ( .A(n28942), .B(n28943), .Z(n28941) );
  XNOR U28767 ( .A(n28940), .B(n28944), .Z(n28942) );
  XOR U28768 ( .A(n28945), .B(n28946), .Z(n28901) );
  NOR U28769 ( .A(n28947), .B(n28948), .Z(n28946) );
  XNOR U28770 ( .A(n28945), .B(n28949), .Z(n28947) );
  XNOR U28771 ( .A(n28846), .B(n28904), .Z(n28906) );
  XNOR U28772 ( .A(n28950), .B(n28951), .Z(n28846) );
  AND U28773 ( .A(n864), .B(n28853), .Z(n28951) );
  XOR U28774 ( .A(n28950), .B(n28851), .Z(n28853) );
  AND U28775 ( .A(n28854), .B(n28857), .Z(n28904) );
  XOR U28776 ( .A(n28952), .B(n28932), .Z(n28857) );
  XNOR U28777 ( .A(p_input[1200]), .B(p_input[2048]), .Z(n28932) );
  XNOR U28778 ( .A(n28919), .B(n28918), .Z(n28952) );
  XNOR U28779 ( .A(n28953), .B(n28926), .Z(n28918) );
  XNOR U28780 ( .A(n28914), .B(n28913), .Z(n28926) );
  XNOR U28781 ( .A(n28954), .B(n28910), .Z(n28913) );
  XNOR U28782 ( .A(p_input[1210]), .B(p_input[2058]), .Z(n28910) );
  XOR U28783 ( .A(p_input[1211]), .B(n16732), .Z(n28954) );
  XOR U28784 ( .A(p_input[1212]), .B(p_input[2060]), .Z(n28914) );
  XOR U28785 ( .A(n28924), .B(n28955), .Z(n28953) );
  IV U28786 ( .A(n28915), .Z(n28955) );
  XOR U28787 ( .A(p_input[1201]), .B(p_input[2049]), .Z(n28915) );
  XNOR U28788 ( .A(n28956), .B(n28931), .Z(n28924) );
  XNOR U28789 ( .A(p_input[1215]), .B(n16735), .Z(n28931) );
  XOR U28790 ( .A(n28921), .B(n28930), .Z(n28956) );
  XOR U28791 ( .A(n28957), .B(n28927), .Z(n28930) );
  XOR U28792 ( .A(p_input[1213]), .B(p_input[2061]), .Z(n28927) );
  XOR U28793 ( .A(p_input[1214]), .B(n16737), .Z(n28957) );
  XOR U28794 ( .A(p_input[1209]), .B(p_input[2057]), .Z(n28921) );
  XOR U28795 ( .A(n28939), .B(n28937), .Z(n28919) );
  XNOR U28796 ( .A(n28958), .B(n28944), .Z(n28937) );
  XOR U28797 ( .A(p_input[1208]), .B(p_input[2056]), .Z(n28944) );
  XOR U28798 ( .A(n28934), .B(n28943), .Z(n28958) );
  XOR U28799 ( .A(n28959), .B(n28940), .Z(n28943) );
  XOR U28800 ( .A(p_input[1206]), .B(p_input[2054]), .Z(n28940) );
  XOR U28801 ( .A(p_input[1207]), .B(n17722), .Z(n28959) );
  XOR U28802 ( .A(p_input[1202]), .B(p_input[2050]), .Z(n28934) );
  XNOR U28803 ( .A(n28949), .B(n28948), .Z(n28939) );
  XOR U28804 ( .A(n28960), .B(n28945), .Z(n28948) );
  XOR U28805 ( .A(p_input[1203]), .B(p_input[2051]), .Z(n28945) );
  XOR U28806 ( .A(p_input[1204]), .B(n17724), .Z(n28960) );
  XOR U28807 ( .A(p_input[1205]), .B(p_input[2053]), .Z(n28949) );
  XNOR U28808 ( .A(n28961), .B(n28962), .Z(n28854) );
  AND U28809 ( .A(n864), .B(n28963), .Z(n28962) );
  XNOR U28810 ( .A(n28964), .B(n28965), .Z(n864) );
  AND U28811 ( .A(n28966), .B(n28967), .Z(n28965) );
  XOR U28812 ( .A(n28964), .B(n28864), .Z(n28967) );
  XNOR U28813 ( .A(n28964), .B(n28818), .Z(n28966) );
  XOR U28814 ( .A(n28968), .B(n28969), .Z(n28964) );
  AND U28815 ( .A(n28970), .B(n28971), .Z(n28969) );
  XOR U28816 ( .A(n28968), .B(n28828), .Z(n28970) );
  XOR U28817 ( .A(n28972), .B(n28973), .Z(n28807) );
  AND U28818 ( .A(n868), .B(n28963), .Z(n28973) );
  XNOR U28819 ( .A(n28961), .B(n28972), .Z(n28963) );
  XNOR U28820 ( .A(n28974), .B(n28975), .Z(n868) );
  AND U28821 ( .A(n28976), .B(n28977), .Z(n28975) );
  XNOR U28822 ( .A(n28978), .B(n28974), .Z(n28977) );
  IV U28823 ( .A(n28864), .Z(n28978) );
  XNOR U28824 ( .A(n28979), .B(n28980), .Z(n28864) );
  AND U28825 ( .A(n871), .B(n28981), .Z(n28980) );
  XNOR U28826 ( .A(n28979), .B(n28982), .Z(n28981) );
  XNOR U28827 ( .A(n28818), .B(n28974), .Z(n28976) );
  XOR U28828 ( .A(n28983), .B(n28984), .Z(n28818) );
  AND U28829 ( .A(n879), .B(n28985), .Z(n28984) );
  XOR U28830 ( .A(n28968), .B(n28986), .Z(n28974) );
  AND U28831 ( .A(n28987), .B(n28971), .Z(n28986) );
  XNOR U28832 ( .A(n28877), .B(n28968), .Z(n28971) );
  XNOR U28833 ( .A(n28988), .B(n28989), .Z(n28877) );
  AND U28834 ( .A(n871), .B(n28990), .Z(n28989) );
  XOR U28835 ( .A(n28991), .B(n28988), .Z(n28990) );
  XNOR U28836 ( .A(n28992), .B(n28968), .Z(n28987) );
  IV U28837 ( .A(n28828), .Z(n28992) );
  XOR U28838 ( .A(n28993), .B(n28994), .Z(n28828) );
  AND U28839 ( .A(n879), .B(n28995), .Z(n28994) );
  XOR U28840 ( .A(n28996), .B(n28997), .Z(n28968) );
  AND U28841 ( .A(n28998), .B(n28999), .Z(n28997) );
  XNOR U28842 ( .A(n28902), .B(n28996), .Z(n28999) );
  XNOR U28843 ( .A(n29000), .B(n29001), .Z(n28902) );
  AND U28844 ( .A(n871), .B(n29002), .Z(n29001) );
  XNOR U28845 ( .A(n29003), .B(n29000), .Z(n29002) );
  XOR U28846 ( .A(n28996), .B(n28839), .Z(n28998) );
  XOR U28847 ( .A(n29004), .B(n29005), .Z(n28839) );
  AND U28848 ( .A(n879), .B(n29006), .Z(n29005) );
  XOR U28849 ( .A(n29007), .B(n29008), .Z(n28996) );
  AND U28850 ( .A(n29009), .B(n29010), .Z(n29008) );
  XNOR U28851 ( .A(n29007), .B(n28950), .Z(n29010) );
  XNOR U28852 ( .A(n29011), .B(n29012), .Z(n28950) );
  AND U28853 ( .A(n871), .B(n29013), .Z(n29012) );
  XOR U28854 ( .A(n29014), .B(n29011), .Z(n29013) );
  XNOR U28855 ( .A(n29015), .B(n29007), .Z(n29009) );
  IV U28856 ( .A(n28851), .Z(n29015) );
  XOR U28857 ( .A(n29016), .B(n29017), .Z(n28851) );
  AND U28858 ( .A(n879), .B(n29018), .Z(n29017) );
  AND U28859 ( .A(n28972), .B(n28961), .Z(n29007) );
  XNOR U28860 ( .A(n29019), .B(n29020), .Z(n28961) );
  AND U28861 ( .A(n871), .B(n29021), .Z(n29020) );
  XNOR U28862 ( .A(n29022), .B(n29019), .Z(n29021) );
  XNOR U28863 ( .A(n29023), .B(n29024), .Z(n871) );
  AND U28864 ( .A(n29025), .B(n29026), .Z(n29024) );
  XOR U28865 ( .A(n28982), .B(n29023), .Z(n29026) );
  AND U28866 ( .A(n29027), .B(n29028), .Z(n28982) );
  XOR U28867 ( .A(n29023), .B(n28979), .Z(n29025) );
  XNOR U28868 ( .A(n29029), .B(n29030), .Z(n28979) );
  AND U28869 ( .A(n875), .B(n28985), .Z(n29030) );
  XOR U28870 ( .A(n28983), .B(n29029), .Z(n28985) );
  XOR U28871 ( .A(n29031), .B(n29032), .Z(n29023) );
  AND U28872 ( .A(n29033), .B(n29034), .Z(n29032) );
  XNOR U28873 ( .A(n29031), .B(n29027), .Z(n29034) );
  IV U28874 ( .A(n28991), .Z(n29027) );
  XOR U28875 ( .A(n29035), .B(n29036), .Z(n28991) );
  XOR U28876 ( .A(n29037), .B(n29028), .Z(n29036) );
  AND U28877 ( .A(n29003), .B(n29038), .Z(n29028) );
  AND U28878 ( .A(n29039), .B(n29040), .Z(n29037) );
  XOR U28879 ( .A(n29041), .B(n29035), .Z(n29039) );
  XNOR U28880 ( .A(n28988), .B(n29031), .Z(n29033) );
  XNOR U28881 ( .A(n29042), .B(n29043), .Z(n28988) );
  AND U28882 ( .A(n875), .B(n28995), .Z(n29043) );
  XOR U28883 ( .A(n29042), .B(n28993), .Z(n28995) );
  XOR U28884 ( .A(n29044), .B(n29045), .Z(n29031) );
  AND U28885 ( .A(n29046), .B(n29047), .Z(n29045) );
  XNOR U28886 ( .A(n29044), .B(n29003), .Z(n29047) );
  XOR U28887 ( .A(n29048), .B(n29040), .Z(n29003) );
  XNOR U28888 ( .A(n29049), .B(n29035), .Z(n29040) );
  XOR U28889 ( .A(n29050), .B(n29051), .Z(n29035) );
  AND U28890 ( .A(n29052), .B(n29053), .Z(n29051) );
  XOR U28891 ( .A(n29054), .B(n29050), .Z(n29052) );
  XNOR U28892 ( .A(n29055), .B(n29056), .Z(n29049) );
  AND U28893 ( .A(n29057), .B(n29058), .Z(n29056) );
  XOR U28894 ( .A(n29055), .B(n29059), .Z(n29057) );
  XNOR U28895 ( .A(n29041), .B(n29038), .Z(n29048) );
  AND U28896 ( .A(n29060), .B(n29061), .Z(n29038) );
  XOR U28897 ( .A(n29062), .B(n29063), .Z(n29041) );
  AND U28898 ( .A(n29064), .B(n29065), .Z(n29063) );
  XOR U28899 ( .A(n29062), .B(n29066), .Z(n29064) );
  XNOR U28900 ( .A(n29000), .B(n29044), .Z(n29046) );
  XNOR U28901 ( .A(n29067), .B(n29068), .Z(n29000) );
  AND U28902 ( .A(n875), .B(n29006), .Z(n29068) );
  XOR U28903 ( .A(n29067), .B(n29004), .Z(n29006) );
  XOR U28904 ( .A(n29069), .B(n29070), .Z(n29044) );
  AND U28905 ( .A(n29071), .B(n29072), .Z(n29070) );
  XNOR U28906 ( .A(n29069), .B(n29060), .Z(n29072) );
  IV U28907 ( .A(n29014), .Z(n29060) );
  XNOR U28908 ( .A(n29073), .B(n29053), .Z(n29014) );
  XNOR U28909 ( .A(n29074), .B(n29059), .Z(n29053) );
  XNOR U28910 ( .A(n29075), .B(n29076), .Z(n29059) );
  NOR U28911 ( .A(n29077), .B(n29078), .Z(n29076) );
  XOR U28912 ( .A(n29075), .B(n29079), .Z(n29077) );
  XNOR U28913 ( .A(n29058), .B(n29050), .Z(n29074) );
  XOR U28914 ( .A(n29080), .B(n29081), .Z(n29050) );
  AND U28915 ( .A(n29082), .B(n29083), .Z(n29081) );
  XOR U28916 ( .A(n29080), .B(n29084), .Z(n29082) );
  XNOR U28917 ( .A(n29085), .B(n29055), .Z(n29058) );
  XOR U28918 ( .A(n29086), .B(n29087), .Z(n29055) );
  AND U28919 ( .A(n29088), .B(n29089), .Z(n29087) );
  XNOR U28920 ( .A(n29090), .B(n29091), .Z(n29088) );
  IV U28921 ( .A(n29086), .Z(n29090) );
  XNOR U28922 ( .A(n29092), .B(n29093), .Z(n29085) );
  NOR U28923 ( .A(n29094), .B(n29095), .Z(n29093) );
  XNOR U28924 ( .A(n29092), .B(n29096), .Z(n29094) );
  XNOR U28925 ( .A(n29054), .B(n29061), .Z(n29073) );
  NOR U28926 ( .A(n29022), .B(n29097), .Z(n29061) );
  XOR U28927 ( .A(n29066), .B(n29065), .Z(n29054) );
  XNOR U28928 ( .A(n29098), .B(n29062), .Z(n29065) );
  XOR U28929 ( .A(n29099), .B(n29100), .Z(n29062) );
  AND U28930 ( .A(n29101), .B(n29102), .Z(n29100) );
  XNOR U28931 ( .A(n29103), .B(n29104), .Z(n29101) );
  IV U28932 ( .A(n29099), .Z(n29103) );
  XNOR U28933 ( .A(n29105), .B(n29106), .Z(n29098) );
  NOR U28934 ( .A(n29107), .B(n29108), .Z(n29106) );
  XNOR U28935 ( .A(n29105), .B(n29109), .Z(n29107) );
  XOR U28936 ( .A(n29110), .B(n29111), .Z(n29066) );
  NOR U28937 ( .A(n29112), .B(n29113), .Z(n29111) );
  XNOR U28938 ( .A(n29110), .B(n29114), .Z(n29112) );
  XNOR U28939 ( .A(n29011), .B(n29069), .Z(n29071) );
  XNOR U28940 ( .A(n29115), .B(n29116), .Z(n29011) );
  AND U28941 ( .A(n875), .B(n29018), .Z(n29116) );
  XOR U28942 ( .A(n29115), .B(n29016), .Z(n29018) );
  AND U28943 ( .A(n29019), .B(n29022), .Z(n29069) );
  XOR U28944 ( .A(n29117), .B(n29097), .Z(n29022) );
  XNOR U28945 ( .A(p_input[1216]), .B(p_input[2048]), .Z(n29097) );
  XNOR U28946 ( .A(n29084), .B(n29083), .Z(n29117) );
  XNOR U28947 ( .A(n29118), .B(n29091), .Z(n29083) );
  XNOR U28948 ( .A(n29079), .B(n29078), .Z(n29091) );
  XNOR U28949 ( .A(n29119), .B(n29075), .Z(n29078) );
  XNOR U28950 ( .A(p_input[1226]), .B(p_input[2058]), .Z(n29075) );
  XOR U28951 ( .A(p_input[1227]), .B(n16732), .Z(n29119) );
  XOR U28952 ( .A(p_input[1228]), .B(p_input[2060]), .Z(n29079) );
  XOR U28953 ( .A(n29089), .B(n29120), .Z(n29118) );
  IV U28954 ( .A(n29080), .Z(n29120) );
  XOR U28955 ( .A(p_input[1217]), .B(p_input[2049]), .Z(n29080) );
  XNOR U28956 ( .A(n29121), .B(n29096), .Z(n29089) );
  XNOR U28957 ( .A(p_input[1231]), .B(n16735), .Z(n29096) );
  XOR U28958 ( .A(n29086), .B(n29095), .Z(n29121) );
  XOR U28959 ( .A(n29122), .B(n29092), .Z(n29095) );
  XOR U28960 ( .A(p_input[1229]), .B(p_input[2061]), .Z(n29092) );
  XOR U28961 ( .A(p_input[1230]), .B(n16737), .Z(n29122) );
  XOR U28962 ( .A(p_input[1225]), .B(p_input[2057]), .Z(n29086) );
  XOR U28963 ( .A(n29104), .B(n29102), .Z(n29084) );
  XNOR U28964 ( .A(n29123), .B(n29109), .Z(n29102) );
  XOR U28965 ( .A(p_input[1224]), .B(p_input[2056]), .Z(n29109) );
  XOR U28966 ( .A(n29099), .B(n29108), .Z(n29123) );
  XOR U28967 ( .A(n29124), .B(n29105), .Z(n29108) );
  XOR U28968 ( .A(p_input[1222]), .B(p_input[2054]), .Z(n29105) );
  XOR U28969 ( .A(p_input[1223]), .B(n17722), .Z(n29124) );
  XOR U28970 ( .A(p_input[1218]), .B(p_input[2050]), .Z(n29099) );
  XNOR U28971 ( .A(n29114), .B(n29113), .Z(n29104) );
  XOR U28972 ( .A(n29125), .B(n29110), .Z(n29113) );
  XOR U28973 ( .A(p_input[1219]), .B(p_input[2051]), .Z(n29110) );
  XOR U28974 ( .A(p_input[1220]), .B(n17724), .Z(n29125) );
  XOR U28975 ( .A(p_input[1221]), .B(p_input[2053]), .Z(n29114) );
  XNOR U28976 ( .A(n29126), .B(n29127), .Z(n29019) );
  AND U28977 ( .A(n875), .B(n29128), .Z(n29127) );
  XNOR U28978 ( .A(n29129), .B(n29130), .Z(n875) );
  AND U28979 ( .A(n29131), .B(n29132), .Z(n29130) );
  XOR U28980 ( .A(n29129), .B(n29029), .Z(n29132) );
  XNOR U28981 ( .A(n29129), .B(n28983), .Z(n29131) );
  XOR U28982 ( .A(n29133), .B(n29134), .Z(n29129) );
  AND U28983 ( .A(n29135), .B(n29136), .Z(n29134) );
  XOR U28984 ( .A(n29133), .B(n28993), .Z(n29135) );
  XOR U28985 ( .A(n29137), .B(n29138), .Z(n28972) );
  AND U28986 ( .A(n879), .B(n29128), .Z(n29138) );
  XNOR U28987 ( .A(n29126), .B(n29137), .Z(n29128) );
  XNOR U28988 ( .A(n29139), .B(n29140), .Z(n879) );
  AND U28989 ( .A(n29141), .B(n29142), .Z(n29140) );
  XNOR U28990 ( .A(n29143), .B(n29139), .Z(n29142) );
  IV U28991 ( .A(n29029), .Z(n29143) );
  XNOR U28992 ( .A(n29144), .B(n29145), .Z(n29029) );
  AND U28993 ( .A(n882), .B(n29146), .Z(n29145) );
  XNOR U28994 ( .A(n29144), .B(n29147), .Z(n29146) );
  XNOR U28995 ( .A(n28983), .B(n29139), .Z(n29141) );
  XOR U28996 ( .A(n29148), .B(n29149), .Z(n28983) );
  AND U28997 ( .A(n890), .B(n29150), .Z(n29149) );
  XOR U28998 ( .A(n29133), .B(n29151), .Z(n29139) );
  AND U28999 ( .A(n29152), .B(n29136), .Z(n29151) );
  XNOR U29000 ( .A(n29042), .B(n29133), .Z(n29136) );
  XNOR U29001 ( .A(n29153), .B(n29154), .Z(n29042) );
  AND U29002 ( .A(n882), .B(n29155), .Z(n29154) );
  XOR U29003 ( .A(n29156), .B(n29153), .Z(n29155) );
  XNOR U29004 ( .A(n29157), .B(n29133), .Z(n29152) );
  IV U29005 ( .A(n28993), .Z(n29157) );
  XOR U29006 ( .A(n29158), .B(n29159), .Z(n28993) );
  AND U29007 ( .A(n890), .B(n29160), .Z(n29159) );
  XOR U29008 ( .A(n29161), .B(n29162), .Z(n29133) );
  AND U29009 ( .A(n29163), .B(n29164), .Z(n29162) );
  XNOR U29010 ( .A(n29067), .B(n29161), .Z(n29164) );
  XNOR U29011 ( .A(n29165), .B(n29166), .Z(n29067) );
  AND U29012 ( .A(n882), .B(n29167), .Z(n29166) );
  XNOR U29013 ( .A(n29168), .B(n29165), .Z(n29167) );
  XOR U29014 ( .A(n29161), .B(n29004), .Z(n29163) );
  XOR U29015 ( .A(n29169), .B(n29170), .Z(n29004) );
  AND U29016 ( .A(n890), .B(n29171), .Z(n29170) );
  XOR U29017 ( .A(n29172), .B(n29173), .Z(n29161) );
  AND U29018 ( .A(n29174), .B(n29175), .Z(n29173) );
  XNOR U29019 ( .A(n29172), .B(n29115), .Z(n29175) );
  XNOR U29020 ( .A(n29176), .B(n29177), .Z(n29115) );
  AND U29021 ( .A(n882), .B(n29178), .Z(n29177) );
  XOR U29022 ( .A(n29179), .B(n29176), .Z(n29178) );
  XNOR U29023 ( .A(n29180), .B(n29172), .Z(n29174) );
  IV U29024 ( .A(n29016), .Z(n29180) );
  XOR U29025 ( .A(n29181), .B(n29182), .Z(n29016) );
  AND U29026 ( .A(n890), .B(n29183), .Z(n29182) );
  AND U29027 ( .A(n29137), .B(n29126), .Z(n29172) );
  XNOR U29028 ( .A(n29184), .B(n29185), .Z(n29126) );
  AND U29029 ( .A(n882), .B(n29186), .Z(n29185) );
  XNOR U29030 ( .A(n29187), .B(n29184), .Z(n29186) );
  XNOR U29031 ( .A(n29188), .B(n29189), .Z(n882) );
  AND U29032 ( .A(n29190), .B(n29191), .Z(n29189) );
  XOR U29033 ( .A(n29147), .B(n29188), .Z(n29191) );
  AND U29034 ( .A(n29192), .B(n29193), .Z(n29147) );
  XOR U29035 ( .A(n29188), .B(n29144), .Z(n29190) );
  XNOR U29036 ( .A(n29194), .B(n29195), .Z(n29144) );
  AND U29037 ( .A(n886), .B(n29150), .Z(n29195) );
  XOR U29038 ( .A(n29148), .B(n29194), .Z(n29150) );
  XOR U29039 ( .A(n29196), .B(n29197), .Z(n29188) );
  AND U29040 ( .A(n29198), .B(n29199), .Z(n29197) );
  XNOR U29041 ( .A(n29196), .B(n29192), .Z(n29199) );
  IV U29042 ( .A(n29156), .Z(n29192) );
  XOR U29043 ( .A(n29200), .B(n29201), .Z(n29156) );
  XOR U29044 ( .A(n29202), .B(n29193), .Z(n29201) );
  AND U29045 ( .A(n29168), .B(n29203), .Z(n29193) );
  AND U29046 ( .A(n29204), .B(n29205), .Z(n29202) );
  XOR U29047 ( .A(n29206), .B(n29200), .Z(n29204) );
  XNOR U29048 ( .A(n29153), .B(n29196), .Z(n29198) );
  XNOR U29049 ( .A(n29207), .B(n29208), .Z(n29153) );
  AND U29050 ( .A(n886), .B(n29160), .Z(n29208) );
  XOR U29051 ( .A(n29207), .B(n29158), .Z(n29160) );
  XOR U29052 ( .A(n29209), .B(n29210), .Z(n29196) );
  AND U29053 ( .A(n29211), .B(n29212), .Z(n29210) );
  XNOR U29054 ( .A(n29209), .B(n29168), .Z(n29212) );
  XOR U29055 ( .A(n29213), .B(n29205), .Z(n29168) );
  XNOR U29056 ( .A(n29214), .B(n29200), .Z(n29205) );
  XOR U29057 ( .A(n29215), .B(n29216), .Z(n29200) );
  AND U29058 ( .A(n29217), .B(n29218), .Z(n29216) );
  XOR U29059 ( .A(n29219), .B(n29215), .Z(n29217) );
  XNOR U29060 ( .A(n29220), .B(n29221), .Z(n29214) );
  AND U29061 ( .A(n29222), .B(n29223), .Z(n29221) );
  XOR U29062 ( .A(n29220), .B(n29224), .Z(n29222) );
  XNOR U29063 ( .A(n29206), .B(n29203), .Z(n29213) );
  AND U29064 ( .A(n29225), .B(n29226), .Z(n29203) );
  XOR U29065 ( .A(n29227), .B(n29228), .Z(n29206) );
  AND U29066 ( .A(n29229), .B(n29230), .Z(n29228) );
  XOR U29067 ( .A(n29227), .B(n29231), .Z(n29229) );
  XNOR U29068 ( .A(n29165), .B(n29209), .Z(n29211) );
  XNOR U29069 ( .A(n29232), .B(n29233), .Z(n29165) );
  AND U29070 ( .A(n886), .B(n29171), .Z(n29233) );
  XOR U29071 ( .A(n29232), .B(n29169), .Z(n29171) );
  XOR U29072 ( .A(n29234), .B(n29235), .Z(n29209) );
  AND U29073 ( .A(n29236), .B(n29237), .Z(n29235) );
  XNOR U29074 ( .A(n29234), .B(n29225), .Z(n29237) );
  IV U29075 ( .A(n29179), .Z(n29225) );
  XNOR U29076 ( .A(n29238), .B(n29218), .Z(n29179) );
  XNOR U29077 ( .A(n29239), .B(n29224), .Z(n29218) );
  XNOR U29078 ( .A(n29240), .B(n29241), .Z(n29224) );
  NOR U29079 ( .A(n29242), .B(n29243), .Z(n29241) );
  XOR U29080 ( .A(n29240), .B(n29244), .Z(n29242) );
  XNOR U29081 ( .A(n29223), .B(n29215), .Z(n29239) );
  XOR U29082 ( .A(n29245), .B(n29246), .Z(n29215) );
  AND U29083 ( .A(n29247), .B(n29248), .Z(n29246) );
  XOR U29084 ( .A(n29245), .B(n29249), .Z(n29247) );
  XNOR U29085 ( .A(n29250), .B(n29220), .Z(n29223) );
  XOR U29086 ( .A(n29251), .B(n29252), .Z(n29220) );
  AND U29087 ( .A(n29253), .B(n29254), .Z(n29252) );
  XNOR U29088 ( .A(n29255), .B(n29256), .Z(n29253) );
  IV U29089 ( .A(n29251), .Z(n29255) );
  XNOR U29090 ( .A(n29257), .B(n29258), .Z(n29250) );
  NOR U29091 ( .A(n29259), .B(n29260), .Z(n29258) );
  XNOR U29092 ( .A(n29257), .B(n29261), .Z(n29259) );
  XNOR U29093 ( .A(n29219), .B(n29226), .Z(n29238) );
  NOR U29094 ( .A(n29187), .B(n29262), .Z(n29226) );
  XOR U29095 ( .A(n29231), .B(n29230), .Z(n29219) );
  XNOR U29096 ( .A(n29263), .B(n29227), .Z(n29230) );
  XOR U29097 ( .A(n29264), .B(n29265), .Z(n29227) );
  AND U29098 ( .A(n29266), .B(n29267), .Z(n29265) );
  XNOR U29099 ( .A(n29268), .B(n29269), .Z(n29266) );
  IV U29100 ( .A(n29264), .Z(n29268) );
  XNOR U29101 ( .A(n29270), .B(n29271), .Z(n29263) );
  NOR U29102 ( .A(n29272), .B(n29273), .Z(n29271) );
  XNOR U29103 ( .A(n29270), .B(n29274), .Z(n29272) );
  XOR U29104 ( .A(n29275), .B(n29276), .Z(n29231) );
  NOR U29105 ( .A(n29277), .B(n29278), .Z(n29276) );
  XNOR U29106 ( .A(n29275), .B(n29279), .Z(n29277) );
  XNOR U29107 ( .A(n29176), .B(n29234), .Z(n29236) );
  XNOR U29108 ( .A(n29280), .B(n29281), .Z(n29176) );
  AND U29109 ( .A(n886), .B(n29183), .Z(n29281) );
  XOR U29110 ( .A(n29280), .B(n29181), .Z(n29183) );
  AND U29111 ( .A(n29184), .B(n29187), .Z(n29234) );
  XOR U29112 ( .A(n29282), .B(n29262), .Z(n29187) );
  XNOR U29113 ( .A(p_input[1232]), .B(p_input[2048]), .Z(n29262) );
  XNOR U29114 ( .A(n29249), .B(n29248), .Z(n29282) );
  XNOR U29115 ( .A(n29283), .B(n29256), .Z(n29248) );
  XNOR U29116 ( .A(n29244), .B(n29243), .Z(n29256) );
  XNOR U29117 ( .A(n29284), .B(n29240), .Z(n29243) );
  XNOR U29118 ( .A(p_input[1242]), .B(p_input[2058]), .Z(n29240) );
  XOR U29119 ( .A(p_input[1243]), .B(n16732), .Z(n29284) );
  XOR U29120 ( .A(p_input[1244]), .B(p_input[2060]), .Z(n29244) );
  XOR U29121 ( .A(n29254), .B(n29285), .Z(n29283) );
  IV U29122 ( .A(n29245), .Z(n29285) );
  XOR U29123 ( .A(p_input[1233]), .B(p_input[2049]), .Z(n29245) );
  XNOR U29124 ( .A(n29286), .B(n29261), .Z(n29254) );
  XNOR U29125 ( .A(p_input[1247]), .B(n16735), .Z(n29261) );
  XOR U29126 ( .A(n29251), .B(n29260), .Z(n29286) );
  XOR U29127 ( .A(n29287), .B(n29257), .Z(n29260) );
  XOR U29128 ( .A(p_input[1245]), .B(p_input[2061]), .Z(n29257) );
  XOR U29129 ( .A(p_input[1246]), .B(n16737), .Z(n29287) );
  XOR U29130 ( .A(p_input[1241]), .B(p_input[2057]), .Z(n29251) );
  XOR U29131 ( .A(n29269), .B(n29267), .Z(n29249) );
  XNOR U29132 ( .A(n29288), .B(n29274), .Z(n29267) );
  XOR U29133 ( .A(p_input[1240]), .B(p_input[2056]), .Z(n29274) );
  XOR U29134 ( .A(n29264), .B(n29273), .Z(n29288) );
  XOR U29135 ( .A(n29289), .B(n29270), .Z(n29273) );
  XOR U29136 ( .A(p_input[1238]), .B(p_input[2054]), .Z(n29270) );
  XOR U29137 ( .A(p_input[1239]), .B(n17722), .Z(n29289) );
  XOR U29138 ( .A(p_input[1234]), .B(p_input[2050]), .Z(n29264) );
  XNOR U29139 ( .A(n29279), .B(n29278), .Z(n29269) );
  XOR U29140 ( .A(n29290), .B(n29275), .Z(n29278) );
  XOR U29141 ( .A(p_input[1235]), .B(p_input[2051]), .Z(n29275) );
  XOR U29142 ( .A(p_input[1236]), .B(n17724), .Z(n29290) );
  XOR U29143 ( .A(p_input[1237]), .B(p_input[2053]), .Z(n29279) );
  XNOR U29144 ( .A(n29291), .B(n29292), .Z(n29184) );
  AND U29145 ( .A(n886), .B(n29293), .Z(n29292) );
  XNOR U29146 ( .A(n29294), .B(n29295), .Z(n886) );
  AND U29147 ( .A(n29296), .B(n29297), .Z(n29295) );
  XOR U29148 ( .A(n29294), .B(n29194), .Z(n29297) );
  XNOR U29149 ( .A(n29294), .B(n29148), .Z(n29296) );
  XOR U29150 ( .A(n29298), .B(n29299), .Z(n29294) );
  AND U29151 ( .A(n29300), .B(n29301), .Z(n29299) );
  XOR U29152 ( .A(n29298), .B(n29158), .Z(n29300) );
  XOR U29153 ( .A(n29302), .B(n29303), .Z(n29137) );
  AND U29154 ( .A(n890), .B(n29293), .Z(n29303) );
  XNOR U29155 ( .A(n29291), .B(n29302), .Z(n29293) );
  XNOR U29156 ( .A(n29304), .B(n29305), .Z(n890) );
  AND U29157 ( .A(n29306), .B(n29307), .Z(n29305) );
  XNOR U29158 ( .A(n29308), .B(n29304), .Z(n29307) );
  IV U29159 ( .A(n29194), .Z(n29308) );
  XNOR U29160 ( .A(n29309), .B(n29310), .Z(n29194) );
  AND U29161 ( .A(n893), .B(n29311), .Z(n29310) );
  XNOR U29162 ( .A(n29309), .B(n29312), .Z(n29311) );
  XNOR U29163 ( .A(n29148), .B(n29304), .Z(n29306) );
  XOR U29164 ( .A(n29313), .B(n29314), .Z(n29148) );
  AND U29165 ( .A(n901), .B(n29315), .Z(n29314) );
  XOR U29166 ( .A(n29298), .B(n29316), .Z(n29304) );
  AND U29167 ( .A(n29317), .B(n29301), .Z(n29316) );
  XNOR U29168 ( .A(n29207), .B(n29298), .Z(n29301) );
  XNOR U29169 ( .A(n29318), .B(n29319), .Z(n29207) );
  AND U29170 ( .A(n893), .B(n29320), .Z(n29319) );
  XOR U29171 ( .A(n29321), .B(n29318), .Z(n29320) );
  XNOR U29172 ( .A(n29322), .B(n29298), .Z(n29317) );
  IV U29173 ( .A(n29158), .Z(n29322) );
  XOR U29174 ( .A(n29323), .B(n29324), .Z(n29158) );
  AND U29175 ( .A(n901), .B(n29325), .Z(n29324) );
  XOR U29176 ( .A(n29326), .B(n29327), .Z(n29298) );
  AND U29177 ( .A(n29328), .B(n29329), .Z(n29327) );
  XNOR U29178 ( .A(n29232), .B(n29326), .Z(n29329) );
  XNOR U29179 ( .A(n29330), .B(n29331), .Z(n29232) );
  AND U29180 ( .A(n893), .B(n29332), .Z(n29331) );
  XNOR U29181 ( .A(n29333), .B(n29330), .Z(n29332) );
  XOR U29182 ( .A(n29326), .B(n29169), .Z(n29328) );
  XOR U29183 ( .A(n29334), .B(n29335), .Z(n29169) );
  AND U29184 ( .A(n901), .B(n29336), .Z(n29335) );
  XOR U29185 ( .A(n29337), .B(n29338), .Z(n29326) );
  AND U29186 ( .A(n29339), .B(n29340), .Z(n29338) );
  XNOR U29187 ( .A(n29337), .B(n29280), .Z(n29340) );
  XNOR U29188 ( .A(n29341), .B(n29342), .Z(n29280) );
  AND U29189 ( .A(n893), .B(n29343), .Z(n29342) );
  XOR U29190 ( .A(n29344), .B(n29341), .Z(n29343) );
  XNOR U29191 ( .A(n29345), .B(n29337), .Z(n29339) );
  IV U29192 ( .A(n29181), .Z(n29345) );
  XOR U29193 ( .A(n29346), .B(n29347), .Z(n29181) );
  AND U29194 ( .A(n901), .B(n29348), .Z(n29347) );
  AND U29195 ( .A(n29302), .B(n29291), .Z(n29337) );
  XNOR U29196 ( .A(n29349), .B(n29350), .Z(n29291) );
  AND U29197 ( .A(n893), .B(n29351), .Z(n29350) );
  XNOR U29198 ( .A(n29352), .B(n29349), .Z(n29351) );
  XNOR U29199 ( .A(n29353), .B(n29354), .Z(n893) );
  AND U29200 ( .A(n29355), .B(n29356), .Z(n29354) );
  XOR U29201 ( .A(n29312), .B(n29353), .Z(n29356) );
  AND U29202 ( .A(n29357), .B(n29358), .Z(n29312) );
  XOR U29203 ( .A(n29353), .B(n29309), .Z(n29355) );
  XNOR U29204 ( .A(n29359), .B(n29360), .Z(n29309) );
  AND U29205 ( .A(n897), .B(n29315), .Z(n29360) );
  XOR U29206 ( .A(n29313), .B(n29359), .Z(n29315) );
  XOR U29207 ( .A(n29361), .B(n29362), .Z(n29353) );
  AND U29208 ( .A(n29363), .B(n29364), .Z(n29362) );
  XNOR U29209 ( .A(n29361), .B(n29357), .Z(n29364) );
  IV U29210 ( .A(n29321), .Z(n29357) );
  XOR U29211 ( .A(n29365), .B(n29366), .Z(n29321) );
  XOR U29212 ( .A(n29367), .B(n29358), .Z(n29366) );
  AND U29213 ( .A(n29333), .B(n29368), .Z(n29358) );
  AND U29214 ( .A(n29369), .B(n29370), .Z(n29367) );
  XOR U29215 ( .A(n29371), .B(n29365), .Z(n29369) );
  XNOR U29216 ( .A(n29318), .B(n29361), .Z(n29363) );
  XNOR U29217 ( .A(n29372), .B(n29373), .Z(n29318) );
  AND U29218 ( .A(n897), .B(n29325), .Z(n29373) );
  XOR U29219 ( .A(n29372), .B(n29323), .Z(n29325) );
  XOR U29220 ( .A(n29374), .B(n29375), .Z(n29361) );
  AND U29221 ( .A(n29376), .B(n29377), .Z(n29375) );
  XNOR U29222 ( .A(n29374), .B(n29333), .Z(n29377) );
  XOR U29223 ( .A(n29378), .B(n29370), .Z(n29333) );
  XNOR U29224 ( .A(n29379), .B(n29365), .Z(n29370) );
  XOR U29225 ( .A(n29380), .B(n29381), .Z(n29365) );
  AND U29226 ( .A(n29382), .B(n29383), .Z(n29381) );
  XOR U29227 ( .A(n29384), .B(n29380), .Z(n29382) );
  XNOR U29228 ( .A(n29385), .B(n29386), .Z(n29379) );
  AND U29229 ( .A(n29387), .B(n29388), .Z(n29386) );
  XOR U29230 ( .A(n29385), .B(n29389), .Z(n29387) );
  XNOR U29231 ( .A(n29371), .B(n29368), .Z(n29378) );
  AND U29232 ( .A(n29390), .B(n29391), .Z(n29368) );
  XOR U29233 ( .A(n29392), .B(n29393), .Z(n29371) );
  AND U29234 ( .A(n29394), .B(n29395), .Z(n29393) );
  XOR U29235 ( .A(n29392), .B(n29396), .Z(n29394) );
  XNOR U29236 ( .A(n29330), .B(n29374), .Z(n29376) );
  XNOR U29237 ( .A(n29397), .B(n29398), .Z(n29330) );
  AND U29238 ( .A(n897), .B(n29336), .Z(n29398) );
  XOR U29239 ( .A(n29397), .B(n29334), .Z(n29336) );
  XOR U29240 ( .A(n29399), .B(n29400), .Z(n29374) );
  AND U29241 ( .A(n29401), .B(n29402), .Z(n29400) );
  XNOR U29242 ( .A(n29399), .B(n29390), .Z(n29402) );
  IV U29243 ( .A(n29344), .Z(n29390) );
  XNOR U29244 ( .A(n29403), .B(n29383), .Z(n29344) );
  XNOR U29245 ( .A(n29404), .B(n29389), .Z(n29383) );
  XNOR U29246 ( .A(n29405), .B(n29406), .Z(n29389) );
  NOR U29247 ( .A(n29407), .B(n29408), .Z(n29406) );
  XOR U29248 ( .A(n29405), .B(n29409), .Z(n29407) );
  XNOR U29249 ( .A(n29388), .B(n29380), .Z(n29404) );
  XOR U29250 ( .A(n29410), .B(n29411), .Z(n29380) );
  AND U29251 ( .A(n29412), .B(n29413), .Z(n29411) );
  XOR U29252 ( .A(n29410), .B(n29414), .Z(n29412) );
  XNOR U29253 ( .A(n29415), .B(n29385), .Z(n29388) );
  XOR U29254 ( .A(n29416), .B(n29417), .Z(n29385) );
  AND U29255 ( .A(n29418), .B(n29419), .Z(n29417) );
  XNOR U29256 ( .A(n29420), .B(n29421), .Z(n29418) );
  IV U29257 ( .A(n29416), .Z(n29420) );
  XNOR U29258 ( .A(n29422), .B(n29423), .Z(n29415) );
  NOR U29259 ( .A(n29424), .B(n29425), .Z(n29423) );
  XNOR U29260 ( .A(n29422), .B(n29426), .Z(n29424) );
  XNOR U29261 ( .A(n29384), .B(n29391), .Z(n29403) );
  NOR U29262 ( .A(n29352), .B(n29427), .Z(n29391) );
  XOR U29263 ( .A(n29396), .B(n29395), .Z(n29384) );
  XNOR U29264 ( .A(n29428), .B(n29392), .Z(n29395) );
  XOR U29265 ( .A(n29429), .B(n29430), .Z(n29392) );
  AND U29266 ( .A(n29431), .B(n29432), .Z(n29430) );
  XNOR U29267 ( .A(n29433), .B(n29434), .Z(n29431) );
  IV U29268 ( .A(n29429), .Z(n29433) );
  XNOR U29269 ( .A(n29435), .B(n29436), .Z(n29428) );
  NOR U29270 ( .A(n29437), .B(n29438), .Z(n29436) );
  XNOR U29271 ( .A(n29435), .B(n29439), .Z(n29437) );
  XOR U29272 ( .A(n29440), .B(n29441), .Z(n29396) );
  NOR U29273 ( .A(n29442), .B(n29443), .Z(n29441) );
  XNOR U29274 ( .A(n29440), .B(n29444), .Z(n29442) );
  XNOR U29275 ( .A(n29341), .B(n29399), .Z(n29401) );
  XNOR U29276 ( .A(n29445), .B(n29446), .Z(n29341) );
  AND U29277 ( .A(n897), .B(n29348), .Z(n29446) );
  XOR U29278 ( .A(n29445), .B(n29346), .Z(n29348) );
  AND U29279 ( .A(n29349), .B(n29352), .Z(n29399) );
  XOR U29280 ( .A(n29447), .B(n29427), .Z(n29352) );
  XNOR U29281 ( .A(p_input[1248]), .B(p_input[2048]), .Z(n29427) );
  XNOR U29282 ( .A(n29414), .B(n29413), .Z(n29447) );
  XNOR U29283 ( .A(n29448), .B(n29421), .Z(n29413) );
  XNOR U29284 ( .A(n29409), .B(n29408), .Z(n29421) );
  XNOR U29285 ( .A(n29449), .B(n29405), .Z(n29408) );
  XNOR U29286 ( .A(p_input[1258]), .B(p_input[2058]), .Z(n29405) );
  XOR U29287 ( .A(p_input[1259]), .B(n16732), .Z(n29449) );
  XOR U29288 ( .A(p_input[1260]), .B(p_input[2060]), .Z(n29409) );
  XOR U29289 ( .A(n29419), .B(n29450), .Z(n29448) );
  IV U29290 ( .A(n29410), .Z(n29450) );
  XOR U29291 ( .A(p_input[1249]), .B(p_input[2049]), .Z(n29410) );
  XNOR U29292 ( .A(n29451), .B(n29426), .Z(n29419) );
  XNOR U29293 ( .A(p_input[1263]), .B(n16735), .Z(n29426) );
  XOR U29294 ( .A(n29416), .B(n29425), .Z(n29451) );
  XOR U29295 ( .A(n29452), .B(n29422), .Z(n29425) );
  XOR U29296 ( .A(p_input[1261]), .B(p_input[2061]), .Z(n29422) );
  XOR U29297 ( .A(p_input[1262]), .B(n16737), .Z(n29452) );
  XOR U29298 ( .A(p_input[1257]), .B(p_input[2057]), .Z(n29416) );
  XOR U29299 ( .A(n29434), .B(n29432), .Z(n29414) );
  XNOR U29300 ( .A(n29453), .B(n29439), .Z(n29432) );
  XOR U29301 ( .A(p_input[1256]), .B(p_input[2056]), .Z(n29439) );
  XOR U29302 ( .A(n29429), .B(n29438), .Z(n29453) );
  XOR U29303 ( .A(n29454), .B(n29435), .Z(n29438) );
  XOR U29304 ( .A(p_input[1254]), .B(p_input[2054]), .Z(n29435) );
  XOR U29305 ( .A(p_input[1255]), .B(n17722), .Z(n29454) );
  XOR U29306 ( .A(p_input[1250]), .B(p_input[2050]), .Z(n29429) );
  XNOR U29307 ( .A(n29444), .B(n29443), .Z(n29434) );
  XOR U29308 ( .A(n29455), .B(n29440), .Z(n29443) );
  XOR U29309 ( .A(p_input[1251]), .B(p_input[2051]), .Z(n29440) );
  XOR U29310 ( .A(p_input[1252]), .B(n17724), .Z(n29455) );
  XOR U29311 ( .A(p_input[1253]), .B(p_input[2053]), .Z(n29444) );
  XNOR U29312 ( .A(n29456), .B(n29457), .Z(n29349) );
  AND U29313 ( .A(n897), .B(n29458), .Z(n29457) );
  XNOR U29314 ( .A(n29459), .B(n29460), .Z(n897) );
  AND U29315 ( .A(n29461), .B(n29462), .Z(n29460) );
  XOR U29316 ( .A(n29459), .B(n29359), .Z(n29462) );
  XNOR U29317 ( .A(n29459), .B(n29313), .Z(n29461) );
  XOR U29318 ( .A(n29463), .B(n29464), .Z(n29459) );
  AND U29319 ( .A(n29465), .B(n29466), .Z(n29464) );
  XOR U29320 ( .A(n29463), .B(n29323), .Z(n29465) );
  XOR U29321 ( .A(n29467), .B(n29468), .Z(n29302) );
  AND U29322 ( .A(n901), .B(n29458), .Z(n29468) );
  XNOR U29323 ( .A(n29456), .B(n29467), .Z(n29458) );
  XNOR U29324 ( .A(n29469), .B(n29470), .Z(n901) );
  AND U29325 ( .A(n29471), .B(n29472), .Z(n29470) );
  XNOR U29326 ( .A(n29473), .B(n29469), .Z(n29472) );
  IV U29327 ( .A(n29359), .Z(n29473) );
  XNOR U29328 ( .A(n29474), .B(n29475), .Z(n29359) );
  AND U29329 ( .A(n904), .B(n29476), .Z(n29475) );
  XNOR U29330 ( .A(n29474), .B(n29477), .Z(n29476) );
  XNOR U29331 ( .A(n29313), .B(n29469), .Z(n29471) );
  XOR U29332 ( .A(n29478), .B(n29479), .Z(n29313) );
  AND U29333 ( .A(n912), .B(n29480), .Z(n29479) );
  XOR U29334 ( .A(n29463), .B(n29481), .Z(n29469) );
  AND U29335 ( .A(n29482), .B(n29466), .Z(n29481) );
  XNOR U29336 ( .A(n29372), .B(n29463), .Z(n29466) );
  XNOR U29337 ( .A(n29483), .B(n29484), .Z(n29372) );
  AND U29338 ( .A(n904), .B(n29485), .Z(n29484) );
  XOR U29339 ( .A(n29486), .B(n29483), .Z(n29485) );
  XNOR U29340 ( .A(n29487), .B(n29463), .Z(n29482) );
  IV U29341 ( .A(n29323), .Z(n29487) );
  XOR U29342 ( .A(n29488), .B(n29489), .Z(n29323) );
  AND U29343 ( .A(n912), .B(n29490), .Z(n29489) );
  XOR U29344 ( .A(n29491), .B(n29492), .Z(n29463) );
  AND U29345 ( .A(n29493), .B(n29494), .Z(n29492) );
  XNOR U29346 ( .A(n29397), .B(n29491), .Z(n29494) );
  XNOR U29347 ( .A(n29495), .B(n29496), .Z(n29397) );
  AND U29348 ( .A(n904), .B(n29497), .Z(n29496) );
  XNOR U29349 ( .A(n29498), .B(n29495), .Z(n29497) );
  XOR U29350 ( .A(n29491), .B(n29334), .Z(n29493) );
  XOR U29351 ( .A(n29499), .B(n29500), .Z(n29334) );
  AND U29352 ( .A(n912), .B(n29501), .Z(n29500) );
  XOR U29353 ( .A(n29502), .B(n29503), .Z(n29491) );
  AND U29354 ( .A(n29504), .B(n29505), .Z(n29503) );
  XNOR U29355 ( .A(n29502), .B(n29445), .Z(n29505) );
  XNOR U29356 ( .A(n29506), .B(n29507), .Z(n29445) );
  AND U29357 ( .A(n904), .B(n29508), .Z(n29507) );
  XOR U29358 ( .A(n29509), .B(n29506), .Z(n29508) );
  XNOR U29359 ( .A(n29510), .B(n29502), .Z(n29504) );
  IV U29360 ( .A(n29346), .Z(n29510) );
  XOR U29361 ( .A(n29511), .B(n29512), .Z(n29346) );
  AND U29362 ( .A(n912), .B(n29513), .Z(n29512) );
  AND U29363 ( .A(n29467), .B(n29456), .Z(n29502) );
  XNOR U29364 ( .A(n29514), .B(n29515), .Z(n29456) );
  AND U29365 ( .A(n904), .B(n29516), .Z(n29515) );
  XNOR U29366 ( .A(n29517), .B(n29514), .Z(n29516) );
  XNOR U29367 ( .A(n29518), .B(n29519), .Z(n904) );
  AND U29368 ( .A(n29520), .B(n29521), .Z(n29519) );
  XOR U29369 ( .A(n29477), .B(n29518), .Z(n29521) );
  AND U29370 ( .A(n29522), .B(n29523), .Z(n29477) );
  XOR U29371 ( .A(n29518), .B(n29474), .Z(n29520) );
  XNOR U29372 ( .A(n29524), .B(n29525), .Z(n29474) );
  AND U29373 ( .A(n908), .B(n29480), .Z(n29525) );
  XOR U29374 ( .A(n29478), .B(n29524), .Z(n29480) );
  XOR U29375 ( .A(n29526), .B(n29527), .Z(n29518) );
  AND U29376 ( .A(n29528), .B(n29529), .Z(n29527) );
  XNOR U29377 ( .A(n29526), .B(n29522), .Z(n29529) );
  IV U29378 ( .A(n29486), .Z(n29522) );
  XOR U29379 ( .A(n29530), .B(n29531), .Z(n29486) );
  XOR U29380 ( .A(n29532), .B(n29523), .Z(n29531) );
  AND U29381 ( .A(n29498), .B(n29533), .Z(n29523) );
  AND U29382 ( .A(n29534), .B(n29535), .Z(n29532) );
  XOR U29383 ( .A(n29536), .B(n29530), .Z(n29534) );
  XNOR U29384 ( .A(n29483), .B(n29526), .Z(n29528) );
  XNOR U29385 ( .A(n29537), .B(n29538), .Z(n29483) );
  AND U29386 ( .A(n908), .B(n29490), .Z(n29538) );
  XOR U29387 ( .A(n29537), .B(n29488), .Z(n29490) );
  XOR U29388 ( .A(n29539), .B(n29540), .Z(n29526) );
  AND U29389 ( .A(n29541), .B(n29542), .Z(n29540) );
  XNOR U29390 ( .A(n29539), .B(n29498), .Z(n29542) );
  XOR U29391 ( .A(n29543), .B(n29535), .Z(n29498) );
  XNOR U29392 ( .A(n29544), .B(n29530), .Z(n29535) );
  XOR U29393 ( .A(n29545), .B(n29546), .Z(n29530) );
  AND U29394 ( .A(n29547), .B(n29548), .Z(n29546) );
  XOR U29395 ( .A(n29549), .B(n29545), .Z(n29547) );
  XNOR U29396 ( .A(n29550), .B(n29551), .Z(n29544) );
  AND U29397 ( .A(n29552), .B(n29553), .Z(n29551) );
  XOR U29398 ( .A(n29550), .B(n29554), .Z(n29552) );
  XNOR U29399 ( .A(n29536), .B(n29533), .Z(n29543) );
  AND U29400 ( .A(n29555), .B(n29556), .Z(n29533) );
  XOR U29401 ( .A(n29557), .B(n29558), .Z(n29536) );
  AND U29402 ( .A(n29559), .B(n29560), .Z(n29558) );
  XOR U29403 ( .A(n29557), .B(n29561), .Z(n29559) );
  XNOR U29404 ( .A(n29495), .B(n29539), .Z(n29541) );
  XNOR U29405 ( .A(n29562), .B(n29563), .Z(n29495) );
  AND U29406 ( .A(n908), .B(n29501), .Z(n29563) );
  XOR U29407 ( .A(n29562), .B(n29499), .Z(n29501) );
  XOR U29408 ( .A(n29564), .B(n29565), .Z(n29539) );
  AND U29409 ( .A(n29566), .B(n29567), .Z(n29565) );
  XNOR U29410 ( .A(n29564), .B(n29555), .Z(n29567) );
  IV U29411 ( .A(n29509), .Z(n29555) );
  XNOR U29412 ( .A(n29568), .B(n29548), .Z(n29509) );
  XNOR U29413 ( .A(n29569), .B(n29554), .Z(n29548) );
  XNOR U29414 ( .A(n29570), .B(n29571), .Z(n29554) );
  NOR U29415 ( .A(n29572), .B(n29573), .Z(n29571) );
  XOR U29416 ( .A(n29570), .B(n29574), .Z(n29572) );
  XNOR U29417 ( .A(n29553), .B(n29545), .Z(n29569) );
  XOR U29418 ( .A(n29575), .B(n29576), .Z(n29545) );
  AND U29419 ( .A(n29577), .B(n29578), .Z(n29576) );
  XOR U29420 ( .A(n29575), .B(n29579), .Z(n29577) );
  XNOR U29421 ( .A(n29580), .B(n29550), .Z(n29553) );
  XOR U29422 ( .A(n29581), .B(n29582), .Z(n29550) );
  AND U29423 ( .A(n29583), .B(n29584), .Z(n29582) );
  XNOR U29424 ( .A(n29585), .B(n29586), .Z(n29583) );
  IV U29425 ( .A(n29581), .Z(n29585) );
  XNOR U29426 ( .A(n29587), .B(n29588), .Z(n29580) );
  NOR U29427 ( .A(n29589), .B(n29590), .Z(n29588) );
  XNOR U29428 ( .A(n29587), .B(n29591), .Z(n29589) );
  XNOR U29429 ( .A(n29549), .B(n29556), .Z(n29568) );
  NOR U29430 ( .A(n29517), .B(n29592), .Z(n29556) );
  XOR U29431 ( .A(n29561), .B(n29560), .Z(n29549) );
  XNOR U29432 ( .A(n29593), .B(n29557), .Z(n29560) );
  XOR U29433 ( .A(n29594), .B(n29595), .Z(n29557) );
  AND U29434 ( .A(n29596), .B(n29597), .Z(n29595) );
  XNOR U29435 ( .A(n29598), .B(n29599), .Z(n29596) );
  IV U29436 ( .A(n29594), .Z(n29598) );
  XNOR U29437 ( .A(n29600), .B(n29601), .Z(n29593) );
  NOR U29438 ( .A(n29602), .B(n29603), .Z(n29601) );
  XNOR U29439 ( .A(n29600), .B(n29604), .Z(n29602) );
  XOR U29440 ( .A(n29605), .B(n29606), .Z(n29561) );
  NOR U29441 ( .A(n29607), .B(n29608), .Z(n29606) );
  XNOR U29442 ( .A(n29605), .B(n29609), .Z(n29607) );
  XNOR U29443 ( .A(n29506), .B(n29564), .Z(n29566) );
  XNOR U29444 ( .A(n29610), .B(n29611), .Z(n29506) );
  AND U29445 ( .A(n908), .B(n29513), .Z(n29611) );
  XOR U29446 ( .A(n29610), .B(n29511), .Z(n29513) );
  AND U29447 ( .A(n29514), .B(n29517), .Z(n29564) );
  XOR U29448 ( .A(n29612), .B(n29592), .Z(n29517) );
  XNOR U29449 ( .A(p_input[1264]), .B(p_input[2048]), .Z(n29592) );
  XNOR U29450 ( .A(n29579), .B(n29578), .Z(n29612) );
  XNOR U29451 ( .A(n29613), .B(n29586), .Z(n29578) );
  XNOR U29452 ( .A(n29574), .B(n29573), .Z(n29586) );
  XNOR U29453 ( .A(n29614), .B(n29570), .Z(n29573) );
  XNOR U29454 ( .A(p_input[1274]), .B(p_input[2058]), .Z(n29570) );
  XOR U29455 ( .A(p_input[1275]), .B(n16732), .Z(n29614) );
  XOR U29456 ( .A(p_input[1276]), .B(p_input[2060]), .Z(n29574) );
  XOR U29457 ( .A(n29584), .B(n29615), .Z(n29613) );
  IV U29458 ( .A(n29575), .Z(n29615) );
  XOR U29459 ( .A(p_input[1265]), .B(p_input[2049]), .Z(n29575) );
  XNOR U29460 ( .A(n29616), .B(n29591), .Z(n29584) );
  XNOR U29461 ( .A(p_input[1279]), .B(n16735), .Z(n29591) );
  XOR U29462 ( .A(n29581), .B(n29590), .Z(n29616) );
  XOR U29463 ( .A(n29617), .B(n29587), .Z(n29590) );
  XOR U29464 ( .A(p_input[1277]), .B(p_input[2061]), .Z(n29587) );
  XOR U29465 ( .A(p_input[1278]), .B(n16737), .Z(n29617) );
  XOR U29466 ( .A(p_input[1273]), .B(p_input[2057]), .Z(n29581) );
  XOR U29467 ( .A(n29599), .B(n29597), .Z(n29579) );
  XNOR U29468 ( .A(n29618), .B(n29604), .Z(n29597) );
  XOR U29469 ( .A(p_input[1272]), .B(p_input[2056]), .Z(n29604) );
  XOR U29470 ( .A(n29594), .B(n29603), .Z(n29618) );
  XOR U29471 ( .A(n29619), .B(n29600), .Z(n29603) );
  XOR U29472 ( .A(p_input[1270]), .B(p_input[2054]), .Z(n29600) );
  XOR U29473 ( .A(p_input[1271]), .B(n17722), .Z(n29619) );
  XOR U29474 ( .A(p_input[1266]), .B(p_input[2050]), .Z(n29594) );
  XNOR U29475 ( .A(n29609), .B(n29608), .Z(n29599) );
  XOR U29476 ( .A(n29620), .B(n29605), .Z(n29608) );
  XOR U29477 ( .A(p_input[1267]), .B(p_input[2051]), .Z(n29605) );
  XOR U29478 ( .A(p_input[1268]), .B(n17724), .Z(n29620) );
  XOR U29479 ( .A(p_input[1269]), .B(p_input[2053]), .Z(n29609) );
  XNOR U29480 ( .A(n29621), .B(n29622), .Z(n29514) );
  AND U29481 ( .A(n908), .B(n29623), .Z(n29622) );
  XNOR U29482 ( .A(n29624), .B(n29625), .Z(n908) );
  AND U29483 ( .A(n29626), .B(n29627), .Z(n29625) );
  XOR U29484 ( .A(n29624), .B(n29524), .Z(n29627) );
  XNOR U29485 ( .A(n29624), .B(n29478), .Z(n29626) );
  XOR U29486 ( .A(n29628), .B(n29629), .Z(n29624) );
  AND U29487 ( .A(n29630), .B(n29631), .Z(n29629) );
  XOR U29488 ( .A(n29628), .B(n29488), .Z(n29630) );
  XOR U29489 ( .A(n29632), .B(n29633), .Z(n29467) );
  AND U29490 ( .A(n912), .B(n29623), .Z(n29633) );
  XNOR U29491 ( .A(n29621), .B(n29632), .Z(n29623) );
  XNOR U29492 ( .A(n29634), .B(n29635), .Z(n912) );
  AND U29493 ( .A(n29636), .B(n29637), .Z(n29635) );
  XNOR U29494 ( .A(n29638), .B(n29634), .Z(n29637) );
  IV U29495 ( .A(n29524), .Z(n29638) );
  XNOR U29496 ( .A(n29639), .B(n29640), .Z(n29524) );
  AND U29497 ( .A(n915), .B(n29641), .Z(n29640) );
  XNOR U29498 ( .A(n29639), .B(n29642), .Z(n29641) );
  XNOR U29499 ( .A(n29478), .B(n29634), .Z(n29636) );
  XOR U29500 ( .A(n29643), .B(n29644), .Z(n29478) );
  AND U29501 ( .A(n923), .B(n29645), .Z(n29644) );
  XOR U29502 ( .A(n29628), .B(n29646), .Z(n29634) );
  AND U29503 ( .A(n29647), .B(n29631), .Z(n29646) );
  XNOR U29504 ( .A(n29537), .B(n29628), .Z(n29631) );
  XNOR U29505 ( .A(n29648), .B(n29649), .Z(n29537) );
  AND U29506 ( .A(n915), .B(n29650), .Z(n29649) );
  XOR U29507 ( .A(n29651), .B(n29648), .Z(n29650) );
  XNOR U29508 ( .A(n29652), .B(n29628), .Z(n29647) );
  IV U29509 ( .A(n29488), .Z(n29652) );
  XOR U29510 ( .A(n29653), .B(n29654), .Z(n29488) );
  AND U29511 ( .A(n923), .B(n29655), .Z(n29654) );
  XOR U29512 ( .A(n29656), .B(n29657), .Z(n29628) );
  AND U29513 ( .A(n29658), .B(n29659), .Z(n29657) );
  XNOR U29514 ( .A(n29562), .B(n29656), .Z(n29659) );
  XNOR U29515 ( .A(n29660), .B(n29661), .Z(n29562) );
  AND U29516 ( .A(n915), .B(n29662), .Z(n29661) );
  XNOR U29517 ( .A(n29663), .B(n29660), .Z(n29662) );
  XOR U29518 ( .A(n29656), .B(n29499), .Z(n29658) );
  XOR U29519 ( .A(n29664), .B(n29665), .Z(n29499) );
  AND U29520 ( .A(n923), .B(n29666), .Z(n29665) );
  XOR U29521 ( .A(n29667), .B(n29668), .Z(n29656) );
  AND U29522 ( .A(n29669), .B(n29670), .Z(n29668) );
  XNOR U29523 ( .A(n29667), .B(n29610), .Z(n29670) );
  XNOR U29524 ( .A(n29671), .B(n29672), .Z(n29610) );
  AND U29525 ( .A(n915), .B(n29673), .Z(n29672) );
  XOR U29526 ( .A(n29674), .B(n29671), .Z(n29673) );
  XNOR U29527 ( .A(n29675), .B(n29667), .Z(n29669) );
  IV U29528 ( .A(n29511), .Z(n29675) );
  XOR U29529 ( .A(n29676), .B(n29677), .Z(n29511) );
  AND U29530 ( .A(n923), .B(n29678), .Z(n29677) );
  AND U29531 ( .A(n29632), .B(n29621), .Z(n29667) );
  XNOR U29532 ( .A(n29679), .B(n29680), .Z(n29621) );
  AND U29533 ( .A(n915), .B(n29681), .Z(n29680) );
  XNOR U29534 ( .A(n29682), .B(n29679), .Z(n29681) );
  XNOR U29535 ( .A(n29683), .B(n29684), .Z(n915) );
  AND U29536 ( .A(n29685), .B(n29686), .Z(n29684) );
  XOR U29537 ( .A(n29642), .B(n29683), .Z(n29686) );
  AND U29538 ( .A(n29687), .B(n29688), .Z(n29642) );
  XOR U29539 ( .A(n29683), .B(n29639), .Z(n29685) );
  XNOR U29540 ( .A(n29689), .B(n29690), .Z(n29639) );
  AND U29541 ( .A(n919), .B(n29645), .Z(n29690) );
  XOR U29542 ( .A(n29643), .B(n29689), .Z(n29645) );
  XOR U29543 ( .A(n29691), .B(n29692), .Z(n29683) );
  AND U29544 ( .A(n29693), .B(n29694), .Z(n29692) );
  XNOR U29545 ( .A(n29691), .B(n29687), .Z(n29694) );
  IV U29546 ( .A(n29651), .Z(n29687) );
  XOR U29547 ( .A(n29695), .B(n29696), .Z(n29651) );
  XOR U29548 ( .A(n29697), .B(n29688), .Z(n29696) );
  AND U29549 ( .A(n29663), .B(n29698), .Z(n29688) );
  AND U29550 ( .A(n29699), .B(n29700), .Z(n29697) );
  XOR U29551 ( .A(n29701), .B(n29695), .Z(n29699) );
  XNOR U29552 ( .A(n29648), .B(n29691), .Z(n29693) );
  XNOR U29553 ( .A(n29702), .B(n29703), .Z(n29648) );
  AND U29554 ( .A(n919), .B(n29655), .Z(n29703) );
  XOR U29555 ( .A(n29702), .B(n29653), .Z(n29655) );
  XOR U29556 ( .A(n29704), .B(n29705), .Z(n29691) );
  AND U29557 ( .A(n29706), .B(n29707), .Z(n29705) );
  XNOR U29558 ( .A(n29704), .B(n29663), .Z(n29707) );
  XOR U29559 ( .A(n29708), .B(n29700), .Z(n29663) );
  XNOR U29560 ( .A(n29709), .B(n29695), .Z(n29700) );
  XOR U29561 ( .A(n29710), .B(n29711), .Z(n29695) );
  AND U29562 ( .A(n29712), .B(n29713), .Z(n29711) );
  XOR U29563 ( .A(n29714), .B(n29710), .Z(n29712) );
  XNOR U29564 ( .A(n29715), .B(n29716), .Z(n29709) );
  AND U29565 ( .A(n29717), .B(n29718), .Z(n29716) );
  XOR U29566 ( .A(n29715), .B(n29719), .Z(n29717) );
  XNOR U29567 ( .A(n29701), .B(n29698), .Z(n29708) );
  AND U29568 ( .A(n29720), .B(n29721), .Z(n29698) );
  XOR U29569 ( .A(n29722), .B(n29723), .Z(n29701) );
  AND U29570 ( .A(n29724), .B(n29725), .Z(n29723) );
  XOR U29571 ( .A(n29722), .B(n29726), .Z(n29724) );
  XNOR U29572 ( .A(n29660), .B(n29704), .Z(n29706) );
  XNOR U29573 ( .A(n29727), .B(n29728), .Z(n29660) );
  AND U29574 ( .A(n919), .B(n29666), .Z(n29728) );
  XOR U29575 ( .A(n29727), .B(n29664), .Z(n29666) );
  XOR U29576 ( .A(n29729), .B(n29730), .Z(n29704) );
  AND U29577 ( .A(n29731), .B(n29732), .Z(n29730) );
  XNOR U29578 ( .A(n29729), .B(n29720), .Z(n29732) );
  IV U29579 ( .A(n29674), .Z(n29720) );
  XNOR U29580 ( .A(n29733), .B(n29713), .Z(n29674) );
  XNOR U29581 ( .A(n29734), .B(n29719), .Z(n29713) );
  XNOR U29582 ( .A(n29735), .B(n29736), .Z(n29719) );
  NOR U29583 ( .A(n29737), .B(n29738), .Z(n29736) );
  XOR U29584 ( .A(n29735), .B(n29739), .Z(n29737) );
  XNOR U29585 ( .A(n29718), .B(n29710), .Z(n29734) );
  XOR U29586 ( .A(n29740), .B(n29741), .Z(n29710) );
  AND U29587 ( .A(n29742), .B(n29743), .Z(n29741) );
  XOR U29588 ( .A(n29740), .B(n29744), .Z(n29742) );
  XNOR U29589 ( .A(n29745), .B(n29715), .Z(n29718) );
  XOR U29590 ( .A(n29746), .B(n29747), .Z(n29715) );
  AND U29591 ( .A(n29748), .B(n29749), .Z(n29747) );
  XNOR U29592 ( .A(n29750), .B(n29751), .Z(n29748) );
  IV U29593 ( .A(n29746), .Z(n29750) );
  XNOR U29594 ( .A(n29752), .B(n29753), .Z(n29745) );
  NOR U29595 ( .A(n29754), .B(n29755), .Z(n29753) );
  XNOR U29596 ( .A(n29752), .B(n29756), .Z(n29754) );
  XNOR U29597 ( .A(n29714), .B(n29721), .Z(n29733) );
  NOR U29598 ( .A(n29682), .B(n29757), .Z(n29721) );
  XOR U29599 ( .A(n29726), .B(n29725), .Z(n29714) );
  XNOR U29600 ( .A(n29758), .B(n29722), .Z(n29725) );
  XOR U29601 ( .A(n29759), .B(n29760), .Z(n29722) );
  AND U29602 ( .A(n29761), .B(n29762), .Z(n29760) );
  XNOR U29603 ( .A(n29763), .B(n29764), .Z(n29761) );
  IV U29604 ( .A(n29759), .Z(n29763) );
  XNOR U29605 ( .A(n29765), .B(n29766), .Z(n29758) );
  NOR U29606 ( .A(n29767), .B(n29768), .Z(n29766) );
  XNOR U29607 ( .A(n29765), .B(n29769), .Z(n29767) );
  XOR U29608 ( .A(n29770), .B(n29771), .Z(n29726) );
  NOR U29609 ( .A(n29772), .B(n29773), .Z(n29771) );
  XNOR U29610 ( .A(n29770), .B(n29774), .Z(n29772) );
  XNOR U29611 ( .A(n29671), .B(n29729), .Z(n29731) );
  XNOR U29612 ( .A(n29775), .B(n29776), .Z(n29671) );
  AND U29613 ( .A(n919), .B(n29678), .Z(n29776) );
  XOR U29614 ( .A(n29775), .B(n29676), .Z(n29678) );
  AND U29615 ( .A(n29679), .B(n29682), .Z(n29729) );
  XOR U29616 ( .A(n29777), .B(n29757), .Z(n29682) );
  XNOR U29617 ( .A(p_input[1280]), .B(p_input[2048]), .Z(n29757) );
  XNOR U29618 ( .A(n29744), .B(n29743), .Z(n29777) );
  XNOR U29619 ( .A(n29778), .B(n29751), .Z(n29743) );
  XNOR U29620 ( .A(n29739), .B(n29738), .Z(n29751) );
  XNOR U29621 ( .A(n29779), .B(n29735), .Z(n29738) );
  XNOR U29622 ( .A(p_input[1290]), .B(p_input[2058]), .Z(n29735) );
  XOR U29623 ( .A(p_input[1291]), .B(n16732), .Z(n29779) );
  XOR U29624 ( .A(p_input[1292]), .B(p_input[2060]), .Z(n29739) );
  XOR U29625 ( .A(n29749), .B(n29780), .Z(n29778) );
  IV U29626 ( .A(n29740), .Z(n29780) );
  XOR U29627 ( .A(p_input[1281]), .B(p_input[2049]), .Z(n29740) );
  XNOR U29628 ( .A(n29781), .B(n29756), .Z(n29749) );
  XNOR U29629 ( .A(p_input[1295]), .B(n16735), .Z(n29756) );
  XOR U29630 ( .A(n29746), .B(n29755), .Z(n29781) );
  XOR U29631 ( .A(n29782), .B(n29752), .Z(n29755) );
  XOR U29632 ( .A(p_input[1293]), .B(p_input[2061]), .Z(n29752) );
  XOR U29633 ( .A(p_input[1294]), .B(n16737), .Z(n29782) );
  XOR U29634 ( .A(p_input[1289]), .B(p_input[2057]), .Z(n29746) );
  XOR U29635 ( .A(n29764), .B(n29762), .Z(n29744) );
  XNOR U29636 ( .A(n29783), .B(n29769), .Z(n29762) );
  XOR U29637 ( .A(p_input[1288]), .B(p_input[2056]), .Z(n29769) );
  XOR U29638 ( .A(n29759), .B(n29768), .Z(n29783) );
  XOR U29639 ( .A(n29784), .B(n29765), .Z(n29768) );
  XOR U29640 ( .A(p_input[1286]), .B(p_input[2054]), .Z(n29765) );
  XOR U29641 ( .A(p_input[1287]), .B(n17722), .Z(n29784) );
  XOR U29642 ( .A(p_input[1282]), .B(p_input[2050]), .Z(n29759) );
  XNOR U29643 ( .A(n29774), .B(n29773), .Z(n29764) );
  XOR U29644 ( .A(n29785), .B(n29770), .Z(n29773) );
  XOR U29645 ( .A(p_input[1283]), .B(p_input[2051]), .Z(n29770) );
  XOR U29646 ( .A(p_input[1284]), .B(n17724), .Z(n29785) );
  XOR U29647 ( .A(p_input[1285]), .B(p_input[2053]), .Z(n29774) );
  XNOR U29648 ( .A(n29786), .B(n29787), .Z(n29679) );
  AND U29649 ( .A(n919), .B(n29788), .Z(n29787) );
  XNOR U29650 ( .A(n29789), .B(n29790), .Z(n919) );
  AND U29651 ( .A(n29791), .B(n29792), .Z(n29790) );
  XOR U29652 ( .A(n29789), .B(n29689), .Z(n29792) );
  XNOR U29653 ( .A(n29789), .B(n29643), .Z(n29791) );
  XOR U29654 ( .A(n29793), .B(n29794), .Z(n29789) );
  AND U29655 ( .A(n29795), .B(n29796), .Z(n29794) );
  XOR U29656 ( .A(n29793), .B(n29653), .Z(n29795) );
  XOR U29657 ( .A(n29797), .B(n29798), .Z(n29632) );
  AND U29658 ( .A(n923), .B(n29788), .Z(n29798) );
  XNOR U29659 ( .A(n29786), .B(n29797), .Z(n29788) );
  XNOR U29660 ( .A(n29799), .B(n29800), .Z(n923) );
  AND U29661 ( .A(n29801), .B(n29802), .Z(n29800) );
  XNOR U29662 ( .A(n29803), .B(n29799), .Z(n29802) );
  IV U29663 ( .A(n29689), .Z(n29803) );
  XNOR U29664 ( .A(n29804), .B(n29805), .Z(n29689) );
  AND U29665 ( .A(n926), .B(n29806), .Z(n29805) );
  XNOR U29666 ( .A(n29804), .B(n29807), .Z(n29806) );
  XNOR U29667 ( .A(n29643), .B(n29799), .Z(n29801) );
  XOR U29668 ( .A(n29808), .B(n29809), .Z(n29643) );
  AND U29669 ( .A(n934), .B(n29810), .Z(n29809) );
  XOR U29670 ( .A(n29793), .B(n29811), .Z(n29799) );
  AND U29671 ( .A(n29812), .B(n29796), .Z(n29811) );
  XNOR U29672 ( .A(n29702), .B(n29793), .Z(n29796) );
  XNOR U29673 ( .A(n29813), .B(n29814), .Z(n29702) );
  AND U29674 ( .A(n926), .B(n29815), .Z(n29814) );
  XOR U29675 ( .A(n29816), .B(n29813), .Z(n29815) );
  XNOR U29676 ( .A(n29817), .B(n29793), .Z(n29812) );
  IV U29677 ( .A(n29653), .Z(n29817) );
  XOR U29678 ( .A(n29818), .B(n29819), .Z(n29653) );
  AND U29679 ( .A(n934), .B(n29820), .Z(n29819) );
  XOR U29680 ( .A(n29821), .B(n29822), .Z(n29793) );
  AND U29681 ( .A(n29823), .B(n29824), .Z(n29822) );
  XNOR U29682 ( .A(n29727), .B(n29821), .Z(n29824) );
  XNOR U29683 ( .A(n29825), .B(n29826), .Z(n29727) );
  AND U29684 ( .A(n926), .B(n29827), .Z(n29826) );
  XNOR U29685 ( .A(n29828), .B(n29825), .Z(n29827) );
  XOR U29686 ( .A(n29821), .B(n29664), .Z(n29823) );
  XOR U29687 ( .A(n29829), .B(n29830), .Z(n29664) );
  AND U29688 ( .A(n934), .B(n29831), .Z(n29830) );
  XOR U29689 ( .A(n29832), .B(n29833), .Z(n29821) );
  AND U29690 ( .A(n29834), .B(n29835), .Z(n29833) );
  XNOR U29691 ( .A(n29832), .B(n29775), .Z(n29835) );
  XNOR U29692 ( .A(n29836), .B(n29837), .Z(n29775) );
  AND U29693 ( .A(n926), .B(n29838), .Z(n29837) );
  XOR U29694 ( .A(n29839), .B(n29836), .Z(n29838) );
  XNOR U29695 ( .A(n29840), .B(n29832), .Z(n29834) );
  IV U29696 ( .A(n29676), .Z(n29840) );
  XOR U29697 ( .A(n29841), .B(n29842), .Z(n29676) );
  AND U29698 ( .A(n934), .B(n29843), .Z(n29842) );
  AND U29699 ( .A(n29797), .B(n29786), .Z(n29832) );
  XNOR U29700 ( .A(n29844), .B(n29845), .Z(n29786) );
  AND U29701 ( .A(n926), .B(n29846), .Z(n29845) );
  XNOR U29702 ( .A(n29847), .B(n29844), .Z(n29846) );
  XNOR U29703 ( .A(n29848), .B(n29849), .Z(n926) );
  AND U29704 ( .A(n29850), .B(n29851), .Z(n29849) );
  XOR U29705 ( .A(n29807), .B(n29848), .Z(n29851) );
  AND U29706 ( .A(n29852), .B(n29853), .Z(n29807) );
  XOR U29707 ( .A(n29848), .B(n29804), .Z(n29850) );
  XNOR U29708 ( .A(n29854), .B(n29855), .Z(n29804) );
  AND U29709 ( .A(n930), .B(n29810), .Z(n29855) );
  XOR U29710 ( .A(n29808), .B(n29854), .Z(n29810) );
  XOR U29711 ( .A(n29856), .B(n29857), .Z(n29848) );
  AND U29712 ( .A(n29858), .B(n29859), .Z(n29857) );
  XNOR U29713 ( .A(n29856), .B(n29852), .Z(n29859) );
  IV U29714 ( .A(n29816), .Z(n29852) );
  XOR U29715 ( .A(n29860), .B(n29861), .Z(n29816) );
  XOR U29716 ( .A(n29862), .B(n29853), .Z(n29861) );
  AND U29717 ( .A(n29828), .B(n29863), .Z(n29853) );
  AND U29718 ( .A(n29864), .B(n29865), .Z(n29862) );
  XOR U29719 ( .A(n29866), .B(n29860), .Z(n29864) );
  XNOR U29720 ( .A(n29813), .B(n29856), .Z(n29858) );
  XNOR U29721 ( .A(n29867), .B(n29868), .Z(n29813) );
  AND U29722 ( .A(n930), .B(n29820), .Z(n29868) );
  XOR U29723 ( .A(n29867), .B(n29818), .Z(n29820) );
  XOR U29724 ( .A(n29869), .B(n29870), .Z(n29856) );
  AND U29725 ( .A(n29871), .B(n29872), .Z(n29870) );
  XNOR U29726 ( .A(n29869), .B(n29828), .Z(n29872) );
  XOR U29727 ( .A(n29873), .B(n29865), .Z(n29828) );
  XNOR U29728 ( .A(n29874), .B(n29860), .Z(n29865) );
  XOR U29729 ( .A(n29875), .B(n29876), .Z(n29860) );
  AND U29730 ( .A(n29877), .B(n29878), .Z(n29876) );
  XOR U29731 ( .A(n29879), .B(n29875), .Z(n29877) );
  XNOR U29732 ( .A(n29880), .B(n29881), .Z(n29874) );
  AND U29733 ( .A(n29882), .B(n29883), .Z(n29881) );
  XOR U29734 ( .A(n29880), .B(n29884), .Z(n29882) );
  XNOR U29735 ( .A(n29866), .B(n29863), .Z(n29873) );
  AND U29736 ( .A(n29885), .B(n29886), .Z(n29863) );
  XOR U29737 ( .A(n29887), .B(n29888), .Z(n29866) );
  AND U29738 ( .A(n29889), .B(n29890), .Z(n29888) );
  XOR U29739 ( .A(n29887), .B(n29891), .Z(n29889) );
  XNOR U29740 ( .A(n29825), .B(n29869), .Z(n29871) );
  XNOR U29741 ( .A(n29892), .B(n29893), .Z(n29825) );
  AND U29742 ( .A(n930), .B(n29831), .Z(n29893) );
  XOR U29743 ( .A(n29892), .B(n29829), .Z(n29831) );
  XOR U29744 ( .A(n29894), .B(n29895), .Z(n29869) );
  AND U29745 ( .A(n29896), .B(n29897), .Z(n29895) );
  XNOR U29746 ( .A(n29894), .B(n29885), .Z(n29897) );
  IV U29747 ( .A(n29839), .Z(n29885) );
  XNOR U29748 ( .A(n29898), .B(n29878), .Z(n29839) );
  XNOR U29749 ( .A(n29899), .B(n29884), .Z(n29878) );
  XNOR U29750 ( .A(n29900), .B(n29901), .Z(n29884) );
  NOR U29751 ( .A(n29902), .B(n29903), .Z(n29901) );
  XOR U29752 ( .A(n29900), .B(n29904), .Z(n29902) );
  XNOR U29753 ( .A(n29883), .B(n29875), .Z(n29899) );
  XOR U29754 ( .A(n29905), .B(n29906), .Z(n29875) );
  AND U29755 ( .A(n29907), .B(n29908), .Z(n29906) );
  XOR U29756 ( .A(n29905), .B(n29909), .Z(n29907) );
  XNOR U29757 ( .A(n29910), .B(n29880), .Z(n29883) );
  XOR U29758 ( .A(n29911), .B(n29912), .Z(n29880) );
  AND U29759 ( .A(n29913), .B(n29914), .Z(n29912) );
  XNOR U29760 ( .A(n29915), .B(n29916), .Z(n29913) );
  IV U29761 ( .A(n29911), .Z(n29915) );
  XNOR U29762 ( .A(n29917), .B(n29918), .Z(n29910) );
  NOR U29763 ( .A(n29919), .B(n29920), .Z(n29918) );
  XNOR U29764 ( .A(n29917), .B(n29921), .Z(n29919) );
  XNOR U29765 ( .A(n29879), .B(n29886), .Z(n29898) );
  NOR U29766 ( .A(n29847), .B(n29922), .Z(n29886) );
  XOR U29767 ( .A(n29891), .B(n29890), .Z(n29879) );
  XNOR U29768 ( .A(n29923), .B(n29887), .Z(n29890) );
  XOR U29769 ( .A(n29924), .B(n29925), .Z(n29887) );
  AND U29770 ( .A(n29926), .B(n29927), .Z(n29925) );
  XNOR U29771 ( .A(n29928), .B(n29929), .Z(n29926) );
  IV U29772 ( .A(n29924), .Z(n29928) );
  XNOR U29773 ( .A(n29930), .B(n29931), .Z(n29923) );
  NOR U29774 ( .A(n29932), .B(n29933), .Z(n29931) );
  XNOR U29775 ( .A(n29930), .B(n29934), .Z(n29932) );
  XOR U29776 ( .A(n29935), .B(n29936), .Z(n29891) );
  NOR U29777 ( .A(n29937), .B(n29938), .Z(n29936) );
  XNOR U29778 ( .A(n29935), .B(n29939), .Z(n29937) );
  XNOR U29779 ( .A(n29836), .B(n29894), .Z(n29896) );
  XNOR U29780 ( .A(n29940), .B(n29941), .Z(n29836) );
  AND U29781 ( .A(n930), .B(n29843), .Z(n29941) );
  XOR U29782 ( .A(n29940), .B(n29841), .Z(n29843) );
  AND U29783 ( .A(n29844), .B(n29847), .Z(n29894) );
  XOR U29784 ( .A(n29942), .B(n29922), .Z(n29847) );
  XNOR U29785 ( .A(p_input[1296]), .B(p_input[2048]), .Z(n29922) );
  XNOR U29786 ( .A(n29909), .B(n29908), .Z(n29942) );
  XNOR U29787 ( .A(n29943), .B(n29916), .Z(n29908) );
  XNOR U29788 ( .A(n29904), .B(n29903), .Z(n29916) );
  XNOR U29789 ( .A(n29944), .B(n29900), .Z(n29903) );
  XNOR U29790 ( .A(p_input[1306]), .B(p_input[2058]), .Z(n29900) );
  XOR U29791 ( .A(p_input[1307]), .B(n16732), .Z(n29944) );
  XOR U29792 ( .A(p_input[1308]), .B(p_input[2060]), .Z(n29904) );
  XOR U29793 ( .A(n29914), .B(n29945), .Z(n29943) );
  IV U29794 ( .A(n29905), .Z(n29945) );
  XOR U29795 ( .A(p_input[1297]), .B(p_input[2049]), .Z(n29905) );
  XNOR U29796 ( .A(n29946), .B(n29921), .Z(n29914) );
  XNOR U29797 ( .A(p_input[1311]), .B(n16735), .Z(n29921) );
  XOR U29798 ( .A(n29911), .B(n29920), .Z(n29946) );
  XOR U29799 ( .A(n29947), .B(n29917), .Z(n29920) );
  XOR U29800 ( .A(p_input[1309]), .B(p_input[2061]), .Z(n29917) );
  XOR U29801 ( .A(p_input[1310]), .B(n16737), .Z(n29947) );
  XOR U29802 ( .A(p_input[1305]), .B(p_input[2057]), .Z(n29911) );
  XOR U29803 ( .A(n29929), .B(n29927), .Z(n29909) );
  XNOR U29804 ( .A(n29948), .B(n29934), .Z(n29927) );
  XOR U29805 ( .A(p_input[1304]), .B(p_input[2056]), .Z(n29934) );
  XOR U29806 ( .A(n29924), .B(n29933), .Z(n29948) );
  XOR U29807 ( .A(n29949), .B(n29930), .Z(n29933) );
  XOR U29808 ( .A(p_input[1302]), .B(p_input[2054]), .Z(n29930) );
  XOR U29809 ( .A(p_input[1303]), .B(n17722), .Z(n29949) );
  XOR U29810 ( .A(p_input[1298]), .B(p_input[2050]), .Z(n29924) );
  XNOR U29811 ( .A(n29939), .B(n29938), .Z(n29929) );
  XOR U29812 ( .A(n29950), .B(n29935), .Z(n29938) );
  XOR U29813 ( .A(p_input[1299]), .B(p_input[2051]), .Z(n29935) );
  XOR U29814 ( .A(p_input[1300]), .B(n17724), .Z(n29950) );
  XOR U29815 ( .A(p_input[1301]), .B(p_input[2053]), .Z(n29939) );
  XNOR U29816 ( .A(n29951), .B(n29952), .Z(n29844) );
  AND U29817 ( .A(n930), .B(n29953), .Z(n29952) );
  XNOR U29818 ( .A(n29954), .B(n29955), .Z(n930) );
  AND U29819 ( .A(n29956), .B(n29957), .Z(n29955) );
  XOR U29820 ( .A(n29954), .B(n29854), .Z(n29957) );
  XNOR U29821 ( .A(n29954), .B(n29808), .Z(n29956) );
  XOR U29822 ( .A(n29958), .B(n29959), .Z(n29954) );
  AND U29823 ( .A(n29960), .B(n29961), .Z(n29959) );
  XOR U29824 ( .A(n29958), .B(n29818), .Z(n29960) );
  XOR U29825 ( .A(n29962), .B(n29963), .Z(n29797) );
  AND U29826 ( .A(n934), .B(n29953), .Z(n29963) );
  XNOR U29827 ( .A(n29951), .B(n29962), .Z(n29953) );
  XNOR U29828 ( .A(n29964), .B(n29965), .Z(n934) );
  AND U29829 ( .A(n29966), .B(n29967), .Z(n29965) );
  XNOR U29830 ( .A(n29968), .B(n29964), .Z(n29967) );
  IV U29831 ( .A(n29854), .Z(n29968) );
  XNOR U29832 ( .A(n29969), .B(n29970), .Z(n29854) );
  AND U29833 ( .A(n937), .B(n29971), .Z(n29970) );
  XNOR U29834 ( .A(n29969), .B(n29972), .Z(n29971) );
  XNOR U29835 ( .A(n29808), .B(n29964), .Z(n29966) );
  XOR U29836 ( .A(n29973), .B(n29974), .Z(n29808) );
  AND U29837 ( .A(n945), .B(n29975), .Z(n29974) );
  XOR U29838 ( .A(n29958), .B(n29976), .Z(n29964) );
  AND U29839 ( .A(n29977), .B(n29961), .Z(n29976) );
  XNOR U29840 ( .A(n29867), .B(n29958), .Z(n29961) );
  XNOR U29841 ( .A(n29978), .B(n29979), .Z(n29867) );
  AND U29842 ( .A(n937), .B(n29980), .Z(n29979) );
  XOR U29843 ( .A(n29981), .B(n29978), .Z(n29980) );
  XNOR U29844 ( .A(n29982), .B(n29958), .Z(n29977) );
  IV U29845 ( .A(n29818), .Z(n29982) );
  XOR U29846 ( .A(n29983), .B(n29984), .Z(n29818) );
  AND U29847 ( .A(n945), .B(n29985), .Z(n29984) );
  XOR U29848 ( .A(n29986), .B(n29987), .Z(n29958) );
  AND U29849 ( .A(n29988), .B(n29989), .Z(n29987) );
  XNOR U29850 ( .A(n29892), .B(n29986), .Z(n29989) );
  XNOR U29851 ( .A(n29990), .B(n29991), .Z(n29892) );
  AND U29852 ( .A(n937), .B(n29992), .Z(n29991) );
  XNOR U29853 ( .A(n29993), .B(n29990), .Z(n29992) );
  XOR U29854 ( .A(n29986), .B(n29829), .Z(n29988) );
  XOR U29855 ( .A(n29994), .B(n29995), .Z(n29829) );
  AND U29856 ( .A(n945), .B(n29996), .Z(n29995) );
  XOR U29857 ( .A(n29997), .B(n29998), .Z(n29986) );
  AND U29858 ( .A(n29999), .B(n30000), .Z(n29998) );
  XNOR U29859 ( .A(n29997), .B(n29940), .Z(n30000) );
  XNOR U29860 ( .A(n30001), .B(n30002), .Z(n29940) );
  AND U29861 ( .A(n937), .B(n30003), .Z(n30002) );
  XOR U29862 ( .A(n30004), .B(n30001), .Z(n30003) );
  XNOR U29863 ( .A(n30005), .B(n29997), .Z(n29999) );
  IV U29864 ( .A(n29841), .Z(n30005) );
  XOR U29865 ( .A(n30006), .B(n30007), .Z(n29841) );
  AND U29866 ( .A(n945), .B(n30008), .Z(n30007) );
  AND U29867 ( .A(n29962), .B(n29951), .Z(n29997) );
  XNOR U29868 ( .A(n30009), .B(n30010), .Z(n29951) );
  AND U29869 ( .A(n937), .B(n30011), .Z(n30010) );
  XNOR U29870 ( .A(n30012), .B(n30009), .Z(n30011) );
  XNOR U29871 ( .A(n30013), .B(n30014), .Z(n937) );
  AND U29872 ( .A(n30015), .B(n30016), .Z(n30014) );
  XOR U29873 ( .A(n29972), .B(n30013), .Z(n30016) );
  AND U29874 ( .A(n30017), .B(n30018), .Z(n29972) );
  XOR U29875 ( .A(n30013), .B(n29969), .Z(n30015) );
  XNOR U29876 ( .A(n30019), .B(n30020), .Z(n29969) );
  AND U29877 ( .A(n941), .B(n29975), .Z(n30020) );
  XOR U29878 ( .A(n29973), .B(n30019), .Z(n29975) );
  XOR U29879 ( .A(n30021), .B(n30022), .Z(n30013) );
  AND U29880 ( .A(n30023), .B(n30024), .Z(n30022) );
  XNOR U29881 ( .A(n30021), .B(n30017), .Z(n30024) );
  IV U29882 ( .A(n29981), .Z(n30017) );
  XOR U29883 ( .A(n30025), .B(n30026), .Z(n29981) );
  XOR U29884 ( .A(n30027), .B(n30018), .Z(n30026) );
  AND U29885 ( .A(n29993), .B(n30028), .Z(n30018) );
  AND U29886 ( .A(n30029), .B(n30030), .Z(n30027) );
  XOR U29887 ( .A(n30031), .B(n30025), .Z(n30029) );
  XNOR U29888 ( .A(n29978), .B(n30021), .Z(n30023) );
  XNOR U29889 ( .A(n30032), .B(n30033), .Z(n29978) );
  AND U29890 ( .A(n941), .B(n29985), .Z(n30033) );
  XOR U29891 ( .A(n30032), .B(n29983), .Z(n29985) );
  XOR U29892 ( .A(n30034), .B(n30035), .Z(n30021) );
  AND U29893 ( .A(n30036), .B(n30037), .Z(n30035) );
  XNOR U29894 ( .A(n30034), .B(n29993), .Z(n30037) );
  XOR U29895 ( .A(n30038), .B(n30030), .Z(n29993) );
  XNOR U29896 ( .A(n30039), .B(n30025), .Z(n30030) );
  XOR U29897 ( .A(n30040), .B(n30041), .Z(n30025) );
  AND U29898 ( .A(n30042), .B(n30043), .Z(n30041) );
  XOR U29899 ( .A(n30044), .B(n30040), .Z(n30042) );
  XNOR U29900 ( .A(n30045), .B(n30046), .Z(n30039) );
  AND U29901 ( .A(n30047), .B(n30048), .Z(n30046) );
  XOR U29902 ( .A(n30045), .B(n30049), .Z(n30047) );
  XNOR U29903 ( .A(n30031), .B(n30028), .Z(n30038) );
  AND U29904 ( .A(n30050), .B(n30051), .Z(n30028) );
  XOR U29905 ( .A(n30052), .B(n30053), .Z(n30031) );
  AND U29906 ( .A(n30054), .B(n30055), .Z(n30053) );
  XOR U29907 ( .A(n30052), .B(n30056), .Z(n30054) );
  XNOR U29908 ( .A(n29990), .B(n30034), .Z(n30036) );
  XNOR U29909 ( .A(n30057), .B(n30058), .Z(n29990) );
  AND U29910 ( .A(n941), .B(n29996), .Z(n30058) );
  XOR U29911 ( .A(n30057), .B(n29994), .Z(n29996) );
  XOR U29912 ( .A(n30059), .B(n30060), .Z(n30034) );
  AND U29913 ( .A(n30061), .B(n30062), .Z(n30060) );
  XNOR U29914 ( .A(n30059), .B(n30050), .Z(n30062) );
  IV U29915 ( .A(n30004), .Z(n30050) );
  XNOR U29916 ( .A(n30063), .B(n30043), .Z(n30004) );
  XNOR U29917 ( .A(n30064), .B(n30049), .Z(n30043) );
  XNOR U29918 ( .A(n30065), .B(n30066), .Z(n30049) );
  NOR U29919 ( .A(n30067), .B(n30068), .Z(n30066) );
  XOR U29920 ( .A(n30065), .B(n30069), .Z(n30067) );
  XNOR U29921 ( .A(n30048), .B(n30040), .Z(n30064) );
  XOR U29922 ( .A(n30070), .B(n30071), .Z(n30040) );
  AND U29923 ( .A(n30072), .B(n30073), .Z(n30071) );
  XOR U29924 ( .A(n30070), .B(n30074), .Z(n30072) );
  XNOR U29925 ( .A(n30075), .B(n30045), .Z(n30048) );
  XOR U29926 ( .A(n30076), .B(n30077), .Z(n30045) );
  AND U29927 ( .A(n30078), .B(n30079), .Z(n30077) );
  XNOR U29928 ( .A(n30080), .B(n30081), .Z(n30078) );
  IV U29929 ( .A(n30076), .Z(n30080) );
  XNOR U29930 ( .A(n30082), .B(n30083), .Z(n30075) );
  NOR U29931 ( .A(n30084), .B(n30085), .Z(n30083) );
  XNOR U29932 ( .A(n30082), .B(n30086), .Z(n30084) );
  XNOR U29933 ( .A(n30044), .B(n30051), .Z(n30063) );
  NOR U29934 ( .A(n30012), .B(n30087), .Z(n30051) );
  XOR U29935 ( .A(n30056), .B(n30055), .Z(n30044) );
  XNOR U29936 ( .A(n30088), .B(n30052), .Z(n30055) );
  XOR U29937 ( .A(n30089), .B(n30090), .Z(n30052) );
  AND U29938 ( .A(n30091), .B(n30092), .Z(n30090) );
  XNOR U29939 ( .A(n30093), .B(n30094), .Z(n30091) );
  IV U29940 ( .A(n30089), .Z(n30093) );
  XNOR U29941 ( .A(n30095), .B(n30096), .Z(n30088) );
  NOR U29942 ( .A(n30097), .B(n30098), .Z(n30096) );
  XNOR U29943 ( .A(n30095), .B(n30099), .Z(n30097) );
  XOR U29944 ( .A(n30100), .B(n30101), .Z(n30056) );
  NOR U29945 ( .A(n30102), .B(n30103), .Z(n30101) );
  XNOR U29946 ( .A(n30100), .B(n30104), .Z(n30102) );
  XNOR U29947 ( .A(n30001), .B(n30059), .Z(n30061) );
  XNOR U29948 ( .A(n30105), .B(n30106), .Z(n30001) );
  AND U29949 ( .A(n941), .B(n30008), .Z(n30106) );
  XOR U29950 ( .A(n30105), .B(n30006), .Z(n30008) );
  AND U29951 ( .A(n30009), .B(n30012), .Z(n30059) );
  XOR U29952 ( .A(n30107), .B(n30087), .Z(n30012) );
  XNOR U29953 ( .A(p_input[1312]), .B(p_input[2048]), .Z(n30087) );
  XNOR U29954 ( .A(n30074), .B(n30073), .Z(n30107) );
  XNOR U29955 ( .A(n30108), .B(n30081), .Z(n30073) );
  XNOR U29956 ( .A(n30069), .B(n30068), .Z(n30081) );
  XNOR U29957 ( .A(n30109), .B(n30065), .Z(n30068) );
  XNOR U29958 ( .A(p_input[1322]), .B(p_input[2058]), .Z(n30065) );
  XOR U29959 ( .A(p_input[1323]), .B(n16732), .Z(n30109) );
  XOR U29960 ( .A(p_input[1324]), .B(p_input[2060]), .Z(n30069) );
  XOR U29961 ( .A(n30079), .B(n30110), .Z(n30108) );
  IV U29962 ( .A(n30070), .Z(n30110) );
  XOR U29963 ( .A(p_input[1313]), .B(p_input[2049]), .Z(n30070) );
  XNOR U29964 ( .A(n30111), .B(n30086), .Z(n30079) );
  XNOR U29965 ( .A(p_input[1327]), .B(n16735), .Z(n30086) );
  XOR U29966 ( .A(n30076), .B(n30085), .Z(n30111) );
  XOR U29967 ( .A(n30112), .B(n30082), .Z(n30085) );
  XOR U29968 ( .A(p_input[1325]), .B(p_input[2061]), .Z(n30082) );
  XOR U29969 ( .A(p_input[1326]), .B(n16737), .Z(n30112) );
  XOR U29970 ( .A(p_input[1321]), .B(p_input[2057]), .Z(n30076) );
  XOR U29971 ( .A(n30094), .B(n30092), .Z(n30074) );
  XNOR U29972 ( .A(n30113), .B(n30099), .Z(n30092) );
  XOR U29973 ( .A(p_input[1320]), .B(p_input[2056]), .Z(n30099) );
  XOR U29974 ( .A(n30089), .B(n30098), .Z(n30113) );
  XOR U29975 ( .A(n30114), .B(n30095), .Z(n30098) );
  XOR U29976 ( .A(p_input[1318]), .B(p_input[2054]), .Z(n30095) );
  XOR U29977 ( .A(p_input[1319]), .B(n17722), .Z(n30114) );
  XOR U29978 ( .A(p_input[1314]), .B(p_input[2050]), .Z(n30089) );
  XNOR U29979 ( .A(n30104), .B(n30103), .Z(n30094) );
  XOR U29980 ( .A(n30115), .B(n30100), .Z(n30103) );
  XOR U29981 ( .A(p_input[1315]), .B(p_input[2051]), .Z(n30100) );
  XOR U29982 ( .A(p_input[1316]), .B(n17724), .Z(n30115) );
  XOR U29983 ( .A(p_input[1317]), .B(p_input[2053]), .Z(n30104) );
  XNOR U29984 ( .A(n30116), .B(n30117), .Z(n30009) );
  AND U29985 ( .A(n941), .B(n30118), .Z(n30117) );
  XNOR U29986 ( .A(n30119), .B(n30120), .Z(n941) );
  AND U29987 ( .A(n30121), .B(n30122), .Z(n30120) );
  XOR U29988 ( .A(n30119), .B(n30019), .Z(n30122) );
  XNOR U29989 ( .A(n30119), .B(n29973), .Z(n30121) );
  XOR U29990 ( .A(n30123), .B(n30124), .Z(n30119) );
  AND U29991 ( .A(n30125), .B(n30126), .Z(n30124) );
  XOR U29992 ( .A(n30123), .B(n29983), .Z(n30125) );
  XOR U29993 ( .A(n30127), .B(n30128), .Z(n29962) );
  AND U29994 ( .A(n945), .B(n30118), .Z(n30128) );
  XNOR U29995 ( .A(n30116), .B(n30127), .Z(n30118) );
  XNOR U29996 ( .A(n30129), .B(n30130), .Z(n945) );
  AND U29997 ( .A(n30131), .B(n30132), .Z(n30130) );
  XNOR U29998 ( .A(n30133), .B(n30129), .Z(n30132) );
  IV U29999 ( .A(n30019), .Z(n30133) );
  XNOR U30000 ( .A(n30134), .B(n30135), .Z(n30019) );
  AND U30001 ( .A(n948), .B(n30136), .Z(n30135) );
  XNOR U30002 ( .A(n30134), .B(n30137), .Z(n30136) );
  XNOR U30003 ( .A(n29973), .B(n30129), .Z(n30131) );
  XOR U30004 ( .A(n30138), .B(n30139), .Z(n29973) );
  AND U30005 ( .A(n956), .B(n30140), .Z(n30139) );
  XOR U30006 ( .A(n30123), .B(n30141), .Z(n30129) );
  AND U30007 ( .A(n30142), .B(n30126), .Z(n30141) );
  XNOR U30008 ( .A(n30032), .B(n30123), .Z(n30126) );
  XNOR U30009 ( .A(n30143), .B(n30144), .Z(n30032) );
  AND U30010 ( .A(n948), .B(n30145), .Z(n30144) );
  XOR U30011 ( .A(n30146), .B(n30143), .Z(n30145) );
  XNOR U30012 ( .A(n30147), .B(n30123), .Z(n30142) );
  IV U30013 ( .A(n29983), .Z(n30147) );
  XOR U30014 ( .A(n30148), .B(n30149), .Z(n29983) );
  AND U30015 ( .A(n956), .B(n30150), .Z(n30149) );
  XOR U30016 ( .A(n30151), .B(n30152), .Z(n30123) );
  AND U30017 ( .A(n30153), .B(n30154), .Z(n30152) );
  XNOR U30018 ( .A(n30057), .B(n30151), .Z(n30154) );
  XNOR U30019 ( .A(n30155), .B(n30156), .Z(n30057) );
  AND U30020 ( .A(n948), .B(n30157), .Z(n30156) );
  XNOR U30021 ( .A(n30158), .B(n30155), .Z(n30157) );
  XOR U30022 ( .A(n30151), .B(n29994), .Z(n30153) );
  XOR U30023 ( .A(n30159), .B(n30160), .Z(n29994) );
  AND U30024 ( .A(n956), .B(n30161), .Z(n30160) );
  XOR U30025 ( .A(n30162), .B(n30163), .Z(n30151) );
  AND U30026 ( .A(n30164), .B(n30165), .Z(n30163) );
  XNOR U30027 ( .A(n30162), .B(n30105), .Z(n30165) );
  XNOR U30028 ( .A(n30166), .B(n30167), .Z(n30105) );
  AND U30029 ( .A(n948), .B(n30168), .Z(n30167) );
  XOR U30030 ( .A(n30169), .B(n30166), .Z(n30168) );
  XNOR U30031 ( .A(n30170), .B(n30162), .Z(n30164) );
  IV U30032 ( .A(n30006), .Z(n30170) );
  XOR U30033 ( .A(n30171), .B(n30172), .Z(n30006) );
  AND U30034 ( .A(n956), .B(n30173), .Z(n30172) );
  AND U30035 ( .A(n30127), .B(n30116), .Z(n30162) );
  XNOR U30036 ( .A(n30174), .B(n30175), .Z(n30116) );
  AND U30037 ( .A(n948), .B(n30176), .Z(n30175) );
  XNOR U30038 ( .A(n30177), .B(n30174), .Z(n30176) );
  XNOR U30039 ( .A(n30178), .B(n30179), .Z(n948) );
  AND U30040 ( .A(n30180), .B(n30181), .Z(n30179) );
  XOR U30041 ( .A(n30137), .B(n30178), .Z(n30181) );
  AND U30042 ( .A(n30182), .B(n30183), .Z(n30137) );
  XOR U30043 ( .A(n30178), .B(n30134), .Z(n30180) );
  XNOR U30044 ( .A(n30184), .B(n30185), .Z(n30134) );
  AND U30045 ( .A(n952), .B(n30140), .Z(n30185) );
  XOR U30046 ( .A(n30138), .B(n30184), .Z(n30140) );
  XOR U30047 ( .A(n30186), .B(n30187), .Z(n30178) );
  AND U30048 ( .A(n30188), .B(n30189), .Z(n30187) );
  XNOR U30049 ( .A(n30186), .B(n30182), .Z(n30189) );
  IV U30050 ( .A(n30146), .Z(n30182) );
  XOR U30051 ( .A(n30190), .B(n30191), .Z(n30146) );
  XOR U30052 ( .A(n30192), .B(n30183), .Z(n30191) );
  AND U30053 ( .A(n30158), .B(n30193), .Z(n30183) );
  AND U30054 ( .A(n30194), .B(n30195), .Z(n30192) );
  XOR U30055 ( .A(n30196), .B(n30190), .Z(n30194) );
  XNOR U30056 ( .A(n30143), .B(n30186), .Z(n30188) );
  XNOR U30057 ( .A(n30197), .B(n30198), .Z(n30143) );
  AND U30058 ( .A(n952), .B(n30150), .Z(n30198) );
  XOR U30059 ( .A(n30197), .B(n30148), .Z(n30150) );
  XOR U30060 ( .A(n30199), .B(n30200), .Z(n30186) );
  AND U30061 ( .A(n30201), .B(n30202), .Z(n30200) );
  XNOR U30062 ( .A(n30199), .B(n30158), .Z(n30202) );
  XOR U30063 ( .A(n30203), .B(n30195), .Z(n30158) );
  XNOR U30064 ( .A(n30204), .B(n30190), .Z(n30195) );
  XOR U30065 ( .A(n30205), .B(n30206), .Z(n30190) );
  AND U30066 ( .A(n30207), .B(n30208), .Z(n30206) );
  XOR U30067 ( .A(n30209), .B(n30205), .Z(n30207) );
  XNOR U30068 ( .A(n30210), .B(n30211), .Z(n30204) );
  AND U30069 ( .A(n30212), .B(n30213), .Z(n30211) );
  XOR U30070 ( .A(n30210), .B(n30214), .Z(n30212) );
  XNOR U30071 ( .A(n30196), .B(n30193), .Z(n30203) );
  AND U30072 ( .A(n30215), .B(n30216), .Z(n30193) );
  XOR U30073 ( .A(n30217), .B(n30218), .Z(n30196) );
  AND U30074 ( .A(n30219), .B(n30220), .Z(n30218) );
  XOR U30075 ( .A(n30217), .B(n30221), .Z(n30219) );
  XNOR U30076 ( .A(n30155), .B(n30199), .Z(n30201) );
  XNOR U30077 ( .A(n30222), .B(n30223), .Z(n30155) );
  AND U30078 ( .A(n952), .B(n30161), .Z(n30223) );
  XOR U30079 ( .A(n30222), .B(n30159), .Z(n30161) );
  XOR U30080 ( .A(n30224), .B(n30225), .Z(n30199) );
  AND U30081 ( .A(n30226), .B(n30227), .Z(n30225) );
  XNOR U30082 ( .A(n30224), .B(n30215), .Z(n30227) );
  IV U30083 ( .A(n30169), .Z(n30215) );
  XNOR U30084 ( .A(n30228), .B(n30208), .Z(n30169) );
  XNOR U30085 ( .A(n30229), .B(n30214), .Z(n30208) );
  XNOR U30086 ( .A(n30230), .B(n30231), .Z(n30214) );
  NOR U30087 ( .A(n30232), .B(n30233), .Z(n30231) );
  XOR U30088 ( .A(n30230), .B(n30234), .Z(n30232) );
  XNOR U30089 ( .A(n30213), .B(n30205), .Z(n30229) );
  XOR U30090 ( .A(n30235), .B(n30236), .Z(n30205) );
  AND U30091 ( .A(n30237), .B(n30238), .Z(n30236) );
  XOR U30092 ( .A(n30235), .B(n30239), .Z(n30237) );
  XNOR U30093 ( .A(n30240), .B(n30210), .Z(n30213) );
  XOR U30094 ( .A(n30241), .B(n30242), .Z(n30210) );
  AND U30095 ( .A(n30243), .B(n30244), .Z(n30242) );
  XNOR U30096 ( .A(n30245), .B(n30246), .Z(n30243) );
  IV U30097 ( .A(n30241), .Z(n30245) );
  XNOR U30098 ( .A(n30247), .B(n30248), .Z(n30240) );
  NOR U30099 ( .A(n30249), .B(n30250), .Z(n30248) );
  XNOR U30100 ( .A(n30247), .B(n30251), .Z(n30249) );
  XNOR U30101 ( .A(n30209), .B(n30216), .Z(n30228) );
  NOR U30102 ( .A(n30177), .B(n30252), .Z(n30216) );
  XOR U30103 ( .A(n30221), .B(n30220), .Z(n30209) );
  XNOR U30104 ( .A(n30253), .B(n30217), .Z(n30220) );
  XOR U30105 ( .A(n30254), .B(n30255), .Z(n30217) );
  AND U30106 ( .A(n30256), .B(n30257), .Z(n30255) );
  XNOR U30107 ( .A(n30258), .B(n30259), .Z(n30256) );
  IV U30108 ( .A(n30254), .Z(n30258) );
  XNOR U30109 ( .A(n30260), .B(n30261), .Z(n30253) );
  NOR U30110 ( .A(n30262), .B(n30263), .Z(n30261) );
  XNOR U30111 ( .A(n30260), .B(n30264), .Z(n30262) );
  XOR U30112 ( .A(n30265), .B(n30266), .Z(n30221) );
  NOR U30113 ( .A(n30267), .B(n30268), .Z(n30266) );
  XNOR U30114 ( .A(n30265), .B(n30269), .Z(n30267) );
  XNOR U30115 ( .A(n30166), .B(n30224), .Z(n30226) );
  XNOR U30116 ( .A(n30270), .B(n30271), .Z(n30166) );
  AND U30117 ( .A(n952), .B(n30173), .Z(n30271) );
  XOR U30118 ( .A(n30270), .B(n30171), .Z(n30173) );
  AND U30119 ( .A(n30174), .B(n30177), .Z(n30224) );
  XOR U30120 ( .A(n30272), .B(n30252), .Z(n30177) );
  XNOR U30121 ( .A(p_input[1328]), .B(p_input[2048]), .Z(n30252) );
  XNOR U30122 ( .A(n30239), .B(n30238), .Z(n30272) );
  XNOR U30123 ( .A(n30273), .B(n30246), .Z(n30238) );
  XNOR U30124 ( .A(n30234), .B(n30233), .Z(n30246) );
  XNOR U30125 ( .A(n30274), .B(n30230), .Z(n30233) );
  XNOR U30126 ( .A(p_input[1338]), .B(p_input[2058]), .Z(n30230) );
  XOR U30127 ( .A(p_input[1339]), .B(n16732), .Z(n30274) );
  XOR U30128 ( .A(p_input[1340]), .B(p_input[2060]), .Z(n30234) );
  XOR U30129 ( .A(n30244), .B(n30275), .Z(n30273) );
  IV U30130 ( .A(n30235), .Z(n30275) );
  XOR U30131 ( .A(p_input[1329]), .B(p_input[2049]), .Z(n30235) );
  XNOR U30132 ( .A(n30276), .B(n30251), .Z(n30244) );
  XNOR U30133 ( .A(p_input[1343]), .B(n16735), .Z(n30251) );
  XOR U30134 ( .A(n30241), .B(n30250), .Z(n30276) );
  XOR U30135 ( .A(n30277), .B(n30247), .Z(n30250) );
  XOR U30136 ( .A(p_input[1341]), .B(p_input[2061]), .Z(n30247) );
  XOR U30137 ( .A(p_input[1342]), .B(n16737), .Z(n30277) );
  XOR U30138 ( .A(p_input[1337]), .B(p_input[2057]), .Z(n30241) );
  XOR U30139 ( .A(n30259), .B(n30257), .Z(n30239) );
  XNOR U30140 ( .A(n30278), .B(n30264), .Z(n30257) );
  XOR U30141 ( .A(p_input[1336]), .B(p_input[2056]), .Z(n30264) );
  XOR U30142 ( .A(n30254), .B(n30263), .Z(n30278) );
  XOR U30143 ( .A(n30279), .B(n30260), .Z(n30263) );
  XOR U30144 ( .A(p_input[1334]), .B(p_input[2054]), .Z(n30260) );
  XOR U30145 ( .A(p_input[1335]), .B(n17722), .Z(n30279) );
  XOR U30146 ( .A(p_input[1330]), .B(p_input[2050]), .Z(n30254) );
  XNOR U30147 ( .A(n30269), .B(n30268), .Z(n30259) );
  XOR U30148 ( .A(n30280), .B(n30265), .Z(n30268) );
  XOR U30149 ( .A(p_input[1331]), .B(p_input[2051]), .Z(n30265) );
  XOR U30150 ( .A(p_input[1332]), .B(n17724), .Z(n30280) );
  XOR U30151 ( .A(p_input[1333]), .B(p_input[2053]), .Z(n30269) );
  XNOR U30152 ( .A(n30281), .B(n30282), .Z(n30174) );
  AND U30153 ( .A(n952), .B(n30283), .Z(n30282) );
  XNOR U30154 ( .A(n30284), .B(n30285), .Z(n952) );
  AND U30155 ( .A(n30286), .B(n30287), .Z(n30285) );
  XOR U30156 ( .A(n30284), .B(n30184), .Z(n30287) );
  XNOR U30157 ( .A(n30284), .B(n30138), .Z(n30286) );
  XOR U30158 ( .A(n30288), .B(n30289), .Z(n30284) );
  AND U30159 ( .A(n30290), .B(n30291), .Z(n30289) );
  XOR U30160 ( .A(n30288), .B(n30148), .Z(n30290) );
  XOR U30161 ( .A(n30292), .B(n30293), .Z(n30127) );
  AND U30162 ( .A(n956), .B(n30283), .Z(n30293) );
  XNOR U30163 ( .A(n30281), .B(n30292), .Z(n30283) );
  XNOR U30164 ( .A(n30294), .B(n30295), .Z(n956) );
  AND U30165 ( .A(n30296), .B(n30297), .Z(n30295) );
  XNOR U30166 ( .A(n30298), .B(n30294), .Z(n30297) );
  IV U30167 ( .A(n30184), .Z(n30298) );
  XNOR U30168 ( .A(n30299), .B(n30300), .Z(n30184) );
  AND U30169 ( .A(n959), .B(n30301), .Z(n30300) );
  XNOR U30170 ( .A(n30299), .B(n30302), .Z(n30301) );
  XNOR U30171 ( .A(n30138), .B(n30294), .Z(n30296) );
  XOR U30172 ( .A(n30303), .B(n30304), .Z(n30138) );
  AND U30173 ( .A(n967), .B(n30305), .Z(n30304) );
  XOR U30174 ( .A(n30288), .B(n30306), .Z(n30294) );
  AND U30175 ( .A(n30307), .B(n30291), .Z(n30306) );
  XNOR U30176 ( .A(n30197), .B(n30288), .Z(n30291) );
  XNOR U30177 ( .A(n30308), .B(n30309), .Z(n30197) );
  AND U30178 ( .A(n959), .B(n30310), .Z(n30309) );
  XOR U30179 ( .A(n30311), .B(n30308), .Z(n30310) );
  XNOR U30180 ( .A(n30312), .B(n30288), .Z(n30307) );
  IV U30181 ( .A(n30148), .Z(n30312) );
  XOR U30182 ( .A(n30313), .B(n30314), .Z(n30148) );
  AND U30183 ( .A(n967), .B(n30315), .Z(n30314) );
  XOR U30184 ( .A(n30316), .B(n30317), .Z(n30288) );
  AND U30185 ( .A(n30318), .B(n30319), .Z(n30317) );
  XNOR U30186 ( .A(n30222), .B(n30316), .Z(n30319) );
  XNOR U30187 ( .A(n30320), .B(n30321), .Z(n30222) );
  AND U30188 ( .A(n959), .B(n30322), .Z(n30321) );
  XNOR U30189 ( .A(n30323), .B(n30320), .Z(n30322) );
  XOR U30190 ( .A(n30316), .B(n30159), .Z(n30318) );
  XOR U30191 ( .A(n30324), .B(n30325), .Z(n30159) );
  AND U30192 ( .A(n967), .B(n30326), .Z(n30325) );
  XOR U30193 ( .A(n30327), .B(n30328), .Z(n30316) );
  AND U30194 ( .A(n30329), .B(n30330), .Z(n30328) );
  XNOR U30195 ( .A(n30327), .B(n30270), .Z(n30330) );
  XNOR U30196 ( .A(n30331), .B(n30332), .Z(n30270) );
  AND U30197 ( .A(n959), .B(n30333), .Z(n30332) );
  XOR U30198 ( .A(n30334), .B(n30331), .Z(n30333) );
  XNOR U30199 ( .A(n30335), .B(n30327), .Z(n30329) );
  IV U30200 ( .A(n30171), .Z(n30335) );
  XOR U30201 ( .A(n30336), .B(n30337), .Z(n30171) );
  AND U30202 ( .A(n967), .B(n30338), .Z(n30337) );
  AND U30203 ( .A(n30292), .B(n30281), .Z(n30327) );
  XNOR U30204 ( .A(n30339), .B(n30340), .Z(n30281) );
  AND U30205 ( .A(n959), .B(n30341), .Z(n30340) );
  XNOR U30206 ( .A(n30342), .B(n30339), .Z(n30341) );
  XNOR U30207 ( .A(n30343), .B(n30344), .Z(n959) );
  AND U30208 ( .A(n30345), .B(n30346), .Z(n30344) );
  XOR U30209 ( .A(n30302), .B(n30343), .Z(n30346) );
  AND U30210 ( .A(n30347), .B(n30348), .Z(n30302) );
  XOR U30211 ( .A(n30343), .B(n30299), .Z(n30345) );
  XNOR U30212 ( .A(n30349), .B(n30350), .Z(n30299) );
  AND U30213 ( .A(n963), .B(n30305), .Z(n30350) );
  XOR U30214 ( .A(n30303), .B(n30349), .Z(n30305) );
  XOR U30215 ( .A(n30351), .B(n30352), .Z(n30343) );
  AND U30216 ( .A(n30353), .B(n30354), .Z(n30352) );
  XNOR U30217 ( .A(n30351), .B(n30347), .Z(n30354) );
  IV U30218 ( .A(n30311), .Z(n30347) );
  XOR U30219 ( .A(n30355), .B(n30356), .Z(n30311) );
  XOR U30220 ( .A(n30357), .B(n30348), .Z(n30356) );
  AND U30221 ( .A(n30323), .B(n30358), .Z(n30348) );
  AND U30222 ( .A(n30359), .B(n30360), .Z(n30357) );
  XOR U30223 ( .A(n30361), .B(n30355), .Z(n30359) );
  XNOR U30224 ( .A(n30308), .B(n30351), .Z(n30353) );
  XNOR U30225 ( .A(n30362), .B(n30363), .Z(n30308) );
  AND U30226 ( .A(n963), .B(n30315), .Z(n30363) );
  XOR U30227 ( .A(n30362), .B(n30313), .Z(n30315) );
  XOR U30228 ( .A(n30364), .B(n30365), .Z(n30351) );
  AND U30229 ( .A(n30366), .B(n30367), .Z(n30365) );
  XNOR U30230 ( .A(n30364), .B(n30323), .Z(n30367) );
  XOR U30231 ( .A(n30368), .B(n30360), .Z(n30323) );
  XNOR U30232 ( .A(n30369), .B(n30355), .Z(n30360) );
  XOR U30233 ( .A(n30370), .B(n30371), .Z(n30355) );
  AND U30234 ( .A(n30372), .B(n30373), .Z(n30371) );
  XOR U30235 ( .A(n30374), .B(n30370), .Z(n30372) );
  XNOR U30236 ( .A(n30375), .B(n30376), .Z(n30369) );
  AND U30237 ( .A(n30377), .B(n30378), .Z(n30376) );
  XOR U30238 ( .A(n30375), .B(n30379), .Z(n30377) );
  XNOR U30239 ( .A(n30361), .B(n30358), .Z(n30368) );
  AND U30240 ( .A(n30380), .B(n30381), .Z(n30358) );
  XOR U30241 ( .A(n30382), .B(n30383), .Z(n30361) );
  AND U30242 ( .A(n30384), .B(n30385), .Z(n30383) );
  XOR U30243 ( .A(n30382), .B(n30386), .Z(n30384) );
  XNOR U30244 ( .A(n30320), .B(n30364), .Z(n30366) );
  XNOR U30245 ( .A(n30387), .B(n30388), .Z(n30320) );
  AND U30246 ( .A(n963), .B(n30326), .Z(n30388) );
  XOR U30247 ( .A(n30387), .B(n30324), .Z(n30326) );
  XOR U30248 ( .A(n30389), .B(n30390), .Z(n30364) );
  AND U30249 ( .A(n30391), .B(n30392), .Z(n30390) );
  XNOR U30250 ( .A(n30389), .B(n30380), .Z(n30392) );
  IV U30251 ( .A(n30334), .Z(n30380) );
  XNOR U30252 ( .A(n30393), .B(n30373), .Z(n30334) );
  XNOR U30253 ( .A(n30394), .B(n30379), .Z(n30373) );
  XNOR U30254 ( .A(n30395), .B(n30396), .Z(n30379) );
  NOR U30255 ( .A(n30397), .B(n30398), .Z(n30396) );
  XOR U30256 ( .A(n30395), .B(n30399), .Z(n30397) );
  XNOR U30257 ( .A(n30378), .B(n30370), .Z(n30394) );
  XOR U30258 ( .A(n30400), .B(n30401), .Z(n30370) );
  AND U30259 ( .A(n30402), .B(n30403), .Z(n30401) );
  XOR U30260 ( .A(n30400), .B(n30404), .Z(n30402) );
  XNOR U30261 ( .A(n30405), .B(n30375), .Z(n30378) );
  XOR U30262 ( .A(n30406), .B(n30407), .Z(n30375) );
  AND U30263 ( .A(n30408), .B(n30409), .Z(n30407) );
  XNOR U30264 ( .A(n30410), .B(n30411), .Z(n30408) );
  IV U30265 ( .A(n30406), .Z(n30410) );
  XNOR U30266 ( .A(n30412), .B(n30413), .Z(n30405) );
  NOR U30267 ( .A(n30414), .B(n30415), .Z(n30413) );
  XNOR U30268 ( .A(n30412), .B(n30416), .Z(n30414) );
  XNOR U30269 ( .A(n30374), .B(n30381), .Z(n30393) );
  NOR U30270 ( .A(n30342), .B(n30417), .Z(n30381) );
  XOR U30271 ( .A(n30386), .B(n30385), .Z(n30374) );
  XNOR U30272 ( .A(n30418), .B(n30382), .Z(n30385) );
  XOR U30273 ( .A(n30419), .B(n30420), .Z(n30382) );
  AND U30274 ( .A(n30421), .B(n30422), .Z(n30420) );
  XNOR U30275 ( .A(n30423), .B(n30424), .Z(n30421) );
  IV U30276 ( .A(n30419), .Z(n30423) );
  XNOR U30277 ( .A(n30425), .B(n30426), .Z(n30418) );
  NOR U30278 ( .A(n30427), .B(n30428), .Z(n30426) );
  XNOR U30279 ( .A(n30425), .B(n30429), .Z(n30427) );
  XOR U30280 ( .A(n30430), .B(n30431), .Z(n30386) );
  NOR U30281 ( .A(n30432), .B(n30433), .Z(n30431) );
  XNOR U30282 ( .A(n30430), .B(n30434), .Z(n30432) );
  XNOR U30283 ( .A(n30331), .B(n30389), .Z(n30391) );
  XNOR U30284 ( .A(n30435), .B(n30436), .Z(n30331) );
  AND U30285 ( .A(n963), .B(n30338), .Z(n30436) );
  XOR U30286 ( .A(n30435), .B(n30336), .Z(n30338) );
  AND U30287 ( .A(n30339), .B(n30342), .Z(n30389) );
  XOR U30288 ( .A(n30437), .B(n30417), .Z(n30342) );
  XNOR U30289 ( .A(p_input[1344]), .B(p_input[2048]), .Z(n30417) );
  XNOR U30290 ( .A(n30404), .B(n30403), .Z(n30437) );
  XNOR U30291 ( .A(n30438), .B(n30411), .Z(n30403) );
  XNOR U30292 ( .A(n30399), .B(n30398), .Z(n30411) );
  XNOR U30293 ( .A(n30439), .B(n30395), .Z(n30398) );
  XNOR U30294 ( .A(p_input[1354]), .B(p_input[2058]), .Z(n30395) );
  XOR U30295 ( .A(p_input[1355]), .B(n16732), .Z(n30439) );
  XOR U30296 ( .A(p_input[1356]), .B(p_input[2060]), .Z(n30399) );
  XOR U30297 ( .A(n30409), .B(n30440), .Z(n30438) );
  IV U30298 ( .A(n30400), .Z(n30440) );
  XOR U30299 ( .A(p_input[1345]), .B(p_input[2049]), .Z(n30400) );
  XNOR U30300 ( .A(n30441), .B(n30416), .Z(n30409) );
  XNOR U30301 ( .A(p_input[1359]), .B(n16735), .Z(n30416) );
  XOR U30302 ( .A(n30406), .B(n30415), .Z(n30441) );
  XOR U30303 ( .A(n30442), .B(n30412), .Z(n30415) );
  XOR U30304 ( .A(p_input[1357]), .B(p_input[2061]), .Z(n30412) );
  XOR U30305 ( .A(p_input[1358]), .B(n16737), .Z(n30442) );
  XOR U30306 ( .A(p_input[1353]), .B(p_input[2057]), .Z(n30406) );
  XOR U30307 ( .A(n30424), .B(n30422), .Z(n30404) );
  XNOR U30308 ( .A(n30443), .B(n30429), .Z(n30422) );
  XOR U30309 ( .A(p_input[1352]), .B(p_input[2056]), .Z(n30429) );
  XOR U30310 ( .A(n30419), .B(n30428), .Z(n30443) );
  XOR U30311 ( .A(n30444), .B(n30425), .Z(n30428) );
  XOR U30312 ( .A(p_input[1350]), .B(p_input[2054]), .Z(n30425) );
  XOR U30313 ( .A(p_input[1351]), .B(n17722), .Z(n30444) );
  XOR U30314 ( .A(p_input[1346]), .B(p_input[2050]), .Z(n30419) );
  XNOR U30315 ( .A(n30434), .B(n30433), .Z(n30424) );
  XOR U30316 ( .A(n30445), .B(n30430), .Z(n30433) );
  XOR U30317 ( .A(p_input[1347]), .B(p_input[2051]), .Z(n30430) );
  XOR U30318 ( .A(p_input[1348]), .B(n17724), .Z(n30445) );
  XOR U30319 ( .A(p_input[1349]), .B(p_input[2053]), .Z(n30434) );
  XNOR U30320 ( .A(n30446), .B(n30447), .Z(n30339) );
  AND U30321 ( .A(n963), .B(n30448), .Z(n30447) );
  XNOR U30322 ( .A(n30449), .B(n30450), .Z(n963) );
  AND U30323 ( .A(n30451), .B(n30452), .Z(n30450) );
  XOR U30324 ( .A(n30449), .B(n30349), .Z(n30452) );
  XNOR U30325 ( .A(n30449), .B(n30303), .Z(n30451) );
  XOR U30326 ( .A(n30453), .B(n30454), .Z(n30449) );
  AND U30327 ( .A(n30455), .B(n30456), .Z(n30454) );
  XOR U30328 ( .A(n30453), .B(n30313), .Z(n30455) );
  XOR U30329 ( .A(n30457), .B(n30458), .Z(n30292) );
  AND U30330 ( .A(n967), .B(n30448), .Z(n30458) );
  XNOR U30331 ( .A(n30446), .B(n30457), .Z(n30448) );
  XNOR U30332 ( .A(n30459), .B(n30460), .Z(n967) );
  AND U30333 ( .A(n30461), .B(n30462), .Z(n30460) );
  XNOR U30334 ( .A(n30463), .B(n30459), .Z(n30462) );
  IV U30335 ( .A(n30349), .Z(n30463) );
  XNOR U30336 ( .A(n30464), .B(n30465), .Z(n30349) );
  AND U30337 ( .A(n970), .B(n30466), .Z(n30465) );
  XNOR U30338 ( .A(n30464), .B(n30467), .Z(n30466) );
  XNOR U30339 ( .A(n30303), .B(n30459), .Z(n30461) );
  XOR U30340 ( .A(n30468), .B(n30469), .Z(n30303) );
  AND U30341 ( .A(n978), .B(n30470), .Z(n30469) );
  XOR U30342 ( .A(n30453), .B(n30471), .Z(n30459) );
  AND U30343 ( .A(n30472), .B(n30456), .Z(n30471) );
  XNOR U30344 ( .A(n30362), .B(n30453), .Z(n30456) );
  XNOR U30345 ( .A(n30473), .B(n30474), .Z(n30362) );
  AND U30346 ( .A(n970), .B(n30475), .Z(n30474) );
  XOR U30347 ( .A(n30476), .B(n30473), .Z(n30475) );
  XNOR U30348 ( .A(n30477), .B(n30453), .Z(n30472) );
  IV U30349 ( .A(n30313), .Z(n30477) );
  XOR U30350 ( .A(n30478), .B(n30479), .Z(n30313) );
  AND U30351 ( .A(n978), .B(n30480), .Z(n30479) );
  XOR U30352 ( .A(n30481), .B(n30482), .Z(n30453) );
  AND U30353 ( .A(n30483), .B(n30484), .Z(n30482) );
  XNOR U30354 ( .A(n30387), .B(n30481), .Z(n30484) );
  XNOR U30355 ( .A(n30485), .B(n30486), .Z(n30387) );
  AND U30356 ( .A(n970), .B(n30487), .Z(n30486) );
  XNOR U30357 ( .A(n30488), .B(n30485), .Z(n30487) );
  XOR U30358 ( .A(n30481), .B(n30324), .Z(n30483) );
  XOR U30359 ( .A(n30489), .B(n30490), .Z(n30324) );
  AND U30360 ( .A(n978), .B(n30491), .Z(n30490) );
  XOR U30361 ( .A(n30492), .B(n30493), .Z(n30481) );
  AND U30362 ( .A(n30494), .B(n30495), .Z(n30493) );
  XNOR U30363 ( .A(n30492), .B(n30435), .Z(n30495) );
  XNOR U30364 ( .A(n30496), .B(n30497), .Z(n30435) );
  AND U30365 ( .A(n970), .B(n30498), .Z(n30497) );
  XOR U30366 ( .A(n30499), .B(n30496), .Z(n30498) );
  XNOR U30367 ( .A(n30500), .B(n30492), .Z(n30494) );
  IV U30368 ( .A(n30336), .Z(n30500) );
  XOR U30369 ( .A(n30501), .B(n30502), .Z(n30336) );
  AND U30370 ( .A(n978), .B(n30503), .Z(n30502) );
  AND U30371 ( .A(n30457), .B(n30446), .Z(n30492) );
  XNOR U30372 ( .A(n30504), .B(n30505), .Z(n30446) );
  AND U30373 ( .A(n970), .B(n30506), .Z(n30505) );
  XNOR U30374 ( .A(n30507), .B(n30504), .Z(n30506) );
  XNOR U30375 ( .A(n30508), .B(n30509), .Z(n970) );
  AND U30376 ( .A(n30510), .B(n30511), .Z(n30509) );
  XOR U30377 ( .A(n30467), .B(n30508), .Z(n30511) );
  AND U30378 ( .A(n30512), .B(n30513), .Z(n30467) );
  XOR U30379 ( .A(n30508), .B(n30464), .Z(n30510) );
  XNOR U30380 ( .A(n30514), .B(n30515), .Z(n30464) );
  AND U30381 ( .A(n974), .B(n30470), .Z(n30515) );
  XOR U30382 ( .A(n30468), .B(n30514), .Z(n30470) );
  XOR U30383 ( .A(n30516), .B(n30517), .Z(n30508) );
  AND U30384 ( .A(n30518), .B(n30519), .Z(n30517) );
  XNOR U30385 ( .A(n30516), .B(n30512), .Z(n30519) );
  IV U30386 ( .A(n30476), .Z(n30512) );
  XOR U30387 ( .A(n30520), .B(n30521), .Z(n30476) );
  XOR U30388 ( .A(n30522), .B(n30513), .Z(n30521) );
  AND U30389 ( .A(n30488), .B(n30523), .Z(n30513) );
  AND U30390 ( .A(n30524), .B(n30525), .Z(n30522) );
  XOR U30391 ( .A(n30526), .B(n30520), .Z(n30524) );
  XNOR U30392 ( .A(n30473), .B(n30516), .Z(n30518) );
  XNOR U30393 ( .A(n30527), .B(n30528), .Z(n30473) );
  AND U30394 ( .A(n974), .B(n30480), .Z(n30528) );
  XOR U30395 ( .A(n30527), .B(n30478), .Z(n30480) );
  XOR U30396 ( .A(n30529), .B(n30530), .Z(n30516) );
  AND U30397 ( .A(n30531), .B(n30532), .Z(n30530) );
  XNOR U30398 ( .A(n30529), .B(n30488), .Z(n30532) );
  XOR U30399 ( .A(n30533), .B(n30525), .Z(n30488) );
  XNOR U30400 ( .A(n30534), .B(n30520), .Z(n30525) );
  XOR U30401 ( .A(n30535), .B(n30536), .Z(n30520) );
  AND U30402 ( .A(n30537), .B(n30538), .Z(n30536) );
  XOR U30403 ( .A(n30539), .B(n30535), .Z(n30537) );
  XNOR U30404 ( .A(n30540), .B(n30541), .Z(n30534) );
  AND U30405 ( .A(n30542), .B(n30543), .Z(n30541) );
  XOR U30406 ( .A(n30540), .B(n30544), .Z(n30542) );
  XNOR U30407 ( .A(n30526), .B(n30523), .Z(n30533) );
  AND U30408 ( .A(n30545), .B(n30546), .Z(n30523) );
  XOR U30409 ( .A(n30547), .B(n30548), .Z(n30526) );
  AND U30410 ( .A(n30549), .B(n30550), .Z(n30548) );
  XOR U30411 ( .A(n30547), .B(n30551), .Z(n30549) );
  XNOR U30412 ( .A(n30485), .B(n30529), .Z(n30531) );
  XNOR U30413 ( .A(n30552), .B(n30553), .Z(n30485) );
  AND U30414 ( .A(n974), .B(n30491), .Z(n30553) );
  XOR U30415 ( .A(n30552), .B(n30489), .Z(n30491) );
  XOR U30416 ( .A(n30554), .B(n30555), .Z(n30529) );
  AND U30417 ( .A(n30556), .B(n30557), .Z(n30555) );
  XNOR U30418 ( .A(n30554), .B(n30545), .Z(n30557) );
  IV U30419 ( .A(n30499), .Z(n30545) );
  XNOR U30420 ( .A(n30558), .B(n30538), .Z(n30499) );
  XNOR U30421 ( .A(n30559), .B(n30544), .Z(n30538) );
  XNOR U30422 ( .A(n30560), .B(n30561), .Z(n30544) );
  NOR U30423 ( .A(n30562), .B(n30563), .Z(n30561) );
  XOR U30424 ( .A(n30560), .B(n30564), .Z(n30562) );
  XNOR U30425 ( .A(n30543), .B(n30535), .Z(n30559) );
  XOR U30426 ( .A(n30565), .B(n30566), .Z(n30535) );
  AND U30427 ( .A(n30567), .B(n30568), .Z(n30566) );
  XOR U30428 ( .A(n30565), .B(n30569), .Z(n30567) );
  XNOR U30429 ( .A(n30570), .B(n30540), .Z(n30543) );
  XOR U30430 ( .A(n30571), .B(n30572), .Z(n30540) );
  AND U30431 ( .A(n30573), .B(n30574), .Z(n30572) );
  XNOR U30432 ( .A(n30575), .B(n30576), .Z(n30573) );
  IV U30433 ( .A(n30571), .Z(n30575) );
  XNOR U30434 ( .A(n30577), .B(n30578), .Z(n30570) );
  NOR U30435 ( .A(n30579), .B(n30580), .Z(n30578) );
  XNOR U30436 ( .A(n30577), .B(n30581), .Z(n30579) );
  XNOR U30437 ( .A(n30539), .B(n30546), .Z(n30558) );
  NOR U30438 ( .A(n30507), .B(n30582), .Z(n30546) );
  XOR U30439 ( .A(n30551), .B(n30550), .Z(n30539) );
  XNOR U30440 ( .A(n30583), .B(n30547), .Z(n30550) );
  XOR U30441 ( .A(n30584), .B(n30585), .Z(n30547) );
  AND U30442 ( .A(n30586), .B(n30587), .Z(n30585) );
  XNOR U30443 ( .A(n30588), .B(n30589), .Z(n30586) );
  IV U30444 ( .A(n30584), .Z(n30588) );
  XNOR U30445 ( .A(n30590), .B(n30591), .Z(n30583) );
  NOR U30446 ( .A(n30592), .B(n30593), .Z(n30591) );
  XNOR U30447 ( .A(n30590), .B(n30594), .Z(n30592) );
  XOR U30448 ( .A(n30595), .B(n30596), .Z(n30551) );
  NOR U30449 ( .A(n30597), .B(n30598), .Z(n30596) );
  XNOR U30450 ( .A(n30595), .B(n30599), .Z(n30597) );
  XNOR U30451 ( .A(n30496), .B(n30554), .Z(n30556) );
  XNOR U30452 ( .A(n30600), .B(n30601), .Z(n30496) );
  AND U30453 ( .A(n974), .B(n30503), .Z(n30601) );
  XOR U30454 ( .A(n30600), .B(n30501), .Z(n30503) );
  AND U30455 ( .A(n30504), .B(n30507), .Z(n30554) );
  XOR U30456 ( .A(n30602), .B(n30582), .Z(n30507) );
  XNOR U30457 ( .A(p_input[1360]), .B(p_input[2048]), .Z(n30582) );
  XNOR U30458 ( .A(n30569), .B(n30568), .Z(n30602) );
  XNOR U30459 ( .A(n30603), .B(n30576), .Z(n30568) );
  XNOR U30460 ( .A(n30564), .B(n30563), .Z(n30576) );
  XNOR U30461 ( .A(n30604), .B(n30560), .Z(n30563) );
  XNOR U30462 ( .A(p_input[1370]), .B(p_input[2058]), .Z(n30560) );
  XOR U30463 ( .A(p_input[1371]), .B(n16732), .Z(n30604) );
  XOR U30464 ( .A(p_input[1372]), .B(p_input[2060]), .Z(n30564) );
  XOR U30465 ( .A(n30574), .B(n30605), .Z(n30603) );
  IV U30466 ( .A(n30565), .Z(n30605) );
  XOR U30467 ( .A(p_input[1361]), .B(p_input[2049]), .Z(n30565) );
  XNOR U30468 ( .A(n30606), .B(n30581), .Z(n30574) );
  XNOR U30469 ( .A(p_input[1375]), .B(n16735), .Z(n30581) );
  XOR U30470 ( .A(n30571), .B(n30580), .Z(n30606) );
  XOR U30471 ( .A(n30607), .B(n30577), .Z(n30580) );
  XOR U30472 ( .A(p_input[1373]), .B(p_input[2061]), .Z(n30577) );
  XOR U30473 ( .A(p_input[1374]), .B(n16737), .Z(n30607) );
  XOR U30474 ( .A(p_input[1369]), .B(p_input[2057]), .Z(n30571) );
  XOR U30475 ( .A(n30589), .B(n30587), .Z(n30569) );
  XNOR U30476 ( .A(n30608), .B(n30594), .Z(n30587) );
  XOR U30477 ( .A(p_input[1368]), .B(p_input[2056]), .Z(n30594) );
  XOR U30478 ( .A(n30584), .B(n30593), .Z(n30608) );
  XOR U30479 ( .A(n30609), .B(n30590), .Z(n30593) );
  XOR U30480 ( .A(p_input[1366]), .B(p_input[2054]), .Z(n30590) );
  XOR U30481 ( .A(p_input[1367]), .B(n17722), .Z(n30609) );
  XOR U30482 ( .A(p_input[1362]), .B(p_input[2050]), .Z(n30584) );
  XNOR U30483 ( .A(n30599), .B(n30598), .Z(n30589) );
  XOR U30484 ( .A(n30610), .B(n30595), .Z(n30598) );
  XOR U30485 ( .A(p_input[1363]), .B(p_input[2051]), .Z(n30595) );
  XOR U30486 ( .A(p_input[1364]), .B(n17724), .Z(n30610) );
  XOR U30487 ( .A(p_input[1365]), .B(p_input[2053]), .Z(n30599) );
  XNOR U30488 ( .A(n30611), .B(n30612), .Z(n30504) );
  AND U30489 ( .A(n974), .B(n30613), .Z(n30612) );
  XNOR U30490 ( .A(n30614), .B(n30615), .Z(n974) );
  AND U30491 ( .A(n30616), .B(n30617), .Z(n30615) );
  XOR U30492 ( .A(n30614), .B(n30514), .Z(n30617) );
  XNOR U30493 ( .A(n30614), .B(n30468), .Z(n30616) );
  XOR U30494 ( .A(n30618), .B(n30619), .Z(n30614) );
  AND U30495 ( .A(n30620), .B(n30621), .Z(n30619) );
  XOR U30496 ( .A(n30618), .B(n30478), .Z(n30620) );
  XOR U30497 ( .A(n30622), .B(n30623), .Z(n30457) );
  AND U30498 ( .A(n978), .B(n30613), .Z(n30623) );
  XNOR U30499 ( .A(n30611), .B(n30622), .Z(n30613) );
  XNOR U30500 ( .A(n30624), .B(n30625), .Z(n978) );
  AND U30501 ( .A(n30626), .B(n30627), .Z(n30625) );
  XNOR U30502 ( .A(n30628), .B(n30624), .Z(n30627) );
  IV U30503 ( .A(n30514), .Z(n30628) );
  XNOR U30504 ( .A(n30629), .B(n30630), .Z(n30514) );
  AND U30505 ( .A(n981), .B(n30631), .Z(n30630) );
  XNOR U30506 ( .A(n30629), .B(n30632), .Z(n30631) );
  XNOR U30507 ( .A(n30468), .B(n30624), .Z(n30626) );
  XOR U30508 ( .A(n30633), .B(n30634), .Z(n30468) );
  AND U30509 ( .A(n989), .B(n30635), .Z(n30634) );
  XOR U30510 ( .A(n30618), .B(n30636), .Z(n30624) );
  AND U30511 ( .A(n30637), .B(n30621), .Z(n30636) );
  XNOR U30512 ( .A(n30527), .B(n30618), .Z(n30621) );
  XNOR U30513 ( .A(n30638), .B(n30639), .Z(n30527) );
  AND U30514 ( .A(n981), .B(n30640), .Z(n30639) );
  XOR U30515 ( .A(n30641), .B(n30638), .Z(n30640) );
  XNOR U30516 ( .A(n30642), .B(n30618), .Z(n30637) );
  IV U30517 ( .A(n30478), .Z(n30642) );
  XOR U30518 ( .A(n30643), .B(n30644), .Z(n30478) );
  AND U30519 ( .A(n989), .B(n30645), .Z(n30644) );
  XOR U30520 ( .A(n30646), .B(n30647), .Z(n30618) );
  AND U30521 ( .A(n30648), .B(n30649), .Z(n30647) );
  XNOR U30522 ( .A(n30552), .B(n30646), .Z(n30649) );
  XNOR U30523 ( .A(n30650), .B(n30651), .Z(n30552) );
  AND U30524 ( .A(n981), .B(n30652), .Z(n30651) );
  XNOR U30525 ( .A(n30653), .B(n30650), .Z(n30652) );
  XOR U30526 ( .A(n30646), .B(n30489), .Z(n30648) );
  XOR U30527 ( .A(n30654), .B(n30655), .Z(n30489) );
  AND U30528 ( .A(n989), .B(n30656), .Z(n30655) );
  XOR U30529 ( .A(n30657), .B(n30658), .Z(n30646) );
  AND U30530 ( .A(n30659), .B(n30660), .Z(n30658) );
  XNOR U30531 ( .A(n30657), .B(n30600), .Z(n30660) );
  XNOR U30532 ( .A(n30661), .B(n30662), .Z(n30600) );
  AND U30533 ( .A(n981), .B(n30663), .Z(n30662) );
  XOR U30534 ( .A(n30664), .B(n30661), .Z(n30663) );
  XNOR U30535 ( .A(n30665), .B(n30657), .Z(n30659) );
  IV U30536 ( .A(n30501), .Z(n30665) );
  XOR U30537 ( .A(n30666), .B(n30667), .Z(n30501) );
  AND U30538 ( .A(n989), .B(n30668), .Z(n30667) );
  AND U30539 ( .A(n30622), .B(n30611), .Z(n30657) );
  XNOR U30540 ( .A(n30669), .B(n30670), .Z(n30611) );
  AND U30541 ( .A(n981), .B(n30671), .Z(n30670) );
  XNOR U30542 ( .A(n30672), .B(n30669), .Z(n30671) );
  XNOR U30543 ( .A(n30673), .B(n30674), .Z(n981) );
  AND U30544 ( .A(n30675), .B(n30676), .Z(n30674) );
  XOR U30545 ( .A(n30632), .B(n30673), .Z(n30676) );
  AND U30546 ( .A(n30677), .B(n30678), .Z(n30632) );
  XOR U30547 ( .A(n30673), .B(n30629), .Z(n30675) );
  XNOR U30548 ( .A(n30679), .B(n30680), .Z(n30629) );
  AND U30549 ( .A(n985), .B(n30635), .Z(n30680) );
  XOR U30550 ( .A(n30633), .B(n30679), .Z(n30635) );
  XOR U30551 ( .A(n30681), .B(n30682), .Z(n30673) );
  AND U30552 ( .A(n30683), .B(n30684), .Z(n30682) );
  XNOR U30553 ( .A(n30681), .B(n30677), .Z(n30684) );
  IV U30554 ( .A(n30641), .Z(n30677) );
  XOR U30555 ( .A(n30685), .B(n30686), .Z(n30641) );
  XOR U30556 ( .A(n30687), .B(n30678), .Z(n30686) );
  AND U30557 ( .A(n30653), .B(n30688), .Z(n30678) );
  AND U30558 ( .A(n30689), .B(n30690), .Z(n30687) );
  XOR U30559 ( .A(n30691), .B(n30685), .Z(n30689) );
  XNOR U30560 ( .A(n30638), .B(n30681), .Z(n30683) );
  XNOR U30561 ( .A(n30692), .B(n30693), .Z(n30638) );
  AND U30562 ( .A(n985), .B(n30645), .Z(n30693) );
  XOR U30563 ( .A(n30692), .B(n30643), .Z(n30645) );
  XOR U30564 ( .A(n30694), .B(n30695), .Z(n30681) );
  AND U30565 ( .A(n30696), .B(n30697), .Z(n30695) );
  XNOR U30566 ( .A(n30694), .B(n30653), .Z(n30697) );
  XOR U30567 ( .A(n30698), .B(n30690), .Z(n30653) );
  XNOR U30568 ( .A(n30699), .B(n30685), .Z(n30690) );
  XOR U30569 ( .A(n30700), .B(n30701), .Z(n30685) );
  AND U30570 ( .A(n30702), .B(n30703), .Z(n30701) );
  XOR U30571 ( .A(n30704), .B(n30700), .Z(n30702) );
  XNOR U30572 ( .A(n30705), .B(n30706), .Z(n30699) );
  AND U30573 ( .A(n30707), .B(n30708), .Z(n30706) );
  XOR U30574 ( .A(n30705), .B(n30709), .Z(n30707) );
  XNOR U30575 ( .A(n30691), .B(n30688), .Z(n30698) );
  AND U30576 ( .A(n30710), .B(n30711), .Z(n30688) );
  XOR U30577 ( .A(n30712), .B(n30713), .Z(n30691) );
  AND U30578 ( .A(n30714), .B(n30715), .Z(n30713) );
  XOR U30579 ( .A(n30712), .B(n30716), .Z(n30714) );
  XNOR U30580 ( .A(n30650), .B(n30694), .Z(n30696) );
  XNOR U30581 ( .A(n30717), .B(n30718), .Z(n30650) );
  AND U30582 ( .A(n985), .B(n30656), .Z(n30718) );
  XOR U30583 ( .A(n30717), .B(n30654), .Z(n30656) );
  XOR U30584 ( .A(n30719), .B(n30720), .Z(n30694) );
  AND U30585 ( .A(n30721), .B(n30722), .Z(n30720) );
  XNOR U30586 ( .A(n30719), .B(n30710), .Z(n30722) );
  IV U30587 ( .A(n30664), .Z(n30710) );
  XNOR U30588 ( .A(n30723), .B(n30703), .Z(n30664) );
  XNOR U30589 ( .A(n30724), .B(n30709), .Z(n30703) );
  XNOR U30590 ( .A(n30725), .B(n30726), .Z(n30709) );
  NOR U30591 ( .A(n30727), .B(n30728), .Z(n30726) );
  XOR U30592 ( .A(n30725), .B(n30729), .Z(n30727) );
  XNOR U30593 ( .A(n30708), .B(n30700), .Z(n30724) );
  XOR U30594 ( .A(n30730), .B(n30731), .Z(n30700) );
  AND U30595 ( .A(n30732), .B(n30733), .Z(n30731) );
  XOR U30596 ( .A(n30730), .B(n30734), .Z(n30732) );
  XNOR U30597 ( .A(n30735), .B(n30705), .Z(n30708) );
  XOR U30598 ( .A(n30736), .B(n30737), .Z(n30705) );
  AND U30599 ( .A(n30738), .B(n30739), .Z(n30737) );
  XNOR U30600 ( .A(n30740), .B(n30741), .Z(n30738) );
  IV U30601 ( .A(n30736), .Z(n30740) );
  XNOR U30602 ( .A(n30742), .B(n30743), .Z(n30735) );
  NOR U30603 ( .A(n30744), .B(n30745), .Z(n30743) );
  XNOR U30604 ( .A(n30742), .B(n30746), .Z(n30744) );
  XNOR U30605 ( .A(n30704), .B(n30711), .Z(n30723) );
  NOR U30606 ( .A(n30672), .B(n30747), .Z(n30711) );
  XOR U30607 ( .A(n30716), .B(n30715), .Z(n30704) );
  XNOR U30608 ( .A(n30748), .B(n30712), .Z(n30715) );
  XOR U30609 ( .A(n30749), .B(n30750), .Z(n30712) );
  AND U30610 ( .A(n30751), .B(n30752), .Z(n30750) );
  XNOR U30611 ( .A(n30753), .B(n30754), .Z(n30751) );
  IV U30612 ( .A(n30749), .Z(n30753) );
  XNOR U30613 ( .A(n30755), .B(n30756), .Z(n30748) );
  NOR U30614 ( .A(n30757), .B(n30758), .Z(n30756) );
  XNOR U30615 ( .A(n30755), .B(n30759), .Z(n30757) );
  XOR U30616 ( .A(n30760), .B(n30761), .Z(n30716) );
  NOR U30617 ( .A(n30762), .B(n30763), .Z(n30761) );
  XNOR U30618 ( .A(n30760), .B(n30764), .Z(n30762) );
  XNOR U30619 ( .A(n30661), .B(n30719), .Z(n30721) );
  XNOR U30620 ( .A(n30765), .B(n30766), .Z(n30661) );
  AND U30621 ( .A(n985), .B(n30668), .Z(n30766) );
  XOR U30622 ( .A(n30765), .B(n30666), .Z(n30668) );
  AND U30623 ( .A(n30669), .B(n30672), .Z(n30719) );
  XOR U30624 ( .A(n30767), .B(n30747), .Z(n30672) );
  XNOR U30625 ( .A(p_input[1376]), .B(p_input[2048]), .Z(n30747) );
  XNOR U30626 ( .A(n30734), .B(n30733), .Z(n30767) );
  XNOR U30627 ( .A(n30768), .B(n30741), .Z(n30733) );
  XNOR U30628 ( .A(n30729), .B(n30728), .Z(n30741) );
  XNOR U30629 ( .A(n30769), .B(n30725), .Z(n30728) );
  XNOR U30630 ( .A(p_input[1386]), .B(p_input[2058]), .Z(n30725) );
  XOR U30631 ( .A(p_input[1387]), .B(n16732), .Z(n30769) );
  XOR U30632 ( .A(p_input[1388]), .B(p_input[2060]), .Z(n30729) );
  XOR U30633 ( .A(n30739), .B(n30770), .Z(n30768) );
  IV U30634 ( .A(n30730), .Z(n30770) );
  XOR U30635 ( .A(p_input[1377]), .B(p_input[2049]), .Z(n30730) );
  XNOR U30636 ( .A(n30771), .B(n30746), .Z(n30739) );
  XNOR U30637 ( .A(p_input[1391]), .B(n16735), .Z(n30746) );
  XOR U30638 ( .A(n30736), .B(n30745), .Z(n30771) );
  XOR U30639 ( .A(n30772), .B(n30742), .Z(n30745) );
  XOR U30640 ( .A(p_input[1389]), .B(p_input[2061]), .Z(n30742) );
  XOR U30641 ( .A(p_input[1390]), .B(n16737), .Z(n30772) );
  XOR U30642 ( .A(p_input[1385]), .B(p_input[2057]), .Z(n30736) );
  XOR U30643 ( .A(n30754), .B(n30752), .Z(n30734) );
  XNOR U30644 ( .A(n30773), .B(n30759), .Z(n30752) );
  XOR U30645 ( .A(p_input[1384]), .B(p_input[2056]), .Z(n30759) );
  XOR U30646 ( .A(n30749), .B(n30758), .Z(n30773) );
  XOR U30647 ( .A(n30774), .B(n30755), .Z(n30758) );
  XOR U30648 ( .A(p_input[1382]), .B(p_input[2054]), .Z(n30755) );
  XOR U30649 ( .A(p_input[1383]), .B(n17722), .Z(n30774) );
  XOR U30650 ( .A(p_input[1378]), .B(p_input[2050]), .Z(n30749) );
  XNOR U30651 ( .A(n30764), .B(n30763), .Z(n30754) );
  XOR U30652 ( .A(n30775), .B(n30760), .Z(n30763) );
  XOR U30653 ( .A(p_input[1379]), .B(p_input[2051]), .Z(n30760) );
  XOR U30654 ( .A(p_input[1380]), .B(n17724), .Z(n30775) );
  XOR U30655 ( .A(p_input[1381]), .B(p_input[2053]), .Z(n30764) );
  XNOR U30656 ( .A(n30776), .B(n30777), .Z(n30669) );
  AND U30657 ( .A(n985), .B(n30778), .Z(n30777) );
  XNOR U30658 ( .A(n30779), .B(n30780), .Z(n985) );
  AND U30659 ( .A(n30781), .B(n30782), .Z(n30780) );
  XOR U30660 ( .A(n30779), .B(n30679), .Z(n30782) );
  XNOR U30661 ( .A(n30779), .B(n30633), .Z(n30781) );
  XOR U30662 ( .A(n30783), .B(n30784), .Z(n30779) );
  AND U30663 ( .A(n30785), .B(n30786), .Z(n30784) );
  XOR U30664 ( .A(n30783), .B(n30643), .Z(n30785) );
  XOR U30665 ( .A(n30787), .B(n30788), .Z(n30622) );
  AND U30666 ( .A(n989), .B(n30778), .Z(n30788) );
  XNOR U30667 ( .A(n30776), .B(n30787), .Z(n30778) );
  XNOR U30668 ( .A(n30789), .B(n30790), .Z(n989) );
  AND U30669 ( .A(n30791), .B(n30792), .Z(n30790) );
  XNOR U30670 ( .A(n30793), .B(n30789), .Z(n30792) );
  IV U30671 ( .A(n30679), .Z(n30793) );
  XNOR U30672 ( .A(n30794), .B(n30795), .Z(n30679) );
  AND U30673 ( .A(n992), .B(n30796), .Z(n30795) );
  XNOR U30674 ( .A(n30794), .B(n30797), .Z(n30796) );
  XNOR U30675 ( .A(n30633), .B(n30789), .Z(n30791) );
  XOR U30676 ( .A(n30798), .B(n30799), .Z(n30633) );
  AND U30677 ( .A(n1000), .B(n30800), .Z(n30799) );
  XOR U30678 ( .A(n30783), .B(n30801), .Z(n30789) );
  AND U30679 ( .A(n30802), .B(n30786), .Z(n30801) );
  XNOR U30680 ( .A(n30692), .B(n30783), .Z(n30786) );
  XNOR U30681 ( .A(n30803), .B(n30804), .Z(n30692) );
  AND U30682 ( .A(n992), .B(n30805), .Z(n30804) );
  XOR U30683 ( .A(n30806), .B(n30803), .Z(n30805) );
  XNOR U30684 ( .A(n30807), .B(n30783), .Z(n30802) );
  IV U30685 ( .A(n30643), .Z(n30807) );
  XOR U30686 ( .A(n30808), .B(n30809), .Z(n30643) );
  AND U30687 ( .A(n1000), .B(n30810), .Z(n30809) );
  XOR U30688 ( .A(n30811), .B(n30812), .Z(n30783) );
  AND U30689 ( .A(n30813), .B(n30814), .Z(n30812) );
  XNOR U30690 ( .A(n30717), .B(n30811), .Z(n30814) );
  XNOR U30691 ( .A(n30815), .B(n30816), .Z(n30717) );
  AND U30692 ( .A(n992), .B(n30817), .Z(n30816) );
  XNOR U30693 ( .A(n30818), .B(n30815), .Z(n30817) );
  XOR U30694 ( .A(n30811), .B(n30654), .Z(n30813) );
  XOR U30695 ( .A(n30819), .B(n30820), .Z(n30654) );
  AND U30696 ( .A(n1000), .B(n30821), .Z(n30820) );
  XOR U30697 ( .A(n30822), .B(n30823), .Z(n30811) );
  AND U30698 ( .A(n30824), .B(n30825), .Z(n30823) );
  XNOR U30699 ( .A(n30822), .B(n30765), .Z(n30825) );
  XNOR U30700 ( .A(n30826), .B(n30827), .Z(n30765) );
  AND U30701 ( .A(n992), .B(n30828), .Z(n30827) );
  XOR U30702 ( .A(n30829), .B(n30826), .Z(n30828) );
  XNOR U30703 ( .A(n30830), .B(n30822), .Z(n30824) );
  IV U30704 ( .A(n30666), .Z(n30830) );
  XOR U30705 ( .A(n30831), .B(n30832), .Z(n30666) );
  AND U30706 ( .A(n1000), .B(n30833), .Z(n30832) );
  AND U30707 ( .A(n30787), .B(n30776), .Z(n30822) );
  XNOR U30708 ( .A(n30834), .B(n30835), .Z(n30776) );
  AND U30709 ( .A(n992), .B(n30836), .Z(n30835) );
  XNOR U30710 ( .A(n30837), .B(n30834), .Z(n30836) );
  XNOR U30711 ( .A(n30838), .B(n30839), .Z(n992) );
  AND U30712 ( .A(n30840), .B(n30841), .Z(n30839) );
  XOR U30713 ( .A(n30797), .B(n30838), .Z(n30841) );
  AND U30714 ( .A(n30842), .B(n30843), .Z(n30797) );
  XOR U30715 ( .A(n30838), .B(n30794), .Z(n30840) );
  XNOR U30716 ( .A(n30844), .B(n30845), .Z(n30794) );
  AND U30717 ( .A(n996), .B(n30800), .Z(n30845) );
  XOR U30718 ( .A(n30798), .B(n30844), .Z(n30800) );
  XOR U30719 ( .A(n30846), .B(n30847), .Z(n30838) );
  AND U30720 ( .A(n30848), .B(n30849), .Z(n30847) );
  XNOR U30721 ( .A(n30846), .B(n30842), .Z(n30849) );
  IV U30722 ( .A(n30806), .Z(n30842) );
  XOR U30723 ( .A(n30850), .B(n30851), .Z(n30806) );
  XOR U30724 ( .A(n30852), .B(n30843), .Z(n30851) );
  AND U30725 ( .A(n30818), .B(n30853), .Z(n30843) );
  AND U30726 ( .A(n30854), .B(n30855), .Z(n30852) );
  XOR U30727 ( .A(n30856), .B(n30850), .Z(n30854) );
  XNOR U30728 ( .A(n30803), .B(n30846), .Z(n30848) );
  XNOR U30729 ( .A(n30857), .B(n30858), .Z(n30803) );
  AND U30730 ( .A(n996), .B(n30810), .Z(n30858) );
  XOR U30731 ( .A(n30857), .B(n30808), .Z(n30810) );
  XOR U30732 ( .A(n30859), .B(n30860), .Z(n30846) );
  AND U30733 ( .A(n30861), .B(n30862), .Z(n30860) );
  XNOR U30734 ( .A(n30859), .B(n30818), .Z(n30862) );
  XOR U30735 ( .A(n30863), .B(n30855), .Z(n30818) );
  XNOR U30736 ( .A(n30864), .B(n30850), .Z(n30855) );
  XOR U30737 ( .A(n30865), .B(n30866), .Z(n30850) );
  AND U30738 ( .A(n30867), .B(n30868), .Z(n30866) );
  XOR U30739 ( .A(n30869), .B(n30865), .Z(n30867) );
  XNOR U30740 ( .A(n30870), .B(n30871), .Z(n30864) );
  AND U30741 ( .A(n30872), .B(n30873), .Z(n30871) );
  XOR U30742 ( .A(n30870), .B(n30874), .Z(n30872) );
  XNOR U30743 ( .A(n30856), .B(n30853), .Z(n30863) );
  AND U30744 ( .A(n30875), .B(n30876), .Z(n30853) );
  XOR U30745 ( .A(n30877), .B(n30878), .Z(n30856) );
  AND U30746 ( .A(n30879), .B(n30880), .Z(n30878) );
  XOR U30747 ( .A(n30877), .B(n30881), .Z(n30879) );
  XNOR U30748 ( .A(n30815), .B(n30859), .Z(n30861) );
  XNOR U30749 ( .A(n30882), .B(n30883), .Z(n30815) );
  AND U30750 ( .A(n996), .B(n30821), .Z(n30883) );
  XOR U30751 ( .A(n30882), .B(n30819), .Z(n30821) );
  XOR U30752 ( .A(n30884), .B(n30885), .Z(n30859) );
  AND U30753 ( .A(n30886), .B(n30887), .Z(n30885) );
  XNOR U30754 ( .A(n30884), .B(n30875), .Z(n30887) );
  IV U30755 ( .A(n30829), .Z(n30875) );
  XNOR U30756 ( .A(n30888), .B(n30868), .Z(n30829) );
  XNOR U30757 ( .A(n30889), .B(n30874), .Z(n30868) );
  XNOR U30758 ( .A(n30890), .B(n30891), .Z(n30874) );
  NOR U30759 ( .A(n30892), .B(n30893), .Z(n30891) );
  XOR U30760 ( .A(n30890), .B(n30894), .Z(n30892) );
  XNOR U30761 ( .A(n30873), .B(n30865), .Z(n30889) );
  XOR U30762 ( .A(n30895), .B(n30896), .Z(n30865) );
  AND U30763 ( .A(n30897), .B(n30898), .Z(n30896) );
  XOR U30764 ( .A(n30895), .B(n30899), .Z(n30897) );
  XNOR U30765 ( .A(n30900), .B(n30870), .Z(n30873) );
  XOR U30766 ( .A(n30901), .B(n30902), .Z(n30870) );
  AND U30767 ( .A(n30903), .B(n30904), .Z(n30902) );
  XNOR U30768 ( .A(n30905), .B(n30906), .Z(n30903) );
  IV U30769 ( .A(n30901), .Z(n30905) );
  XNOR U30770 ( .A(n30907), .B(n30908), .Z(n30900) );
  NOR U30771 ( .A(n30909), .B(n30910), .Z(n30908) );
  XNOR U30772 ( .A(n30907), .B(n30911), .Z(n30909) );
  XNOR U30773 ( .A(n30869), .B(n30876), .Z(n30888) );
  NOR U30774 ( .A(n30837), .B(n30912), .Z(n30876) );
  XOR U30775 ( .A(n30881), .B(n30880), .Z(n30869) );
  XNOR U30776 ( .A(n30913), .B(n30877), .Z(n30880) );
  XOR U30777 ( .A(n30914), .B(n30915), .Z(n30877) );
  AND U30778 ( .A(n30916), .B(n30917), .Z(n30915) );
  XNOR U30779 ( .A(n30918), .B(n30919), .Z(n30916) );
  IV U30780 ( .A(n30914), .Z(n30918) );
  XNOR U30781 ( .A(n30920), .B(n30921), .Z(n30913) );
  NOR U30782 ( .A(n30922), .B(n30923), .Z(n30921) );
  XNOR U30783 ( .A(n30920), .B(n30924), .Z(n30922) );
  XOR U30784 ( .A(n30925), .B(n30926), .Z(n30881) );
  NOR U30785 ( .A(n30927), .B(n30928), .Z(n30926) );
  XNOR U30786 ( .A(n30925), .B(n30929), .Z(n30927) );
  XNOR U30787 ( .A(n30826), .B(n30884), .Z(n30886) );
  XNOR U30788 ( .A(n30930), .B(n30931), .Z(n30826) );
  AND U30789 ( .A(n996), .B(n30833), .Z(n30931) );
  XOR U30790 ( .A(n30930), .B(n30831), .Z(n30833) );
  AND U30791 ( .A(n30834), .B(n30837), .Z(n30884) );
  XOR U30792 ( .A(n30932), .B(n30912), .Z(n30837) );
  XNOR U30793 ( .A(p_input[1392]), .B(p_input[2048]), .Z(n30912) );
  XNOR U30794 ( .A(n30899), .B(n30898), .Z(n30932) );
  XNOR U30795 ( .A(n30933), .B(n30906), .Z(n30898) );
  XNOR U30796 ( .A(n30894), .B(n30893), .Z(n30906) );
  XNOR U30797 ( .A(n30934), .B(n30890), .Z(n30893) );
  XNOR U30798 ( .A(p_input[1402]), .B(p_input[2058]), .Z(n30890) );
  XOR U30799 ( .A(p_input[1403]), .B(n16732), .Z(n30934) );
  XOR U30800 ( .A(p_input[1404]), .B(p_input[2060]), .Z(n30894) );
  XOR U30801 ( .A(n30904), .B(n30935), .Z(n30933) );
  IV U30802 ( .A(n30895), .Z(n30935) );
  XOR U30803 ( .A(p_input[1393]), .B(p_input[2049]), .Z(n30895) );
  XNOR U30804 ( .A(n30936), .B(n30911), .Z(n30904) );
  XNOR U30805 ( .A(p_input[1407]), .B(n16735), .Z(n30911) );
  XOR U30806 ( .A(n30901), .B(n30910), .Z(n30936) );
  XOR U30807 ( .A(n30937), .B(n30907), .Z(n30910) );
  XOR U30808 ( .A(p_input[1405]), .B(p_input[2061]), .Z(n30907) );
  XOR U30809 ( .A(p_input[1406]), .B(n16737), .Z(n30937) );
  XOR U30810 ( .A(p_input[1401]), .B(p_input[2057]), .Z(n30901) );
  XOR U30811 ( .A(n30919), .B(n30917), .Z(n30899) );
  XNOR U30812 ( .A(n30938), .B(n30924), .Z(n30917) );
  XOR U30813 ( .A(p_input[1400]), .B(p_input[2056]), .Z(n30924) );
  XOR U30814 ( .A(n30914), .B(n30923), .Z(n30938) );
  XOR U30815 ( .A(n30939), .B(n30920), .Z(n30923) );
  XOR U30816 ( .A(p_input[1398]), .B(p_input[2054]), .Z(n30920) );
  XOR U30817 ( .A(p_input[1399]), .B(n17722), .Z(n30939) );
  XOR U30818 ( .A(p_input[1394]), .B(p_input[2050]), .Z(n30914) );
  XNOR U30819 ( .A(n30929), .B(n30928), .Z(n30919) );
  XOR U30820 ( .A(n30940), .B(n30925), .Z(n30928) );
  XOR U30821 ( .A(p_input[1395]), .B(p_input[2051]), .Z(n30925) );
  XOR U30822 ( .A(p_input[1396]), .B(n17724), .Z(n30940) );
  XOR U30823 ( .A(p_input[1397]), .B(p_input[2053]), .Z(n30929) );
  XNOR U30824 ( .A(n30941), .B(n30942), .Z(n30834) );
  AND U30825 ( .A(n996), .B(n30943), .Z(n30942) );
  XNOR U30826 ( .A(n30944), .B(n30945), .Z(n996) );
  AND U30827 ( .A(n30946), .B(n30947), .Z(n30945) );
  XOR U30828 ( .A(n30944), .B(n30844), .Z(n30947) );
  XNOR U30829 ( .A(n30944), .B(n30798), .Z(n30946) );
  XOR U30830 ( .A(n30948), .B(n30949), .Z(n30944) );
  AND U30831 ( .A(n30950), .B(n30951), .Z(n30949) );
  XOR U30832 ( .A(n30948), .B(n30808), .Z(n30950) );
  XOR U30833 ( .A(n30952), .B(n30953), .Z(n30787) );
  AND U30834 ( .A(n1000), .B(n30943), .Z(n30953) );
  XNOR U30835 ( .A(n30941), .B(n30952), .Z(n30943) );
  XNOR U30836 ( .A(n30954), .B(n30955), .Z(n1000) );
  AND U30837 ( .A(n30956), .B(n30957), .Z(n30955) );
  XNOR U30838 ( .A(n30958), .B(n30954), .Z(n30957) );
  IV U30839 ( .A(n30844), .Z(n30958) );
  XNOR U30840 ( .A(n30959), .B(n30960), .Z(n30844) );
  AND U30841 ( .A(n1003), .B(n30961), .Z(n30960) );
  XNOR U30842 ( .A(n30959), .B(n30962), .Z(n30961) );
  XNOR U30843 ( .A(n30798), .B(n30954), .Z(n30956) );
  XOR U30844 ( .A(n30963), .B(n30964), .Z(n30798) );
  AND U30845 ( .A(n1011), .B(n30965), .Z(n30964) );
  XOR U30846 ( .A(n30948), .B(n30966), .Z(n30954) );
  AND U30847 ( .A(n30967), .B(n30951), .Z(n30966) );
  XNOR U30848 ( .A(n30857), .B(n30948), .Z(n30951) );
  XNOR U30849 ( .A(n30968), .B(n30969), .Z(n30857) );
  AND U30850 ( .A(n1003), .B(n30970), .Z(n30969) );
  XOR U30851 ( .A(n30971), .B(n30968), .Z(n30970) );
  XNOR U30852 ( .A(n30972), .B(n30948), .Z(n30967) );
  IV U30853 ( .A(n30808), .Z(n30972) );
  XOR U30854 ( .A(n30973), .B(n30974), .Z(n30808) );
  AND U30855 ( .A(n1011), .B(n30975), .Z(n30974) );
  XOR U30856 ( .A(n30976), .B(n30977), .Z(n30948) );
  AND U30857 ( .A(n30978), .B(n30979), .Z(n30977) );
  XNOR U30858 ( .A(n30882), .B(n30976), .Z(n30979) );
  XNOR U30859 ( .A(n30980), .B(n30981), .Z(n30882) );
  AND U30860 ( .A(n1003), .B(n30982), .Z(n30981) );
  XNOR U30861 ( .A(n30983), .B(n30980), .Z(n30982) );
  XOR U30862 ( .A(n30976), .B(n30819), .Z(n30978) );
  XOR U30863 ( .A(n30984), .B(n30985), .Z(n30819) );
  AND U30864 ( .A(n1011), .B(n30986), .Z(n30985) );
  XOR U30865 ( .A(n30987), .B(n30988), .Z(n30976) );
  AND U30866 ( .A(n30989), .B(n30990), .Z(n30988) );
  XNOR U30867 ( .A(n30987), .B(n30930), .Z(n30990) );
  XNOR U30868 ( .A(n30991), .B(n30992), .Z(n30930) );
  AND U30869 ( .A(n1003), .B(n30993), .Z(n30992) );
  XOR U30870 ( .A(n30994), .B(n30991), .Z(n30993) );
  XNOR U30871 ( .A(n30995), .B(n30987), .Z(n30989) );
  IV U30872 ( .A(n30831), .Z(n30995) );
  XOR U30873 ( .A(n30996), .B(n30997), .Z(n30831) );
  AND U30874 ( .A(n1011), .B(n30998), .Z(n30997) );
  AND U30875 ( .A(n30952), .B(n30941), .Z(n30987) );
  XNOR U30876 ( .A(n30999), .B(n31000), .Z(n30941) );
  AND U30877 ( .A(n1003), .B(n31001), .Z(n31000) );
  XNOR U30878 ( .A(n31002), .B(n30999), .Z(n31001) );
  XNOR U30879 ( .A(n31003), .B(n31004), .Z(n1003) );
  AND U30880 ( .A(n31005), .B(n31006), .Z(n31004) );
  XOR U30881 ( .A(n30962), .B(n31003), .Z(n31006) );
  AND U30882 ( .A(n31007), .B(n31008), .Z(n30962) );
  XOR U30883 ( .A(n31003), .B(n30959), .Z(n31005) );
  XNOR U30884 ( .A(n31009), .B(n31010), .Z(n30959) );
  AND U30885 ( .A(n1007), .B(n30965), .Z(n31010) );
  XOR U30886 ( .A(n30963), .B(n31009), .Z(n30965) );
  XOR U30887 ( .A(n31011), .B(n31012), .Z(n31003) );
  AND U30888 ( .A(n31013), .B(n31014), .Z(n31012) );
  XNOR U30889 ( .A(n31011), .B(n31007), .Z(n31014) );
  IV U30890 ( .A(n30971), .Z(n31007) );
  XOR U30891 ( .A(n31015), .B(n31016), .Z(n30971) );
  XOR U30892 ( .A(n31017), .B(n31008), .Z(n31016) );
  AND U30893 ( .A(n30983), .B(n31018), .Z(n31008) );
  AND U30894 ( .A(n31019), .B(n31020), .Z(n31017) );
  XOR U30895 ( .A(n31021), .B(n31015), .Z(n31019) );
  XNOR U30896 ( .A(n30968), .B(n31011), .Z(n31013) );
  XNOR U30897 ( .A(n31022), .B(n31023), .Z(n30968) );
  AND U30898 ( .A(n1007), .B(n30975), .Z(n31023) );
  XOR U30899 ( .A(n31022), .B(n30973), .Z(n30975) );
  XOR U30900 ( .A(n31024), .B(n31025), .Z(n31011) );
  AND U30901 ( .A(n31026), .B(n31027), .Z(n31025) );
  XNOR U30902 ( .A(n31024), .B(n30983), .Z(n31027) );
  XOR U30903 ( .A(n31028), .B(n31020), .Z(n30983) );
  XNOR U30904 ( .A(n31029), .B(n31015), .Z(n31020) );
  XOR U30905 ( .A(n31030), .B(n31031), .Z(n31015) );
  AND U30906 ( .A(n31032), .B(n31033), .Z(n31031) );
  XOR U30907 ( .A(n31034), .B(n31030), .Z(n31032) );
  XNOR U30908 ( .A(n31035), .B(n31036), .Z(n31029) );
  AND U30909 ( .A(n31037), .B(n31038), .Z(n31036) );
  XOR U30910 ( .A(n31035), .B(n31039), .Z(n31037) );
  XNOR U30911 ( .A(n31021), .B(n31018), .Z(n31028) );
  AND U30912 ( .A(n31040), .B(n31041), .Z(n31018) );
  XOR U30913 ( .A(n31042), .B(n31043), .Z(n31021) );
  AND U30914 ( .A(n31044), .B(n31045), .Z(n31043) );
  XOR U30915 ( .A(n31042), .B(n31046), .Z(n31044) );
  XNOR U30916 ( .A(n30980), .B(n31024), .Z(n31026) );
  XNOR U30917 ( .A(n31047), .B(n31048), .Z(n30980) );
  AND U30918 ( .A(n1007), .B(n30986), .Z(n31048) );
  XOR U30919 ( .A(n31047), .B(n30984), .Z(n30986) );
  XOR U30920 ( .A(n31049), .B(n31050), .Z(n31024) );
  AND U30921 ( .A(n31051), .B(n31052), .Z(n31050) );
  XNOR U30922 ( .A(n31049), .B(n31040), .Z(n31052) );
  IV U30923 ( .A(n30994), .Z(n31040) );
  XNOR U30924 ( .A(n31053), .B(n31033), .Z(n30994) );
  XNOR U30925 ( .A(n31054), .B(n31039), .Z(n31033) );
  XNOR U30926 ( .A(n31055), .B(n31056), .Z(n31039) );
  NOR U30927 ( .A(n31057), .B(n31058), .Z(n31056) );
  XOR U30928 ( .A(n31055), .B(n31059), .Z(n31057) );
  XNOR U30929 ( .A(n31038), .B(n31030), .Z(n31054) );
  XOR U30930 ( .A(n31060), .B(n31061), .Z(n31030) );
  AND U30931 ( .A(n31062), .B(n31063), .Z(n31061) );
  XOR U30932 ( .A(n31060), .B(n31064), .Z(n31062) );
  XNOR U30933 ( .A(n31065), .B(n31035), .Z(n31038) );
  XOR U30934 ( .A(n31066), .B(n31067), .Z(n31035) );
  AND U30935 ( .A(n31068), .B(n31069), .Z(n31067) );
  XNOR U30936 ( .A(n31070), .B(n31071), .Z(n31068) );
  IV U30937 ( .A(n31066), .Z(n31070) );
  XNOR U30938 ( .A(n31072), .B(n31073), .Z(n31065) );
  NOR U30939 ( .A(n31074), .B(n31075), .Z(n31073) );
  XNOR U30940 ( .A(n31072), .B(n31076), .Z(n31074) );
  XNOR U30941 ( .A(n31034), .B(n31041), .Z(n31053) );
  NOR U30942 ( .A(n31002), .B(n31077), .Z(n31041) );
  XOR U30943 ( .A(n31046), .B(n31045), .Z(n31034) );
  XNOR U30944 ( .A(n31078), .B(n31042), .Z(n31045) );
  XOR U30945 ( .A(n31079), .B(n31080), .Z(n31042) );
  AND U30946 ( .A(n31081), .B(n31082), .Z(n31080) );
  XNOR U30947 ( .A(n31083), .B(n31084), .Z(n31081) );
  IV U30948 ( .A(n31079), .Z(n31083) );
  XNOR U30949 ( .A(n31085), .B(n31086), .Z(n31078) );
  NOR U30950 ( .A(n31087), .B(n31088), .Z(n31086) );
  XNOR U30951 ( .A(n31085), .B(n31089), .Z(n31087) );
  XOR U30952 ( .A(n31090), .B(n31091), .Z(n31046) );
  NOR U30953 ( .A(n31092), .B(n31093), .Z(n31091) );
  XNOR U30954 ( .A(n31090), .B(n31094), .Z(n31092) );
  XNOR U30955 ( .A(n30991), .B(n31049), .Z(n31051) );
  XNOR U30956 ( .A(n31095), .B(n31096), .Z(n30991) );
  AND U30957 ( .A(n1007), .B(n30998), .Z(n31096) );
  XOR U30958 ( .A(n31095), .B(n30996), .Z(n30998) );
  AND U30959 ( .A(n30999), .B(n31002), .Z(n31049) );
  XOR U30960 ( .A(n31097), .B(n31077), .Z(n31002) );
  XNOR U30961 ( .A(p_input[1408]), .B(p_input[2048]), .Z(n31077) );
  XNOR U30962 ( .A(n31064), .B(n31063), .Z(n31097) );
  XNOR U30963 ( .A(n31098), .B(n31071), .Z(n31063) );
  XNOR U30964 ( .A(n31059), .B(n31058), .Z(n31071) );
  XNOR U30965 ( .A(n31099), .B(n31055), .Z(n31058) );
  XNOR U30966 ( .A(p_input[1418]), .B(p_input[2058]), .Z(n31055) );
  XOR U30967 ( .A(p_input[1419]), .B(n16732), .Z(n31099) );
  XOR U30968 ( .A(p_input[1420]), .B(p_input[2060]), .Z(n31059) );
  XOR U30969 ( .A(n31069), .B(n31100), .Z(n31098) );
  IV U30970 ( .A(n31060), .Z(n31100) );
  XOR U30971 ( .A(p_input[1409]), .B(p_input[2049]), .Z(n31060) );
  XNOR U30972 ( .A(n31101), .B(n31076), .Z(n31069) );
  XNOR U30973 ( .A(p_input[1423]), .B(n16735), .Z(n31076) );
  XOR U30974 ( .A(n31066), .B(n31075), .Z(n31101) );
  XOR U30975 ( .A(n31102), .B(n31072), .Z(n31075) );
  XOR U30976 ( .A(p_input[1421]), .B(p_input[2061]), .Z(n31072) );
  XOR U30977 ( .A(p_input[1422]), .B(n16737), .Z(n31102) );
  XOR U30978 ( .A(p_input[1417]), .B(p_input[2057]), .Z(n31066) );
  XOR U30979 ( .A(n31084), .B(n31082), .Z(n31064) );
  XNOR U30980 ( .A(n31103), .B(n31089), .Z(n31082) );
  XOR U30981 ( .A(p_input[1416]), .B(p_input[2056]), .Z(n31089) );
  XOR U30982 ( .A(n31079), .B(n31088), .Z(n31103) );
  XOR U30983 ( .A(n31104), .B(n31085), .Z(n31088) );
  XOR U30984 ( .A(p_input[1414]), .B(p_input[2054]), .Z(n31085) );
  XOR U30985 ( .A(p_input[1415]), .B(n17722), .Z(n31104) );
  XOR U30986 ( .A(p_input[1410]), .B(p_input[2050]), .Z(n31079) );
  XNOR U30987 ( .A(n31094), .B(n31093), .Z(n31084) );
  XOR U30988 ( .A(n31105), .B(n31090), .Z(n31093) );
  XOR U30989 ( .A(p_input[1411]), .B(p_input[2051]), .Z(n31090) );
  XOR U30990 ( .A(p_input[1412]), .B(n17724), .Z(n31105) );
  XOR U30991 ( .A(p_input[1413]), .B(p_input[2053]), .Z(n31094) );
  XNOR U30992 ( .A(n31106), .B(n31107), .Z(n30999) );
  AND U30993 ( .A(n1007), .B(n31108), .Z(n31107) );
  XNOR U30994 ( .A(n31109), .B(n31110), .Z(n1007) );
  AND U30995 ( .A(n31111), .B(n31112), .Z(n31110) );
  XOR U30996 ( .A(n31109), .B(n31009), .Z(n31112) );
  XNOR U30997 ( .A(n31109), .B(n30963), .Z(n31111) );
  XOR U30998 ( .A(n31113), .B(n31114), .Z(n31109) );
  AND U30999 ( .A(n31115), .B(n31116), .Z(n31114) );
  XOR U31000 ( .A(n31113), .B(n30973), .Z(n31115) );
  XOR U31001 ( .A(n31117), .B(n31118), .Z(n30952) );
  AND U31002 ( .A(n1011), .B(n31108), .Z(n31118) );
  XNOR U31003 ( .A(n31106), .B(n31117), .Z(n31108) );
  XNOR U31004 ( .A(n31119), .B(n31120), .Z(n1011) );
  AND U31005 ( .A(n31121), .B(n31122), .Z(n31120) );
  XNOR U31006 ( .A(n31123), .B(n31119), .Z(n31122) );
  IV U31007 ( .A(n31009), .Z(n31123) );
  XNOR U31008 ( .A(n31124), .B(n31125), .Z(n31009) );
  AND U31009 ( .A(n1014), .B(n31126), .Z(n31125) );
  XNOR U31010 ( .A(n31124), .B(n31127), .Z(n31126) );
  XNOR U31011 ( .A(n30963), .B(n31119), .Z(n31121) );
  XOR U31012 ( .A(n31128), .B(n31129), .Z(n30963) );
  AND U31013 ( .A(n1022), .B(n31130), .Z(n31129) );
  XOR U31014 ( .A(n31113), .B(n31131), .Z(n31119) );
  AND U31015 ( .A(n31132), .B(n31116), .Z(n31131) );
  XNOR U31016 ( .A(n31022), .B(n31113), .Z(n31116) );
  XNOR U31017 ( .A(n31133), .B(n31134), .Z(n31022) );
  AND U31018 ( .A(n1014), .B(n31135), .Z(n31134) );
  XOR U31019 ( .A(n31136), .B(n31133), .Z(n31135) );
  XNOR U31020 ( .A(n31137), .B(n31113), .Z(n31132) );
  IV U31021 ( .A(n30973), .Z(n31137) );
  XOR U31022 ( .A(n31138), .B(n31139), .Z(n30973) );
  AND U31023 ( .A(n1022), .B(n31140), .Z(n31139) );
  XOR U31024 ( .A(n31141), .B(n31142), .Z(n31113) );
  AND U31025 ( .A(n31143), .B(n31144), .Z(n31142) );
  XNOR U31026 ( .A(n31047), .B(n31141), .Z(n31144) );
  XNOR U31027 ( .A(n31145), .B(n31146), .Z(n31047) );
  AND U31028 ( .A(n1014), .B(n31147), .Z(n31146) );
  XNOR U31029 ( .A(n31148), .B(n31145), .Z(n31147) );
  XOR U31030 ( .A(n31141), .B(n30984), .Z(n31143) );
  XOR U31031 ( .A(n31149), .B(n31150), .Z(n30984) );
  AND U31032 ( .A(n1022), .B(n31151), .Z(n31150) );
  XOR U31033 ( .A(n31152), .B(n31153), .Z(n31141) );
  AND U31034 ( .A(n31154), .B(n31155), .Z(n31153) );
  XNOR U31035 ( .A(n31152), .B(n31095), .Z(n31155) );
  XNOR U31036 ( .A(n31156), .B(n31157), .Z(n31095) );
  AND U31037 ( .A(n1014), .B(n31158), .Z(n31157) );
  XOR U31038 ( .A(n31159), .B(n31156), .Z(n31158) );
  XNOR U31039 ( .A(n31160), .B(n31152), .Z(n31154) );
  IV U31040 ( .A(n30996), .Z(n31160) );
  XOR U31041 ( .A(n31161), .B(n31162), .Z(n30996) );
  AND U31042 ( .A(n1022), .B(n31163), .Z(n31162) );
  AND U31043 ( .A(n31117), .B(n31106), .Z(n31152) );
  XNOR U31044 ( .A(n31164), .B(n31165), .Z(n31106) );
  AND U31045 ( .A(n1014), .B(n31166), .Z(n31165) );
  XNOR U31046 ( .A(n31167), .B(n31164), .Z(n31166) );
  XNOR U31047 ( .A(n31168), .B(n31169), .Z(n1014) );
  AND U31048 ( .A(n31170), .B(n31171), .Z(n31169) );
  XOR U31049 ( .A(n31127), .B(n31168), .Z(n31171) );
  AND U31050 ( .A(n31172), .B(n31173), .Z(n31127) );
  XOR U31051 ( .A(n31168), .B(n31124), .Z(n31170) );
  XNOR U31052 ( .A(n31174), .B(n31175), .Z(n31124) );
  AND U31053 ( .A(n1018), .B(n31130), .Z(n31175) );
  XOR U31054 ( .A(n31128), .B(n31174), .Z(n31130) );
  XOR U31055 ( .A(n31176), .B(n31177), .Z(n31168) );
  AND U31056 ( .A(n31178), .B(n31179), .Z(n31177) );
  XNOR U31057 ( .A(n31176), .B(n31172), .Z(n31179) );
  IV U31058 ( .A(n31136), .Z(n31172) );
  XOR U31059 ( .A(n31180), .B(n31181), .Z(n31136) );
  XOR U31060 ( .A(n31182), .B(n31173), .Z(n31181) );
  AND U31061 ( .A(n31148), .B(n31183), .Z(n31173) );
  AND U31062 ( .A(n31184), .B(n31185), .Z(n31182) );
  XOR U31063 ( .A(n31186), .B(n31180), .Z(n31184) );
  XNOR U31064 ( .A(n31133), .B(n31176), .Z(n31178) );
  XNOR U31065 ( .A(n31187), .B(n31188), .Z(n31133) );
  AND U31066 ( .A(n1018), .B(n31140), .Z(n31188) );
  XOR U31067 ( .A(n31187), .B(n31138), .Z(n31140) );
  XOR U31068 ( .A(n31189), .B(n31190), .Z(n31176) );
  AND U31069 ( .A(n31191), .B(n31192), .Z(n31190) );
  XNOR U31070 ( .A(n31189), .B(n31148), .Z(n31192) );
  XOR U31071 ( .A(n31193), .B(n31185), .Z(n31148) );
  XNOR U31072 ( .A(n31194), .B(n31180), .Z(n31185) );
  XOR U31073 ( .A(n31195), .B(n31196), .Z(n31180) );
  AND U31074 ( .A(n31197), .B(n31198), .Z(n31196) );
  XOR U31075 ( .A(n31199), .B(n31195), .Z(n31197) );
  XNOR U31076 ( .A(n31200), .B(n31201), .Z(n31194) );
  AND U31077 ( .A(n31202), .B(n31203), .Z(n31201) );
  XOR U31078 ( .A(n31200), .B(n31204), .Z(n31202) );
  XNOR U31079 ( .A(n31186), .B(n31183), .Z(n31193) );
  AND U31080 ( .A(n31205), .B(n31206), .Z(n31183) );
  XOR U31081 ( .A(n31207), .B(n31208), .Z(n31186) );
  AND U31082 ( .A(n31209), .B(n31210), .Z(n31208) );
  XOR U31083 ( .A(n31207), .B(n31211), .Z(n31209) );
  XNOR U31084 ( .A(n31145), .B(n31189), .Z(n31191) );
  XNOR U31085 ( .A(n31212), .B(n31213), .Z(n31145) );
  AND U31086 ( .A(n1018), .B(n31151), .Z(n31213) );
  XOR U31087 ( .A(n31212), .B(n31149), .Z(n31151) );
  XOR U31088 ( .A(n31214), .B(n31215), .Z(n31189) );
  AND U31089 ( .A(n31216), .B(n31217), .Z(n31215) );
  XNOR U31090 ( .A(n31214), .B(n31205), .Z(n31217) );
  IV U31091 ( .A(n31159), .Z(n31205) );
  XNOR U31092 ( .A(n31218), .B(n31198), .Z(n31159) );
  XNOR U31093 ( .A(n31219), .B(n31204), .Z(n31198) );
  XNOR U31094 ( .A(n31220), .B(n31221), .Z(n31204) );
  NOR U31095 ( .A(n31222), .B(n31223), .Z(n31221) );
  XOR U31096 ( .A(n31220), .B(n31224), .Z(n31222) );
  XNOR U31097 ( .A(n31203), .B(n31195), .Z(n31219) );
  XOR U31098 ( .A(n31225), .B(n31226), .Z(n31195) );
  AND U31099 ( .A(n31227), .B(n31228), .Z(n31226) );
  XOR U31100 ( .A(n31225), .B(n31229), .Z(n31227) );
  XNOR U31101 ( .A(n31230), .B(n31200), .Z(n31203) );
  XOR U31102 ( .A(n31231), .B(n31232), .Z(n31200) );
  AND U31103 ( .A(n31233), .B(n31234), .Z(n31232) );
  XNOR U31104 ( .A(n31235), .B(n31236), .Z(n31233) );
  IV U31105 ( .A(n31231), .Z(n31235) );
  XNOR U31106 ( .A(n31237), .B(n31238), .Z(n31230) );
  NOR U31107 ( .A(n31239), .B(n31240), .Z(n31238) );
  XNOR U31108 ( .A(n31237), .B(n31241), .Z(n31239) );
  XNOR U31109 ( .A(n31199), .B(n31206), .Z(n31218) );
  NOR U31110 ( .A(n31167), .B(n31242), .Z(n31206) );
  XOR U31111 ( .A(n31211), .B(n31210), .Z(n31199) );
  XNOR U31112 ( .A(n31243), .B(n31207), .Z(n31210) );
  XOR U31113 ( .A(n31244), .B(n31245), .Z(n31207) );
  AND U31114 ( .A(n31246), .B(n31247), .Z(n31245) );
  XNOR U31115 ( .A(n31248), .B(n31249), .Z(n31246) );
  IV U31116 ( .A(n31244), .Z(n31248) );
  XNOR U31117 ( .A(n31250), .B(n31251), .Z(n31243) );
  NOR U31118 ( .A(n31252), .B(n31253), .Z(n31251) );
  XNOR U31119 ( .A(n31250), .B(n31254), .Z(n31252) );
  XOR U31120 ( .A(n31255), .B(n31256), .Z(n31211) );
  NOR U31121 ( .A(n31257), .B(n31258), .Z(n31256) );
  XNOR U31122 ( .A(n31255), .B(n31259), .Z(n31257) );
  XNOR U31123 ( .A(n31156), .B(n31214), .Z(n31216) );
  XNOR U31124 ( .A(n31260), .B(n31261), .Z(n31156) );
  AND U31125 ( .A(n1018), .B(n31163), .Z(n31261) );
  XOR U31126 ( .A(n31260), .B(n31161), .Z(n31163) );
  AND U31127 ( .A(n31164), .B(n31167), .Z(n31214) );
  XOR U31128 ( .A(n31262), .B(n31242), .Z(n31167) );
  XNOR U31129 ( .A(p_input[1424]), .B(p_input[2048]), .Z(n31242) );
  XNOR U31130 ( .A(n31229), .B(n31228), .Z(n31262) );
  XNOR U31131 ( .A(n31263), .B(n31236), .Z(n31228) );
  XNOR U31132 ( .A(n31224), .B(n31223), .Z(n31236) );
  XNOR U31133 ( .A(n31264), .B(n31220), .Z(n31223) );
  XNOR U31134 ( .A(p_input[1434]), .B(p_input[2058]), .Z(n31220) );
  XOR U31135 ( .A(p_input[1435]), .B(n16732), .Z(n31264) );
  XOR U31136 ( .A(p_input[1436]), .B(p_input[2060]), .Z(n31224) );
  XOR U31137 ( .A(n31234), .B(n31265), .Z(n31263) );
  IV U31138 ( .A(n31225), .Z(n31265) );
  XOR U31139 ( .A(p_input[1425]), .B(p_input[2049]), .Z(n31225) );
  XNOR U31140 ( .A(n31266), .B(n31241), .Z(n31234) );
  XNOR U31141 ( .A(p_input[1439]), .B(n16735), .Z(n31241) );
  XOR U31142 ( .A(n31231), .B(n31240), .Z(n31266) );
  XOR U31143 ( .A(n31267), .B(n31237), .Z(n31240) );
  XOR U31144 ( .A(p_input[1437]), .B(p_input[2061]), .Z(n31237) );
  XOR U31145 ( .A(p_input[1438]), .B(n16737), .Z(n31267) );
  XOR U31146 ( .A(p_input[1433]), .B(p_input[2057]), .Z(n31231) );
  XOR U31147 ( .A(n31249), .B(n31247), .Z(n31229) );
  XNOR U31148 ( .A(n31268), .B(n31254), .Z(n31247) );
  XOR U31149 ( .A(p_input[1432]), .B(p_input[2056]), .Z(n31254) );
  XOR U31150 ( .A(n31244), .B(n31253), .Z(n31268) );
  XOR U31151 ( .A(n31269), .B(n31250), .Z(n31253) );
  XOR U31152 ( .A(p_input[1430]), .B(p_input[2054]), .Z(n31250) );
  XOR U31153 ( .A(p_input[1431]), .B(n17722), .Z(n31269) );
  XOR U31154 ( .A(p_input[1426]), .B(p_input[2050]), .Z(n31244) );
  XNOR U31155 ( .A(n31259), .B(n31258), .Z(n31249) );
  XOR U31156 ( .A(n31270), .B(n31255), .Z(n31258) );
  XOR U31157 ( .A(p_input[1427]), .B(p_input[2051]), .Z(n31255) );
  XOR U31158 ( .A(p_input[1428]), .B(n17724), .Z(n31270) );
  XOR U31159 ( .A(p_input[1429]), .B(p_input[2053]), .Z(n31259) );
  XNOR U31160 ( .A(n31271), .B(n31272), .Z(n31164) );
  AND U31161 ( .A(n1018), .B(n31273), .Z(n31272) );
  XNOR U31162 ( .A(n31274), .B(n31275), .Z(n1018) );
  AND U31163 ( .A(n31276), .B(n31277), .Z(n31275) );
  XOR U31164 ( .A(n31274), .B(n31174), .Z(n31277) );
  XNOR U31165 ( .A(n31274), .B(n31128), .Z(n31276) );
  XOR U31166 ( .A(n31278), .B(n31279), .Z(n31274) );
  AND U31167 ( .A(n31280), .B(n31281), .Z(n31279) );
  XOR U31168 ( .A(n31278), .B(n31138), .Z(n31280) );
  XOR U31169 ( .A(n31282), .B(n31283), .Z(n31117) );
  AND U31170 ( .A(n1022), .B(n31273), .Z(n31283) );
  XNOR U31171 ( .A(n31271), .B(n31282), .Z(n31273) );
  XNOR U31172 ( .A(n31284), .B(n31285), .Z(n1022) );
  AND U31173 ( .A(n31286), .B(n31287), .Z(n31285) );
  XNOR U31174 ( .A(n31288), .B(n31284), .Z(n31287) );
  IV U31175 ( .A(n31174), .Z(n31288) );
  XNOR U31176 ( .A(n31289), .B(n31290), .Z(n31174) );
  AND U31177 ( .A(n1025), .B(n31291), .Z(n31290) );
  XNOR U31178 ( .A(n31289), .B(n31292), .Z(n31291) );
  XNOR U31179 ( .A(n31128), .B(n31284), .Z(n31286) );
  XOR U31180 ( .A(n31293), .B(n31294), .Z(n31128) );
  AND U31181 ( .A(n1033), .B(n31295), .Z(n31294) );
  XOR U31182 ( .A(n31278), .B(n31296), .Z(n31284) );
  AND U31183 ( .A(n31297), .B(n31281), .Z(n31296) );
  XNOR U31184 ( .A(n31187), .B(n31278), .Z(n31281) );
  XNOR U31185 ( .A(n31298), .B(n31299), .Z(n31187) );
  AND U31186 ( .A(n1025), .B(n31300), .Z(n31299) );
  XOR U31187 ( .A(n31301), .B(n31298), .Z(n31300) );
  XNOR U31188 ( .A(n31302), .B(n31278), .Z(n31297) );
  IV U31189 ( .A(n31138), .Z(n31302) );
  XOR U31190 ( .A(n31303), .B(n31304), .Z(n31138) );
  AND U31191 ( .A(n1033), .B(n31305), .Z(n31304) );
  XOR U31192 ( .A(n31306), .B(n31307), .Z(n31278) );
  AND U31193 ( .A(n31308), .B(n31309), .Z(n31307) );
  XNOR U31194 ( .A(n31212), .B(n31306), .Z(n31309) );
  XNOR U31195 ( .A(n31310), .B(n31311), .Z(n31212) );
  AND U31196 ( .A(n1025), .B(n31312), .Z(n31311) );
  XNOR U31197 ( .A(n31313), .B(n31310), .Z(n31312) );
  XOR U31198 ( .A(n31306), .B(n31149), .Z(n31308) );
  XOR U31199 ( .A(n31314), .B(n31315), .Z(n31149) );
  AND U31200 ( .A(n1033), .B(n31316), .Z(n31315) );
  XOR U31201 ( .A(n31317), .B(n31318), .Z(n31306) );
  AND U31202 ( .A(n31319), .B(n31320), .Z(n31318) );
  XNOR U31203 ( .A(n31317), .B(n31260), .Z(n31320) );
  XNOR U31204 ( .A(n31321), .B(n31322), .Z(n31260) );
  AND U31205 ( .A(n1025), .B(n31323), .Z(n31322) );
  XOR U31206 ( .A(n31324), .B(n31321), .Z(n31323) );
  XNOR U31207 ( .A(n31325), .B(n31317), .Z(n31319) );
  IV U31208 ( .A(n31161), .Z(n31325) );
  XOR U31209 ( .A(n31326), .B(n31327), .Z(n31161) );
  AND U31210 ( .A(n1033), .B(n31328), .Z(n31327) );
  AND U31211 ( .A(n31282), .B(n31271), .Z(n31317) );
  XNOR U31212 ( .A(n31329), .B(n31330), .Z(n31271) );
  AND U31213 ( .A(n1025), .B(n31331), .Z(n31330) );
  XNOR U31214 ( .A(n31332), .B(n31329), .Z(n31331) );
  XNOR U31215 ( .A(n31333), .B(n31334), .Z(n1025) );
  AND U31216 ( .A(n31335), .B(n31336), .Z(n31334) );
  XOR U31217 ( .A(n31292), .B(n31333), .Z(n31336) );
  AND U31218 ( .A(n31337), .B(n31338), .Z(n31292) );
  XOR U31219 ( .A(n31333), .B(n31289), .Z(n31335) );
  XNOR U31220 ( .A(n31339), .B(n31340), .Z(n31289) );
  AND U31221 ( .A(n1029), .B(n31295), .Z(n31340) );
  XOR U31222 ( .A(n31293), .B(n31339), .Z(n31295) );
  XOR U31223 ( .A(n31341), .B(n31342), .Z(n31333) );
  AND U31224 ( .A(n31343), .B(n31344), .Z(n31342) );
  XNOR U31225 ( .A(n31341), .B(n31337), .Z(n31344) );
  IV U31226 ( .A(n31301), .Z(n31337) );
  XOR U31227 ( .A(n31345), .B(n31346), .Z(n31301) );
  XOR U31228 ( .A(n31347), .B(n31338), .Z(n31346) );
  AND U31229 ( .A(n31313), .B(n31348), .Z(n31338) );
  AND U31230 ( .A(n31349), .B(n31350), .Z(n31347) );
  XOR U31231 ( .A(n31351), .B(n31345), .Z(n31349) );
  XNOR U31232 ( .A(n31298), .B(n31341), .Z(n31343) );
  XNOR U31233 ( .A(n31352), .B(n31353), .Z(n31298) );
  AND U31234 ( .A(n1029), .B(n31305), .Z(n31353) );
  XOR U31235 ( .A(n31352), .B(n31303), .Z(n31305) );
  XOR U31236 ( .A(n31354), .B(n31355), .Z(n31341) );
  AND U31237 ( .A(n31356), .B(n31357), .Z(n31355) );
  XNOR U31238 ( .A(n31354), .B(n31313), .Z(n31357) );
  XOR U31239 ( .A(n31358), .B(n31350), .Z(n31313) );
  XNOR U31240 ( .A(n31359), .B(n31345), .Z(n31350) );
  XOR U31241 ( .A(n31360), .B(n31361), .Z(n31345) );
  AND U31242 ( .A(n31362), .B(n31363), .Z(n31361) );
  XOR U31243 ( .A(n31364), .B(n31360), .Z(n31362) );
  XNOR U31244 ( .A(n31365), .B(n31366), .Z(n31359) );
  AND U31245 ( .A(n31367), .B(n31368), .Z(n31366) );
  XOR U31246 ( .A(n31365), .B(n31369), .Z(n31367) );
  XNOR U31247 ( .A(n31351), .B(n31348), .Z(n31358) );
  AND U31248 ( .A(n31370), .B(n31371), .Z(n31348) );
  XOR U31249 ( .A(n31372), .B(n31373), .Z(n31351) );
  AND U31250 ( .A(n31374), .B(n31375), .Z(n31373) );
  XOR U31251 ( .A(n31372), .B(n31376), .Z(n31374) );
  XNOR U31252 ( .A(n31310), .B(n31354), .Z(n31356) );
  XNOR U31253 ( .A(n31377), .B(n31378), .Z(n31310) );
  AND U31254 ( .A(n1029), .B(n31316), .Z(n31378) );
  XOR U31255 ( .A(n31377), .B(n31314), .Z(n31316) );
  XOR U31256 ( .A(n31379), .B(n31380), .Z(n31354) );
  AND U31257 ( .A(n31381), .B(n31382), .Z(n31380) );
  XNOR U31258 ( .A(n31379), .B(n31370), .Z(n31382) );
  IV U31259 ( .A(n31324), .Z(n31370) );
  XNOR U31260 ( .A(n31383), .B(n31363), .Z(n31324) );
  XNOR U31261 ( .A(n31384), .B(n31369), .Z(n31363) );
  XNOR U31262 ( .A(n31385), .B(n31386), .Z(n31369) );
  NOR U31263 ( .A(n31387), .B(n31388), .Z(n31386) );
  XOR U31264 ( .A(n31385), .B(n31389), .Z(n31387) );
  XNOR U31265 ( .A(n31368), .B(n31360), .Z(n31384) );
  XOR U31266 ( .A(n31390), .B(n31391), .Z(n31360) );
  AND U31267 ( .A(n31392), .B(n31393), .Z(n31391) );
  XOR U31268 ( .A(n31390), .B(n31394), .Z(n31392) );
  XNOR U31269 ( .A(n31395), .B(n31365), .Z(n31368) );
  XOR U31270 ( .A(n31396), .B(n31397), .Z(n31365) );
  AND U31271 ( .A(n31398), .B(n31399), .Z(n31397) );
  XNOR U31272 ( .A(n31400), .B(n31401), .Z(n31398) );
  IV U31273 ( .A(n31396), .Z(n31400) );
  XNOR U31274 ( .A(n31402), .B(n31403), .Z(n31395) );
  NOR U31275 ( .A(n31404), .B(n31405), .Z(n31403) );
  XNOR U31276 ( .A(n31402), .B(n31406), .Z(n31404) );
  XNOR U31277 ( .A(n31364), .B(n31371), .Z(n31383) );
  NOR U31278 ( .A(n31332), .B(n31407), .Z(n31371) );
  XOR U31279 ( .A(n31376), .B(n31375), .Z(n31364) );
  XNOR U31280 ( .A(n31408), .B(n31372), .Z(n31375) );
  XOR U31281 ( .A(n31409), .B(n31410), .Z(n31372) );
  AND U31282 ( .A(n31411), .B(n31412), .Z(n31410) );
  XNOR U31283 ( .A(n31413), .B(n31414), .Z(n31411) );
  IV U31284 ( .A(n31409), .Z(n31413) );
  XNOR U31285 ( .A(n31415), .B(n31416), .Z(n31408) );
  NOR U31286 ( .A(n31417), .B(n31418), .Z(n31416) );
  XNOR U31287 ( .A(n31415), .B(n31419), .Z(n31417) );
  XOR U31288 ( .A(n31420), .B(n31421), .Z(n31376) );
  NOR U31289 ( .A(n31422), .B(n31423), .Z(n31421) );
  XNOR U31290 ( .A(n31420), .B(n31424), .Z(n31422) );
  XNOR U31291 ( .A(n31321), .B(n31379), .Z(n31381) );
  XNOR U31292 ( .A(n31425), .B(n31426), .Z(n31321) );
  AND U31293 ( .A(n1029), .B(n31328), .Z(n31426) );
  XOR U31294 ( .A(n31425), .B(n31326), .Z(n31328) );
  AND U31295 ( .A(n31329), .B(n31332), .Z(n31379) );
  XOR U31296 ( .A(n31427), .B(n31407), .Z(n31332) );
  XNOR U31297 ( .A(p_input[1440]), .B(p_input[2048]), .Z(n31407) );
  XNOR U31298 ( .A(n31394), .B(n31393), .Z(n31427) );
  XNOR U31299 ( .A(n31428), .B(n31401), .Z(n31393) );
  XNOR U31300 ( .A(n31389), .B(n31388), .Z(n31401) );
  XNOR U31301 ( .A(n31429), .B(n31385), .Z(n31388) );
  XNOR U31302 ( .A(p_input[1450]), .B(p_input[2058]), .Z(n31385) );
  XOR U31303 ( .A(p_input[1451]), .B(n16732), .Z(n31429) );
  XOR U31304 ( .A(p_input[1452]), .B(p_input[2060]), .Z(n31389) );
  XOR U31305 ( .A(n31399), .B(n31430), .Z(n31428) );
  IV U31306 ( .A(n31390), .Z(n31430) );
  XOR U31307 ( .A(p_input[1441]), .B(p_input[2049]), .Z(n31390) );
  XNOR U31308 ( .A(n31431), .B(n31406), .Z(n31399) );
  XNOR U31309 ( .A(p_input[1455]), .B(n16735), .Z(n31406) );
  XOR U31310 ( .A(n31396), .B(n31405), .Z(n31431) );
  XOR U31311 ( .A(n31432), .B(n31402), .Z(n31405) );
  XOR U31312 ( .A(p_input[1453]), .B(p_input[2061]), .Z(n31402) );
  XOR U31313 ( .A(p_input[1454]), .B(n16737), .Z(n31432) );
  XOR U31314 ( .A(p_input[1449]), .B(p_input[2057]), .Z(n31396) );
  XOR U31315 ( .A(n31414), .B(n31412), .Z(n31394) );
  XNOR U31316 ( .A(n31433), .B(n31419), .Z(n31412) );
  XOR U31317 ( .A(p_input[1448]), .B(p_input[2056]), .Z(n31419) );
  XOR U31318 ( .A(n31409), .B(n31418), .Z(n31433) );
  XOR U31319 ( .A(n31434), .B(n31415), .Z(n31418) );
  XOR U31320 ( .A(p_input[1446]), .B(p_input[2054]), .Z(n31415) );
  XOR U31321 ( .A(p_input[1447]), .B(n17722), .Z(n31434) );
  XOR U31322 ( .A(p_input[1442]), .B(p_input[2050]), .Z(n31409) );
  XNOR U31323 ( .A(n31424), .B(n31423), .Z(n31414) );
  XOR U31324 ( .A(n31435), .B(n31420), .Z(n31423) );
  XOR U31325 ( .A(p_input[1443]), .B(p_input[2051]), .Z(n31420) );
  XOR U31326 ( .A(p_input[1444]), .B(n17724), .Z(n31435) );
  XOR U31327 ( .A(p_input[1445]), .B(p_input[2053]), .Z(n31424) );
  XNOR U31328 ( .A(n31436), .B(n31437), .Z(n31329) );
  AND U31329 ( .A(n1029), .B(n31438), .Z(n31437) );
  XNOR U31330 ( .A(n31439), .B(n31440), .Z(n1029) );
  AND U31331 ( .A(n31441), .B(n31442), .Z(n31440) );
  XOR U31332 ( .A(n31439), .B(n31339), .Z(n31442) );
  XNOR U31333 ( .A(n31439), .B(n31293), .Z(n31441) );
  XOR U31334 ( .A(n31443), .B(n31444), .Z(n31439) );
  AND U31335 ( .A(n31445), .B(n31446), .Z(n31444) );
  XOR U31336 ( .A(n31443), .B(n31303), .Z(n31445) );
  XOR U31337 ( .A(n31447), .B(n31448), .Z(n31282) );
  AND U31338 ( .A(n1033), .B(n31438), .Z(n31448) );
  XNOR U31339 ( .A(n31436), .B(n31447), .Z(n31438) );
  XNOR U31340 ( .A(n31449), .B(n31450), .Z(n1033) );
  AND U31341 ( .A(n31451), .B(n31452), .Z(n31450) );
  XNOR U31342 ( .A(n31453), .B(n31449), .Z(n31452) );
  IV U31343 ( .A(n31339), .Z(n31453) );
  XNOR U31344 ( .A(n31454), .B(n31455), .Z(n31339) );
  AND U31345 ( .A(n1036), .B(n31456), .Z(n31455) );
  XNOR U31346 ( .A(n31454), .B(n31457), .Z(n31456) );
  XNOR U31347 ( .A(n31293), .B(n31449), .Z(n31451) );
  XOR U31348 ( .A(n31458), .B(n31459), .Z(n31293) );
  AND U31349 ( .A(n1044), .B(n31460), .Z(n31459) );
  XOR U31350 ( .A(n31443), .B(n31461), .Z(n31449) );
  AND U31351 ( .A(n31462), .B(n31446), .Z(n31461) );
  XNOR U31352 ( .A(n31352), .B(n31443), .Z(n31446) );
  XNOR U31353 ( .A(n31463), .B(n31464), .Z(n31352) );
  AND U31354 ( .A(n1036), .B(n31465), .Z(n31464) );
  XOR U31355 ( .A(n31466), .B(n31463), .Z(n31465) );
  XNOR U31356 ( .A(n31467), .B(n31443), .Z(n31462) );
  IV U31357 ( .A(n31303), .Z(n31467) );
  XOR U31358 ( .A(n31468), .B(n31469), .Z(n31303) );
  AND U31359 ( .A(n1044), .B(n31470), .Z(n31469) );
  XOR U31360 ( .A(n31471), .B(n31472), .Z(n31443) );
  AND U31361 ( .A(n31473), .B(n31474), .Z(n31472) );
  XNOR U31362 ( .A(n31377), .B(n31471), .Z(n31474) );
  XNOR U31363 ( .A(n31475), .B(n31476), .Z(n31377) );
  AND U31364 ( .A(n1036), .B(n31477), .Z(n31476) );
  XNOR U31365 ( .A(n31478), .B(n31475), .Z(n31477) );
  XOR U31366 ( .A(n31471), .B(n31314), .Z(n31473) );
  XOR U31367 ( .A(n31479), .B(n31480), .Z(n31314) );
  AND U31368 ( .A(n1044), .B(n31481), .Z(n31480) );
  XOR U31369 ( .A(n31482), .B(n31483), .Z(n31471) );
  AND U31370 ( .A(n31484), .B(n31485), .Z(n31483) );
  XNOR U31371 ( .A(n31482), .B(n31425), .Z(n31485) );
  XNOR U31372 ( .A(n31486), .B(n31487), .Z(n31425) );
  AND U31373 ( .A(n1036), .B(n31488), .Z(n31487) );
  XOR U31374 ( .A(n31489), .B(n31486), .Z(n31488) );
  XNOR U31375 ( .A(n31490), .B(n31482), .Z(n31484) );
  IV U31376 ( .A(n31326), .Z(n31490) );
  XOR U31377 ( .A(n31491), .B(n31492), .Z(n31326) );
  AND U31378 ( .A(n1044), .B(n31493), .Z(n31492) );
  AND U31379 ( .A(n31447), .B(n31436), .Z(n31482) );
  XNOR U31380 ( .A(n31494), .B(n31495), .Z(n31436) );
  AND U31381 ( .A(n1036), .B(n31496), .Z(n31495) );
  XNOR U31382 ( .A(n31497), .B(n31494), .Z(n31496) );
  XNOR U31383 ( .A(n31498), .B(n31499), .Z(n1036) );
  AND U31384 ( .A(n31500), .B(n31501), .Z(n31499) );
  XOR U31385 ( .A(n31457), .B(n31498), .Z(n31501) );
  AND U31386 ( .A(n31502), .B(n31503), .Z(n31457) );
  XOR U31387 ( .A(n31498), .B(n31454), .Z(n31500) );
  XNOR U31388 ( .A(n31504), .B(n31505), .Z(n31454) );
  AND U31389 ( .A(n1040), .B(n31460), .Z(n31505) );
  XOR U31390 ( .A(n31458), .B(n31504), .Z(n31460) );
  XOR U31391 ( .A(n31506), .B(n31507), .Z(n31498) );
  AND U31392 ( .A(n31508), .B(n31509), .Z(n31507) );
  XNOR U31393 ( .A(n31506), .B(n31502), .Z(n31509) );
  IV U31394 ( .A(n31466), .Z(n31502) );
  XOR U31395 ( .A(n31510), .B(n31511), .Z(n31466) );
  XOR U31396 ( .A(n31512), .B(n31503), .Z(n31511) );
  AND U31397 ( .A(n31478), .B(n31513), .Z(n31503) );
  AND U31398 ( .A(n31514), .B(n31515), .Z(n31512) );
  XOR U31399 ( .A(n31516), .B(n31510), .Z(n31514) );
  XNOR U31400 ( .A(n31463), .B(n31506), .Z(n31508) );
  XNOR U31401 ( .A(n31517), .B(n31518), .Z(n31463) );
  AND U31402 ( .A(n1040), .B(n31470), .Z(n31518) );
  XOR U31403 ( .A(n31517), .B(n31468), .Z(n31470) );
  XOR U31404 ( .A(n31519), .B(n31520), .Z(n31506) );
  AND U31405 ( .A(n31521), .B(n31522), .Z(n31520) );
  XNOR U31406 ( .A(n31519), .B(n31478), .Z(n31522) );
  XOR U31407 ( .A(n31523), .B(n31515), .Z(n31478) );
  XNOR U31408 ( .A(n31524), .B(n31510), .Z(n31515) );
  XOR U31409 ( .A(n31525), .B(n31526), .Z(n31510) );
  AND U31410 ( .A(n31527), .B(n31528), .Z(n31526) );
  XOR U31411 ( .A(n31529), .B(n31525), .Z(n31527) );
  XNOR U31412 ( .A(n31530), .B(n31531), .Z(n31524) );
  AND U31413 ( .A(n31532), .B(n31533), .Z(n31531) );
  XOR U31414 ( .A(n31530), .B(n31534), .Z(n31532) );
  XNOR U31415 ( .A(n31516), .B(n31513), .Z(n31523) );
  AND U31416 ( .A(n31535), .B(n31536), .Z(n31513) );
  XOR U31417 ( .A(n31537), .B(n31538), .Z(n31516) );
  AND U31418 ( .A(n31539), .B(n31540), .Z(n31538) );
  XOR U31419 ( .A(n31537), .B(n31541), .Z(n31539) );
  XNOR U31420 ( .A(n31475), .B(n31519), .Z(n31521) );
  XNOR U31421 ( .A(n31542), .B(n31543), .Z(n31475) );
  AND U31422 ( .A(n1040), .B(n31481), .Z(n31543) );
  XOR U31423 ( .A(n31542), .B(n31479), .Z(n31481) );
  XOR U31424 ( .A(n31544), .B(n31545), .Z(n31519) );
  AND U31425 ( .A(n31546), .B(n31547), .Z(n31545) );
  XNOR U31426 ( .A(n31544), .B(n31535), .Z(n31547) );
  IV U31427 ( .A(n31489), .Z(n31535) );
  XNOR U31428 ( .A(n31548), .B(n31528), .Z(n31489) );
  XNOR U31429 ( .A(n31549), .B(n31534), .Z(n31528) );
  XNOR U31430 ( .A(n31550), .B(n31551), .Z(n31534) );
  NOR U31431 ( .A(n31552), .B(n31553), .Z(n31551) );
  XOR U31432 ( .A(n31550), .B(n31554), .Z(n31552) );
  XNOR U31433 ( .A(n31533), .B(n31525), .Z(n31549) );
  XOR U31434 ( .A(n31555), .B(n31556), .Z(n31525) );
  AND U31435 ( .A(n31557), .B(n31558), .Z(n31556) );
  XOR U31436 ( .A(n31555), .B(n31559), .Z(n31557) );
  XNOR U31437 ( .A(n31560), .B(n31530), .Z(n31533) );
  XOR U31438 ( .A(n31561), .B(n31562), .Z(n31530) );
  AND U31439 ( .A(n31563), .B(n31564), .Z(n31562) );
  XNOR U31440 ( .A(n31565), .B(n31566), .Z(n31563) );
  IV U31441 ( .A(n31561), .Z(n31565) );
  XNOR U31442 ( .A(n31567), .B(n31568), .Z(n31560) );
  NOR U31443 ( .A(n31569), .B(n31570), .Z(n31568) );
  XNOR U31444 ( .A(n31567), .B(n31571), .Z(n31569) );
  XNOR U31445 ( .A(n31529), .B(n31536), .Z(n31548) );
  NOR U31446 ( .A(n31497), .B(n31572), .Z(n31536) );
  XOR U31447 ( .A(n31541), .B(n31540), .Z(n31529) );
  XNOR U31448 ( .A(n31573), .B(n31537), .Z(n31540) );
  XOR U31449 ( .A(n31574), .B(n31575), .Z(n31537) );
  AND U31450 ( .A(n31576), .B(n31577), .Z(n31575) );
  XNOR U31451 ( .A(n31578), .B(n31579), .Z(n31576) );
  IV U31452 ( .A(n31574), .Z(n31578) );
  XNOR U31453 ( .A(n31580), .B(n31581), .Z(n31573) );
  NOR U31454 ( .A(n31582), .B(n31583), .Z(n31581) );
  XNOR U31455 ( .A(n31580), .B(n31584), .Z(n31582) );
  XOR U31456 ( .A(n31585), .B(n31586), .Z(n31541) );
  NOR U31457 ( .A(n31587), .B(n31588), .Z(n31586) );
  XNOR U31458 ( .A(n31585), .B(n31589), .Z(n31587) );
  XNOR U31459 ( .A(n31486), .B(n31544), .Z(n31546) );
  XNOR U31460 ( .A(n31590), .B(n31591), .Z(n31486) );
  AND U31461 ( .A(n1040), .B(n31493), .Z(n31591) );
  XOR U31462 ( .A(n31590), .B(n31491), .Z(n31493) );
  AND U31463 ( .A(n31494), .B(n31497), .Z(n31544) );
  XOR U31464 ( .A(n31592), .B(n31572), .Z(n31497) );
  XNOR U31465 ( .A(p_input[1456]), .B(p_input[2048]), .Z(n31572) );
  XNOR U31466 ( .A(n31559), .B(n31558), .Z(n31592) );
  XNOR U31467 ( .A(n31593), .B(n31566), .Z(n31558) );
  XNOR U31468 ( .A(n31554), .B(n31553), .Z(n31566) );
  XNOR U31469 ( .A(n31594), .B(n31550), .Z(n31553) );
  XNOR U31470 ( .A(p_input[1466]), .B(p_input[2058]), .Z(n31550) );
  XOR U31471 ( .A(p_input[1467]), .B(n16732), .Z(n31594) );
  XOR U31472 ( .A(p_input[1468]), .B(p_input[2060]), .Z(n31554) );
  XOR U31473 ( .A(n31564), .B(n31595), .Z(n31593) );
  IV U31474 ( .A(n31555), .Z(n31595) );
  XOR U31475 ( .A(p_input[1457]), .B(p_input[2049]), .Z(n31555) );
  XNOR U31476 ( .A(n31596), .B(n31571), .Z(n31564) );
  XNOR U31477 ( .A(p_input[1471]), .B(n16735), .Z(n31571) );
  XOR U31478 ( .A(n31561), .B(n31570), .Z(n31596) );
  XOR U31479 ( .A(n31597), .B(n31567), .Z(n31570) );
  XOR U31480 ( .A(p_input[1469]), .B(p_input[2061]), .Z(n31567) );
  XOR U31481 ( .A(p_input[1470]), .B(n16737), .Z(n31597) );
  XOR U31482 ( .A(p_input[1465]), .B(p_input[2057]), .Z(n31561) );
  XOR U31483 ( .A(n31579), .B(n31577), .Z(n31559) );
  XNOR U31484 ( .A(n31598), .B(n31584), .Z(n31577) );
  XOR U31485 ( .A(p_input[1464]), .B(p_input[2056]), .Z(n31584) );
  XOR U31486 ( .A(n31574), .B(n31583), .Z(n31598) );
  XOR U31487 ( .A(n31599), .B(n31580), .Z(n31583) );
  XOR U31488 ( .A(p_input[1462]), .B(p_input[2054]), .Z(n31580) );
  XOR U31489 ( .A(p_input[1463]), .B(n17722), .Z(n31599) );
  XOR U31490 ( .A(p_input[1458]), .B(p_input[2050]), .Z(n31574) );
  XNOR U31491 ( .A(n31589), .B(n31588), .Z(n31579) );
  XOR U31492 ( .A(n31600), .B(n31585), .Z(n31588) );
  XOR U31493 ( .A(p_input[1459]), .B(p_input[2051]), .Z(n31585) );
  XOR U31494 ( .A(p_input[1460]), .B(n17724), .Z(n31600) );
  XOR U31495 ( .A(p_input[1461]), .B(p_input[2053]), .Z(n31589) );
  XNOR U31496 ( .A(n31601), .B(n31602), .Z(n31494) );
  AND U31497 ( .A(n1040), .B(n31603), .Z(n31602) );
  XNOR U31498 ( .A(n31604), .B(n31605), .Z(n1040) );
  AND U31499 ( .A(n31606), .B(n31607), .Z(n31605) );
  XOR U31500 ( .A(n31604), .B(n31504), .Z(n31607) );
  XNOR U31501 ( .A(n31604), .B(n31458), .Z(n31606) );
  XOR U31502 ( .A(n31608), .B(n31609), .Z(n31604) );
  AND U31503 ( .A(n31610), .B(n31611), .Z(n31609) );
  XOR U31504 ( .A(n31608), .B(n31468), .Z(n31610) );
  XOR U31505 ( .A(n31612), .B(n31613), .Z(n31447) );
  AND U31506 ( .A(n1044), .B(n31603), .Z(n31613) );
  XNOR U31507 ( .A(n31601), .B(n31612), .Z(n31603) );
  XNOR U31508 ( .A(n31614), .B(n31615), .Z(n1044) );
  AND U31509 ( .A(n31616), .B(n31617), .Z(n31615) );
  XNOR U31510 ( .A(n31618), .B(n31614), .Z(n31617) );
  IV U31511 ( .A(n31504), .Z(n31618) );
  XNOR U31512 ( .A(n31619), .B(n31620), .Z(n31504) );
  AND U31513 ( .A(n1047), .B(n31621), .Z(n31620) );
  XNOR U31514 ( .A(n31619), .B(n31622), .Z(n31621) );
  XNOR U31515 ( .A(n31458), .B(n31614), .Z(n31616) );
  XOR U31516 ( .A(n31623), .B(n31624), .Z(n31458) );
  AND U31517 ( .A(n1055), .B(n31625), .Z(n31624) );
  XOR U31518 ( .A(n31608), .B(n31626), .Z(n31614) );
  AND U31519 ( .A(n31627), .B(n31611), .Z(n31626) );
  XNOR U31520 ( .A(n31517), .B(n31608), .Z(n31611) );
  XNOR U31521 ( .A(n31628), .B(n31629), .Z(n31517) );
  AND U31522 ( .A(n1047), .B(n31630), .Z(n31629) );
  XOR U31523 ( .A(n31631), .B(n31628), .Z(n31630) );
  XNOR U31524 ( .A(n31632), .B(n31608), .Z(n31627) );
  IV U31525 ( .A(n31468), .Z(n31632) );
  XOR U31526 ( .A(n31633), .B(n31634), .Z(n31468) );
  AND U31527 ( .A(n1055), .B(n31635), .Z(n31634) );
  XOR U31528 ( .A(n31636), .B(n31637), .Z(n31608) );
  AND U31529 ( .A(n31638), .B(n31639), .Z(n31637) );
  XNOR U31530 ( .A(n31542), .B(n31636), .Z(n31639) );
  XNOR U31531 ( .A(n31640), .B(n31641), .Z(n31542) );
  AND U31532 ( .A(n1047), .B(n31642), .Z(n31641) );
  XNOR U31533 ( .A(n31643), .B(n31640), .Z(n31642) );
  XOR U31534 ( .A(n31636), .B(n31479), .Z(n31638) );
  XOR U31535 ( .A(n31644), .B(n31645), .Z(n31479) );
  AND U31536 ( .A(n1055), .B(n31646), .Z(n31645) );
  XOR U31537 ( .A(n31647), .B(n31648), .Z(n31636) );
  AND U31538 ( .A(n31649), .B(n31650), .Z(n31648) );
  XNOR U31539 ( .A(n31647), .B(n31590), .Z(n31650) );
  XNOR U31540 ( .A(n31651), .B(n31652), .Z(n31590) );
  AND U31541 ( .A(n1047), .B(n31653), .Z(n31652) );
  XOR U31542 ( .A(n31654), .B(n31651), .Z(n31653) );
  XNOR U31543 ( .A(n31655), .B(n31647), .Z(n31649) );
  IV U31544 ( .A(n31491), .Z(n31655) );
  XOR U31545 ( .A(n31656), .B(n31657), .Z(n31491) );
  AND U31546 ( .A(n1055), .B(n31658), .Z(n31657) );
  AND U31547 ( .A(n31612), .B(n31601), .Z(n31647) );
  XNOR U31548 ( .A(n31659), .B(n31660), .Z(n31601) );
  AND U31549 ( .A(n1047), .B(n31661), .Z(n31660) );
  XNOR U31550 ( .A(n31662), .B(n31659), .Z(n31661) );
  XNOR U31551 ( .A(n31663), .B(n31664), .Z(n1047) );
  AND U31552 ( .A(n31665), .B(n31666), .Z(n31664) );
  XOR U31553 ( .A(n31622), .B(n31663), .Z(n31666) );
  AND U31554 ( .A(n31667), .B(n31668), .Z(n31622) );
  XOR U31555 ( .A(n31663), .B(n31619), .Z(n31665) );
  XNOR U31556 ( .A(n31669), .B(n31670), .Z(n31619) );
  AND U31557 ( .A(n1051), .B(n31625), .Z(n31670) );
  XOR U31558 ( .A(n31623), .B(n31669), .Z(n31625) );
  XOR U31559 ( .A(n31671), .B(n31672), .Z(n31663) );
  AND U31560 ( .A(n31673), .B(n31674), .Z(n31672) );
  XNOR U31561 ( .A(n31671), .B(n31667), .Z(n31674) );
  IV U31562 ( .A(n31631), .Z(n31667) );
  XOR U31563 ( .A(n31675), .B(n31676), .Z(n31631) );
  XOR U31564 ( .A(n31677), .B(n31668), .Z(n31676) );
  AND U31565 ( .A(n31643), .B(n31678), .Z(n31668) );
  AND U31566 ( .A(n31679), .B(n31680), .Z(n31677) );
  XOR U31567 ( .A(n31681), .B(n31675), .Z(n31679) );
  XNOR U31568 ( .A(n31628), .B(n31671), .Z(n31673) );
  XNOR U31569 ( .A(n31682), .B(n31683), .Z(n31628) );
  AND U31570 ( .A(n1051), .B(n31635), .Z(n31683) );
  XOR U31571 ( .A(n31682), .B(n31633), .Z(n31635) );
  XOR U31572 ( .A(n31684), .B(n31685), .Z(n31671) );
  AND U31573 ( .A(n31686), .B(n31687), .Z(n31685) );
  XNOR U31574 ( .A(n31684), .B(n31643), .Z(n31687) );
  XOR U31575 ( .A(n31688), .B(n31680), .Z(n31643) );
  XNOR U31576 ( .A(n31689), .B(n31675), .Z(n31680) );
  XOR U31577 ( .A(n31690), .B(n31691), .Z(n31675) );
  AND U31578 ( .A(n31692), .B(n31693), .Z(n31691) );
  XOR U31579 ( .A(n31694), .B(n31690), .Z(n31692) );
  XNOR U31580 ( .A(n31695), .B(n31696), .Z(n31689) );
  AND U31581 ( .A(n31697), .B(n31698), .Z(n31696) );
  XOR U31582 ( .A(n31695), .B(n31699), .Z(n31697) );
  XNOR U31583 ( .A(n31681), .B(n31678), .Z(n31688) );
  AND U31584 ( .A(n31700), .B(n31701), .Z(n31678) );
  XOR U31585 ( .A(n31702), .B(n31703), .Z(n31681) );
  AND U31586 ( .A(n31704), .B(n31705), .Z(n31703) );
  XOR U31587 ( .A(n31702), .B(n31706), .Z(n31704) );
  XNOR U31588 ( .A(n31640), .B(n31684), .Z(n31686) );
  XNOR U31589 ( .A(n31707), .B(n31708), .Z(n31640) );
  AND U31590 ( .A(n1051), .B(n31646), .Z(n31708) );
  XOR U31591 ( .A(n31707), .B(n31644), .Z(n31646) );
  XOR U31592 ( .A(n31709), .B(n31710), .Z(n31684) );
  AND U31593 ( .A(n31711), .B(n31712), .Z(n31710) );
  XNOR U31594 ( .A(n31709), .B(n31700), .Z(n31712) );
  IV U31595 ( .A(n31654), .Z(n31700) );
  XNOR U31596 ( .A(n31713), .B(n31693), .Z(n31654) );
  XNOR U31597 ( .A(n31714), .B(n31699), .Z(n31693) );
  XNOR U31598 ( .A(n31715), .B(n31716), .Z(n31699) );
  NOR U31599 ( .A(n31717), .B(n31718), .Z(n31716) );
  XOR U31600 ( .A(n31715), .B(n31719), .Z(n31717) );
  XNOR U31601 ( .A(n31698), .B(n31690), .Z(n31714) );
  XOR U31602 ( .A(n31720), .B(n31721), .Z(n31690) );
  AND U31603 ( .A(n31722), .B(n31723), .Z(n31721) );
  XOR U31604 ( .A(n31720), .B(n31724), .Z(n31722) );
  XNOR U31605 ( .A(n31725), .B(n31695), .Z(n31698) );
  XOR U31606 ( .A(n31726), .B(n31727), .Z(n31695) );
  AND U31607 ( .A(n31728), .B(n31729), .Z(n31727) );
  XNOR U31608 ( .A(n31730), .B(n31731), .Z(n31728) );
  IV U31609 ( .A(n31726), .Z(n31730) );
  XNOR U31610 ( .A(n31732), .B(n31733), .Z(n31725) );
  NOR U31611 ( .A(n31734), .B(n31735), .Z(n31733) );
  XNOR U31612 ( .A(n31732), .B(n31736), .Z(n31734) );
  XNOR U31613 ( .A(n31694), .B(n31701), .Z(n31713) );
  NOR U31614 ( .A(n31662), .B(n31737), .Z(n31701) );
  XOR U31615 ( .A(n31706), .B(n31705), .Z(n31694) );
  XNOR U31616 ( .A(n31738), .B(n31702), .Z(n31705) );
  XOR U31617 ( .A(n31739), .B(n31740), .Z(n31702) );
  AND U31618 ( .A(n31741), .B(n31742), .Z(n31740) );
  XNOR U31619 ( .A(n31743), .B(n31744), .Z(n31741) );
  IV U31620 ( .A(n31739), .Z(n31743) );
  XNOR U31621 ( .A(n31745), .B(n31746), .Z(n31738) );
  NOR U31622 ( .A(n31747), .B(n31748), .Z(n31746) );
  XNOR U31623 ( .A(n31745), .B(n31749), .Z(n31747) );
  XOR U31624 ( .A(n31750), .B(n31751), .Z(n31706) );
  NOR U31625 ( .A(n31752), .B(n31753), .Z(n31751) );
  XNOR U31626 ( .A(n31750), .B(n31754), .Z(n31752) );
  XNOR U31627 ( .A(n31651), .B(n31709), .Z(n31711) );
  XNOR U31628 ( .A(n31755), .B(n31756), .Z(n31651) );
  AND U31629 ( .A(n1051), .B(n31658), .Z(n31756) );
  XOR U31630 ( .A(n31755), .B(n31656), .Z(n31658) );
  AND U31631 ( .A(n31659), .B(n31662), .Z(n31709) );
  XOR U31632 ( .A(n31757), .B(n31737), .Z(n31662) );
  XNOR U31633 ( .A(p_input[1472]), .B(p_input[2048]), .Z(n31737) );
  XNOR U31634 ( .A(n31724), .B(n31723), .Z(n31757) );
  XNOR U31635 ( .A(n31758), .B(n31731), .Z(n31723) );
  XNOR U31636 ( .A(n31719), .B(n31718), .Z(n31731) );
  XNOR U31637 ( .A(n31759), .B(n31715), .Z(n31718) );
  XNOR U31638 ( .A(p_input[1482]), .B(p_input[2058]), .Z(n31715) );
  XOR U31639 ( .A(p_input[1483]), .B(n16732), .Z(n31759) );
  XOR U31640 ( .A(p_input[1484]), .B(p_input[2060]), .Z(n31719) );
  XOR U31641 ( .A(n31729), .B(n31760), .Z(n31758) );
  IV U31642 ( .A(n31720), .Z(n31760) );
  XOR U31643 ( .A(p_input[1473]), .B(p_input[2049]), .Z(n31720) );
  XNOR U31644 ( .A(n31761), .B(n31736), .Z(n31729) );
  XNOR U31645 ( .A(p_input[1487]), .B(n16735), .Z(n31736) );
  XOR U31646 ( .A(n31726), .B(n31735), .Z(n31761) );
  XOR U31647 ( .A(n31762), .B(n31732), .Z(n31735) );
  XOR U31648 ( .A(p_input[1485]), .B(p_input[2061]), .Z(n31732) );
  XOR U31649 ( .A(p_input[1486]), .B(n16737), .Z(n31762) );
  XOR U31650 ( .A(p_input[1481]), .B(p_input[2057]), .Z(n31726) );
  XOR U31651 ( .A(n31744), .B(n31742), .Z(n31724) );
  XNOR U31652 ( .A(n31763), .B(n31749), .Z(n31742) );
  XOR U31653 ( .A(p_input[1480]), .B(p_input[2056]), .Z(n31749) );
  XOR U31654 ( .A(n31739), .B(n31748), .Z(n31763) );
  XOR U31655 ( .A(n31764), .B(n31745), .Z(n31748) );
  XOR U31656 ( .A(p_input[1478]), .B(p_input[2054]), .Z(n31745) );
  XOR U31657 ( .A(p_input[1479]), .B(n17722), .Z(n31764) );
  XOR U31658 ( .A(p_input[1474]), .B(p_input[2050]), .Z(n31739) );
  XNOR U31659 ( .A(n31754), .B(n31753), .Z(n31744) );
  XOR U31660 ( .A(n31765), .B(n31750), .Z(n31753) );
  XOR U31661 ( .A(p_input[1475]), .B(p_input[2051]), .Z(n31750) );
  XOR U31662 ( .A(p_input[1476]), .B(n17724), .Z(n31765) );
  XOR U31663 ( .A(p_input[1477]), .B(p_input[2053]), .Z(n31754) );
  XNOR U31664 ( .A(n31766), .B(n31767), .Z(n31659) );
  AND U31665 ( .A(n1051), .B(n31768), .Z(n31767) );
  XNOR U31666 ( .A(n31769), .B(n31770), .Z(n1051) );
  AND U31667 ( .A(n31771), .B(n31772), .Z(n31770) );
  XOR U31668 ( .A(n31769), .B(n31669), .Z(n31772) );
  XNOR U31669 ( .A(n31769), .B(n31623), .Z(n31771) );
  XOR U31670 ( .A(n31773), .B(n31774), .Z(n31769) );
  AND U31671 ( .A(n31775), .B(n31776), .Z(n31774) );
  XOR U31672 ( .A(n31773), .B(n31633), .Z(n31775) );
  XOR U31673 ( .A(n31777), .B(n31778), .Z(n31612) );
  AND U31674 ( .A(n1055), .B(n31768), .Z(n31778) );
  XNOR U31675 ( .A(n31766), .B(n31777), .Z(n31768) );
  XNOR U31676 ( .A(n31779), .B(n31780), .Z(n1055) );
  AND U31677 ( .A(n31781), .B(n31782), .Z(n31780) );
  XNOR U31678 ( .A(n31783), .B(n31779), .Z(n31782) );
  IV U31679 ( .A(n31669), .Z(n31783) );
  XNOR U31680 ( .A(n31784), .B(n31785), .Z(n31669) );
  AND U31681 ( .A(n1058), .B(n31786), .Z(n31785) );
  XNOR U31682 ( .A(n31784), .B(n31787), .Z(n31786) );
  XNOR U31683 ( .A(n31623), .B(n31779), .Z(n31781) );
  XOR U31684 ( .A(n31788), .B(n31789), .Z(n31623) );
  AND U31685 ( .A(n1066), .B(n31790), .Z(n31789) );
  XOR U31686 ( .A(n31773), .B(n31791), .Z(n31779) );
  AND U31687 ( .A(n31792), .B(n31776), .Z(n31791) );
  XNOR U31688 ( .A(n31682), .B(n31773), .Z(n31776) );
  XNOR U31689 ( .A(n31793), .B(n31794), .Z(n31682) );
  AND U31690 ( .A(n1058), .B(n31795), .Z(n31794) );
  XOR U31691 ( .A(n31796), .B(n31793), .Z(n31795) );
  XNOR U31692 ( .A(n31797), .B(n31773), .Z(n31792) );
  IV U31693 ( .A(n31633), .Z(n31797) );
  XOR U31694 ( .A(n31798), .B(n31799), .Z(n31633) );
  AND U31695 ( .A(n1066), .B(n31800), .Z(n31799) );
  XOR U31696 ( .A(n31801), .B(n31802), .Z(n31773) );
  AND U31697 ( .A(n31803), .B(n31804), .Z(n31802) );
  XNOR U31698 ( .A(n31707), .B(n31801), .Z(n31804) );
  XNOR U31699 ( .A(n31805), .B(n31806), .Z(n31707) );
  AND U31700 ( .A(n1058), .B(n31807), .Z(n31806) );
  XNOR U31701 ( .A(n31808), .B(n31805), .Z(n31807) );
  XOR U31702 ( .A(n31801), .B(n31644), .Z(n31803) );
  XOR U31703 ( .A(n31809), .B(n31810), .Z(n31644) );
  AND U31704 ( .A(n1066), .B(n31811), .Z(n31810) );
  XOR U31705 ( .A(n31812), .B(n31813), .Z(n31801) );
  AND U31706 ( .A(n31814), .B(n31815), .Z(n31813) );
  XNOR U31707 ( .A(n31812), .B(n31755), .Z(n31815) );
  XNOR U31708 ( .A(n31816), .B(n31817), .Z(n31755) );
  AND U31709 ( .A(n1058), .B(n31818), .Z(n31817) );
  XOR U31710 ( .A(n31819), .B(n31816), .Z(n31818) );
  XNOR U31711 ( .A(n31820), .B(n31812), .Z(n31814) );
  IV U31712 ( .A(n31656), .Z(n31820) );
  XOR U31713 ( .A(n31821), .B(n31822), .Z(n31656) );
  AND U31714 ( .A(n1066), .B(n31823), .Z(n31822) );
  AND U31715 ( .A(n31777), .B(n31766), .Z(n31812) );
  XNOR U31716 ( .A(n31824), .B(n31825), .Z(n31766) );
  AND U31717 ( .A(n1058), .B(n31826), .Z(n31825) );
  XNOR U31718 ( .A(n31827), .B(n31824), .Z(n31826) );
  XNOR U31719 ( .A(n31828), .B(n31829), .Z(n1058) );
  AND U31720 ( .A(n31830), .B(n31831), .Z(n31829) );
  XOR U31721 ( .A(n31787), .B(n31828), .Z(n31831) );
  AND U31722 ( .A(n31832), .B(n31833), .Z(n31787) );
  XOR U31723 ( .A(n31828), .B(n31784), .Z(n31830) );
  XNOR U31724 ( .A(n31834), .B(n31835), .Z(n31784) );
  AND U31725 ( .A(n1062), .B(n31790), .Z(n31835) );
  XOR U31726 ( .A(n31788), .B(n31834), .Z(n31790) );
  XOR U31727 ( .A(n31836), .B(n31837), .Z(n31828) );
  AND U31728 ( .A(n31838), .B(n31839), .Z(n31837) );
  XNOR U31729 ( .A(n31836), .B(n31832), .Z(n31839) );
  IV U31730 ( .A(n31796), .Z(n31832) );
  XOR U31731 ( .A(n31840), .B(n31841), .Z(n31796) );
  XOR U31732 ( .A(n31842), .B(n31833), .Z(n31841) );
  AND U31733 ( .A(n31808), .B(n31843), .Z(n31833) );
  AND U31734 ( .A(n31844), .B(n31845), .Z(n31842) );
  XOR U31735 ( .A(n31846), .B(n31840), .Z(n31844) );
  XNOR U31736 ( .A(n31793), .B(n31836), .Z(n31838) );
  XNOR U31737 ( .A(n31847), .B(n31848), .Z(n31793) );
  AND U31738 ( .A(n1062), .B(n31800), .Z(n31848) );
  XOR U31739 ( .A(n31847), .B(n31798), .Z(n31800) );
  XOR U31740 ( .A(n31849), .B(n31850), .Z(n31836) );
  AND U31741 ( .A(n31851), .B(n31852), .Z(n31850) );
  XNOR U31742 ( .A(n31849), .B(n31808), .Z(n31852) );
  XOR U31743 ( .A(n31853), .B(n31845), .Z(n31808) );
  XNOR U31744 ( .A(n31854), .B(n31840), .Z(n31845) );
  XOR U31745 ( .A(n31855), .B(n31856), .Z(n31840) );
  AND U31746 ( .A(n31857), .B(n31858), .Z(n31856) );
  XOR U31747 ( .A(n31859), .B(n31855), .Z(n31857) );
  XNOR U31748 ( .A(n31860), .B(n31861), .Z(n31854) );
  AND U31749 ( .A(n31862), .B(n31863), .Z(n31861) );
  XOR U31750 ( .A(n31860), .B(n31864), .Z(n31862) );
  XNOR U31751 ( .A(n31846), .B(n31843), .Z(n31853) );
  AND U31752 ( .A(n31865), .B(n31866), .Z(n31843) );
  XOR U31753 ( .A(n31867), .B(n31868), .Z(n31846) );
  AND U31754 ( .A(n31869), .B(n31870), .Z(n31868) );
  XOR U31755 ( .A(n31867), .B(n31871), .Z(n31869) );
  XNOR U31756 ( .A(n31805), .B(n31849), .Z(n31851) );
  XNOR U31757 ( .A(n31872), .B(n31873), .Z(n31805) );
  AND U31758 ( .A(n1062), .B(n31811), .Z(n31873) );
  XOR U31759 ( .A(n31872), .B(n31809), .Z(n31811) );
  XOR U31760 ( .A(n31874), .B(n31875), .Z(n31849) );
  AND U31761 ( .A(n31876), .B(n31877), .Z(n31875) );
  XNOR U31762 ( .A(n31874), .B(n31865), .Z(n31877) );
  IV U31763 ( .A(n31819), .Z(n31865) );
  XNOR U31764 ( .A(n31878), .B(n31858), .Z(n31819) );
  XNOR U31765 ( .A(n31879), .B(n31864), .Z(n31858) );
  XNOR U31766 ( .A(n31880), .B(n31881), .Z(n31864) );
  NOR U31767 ( .A(n31882), .B(n31883), .Z(n31881) );
  XOR U31768 ( .A(n31880), .B(n31884), .Z(n31882) );
  XNOR U31769 ( .A(n31863), .B(n31855), .Z(n31879) );
  XOR U31770 ( .A(n31885), .B(n31886), .Z(n31855) );
  AND U31771 ( .A(n31887), .B(n31888), .Z(n31886) );
  XOR U31772 ( .A(n31885), .B(n31889), .Z(n31887) );
  XNOR U31773 ( .A(n31890), .B(n31860), .Z(n31863) );
  XOR U31774 ( .A(n31891), .B(n31892), .Z(n31860) );
  AND U31775 ( .A(n31893), .B(n31894), .Z(n31892) );
  XNOR U31776 ( .A(n31895), .B(n31896), .Z(n31893) );
  IV U31777 ( .A(n31891), .Z(n31895) );
  XNOR U31778 ( .A(n31897), .B(n31898), .Z(n31890) );
  NOR U31779 ( .A(n31899), .B(n31900), .Z(n31898) );
  XNOR U31780 ( .A(n31897), .B(n31901), .Z(n31899) );
  XNOR U31781 ( .A(n31859), .B(n31866), .Z(n31878) );
  NOR U31782 ( .A(n31827), .B(n31902), .Z(n31866) );
  XOR U31783 ( .A(n31871), .B(n31870), .Z(n31859) );
  XNOR U31784 ( .A(n31903), .B(n31867), .Z(n31870) );
  XOR U31785 ( .A(n31904), .B(n31905), .Z(n31867) );
  AND U31786 ( .A(n31906), .B(n31907), .Z(n31905) );
  XNOR U31787 ( .A(n31908), .B(n31909), .Z(n31906) );
  IV U31788 ( .A(n31904), .Z(n31908) );
  XNOR U31789 ( .A(n31910), .B(n31911), .Z(n31903) );
  NOR U31790 ( .A(n31912), .B(n31913), .Z(n31911) );
  XNOR U31791 ( .A(n31910), .B(n31914), .Z(n31912) );
  XOR U31792 ( .A(n31915), .B(n31916), .Z(n31871) );
  NOR U31793 ( .A(n31917), .B(n31918), .Z(n31916) );
  XNOR U31794 ( .A(n31915), .B(n31919), .Z(n31917) );
  XNOR U31795 ( .A(n31816), .B(n31874), .Z(n31876) );
  XNOR U31796 ( .A(n31920), .B(n31921), .Z(n31816) );
  AND U31797 ( .A(n1062), .B(n31823), .Z(n31921) );
  XOR U31798 ( .A(n31920), .B(n31821), .Z(n31823) );
  AND U31799 ( .A(n31824), .B(n31827), .Z(n31874) );
  XOR U31800 ( .A(n31922), .B(n31902), .Z(n31827) );
  XNOR U31801 ( .A(p_input[1488]), .B(p_input[2048]), .Z(n31902) );
  XNOR U31802 ( .A(n31889), .B(n31888), .Z(n31922) );
  XNOR U31803 ( .A(n31923), .B(n31896), .Z(n31888) );
  XNOR U31804 ( .A(n31884), .B(n31883), .Z(n31896) );
  XNOR U31805 ( .A(n31924), .B(n31880), .Z(n31883) );
  XNOR U31806 ( .A(p_input[1498]), .B(p_input[2058]), .Z(n31880) );
  XOR U31807 ( .A(p_input[1499]), .B(n16732), .Z(n31924) );
  XOR U31808 ( .A(p_input[1500]), .B(p_input[2060]), .Z(n31884) );
  XOR U31809 ( .A(n31894), .B(n31925), .Z(n31923) );
  IV U31810 ( .A(n31885), .Z(n31925) );
  XOR U31811 ( .A(p_input[1489]), .B(p_input[2049]), .Z(n31885) );
  XNOR U31812 ( .A(n31926), .B(n31901), .Z(n31894) );
  XNOR U31813 ( .A(p_input[1503]), .B(n16735), .Z(n31901) );
  XOR U31814 ( .A(n31891), .B(n31900), .Z(n31926) );
  XOR U31815 ( .A(n31927), .B(n31897), .Z(n31900) );
  XOR U31816 ( .A(p_input[1501]), .B(p_input[2061]), .Z(n31897) );
  XOR U31817 ( .A(p_input[1502]), .B(n16737), .Z(n31927) );
  XOR U31818 ( .A(p_input[1497]), .B(p_input[2057]), .Z(n31891) );
  XOR U31819 ( .A(n31909), .B(n31907), .Z(n31889) );
  XNOR U31820 ( .A(n31928), .B(n31914), .Z(n31907) );
  XOR U31821 ( .A(p_input[1496]), .B(p_input[2056]), .Z(n31914) );
  XOR U31822 ( .A(n31904), .B(n31913), .Z(n31928) );
  XOR U31823 ( .A(n31929), .B(n31910), .Z(n31913) );
  XOR U31824 ( .A(p_input[1494]), .B(p_input[2054]), .Z(n31910) );
  XOR U31825 ( .A(p_input[1495]), .B(n17722), .Z(n31929) );
  XOR U31826 ( .A(p_input[1490]), .B(p_input[2050]), .Z(n31904) );
  XNOR U31827 ( .A(n31919), .B(n31918), .Z(n31909) );
  XOR U31828 ( .A(n31930), .B(n31915), .Z(n31918) );
  XOR U31829 ( .A(p_input[1491]), .B(p_input[2051]), .Z(n31915) );
  XOR U31830 ( .A(p_input[1492]), .B(n17724), .Z(n31930) );
  XOR U31831 ( .A(p_input[1493]), .B(p_input[2053]), .Z(n31919) );
  XNOR U31832 ( .A(n31931), .B(n31932), .Z(n31824) );
  AND U31833 ( .A(n1062), .B(n31933), .Z(n31932) );
  XNOR U31834 ( .A(n31934), .B(n31935), .Z(n1062) );
  AND U31835 ( .A(n31936), .B(n31937), .Z(n31935) );
  XOR U31836 ( .A(n31934), .B(n31834), .Z(n31937) );
  XNOR U31837 ( .A(n31934), .B(n31788), .Z(n31936) );
  XOR U31838 ( .A(n31938), .B(n31939), .Z(n31934) );
  AND U31839 ( .A(n31940), .B(n31941), .Z(n31939) );
  XOR U31840 ( .A(n31938), .B(n31798), .Z(n31940) );
  XOR U31841 ( .A(n31942), .B(n31943), .Z(n31777) );
  AND U31842 ( .A(n1066), .B(n31933), .Z(n31943) );
  XNOR U31843 ( .A(n31931), .B(n31942), .Z(n31933) );
  XNOR U31844 ( .A(n31944), .B(n31945), .Z(n1066) );
  AND U31845 ( .A(n31946), .B(n31947), .Z(n31945) );
  XNOR U31846 ( .A(n31948), .B(n31944), .Z(n31947) );
  IV U31847 ( .A(n31834), .Z(n31948) );
  XNOR U31848 ( .A(n31949), .B(n31950), .Z(n31834) );
  AND U31849 ( .A(n1069), .B(n31951), .Z(n31950) );
  XNOR U31850 ( .A(n31949), .B(n31952), .Z(n31951) );
  XNOR U31851 ( .A(n31788), .B(n31944), .Z(n31946) );
  XOR U31852 ( .A(n31953), .B(n31954), .Z(n31788) );
  AND U31853 ( .A(n1077), .B(n31955), .Z(n31954) );
  XOR U31854 ( .A(n31938), .B(n31956), .Z(n31944) );
  AND U31855 ( .A(n31957), .B(n31941), .Z(n31956) );
  XNOR U31856 ( .A(n31847), .B(n31938), .Z(n31941) );
  XNOR U31857 ( .A(n31958), .B(n31959), .Z(n31847) );
  AND U31858 ( .A(n1069), .B(n31960), .Z(n31959) );
  XOR U31859 ( .A(n31961), .B(n31958), .Z(n31960) );
  XNOR U31860 ( .A(n31962), .B(n31938), .Z(n31957) );
  IV U31861 ( .A(n31798), .Z(n31962) );
  XOR U31862 ( .A(n31963), .B(n31964), .Z(n31798) );
  AND U31863 ( .A(n1077), .B(n31965), .Z(n31964) );
  XOR U31864 ( .A(n31966), .B(n31967), .Z(n31938) );
  AND U31865 ( .A(n31968), .B(n31969), .Z(n31967) );
  XNOR U31866 ( .A(n31872), .B(n31966), .Z(n31969) );
  XNOR U31867 ( .A(n31970), .B(n31971), .Z(n31872) );
  AND U31868 ( .A(n1069), .B(n31972), .Z(n31971) );
  XNOR U31869 ( .A(n31973), .B(n31970), .Z(n31972) );
  XOR U31870 ( .A(n31966), .B(n31809), .Z(n31968) );
  XOR U31871 ( .A(n31974), .B(n31975), .Z(n31809) );
  AND U31872 ( .A(n1077), .B(n31976), .Z(n31975) );
  XOR U31873 ( .A(n31977), .B(n31978), .Z(n31966) );
  AND U31874 ( .A(n31979), .B(n31980), .Z(n31978) );
  XNOR U31875 ( .A(n31977), .B(n31920), .Z(n31980) );
  XNOR U31876 ( .A(n31981), .B(n31982), .Z(n31920) );
  AND U31877 ( .A(n1069), .B(n31983), .Z(n31982) );
  XOR U31878 ( .A(n31984), .B(n31981), .Z(n31983) );
  XNOR U31879 ( .A(n31985), .B(n31977), .Z(n31979) );
  IV U31880 ( .A(n31821), .Z(n31985) );
  XOR U31881 ( .A(n31986), .B(n31987), .Z(n31821) );
  AND U31882 ( .A(n1077), .B(n31988), .Z(n31987) );
  AND U31883 ( .A(n31942), .B(n31931), .Z(n31977) );
  XNOR U31884 ( .A(n31989), .B(n31990), .Z(n31931) );
  AND U31885 ( .A(n1069), .B(n31991), .Z(n31990) );
  XNOR U31886 ( .A(n31992), .B(n31989), .Z(n31991) );
  XNOR U31887 ( .A(n31993), .B(n31994), .Z(n1069) );
  AND U31888 ( .A(n31995), .B(n31996), .Z(n31994) );
  XOR U31889 ( .A(n31952), .B(n31993), .Z(n31996) );
  AND U31890 ( .A(n31997), .B(n31998), .Z(n31952) );
  XOR U31891 ( .A(n31993), .B(n31949), .Z(n31995) );
  XNOR U31892 ( .A(n31999), .B(n32000), .Z(n31949) );
  AND U31893 ( .A(n1073), .B(n31955), .Z(n32000) );
  XOR U31894 ( .A(n31953), .B(n31999), .Z(n31955) );
  XOR U31895 ( .A(n32001), .B(n32002), .Z(n31993) );
  AND U31896 ( .A(n32003), .B(n32004), .Z(n32002) );
  XNOR U31897 ( .A(n32001), .B(n31997), .Z(n32004) );
  IV U31898 ( .A(n31961), .Z(n31997) );
  XOR U31899 ( .A(n32005), .B(n32006), .Z(n31961) );
  XOR U31900 ( .A(n32007), .B(n31998), .Z(n32006) );
  AND U31901 ( .A(n31973), .B(n32008), .Z(n31998) );
  AND U31902 ( .A(n32009), .B(n32010), .Z(n32007) );
  XOR U31903 ( .A(n32011), .B(n32005), .Z(n32009) );
  XNOR U31904 ( .A(n31958), .B(n32001), .Z(n32003) );
  XNOR U31905 ( .A(n32012), .B(n32013), .Z(n31958) );
  AND U31906 ( .A(n1073), .B(n31965), .Z(n32013) );
  XOR U31907 ( .A(n32012), .B(n31963), .Z(n31965) );
  XOR U31908 ( .A(n32014), .B(n32015), .Z(n32001) );
  AND U31909 ( .A(n32016), .B(n32017), .Z(n32015) );
  XNOR U31910 ( .A(n32014), .B(n31973), .Z(n32017) );
  XOR U31911 ( .A(n32018), .B(n32010), .Z(n31973) );
  XNOR U31912 ( .A(n32019), .B(n32005), .Z(n32010) );
  XOR U31913 ( .A(n32020), .B(n32021), .Z(n32005) );
  AND U31914 ( .A(n32022), .B(n32023), .Z(n32021) );
  XOR U31915 ( .A(n32024), .B(n32020), .Z(n32022) );
  XNOR U31916 ( .A(n32025), .B(n32026), .Z(n32019) );
  AND U31917 ( .A(n32027), .B(n32028), .Z(n32026) );
  XOR U31918 ( .A(n32025), .B(n32029), .Z(n32027) );
  XNOR U31919 ( .A(n32011), .B(n32008), .Z(n32018) );
  AND U31920 ( .A(n32030), .B(n32031), .Z(n32008) );
  XOR U31921 ( .A(n32032), .B(n32033), .Z(n32011) );
  AND U31922 ( .A(n32034), .B(n32035), .Z(n32033) );
  XOR U31923 ( .A(n32032), .B(n32036), .Z(n32034) );
  XNOR U31924 ( .A(n31970), .B(n32014), .Z(n32016) );
  XNOR U31925 ( .A(n32037), .B(n32038), .Z(n31970) );
  AND U31926 ( .A(n1073), .B(n31976), .Z(n32038) );
  XOR U31927 ( .A(n32037), .B(n31974), .Z(n31976) );
  XOR U31928 ( .A(n32039), .B(n32040), .Z(n32014) );
  AND U31929 ( .A(n32041), .B(n32042), .Z(n32040) );
  XNOR U31930 ( .A(n32039), .B(n32030), .Z(n32042) );
  IV U31931 ( .A(n31984), .Z(n32030) );
  XNOR U31932 ( .A(n32043), .B(n32023), .Z(n31984) );
  XNOR U31933 ( .A(n32044), .B(n32029), .Z(n32023) );
  XNOR U31934 ( .A(n32045), .B(n32046), .Z(n32029) );
  NOR U31935 ( .A(n32047), .B(n32048), .Z(n32046) );
  XOR U31936 ( .A(n32045), .B(n32049), .Z(n32047) );
  XNOR U31937 ( .A(n32028), .B(n32020), .Z(n32044) );
  XOR U31938 ( .A(n32050), .B(n32051), .Z(n32020) );
  AND U31939 ( .A(n32052), .B(n32053), .Z(n32051) );
  XOR U31940 ( .A(n32050), .B(n32054), .Z(n32052) );
  XNOR U31941 ( .A(n32055), .B(n32025), .Z(n32028) );
  XOR U31942 ( .A(n32056), .B(n32057), .Z(n32025) );
  AND U31943 ( .A(n32058), .B(n32059), .Z(n32057) );
  XNOR U31944 ( .A(n32060), .B(n32061), .Z(n32058) );
  IV U31945 ( .A(n32056), .Z(n32060) );
  XNOR U31946 ( .A(n32062), .B(n32063), .Z(n32055) );
  NOR U31947 ( .A(n32064), .B(n32065), .Z(n32063) );
  XNOR U31948 ( .A(n32062), .B(n32066), .Z(n32064) );
  XNOR U31949 ( .A(n32024), .B(n32031), .Z(n32043) );
  NOR U31950 ( .A(n31992), .B(n32067), .Z(n32031) );
  XOR U31951 ( .A(n32036), .B(n32035), .Z(n32024) );
  XNOR U31952 ( .A(n32068), .B(n32032), .Z(n32035) );
  XOR U31953 ( .A(n32069), .B(n32070), .Z(n32032) );
  AND U31954 ( .A(n32071), .B(n32072), .Z(n32070) );
  XNOR U31955 ( .A(n32073), .B(n32074), .Z(n32071) );
  IV U31956 ( .A(n32069), .Z(n32073) );
  XNOR U31957 ( .A(n32075), .B(n32076), .Z(n32068) );
  NOR U31958 ( .A(n32077), .B(n32078), .Z(n32076) );
  XNOR U31959 ( .A(n32075), .B(n32079), .Z(n32077) );
  XOR U31960 ( .A(n32080), .B(n32081), .Z(n32036) );
  NOR U31961 ( .A(n32082), .B(n32083), .Z(n32081) );
  XNOR U31962 ( .A(n32080), .B(n32084), .Z(n32082) );
  XNOR U31963 ( .A(n31981), .B(n32039), .Z(n32041) );
  XNOR U31964 ( .A(n32085), .B(n32086), .Z(n31981) );
  AND U31965 ( .A(n1073), .B(n31988), .Z(n32086) );
  XOR U31966 ( .A(n32085), .B(n31986), .Z(n31988) );
  AND U31967 ( .A(n31989), .B(n31992), .Z(n32039) );
  XOR U31968 ( .A(n32087), .B(n32067), .Z(n31992) );
  XNOR U31969 ( .A(p_input[1504]), .B(p_input[2048]), .Z(n32067) );
  XNOR U31970 ( .A(n32054), .B(n32053), .Z(n32087) );
  XNOR U31971 ( .A(n32088), .B(n32061), .Z(n32053) );
  XNOR U31972 ( .A(n32049), .B(n32048), .Z(n32061) );
  XNOR U31973 ( .A(n32089), .B(n32045), .Z(n32048) );
  XNOR U31974 ( .A(p_input[1514]), .B(p_input[2058]), .Z(n32045) );
  XOR U31975 ( .A(p_input[1515]), .B(n16732), .Z(n32089) );
  XOR U31976 ( .A(p_input[1516]), .B(p_input[2060]), .Z(n32049) );
  XOR U31977 ( .A(n32059), .B(n32090), .Z(n32088) );
  IV U31978 ( .A(n32050), .Z(n32090) );
  XOR U31979 ( .A(p_input[1505]), .B(p_input[2049]), .Z(n32050) );
  XNOR U31980 ( .A(n32091), .B(n32066), .Z(n32059) );
  XNOR U31981 ( .A(p_input[1519]), .B(n16735), .Z(n32066) );
  XOR U31982 ( .A(n32056), .B(n32065), .Z(n32091) );
  XOR U31983 ( .A(n32092), .B(n32062), .Z(n32065) );
  XOR U31984 ( .A(p_input[1517]), .B(p_input[2061]), .Z(n32062) );
  XOR U31985 ( .A(p_input[1518]), .B(n16737), .Z(n32092) );
  XOR U31986 ( .A(p_input[1513]), .B(p_input[2057]), .Z(n32056) );
  XOR U31987 ( .A(n32074), .B(n32072), .Z(n32054) );
  XNOR U31988 ( .A(n32093), .B(n32079), .Z(n32072) );
  XOR U31989 ( .A(p_input[1512]), .B(p_input[2056]), .Z(n32079) );
  XOR U31990 ( .A(n32069), .B(n32078), .Z(n32093) );
  XOR U31991 ( .A(n32094), .B(n32075), .Z(n32078) );
  XOR U31992 ( .A(p_input[1510]), .B(p_input[2054]), .Z(n32075) );
  XOR U31993 ( .A(p_input[1511]), .B(n17722), .Z(n32094) );
  XOR U31994 ( .A(p_input[1506]), .B(p_input[2050]), .Z(n32069) );
  XNOR U31995 ( .A(n32084), .B(n32083), .Z(n32074) );
  XOR U31996 ( .A(n32095), .B(n32080), .Z(n32083) );
  XOR U31997 ( .A(p_input[1507]), .B(p_input[2051]), .Z(n32080) );
  XOR U31998 ( .A(p_input[1508]), .B(n17724), .Z(n32095) );
  XOR U31999 ( .A(p_input[1509]), .B(p_input[2053]), .Z(n32084) );
  XNOR U32000 ( .A(n32096), .B(n32097), .Z(n31989) );
  AND U32001 ( .A(n1073), .B(n32098), .Z(n32097) );
  XNOR U32002 ( .A(n32099), .B(n32100), .Z(n1073) );
  AND U32003 ( .A(n32101), .B(n32102), .Z(n32100) );
  XOR U32004 ( .A(n32099), .B(n31999), .Z(n32102) );
  XNOR U32005 ( .A(n32099), .B(n31953), .Z(n32101) );
  XOR U32006 ( .A(n32103), .B(n32104), .Z(n32099) );
  AND U32007 ( .A(n32105), .B(n32106), .Z(n32104) );
  XOR U32008 ( .A(n32103), .B(n31963), .Z(n32105) );
  XOR U32009 ( .A(n32107), .B(n32108), .Z(n31942) );
  AND U32010 ( .A(n1077), .B(n32098), .Z(n32108) );
  XNOR U32011 ( .A(n32096), .B(n32107), .Z(n32098) );
  XNOR U32012 ( .A(n32109), .B(n32110), .Z(n1077) );
  AND U32013 ( .A(n32111), .B(n32112), .Z(n32110) );
  XNOR U32014 ( .A(n32113), .B(n32109), .Z(n32112) );
  IV U32015 ( .A(n31999), .Z(n32113) );
  XNOR U32016 ( .A(n32114), .B(n32115), .Z(n31999) );
  AND U32017 ( .A(n1080), .B(n32116), .Z(n32115) );
  XNOR U32018 ( .A(n32114), .B(n32117), .Z(n32116) );
  XNOR U32019 ( .A(n31953), .B(n32109), .Z(n32111) );
  XOR U32020 ( .A(n32118), .B(n32119), .Z(n31953) );
  AND U32021 ( .A(n1088), .B(n32120), .Z(n32119) );
  XOR U32022 ( .A(n32103), .B(n32121), .Z(n32109) );
  AND U32023 ( .A(n32122), .B(n32106), .Z(n32121) );
  XNOR U32024 ( .A(n32012), .B(n32103), .Z(n32106) );
  XNOR U32025 ( .A(n32123), .B(n32124), .Z(n32012) );
  AND U32026 ( .A(n1080), .B(n32125), .Z(n32124) );
  XOR U32027 ( .A(n32126), .B(n32123), .Z(n32125) );
  XNOR U32028 ( .A(n32127), .B(n32103), .Z(n32122) );
  IV U32029 ( .A(n31963), .Z(n32127) );
  XOR U32030 ( .A(n32128), .B(n32129), .Z(n31963) );
  AND U32031 ( .A(n1088), .B(n32130), .Z(n32129) );
  XOR U32032 ( .A(n32131), .B(n32132), .Z(n32103) );
  AND U32033 ( .A(n32133), .B(n32134), .Z(n32132) );
  XNOR U32034 ( .A(n32037), .B(n32131), .Z(n32134) );
  XNOR U32035 ( .A(n32135), .B(n32136), .Z(n32037) );
  AND U32036 ( .A(n1080), .B(n32137), .Z(n32136) );
  XNOR U32037 ( .A(n32138), .B(n32135), .Z(n32137) );
  XOR U32038 ( .A(n32131), .B(n31974), .Z(n32133) );
  XOR U32039 ( .A(n32139), .B(n32140), .Z(n31974) );
  AND U32040 ( .A(n1088), .B(n32141), .Z(n32140) );
  XOR U32041 ( .A(n32142), .B(n32143), .Z(n32131) );
  AND U32042 ( .A(n32144), .B(n32145), .Z(n32143) );
  XNOR U32043 ( .A(n32142), .B(n32085), .Z(n32145) );
  XNOR U32044 ( .A(n32146), .B(n32147), .Z(n32085) );
  AND U32045 ( .A(n1080), .B(n32148), .Z(n32147) );
  XOR U32046 ( .A(n32149), .B(n32146), .Z(n32148) );
  XNOR U32047 ( .A(n32150), .B(n32142), .Z(n32144) );
  IV U32048 ( .A(n31986), .Z(n32150) );
  XOR U32049 ( .A(n32151), .B(n32152), .Z(n31986) );
  AND U32050 ( .A(n1088), .B(n32153), .Z(n32152) );
  AND U32051 ( .A(n32107), .B(n32096), .Z(n32142) );
  XNOR U32052 ( .A(n32154), .B(n32155), .Z(n32096) );
  AND U32053 ( .A(n1080), .B(n32156), .Z(n32155) );
  XNOR U32054 ( .A(n32157), .B(n32154), .Z(n32156) );
  XNOR U32055 ( .A(n32158), .B(n32159), .Z(n1080) );
  AND U32056 ( .A(n32160), .B(n32161), .Z(n32159) );
  XOR U32057 ( .A(n32117), .B(n32158), .Z(n32161) );
  AND U32058 ( .A(n32162), .B(n32163), .Z(n32117) );
  XOR U32059 ( .A(n32158), .B(n32114), .Z(n32160) );
  XNOR U32060 ( .A(n32164), .B(n32165), .Z(n32114) );
  AND U32061 ( .A(n1084), .B(n32120), .Z(n32165) );
  XOR U32062 ( .A(n32118), .B(n32164), .Z(n32120) );
  XOR U32063 ( .A(n32166), .B(n32167), .Z(n32158) );
  AND U32064 ( .A(n32168), .B(n32169), .Z(n32167) );
  XNOR U32065 ( .A(n32166), .B(n32162), .Z(n32169) );
  IV U32066 ( .A(n32126), .Z(n32162) );
  XOR U32067 ( .A(n32170), .B(n32171), .Z(n32126) );
  XOR U32068 ( .A(n32172), .B(n32163), .Z(n32171) );
  AND U32069 ( .A(n32138), .B(n32173), .Z(n32163) );
  AND U32070 ( .A(n32174), .B(n32175), .Z(n32172) );
  XOR U32071 ( .A(n32176), .B(n32170), .Z(n32174) );
  XNOR U32072 ( .A(n32123), .B(n32166), .Z(n32168) );
  XNOR U32073 ( .A(n32177), .B(n32178), .Z(n32123) );
  AND U32074 ( .A(n1084), .B(n32130), .Z(n32178) );
  XOR U32075 ( .A(n32177), .B(n32128), .Z(n32130) );
  XOR U32076 ( .A(n32179), .B(n32180), .Z(n32166) );
  AND U32077 ( .A(n32181), .B(n32182), .Z(n32180) );
  XNOR U32078 ( .A(n32179), .B(n32138), .Z(n32182) );
  XOR U32079 ( .A(n32183), .B(n32175), .Z(n32138) );
  XNOR U32080 ( .A(n32184), .B(n32170), .Z(n32175) );
  XOR U32081 ( .A(n32185), .B(n32186), .Z(n32170) );
  AND U32082 ( .A(n32187), .B(n32188), .Z(n32186) );
  XOR U32083 ( .A(n32189), .B(n32185), .Z(n32187) );
  XNOR U32084 ( .A(n32190), .B(n32191), .Z(n32184) );
  AND U32085 ( .A(n32192), .B(n32193), .Z(n32191) );
  XOR U32086 ( .A(n32190), .B(n32194), .Z(n32192) );
  XNOR U32087 ( .A(n32176), .B(n32173), .Z(n32183) );
  AND U32088 ( .A(n32195), .B(n32196), .Z(n32173) );
  XOR U32089 ( .A(n32197), .B(n32198), .Z(n32176) );
  AND U32090 ( .A(n32199), .B(n32200), .Z(n32198) );
  XOR U32091 ( .A(n32197), .B(n32201), .Z(n32199) );
  XNOR U32092 ( .A(n32135), .B(n32179), .Z(n32181) );
  XNOR U32093 ( .A(n32202), .B(n32203), .Z(n32135) );
  AND U32094 ( .A(n1084), .B(n32141), .Z(n32203) );
  XOR U32095 ( .A(n32202), .B(n32139), .Z(n32141) );
  XOR U32096 ( .A(n32204), .B(n32205), .Z(n32179) );
  AND U32097 ( .A(n32206), .B(n32207), .Z(n32205) );
  XNOR U32098 ( .A(n32204), .B(n32195), .Z(n32207) );
  IV U32099 ( .A(n32149), .Z(n32195) );
  XNOR U32100 ( .A(n32208), .B(n32188), .Z(n32149) );
  XNOR U32101 ( .A(n32209), .B(n32194), .Z(n32188) );
  XNOR U32102 ( .A(n32210), .B(n32211), .Z(n32194) );
  NOR U32103 ( .A(n32212), .B(n32213), .Z(n32211) );
  XOR U32104 ( .A(n32210), .B(n32214), .Z(n32212) );
  XNOR U32105 ( .A(n32193), .B(n32185), .Z(n32209) );
  XOR U32106 ( .A(n32215), .B(n32216), .Z(n32185) );
  AND U32107 ( .A(n32217), .B(n32218), .Z(n32216) );
  XOR U32108 ( .A(n32215), .B(n32219), .Z(n32217) );
  XNOR U32109 ( .A(n32220), .B(n32190), .Z(n32193) );
  XOR U32110 ( .A(n32221), .B(n32222), .Z(n32190) );
  AND U32111 ( .A(n32223), .B(n32224), .Z(n32222) );
  XNOR U32112 ( .A(n32225), .B(n32226), .Z(n32223) );
  IV U32113 ( .A(n32221), .Z(n32225) );
  XNOR U32114 ( .A(n32227), .B(n32228), .Z(n32220) );
  NOR U32115 ( .A(n32229), .B(n32230), .Z(n32228) );
  XNOR U32116 ( .A(n32227), .B(n32231), .Z(n32229) );
  XNOR U32117 ( .A(n32189), .B(n32196), .Z(n32208) );
  NOR U32118 ( .A(n32157), .B(n32232), .Z(n32196) );
  XOR U32119 ( .A(n32201), .B(n32200), .Z(n32189) );
  XNOR U32120 ( .A(n32233), .B(n32197), .Z(n32200) );
  XOR U32121 ( .A(n32234), .B(n32235), .Z(n32197) );
  AND U32122 ( .A(n32236), .B(n32237), .Z(n32235) );
  XNOR U32123 ( .A(n32238), .B(n32239), .Z(n32236) );
  IV U32124 ( .A(n32234), .Z(n32238) );
  XNOR U32125 ( .A(n32240), .B(n32241), .Z(n32233) );
  NOR U32126 ( .A(n32242), .B(n32243), .Z(n32241) );
  XNOR U32127 ( .A(n32240), .B(n32244), .Z(n32242) );
  XOR U32128 ( .A(n32245), .B(n32246), .Z(n32201) );
  NOR U32129 ( .A(n32247), .B(n32248), .Z(n32246) );
  XNOR U32130 ( .A(n32245), .B(n32249), .Z(n32247) );
  XNOR U32131 ( .A(n32146), .B(n32204), .Z(n32206) );
  XNOR U32132 ( .A(n32250), .B(n32251), .Z(n32146) );
  AND U32133 ( .A(n1084), .B(n32153), .Z(n32251) );
  XOR U32134 ( .A(n32250), .B(n32151), .Z(n32153) );
  AND U32135 ( .A(n32154), .B(n32157), .Z(n32204) );
  XOR U32136 ( .A(n32252), .B(n32232), .Z(n32157) );
  XNOR U32137 ( .A(p_input[1520]), .B(p_input[2048]), .Z(n32232) );
  XNOR U32138 ( .A(n32219), .B(n32218), .Z(n32252) );
  XNOR U32139 ( .A(n32253), .B(n32226), .Z(n32218) );
  XNOR U32140 ( .A(n32214), .B(n32213), .Z(n32226) );
  XNOR U32141 ( .A(n32254), .B(n32210), .Z(n32213) );
  XNOR U32142 ( .A(p_input[1530]), .B(p_input[2058]), .Z(n32210) );
  XOR U32143 ( .A(p_input[1531]), .B(n16732), .Z(n32254) );
  XOR U32144 ( .A(p_input[1532]), .B(p_input[2060]), .Z(n32214) );
  XOR U32145 ( .A(n32224), .B(n32255), .Z(n32253) );
  IV U32146 ( .A(n32215), .Z(n32255) );
  XOR U32147 ( .A(p_input[1521]), .B(p_input[2049]), .Z(n32215) );
  XNOR U32148 ( .A(n32256), .B(n32231), .Z(n32224) );
  XNOR U32149 ( .A(p_input[1535]), .B(n16735), .Z(n32231) );
  XOR U32150 ( .A(n32221), .B(n32230), .Z(n32256) );
  XOR U32151 ( .A(n32257), .B(n32227), .Z(n32230) );
  XOR U32152 ( .A(p_input[1533]), .B(p_input[2061]), .Z(n32227) );
  XOR U32153 ( .A(p_input[1534]), .B(n16737), .Z(n32257) );
  XOR U32154 ( .A(p_input[1529]), .B(p_input[2057]), .Z(n32221) );
  XOR U32155 ( .A(n32239), .B(n32237), .Z(n32219) );
  XNOR U32156 ( .A(n32258), .B(n32244), .Z(n32237) );
  XOR U32157 ( .A(p_input[1528]), .B(p_input[2056]), .Z(n32244) );
  XOR U32158 ( .A(n32234), .B(n32243), .Z(n32258) );
  XOR U32159 ( .A(n32259), .B(n32240), .Z(n32243) );
  XOR U32160 ( .A(p_input[1526]), .B(p_input[2054]), .Z(n32240) );
  XOR U32161 ( .A(p_input[1527]), .B(n17722), .Z(n32259) );
  XOR U32162 ( .A(p_input[1522]), .B(p_input[2050]), .Z(n32234) );
  XNOR U32163 ( .A(n32249), .B(n32248), .Z(n32239) );
  XOR U32164 ( .A(n32260), .B(n32245), .Z(n32248) );
  XOR U32165 ( .A(p_input[1523]), .B(p_input[2051]), .Z(n32245) );
  XOR U32166 ( .A(p_input[1524]), .B(n17724), .Z(n32260) );
  XOR U32167 ( .A(p_input[1525]), .B(p_input[2053]), .Z(n32249) );
  XNOR U32168 ( .A(n32261), .B(n32262), .Z(n32154) );
  AND U32169 ( .A(n1084), .B(n32263), .Z(n32262) );
  XNOR U32170 ( .A(n32264), .B(n32265), .Z(n1084) );
  AND U32171 ( .A(n32266), .B(n32267), .Z(n32265) );
  XOR U32172 ( .A(n32264), .B(n32164), .Z(n32267) );
  XNOR U32173 ( .A(n32264), .B(n32118), .Z(n32266) );
  XOR U32174 ( .A(n32268), .B(n32269), .Z(n32264) );
  AND U32175 ( .A(n32270), .B(n32271), .Z(n32269) );
  XOR U32176 ( .A(n32268), .B(n32128), .Z(n32270) );
  XOR U32177 ( .A(n32272), .B(n32273), .Z(n32107) );
  AND U32178 ( .A(n1088), .B(n32263), .Z(n32273) );
  XNOR U32179 ( .A(n32261), .B(n32272), .Z(n32263) );
  XNOR U32180 ( .A(n32274), .B(n32275), .Z(n1088) );
  AND U32181 ( .A(n32276), .B(n32277), .Z(n32275) );
  XNOR U32182 ( .A(n32278), .B(n32274), .Z(n32277) );
  IV U32183 ( .A(n32164), .Z(n32278) );
  XNOR U32184 ( .A(n32279), .B(n32280), .Z(n32164) );
  AND U32185 ( .A(n1091), .B(n32281), .Z(n32280) );
  XNOR U32186 ( .A(n32279), .B(n32282), .Z(n32281) );
  XNOR U32187 ( .A(n32118), .B(n32274), .Z(n32276) );
  XOR U32188 ( .A(n32283), .B(n32284), .Z(n32118) );
  AND U32189 ( .A(n1099), .B(n32285), .Z(n32284) );
  XOR U32190 ( .A(n32268), .B(n32286), .Z(n32274) );
  AND U32191 ( .A(n32287), .B(n32271), .Z(n32286) );
  XNOR U32192 ( .A(n32177), .B(n32268), .Z(n32271) );
  XNOR U32193 ( .A(n32288), .B(n32289), .Z(n32177) );
  AND U32194 ( .A(n1091), .B(n32290), .Z(n32289) );
  XOR U32195 ( .A(n32291), .B(n32288), .Z(n32290) );
  XNOR U32196 ( .A(n32292), .B(n32268), .Z(n32287) );
  IV U32197 ( .A(n32128), .Z(n32292) );
  XOR U32198 ( .A(n32293), .B(n32294), .Z(n32128) );
  AND U32199 ( .A(n1099), .B(n32295), .Z(n32294) );
  XOR U32200 ( .A(n32296), .B(n32297), .Z(n32268) );
  AND U32201 ( .A(n32298), .B(n32299), .Z(n32297) );
  XNOR U32202 ( .A(n32202), .B(n32296), .Z(n32299) );
  XNOR U32203 ( .A(n32300), .B(n32301), .Z(n32202) );
  AND U32204 ( .A(n1091), .B(n32302), .Z(n32301) );
  XNOR U32205 ( .A(n32303), .B(n32300), .Z(n32302) );
  XOR U32206 ( .A(n32296), .B(n32139), .Z(n32298) );
  XOR U32207 ( .A(n32304), .B(n32305), .Z(n32139) );
  AND U32208 ( .A(n1099), .B(n32306), .Z(n32305) );
  XOR U32209 ( .A(n32307), .B(n32308), .Z(n32296) );
  AND U32210 ( .A(n32309), .B(n32310), .Z(n32308) );
  XNOR U32211 ( .A(n32307), .B(n32250), .Z(n32310) );
  XNOR U32212 ( .A(n32311), .B(n32312), .Z(n32250) );
  AND U32213 ( .A(n1091), .B(n32313), .Z(n32312) );
  XOR U32214 ( .A(n32314), .B(n32311), .Z(n32313) );
  XNOR U32215 ( .A(n32315), .B(n32307), .Z(n32309) );
  IV U32216 ( .A(n32151), .Z(n32315) );
  XOR U32217 ( .A(n32316), .B(n32317), .Z(n32151) );
  AND U32218 ( .A(n1099), .B(n32318), .Z(n32317) );
  AND U32219 ( .A(n32272), .B(n32261), .Z(n32307) );
  XNOR U32220 ( .A(n32319), .B(n32320), .Z(n32261) );
  AND U32221 ( .A(n1091), .B(n32321), .Z(n32320) );
  XNOR U32222 ( .A(n32322), .B(n32319), .Z(n32321) );
  XNOR U32223 ( .A(n32323), .B(n32324), .Z(n1091) );
  AND U32224 ( .A(n32325), .B(n32326), .Z(n32324) );
  XOR U32225 ( .A(n32282), .B(n32323), .Z(n32326) );
  AND U32226 ( .A(n32327), .B(n32328), .Z(n32282) );
  XOR U32227 ( .A(n32323), .B(n32279), .Z(n32325) );
  XNOR U32228 ( .A(n32329), .B(n32330), .Z(n32279) );
  AND U32229 ( .A(n1095), .B(n32285), .Z(n32330) );
  XOR U32230 ( .A(n32283), .B(n32329), .Z(n32285) );
  XOR U32231 ( .A(n32331), .B(n32332), .Z(n32323) );
  AND U32232 ( .A(n32333), .B(n32334), .Z(n32332) );
  XNOR U32233 ( .A(n32331), .B(n32327), .Z(n32334) );
  IV U32234 ( .A(n32291), .Z(n32327) );
  XOR U32235 ( .A(n32335), .B(n32336), .Z(n32291) );
  XOR U32236 ( .A(n32337), .B(n32328), .Z(n32336) );
  AND U32237 ( .A(n32303), .B(n32338), .Z(n32328) );
  AND U32238 ( .A(n32339), .B(n32340), .Z(n32337) );
  XOR U32239 ( .A(n32341), .B(n32335), .Z(n32339) );
  XNOR U32240 ( .A(n32288), .B(n32331), .Z(n32333) );
  XNOR U32241 ( .A(n32342), .B(n32343), .Z(n32288) );
  AND U32242 ( .A(n1095), .B(n32295), .Z(n32343) );
  XOR U32243 ( .A(n32342), .B(n32293), .Z(n32295) );
  XOR U32244 ( .A(n32344), .B(n32345), .Z(n32331) );
  AND U32245 ( .A(n32346), .B(n32347), .Z(n32345) );
  XNOR U32246 ( .A(n32344), .B(n32303), .Z(n32347) );
  XOR U32247 ( .A(n32348), .B(n32340), .Z(n32303) );
  XNOR U32248 ( .A(n32349), .B(n32335), .Z(n32340) );
  XOR U32249 ( .A(n32350), .B(n32351), .Z(n32335) );
  AND U32250 ( .A(n32352), .B(n32353), .Z(n32351) );
  XOR U32251 ( .A(n32354), .B(n32350), .Z(n32352) );
  XNOR U32252 ( .A(n32355), .B(n32356), .Z(n32349) );
  AND U32253 ( .A(n32357), .B(n32358), .Z(n32356) );
  XOR U32254 ( .A(n32355), .B(n32359), .Z(n32357) );
  XNOR U32255 ( .A(n32341), .B(n32338), .Z(n32348) );
  AND U32256 ( .A(n32360), .B(n32361), .Z(n32338) );
  XOR U32257 ( .A(n32362), .B(n32363), .Z(n32341) );
  AND U32258 ( .A(n32364), .B(n32365), .Z(n32363) );
  XOR U32259 ( .A(n32362), .B(n32366), .Z(n32364) );
  XNOR U32260 ( .A(n32300), .B(n32344), .Z(n32346) );
  XNOR U32261 ( .A(n32367), .B(n32368), .Z(n32300) );
  AND U32262 ( .A(n1095), .B(n32306), .Z(n32368) );
  XOR U32263 ( .A(n32367), .B(n32304), .Z(n32306) );
  XOR U32264 ( .A(n32369), .B(n32370), .Z(n32344) );
  AND U32265 ( .A(n32371), .B(n32372), .Z(n32370) );
  XNOR U32266 ( .A(n32369), .B(n32360), .Z(n32372) );
  IV U32267 ( .A(n32314), .Z(n32360) );
  XNOR U32268 ( .A(n32373), .B(n32353), .Z(n32314) );
  XNOR U32269 ( .A(n32374), .B(n32359), .Z(n32353) );
  XNOR U32270 ( .A(n32375), .B(n32376), .Z(n32359) );
  NOR U32271 ( .A(n32377), .B(n32378), .Z(n32376) );
  XOR U32272 ( .A(n32375), .B(n32379), .Z(n32377) );
  XNOR U32273 ( .A(n32358), .B(n32350), .Z(n32374) );
  XOR U32274 ( .A(n32380), .B(n32381), .Z(n32350) );
  AND U32275 ( .A(n32382), .B(n32383), .Z(n32381) );
  XOR U32276 ( .A(n32380), .B(n32384), .Z(n32382) );
  XNOR U32277 ( .A(n32385), .B(n32355), .Z(n32358) );
  XOR U32278 ( .A(n32386), .B(n32387), .Z(n32355) );
  AND U32279 ( .A(n32388), .B(n32389), .Z(n32387) );
  XNOR U32280 ( .A(n32390), .B(n32391), .Z(n32388) );
  IV U32281 ( .A(n32386), .Z(n32390) );
  XNOR U32282 ( .A(n32392), .B(n32393), .Z(n32385) );
  NOR U32283 ( .A(n32394), .B(n32395), .Z(n32393) );
  XNOR U32284 ( .A(n32392), .B(n32396), .Z(n32394) );
  XNOR U32285 ( .A(n32354), .B(n32361), .Z(n32373) );
  NOR U32286 ( .A(n32322), .B(n32397), .Z(n32361) );
  XOR U32287 ( .A(n32366), .B(n32365), .Z(n32354) );
  XNOR U32288 ( .A(n32398), .B(n32362), .Z(n32365) );
  XOR U32289 ( .A(n32399), .B(n32400), .Z(n32362) );
  AND U32290 ( .A(n32401), .B(n32402), .Z(n32400) );
  XNOR U32291 ( .A(n32403), .B(n32404), .Z(n32401) );
  IV U32292 ( .A(n32399), .Z(n32403) );
  XNOR U32293 ( .A(n32405), .B(n32406), .Z(n32398) );
  NOR U32294 ( .A(n32407), .B(n32408), .Z(n32406) );
  XNOR U32295 ( .A(n32405), .B(n32409), .Z(n32407) );
  XOR U32296 ( .A(n32410), .B(n32411), .Z(n32366) );
  NOR U32297 ( .A(n32412), .B(n32413), .Z(n32411) );
  XNOR U32298 ( .A(n32410), .B(n32414), .Z(n32412) );
  XNOR U32299 ( .A(n32311), .B(n32369), .Z(n32371) );
  XNOR U32300 ( .A(n32415), .B(n32416), .Z(n32311) );
  AND U32301 ( .A(n1095), .B(n32318), .Z(n32416) );
  XOR U32302 ( .A(n32415), .B(n32316), .Z(n32318) );
  AND U32303 ( .A(n32319), .B(n32322), .Z(n32369) );
  XOR U32304 ( .A(n32417), .B(n32397), .Z(n32322) );
  XNOR U32305 ( .A(p_input[1536]), .B(p_input[2048]), .Z(n32397) );
  XNOR U32306 ( .A(n32384), .B(n32383), .Z(n32417) );
  XNOR U32307 ( .A(n32418), .B(n32391), .Z(n32383) );
  XNOR U32308 ( .A(n32379), .B(n32378), .Z(n32391) );
  XNOR U32309 ( .A(n32419), .B(n32375), .Z(n32378) );
  XNOR U32310 ( .A(p_input[1546]), .B(p_input[2058]), .Z(n32375) );
  XOR U32311 ( .A(p_input[1547]), .B(n16732), .Z(n32419) );
  XOR U32312 ( .A(p_input[1548]), .B(p_input[2060]), .Z(n32379) );
  XOR U32313 ( .A(n32389), .B(n32420), .Z(n32418) );
  IV U32314 ( .A(n32380), .Z(n32420) );
  XOR U32315 ( .A(p_input[1537]), .B(p_input[2049]), .Z(n32380) );
  XNOR U32316 ( .A(n32421), .B(n32396), .Z(n32389) );
  XNOR U32317 ( .A(p_input[1551]), .B(n16735), .Z(n32396) );
  XOR U32318 ( .A(n32386), .B(n32395), .Z(n32421) );
  XOR U32319 ( .A(n32422), .B(n32392), .Z(n32395) );
  XOR U32320 ( .A(p_input[1549]), .B(p_input[2061]), .Z(n32392) );
  XOR U32321 ( .A(p_input[1550]), .B(n16737), .Z(n32422) );
  XOR U32322 ( .A(p_input[1545]), .B(p_input[2057]), .Z(n32386) );
  XOR U32323 ( .A(n32404), .B(n32402), .Z(n32384) );
  XNOR U32324 ( .A(n32423), .B(n32409), .Z(n32402) );
  XOR U32325 ( .A(p_input[1544]), .B(p_input[2056]), .Z(n32409) );
  XOR U32326 ( .A(n32399), .B(n32408), .Z(n32423) );
  XOR U32327 ( .A(n32424), .B(n32405), .Z(n32408) );
  XOR U32328 ( .A(p_input[1542]), .B(p_input[2054]), .Z(n32405) );
  XOR U32329 ( .A(p_input[1543]), .B(n17722), .Z(n32424) );
  XOR U32330 ( .A(p_input[1538]), .B(p_input[2050]), .Z(n32399) );
  XNOR U32331 ( .A(n32414), .B(n32413), .Z(n32404) );
  XOR U32332 ( .A(n32425), .B(n32410), .Z(n32413) );
  XOR U32333 ( .A(p_input[1539]), .B(p_input[2051]), .Z(n32410) );
  XOR U32334 ( .A(p_input[1540]), .B(n17724), .Z(n32425) );
  XOR U32335 ( .A(p_input[1541]), .B(p_input[2053]), .Z(n32414) );
  XNOR U32336 ( .A(n32426), .B(n32427), .Z(n32319) );
  AND U32337 ( .A(n1095), .B(n32428), .Z(n32427) );
  XNOR U32338 ( .A(n32429), .B(n32430), .Z(n1095) );
  AND U32339 ( .A(n32431), .B(n32432), .Z(n32430) );
  XOR U32340 ( .A(n32429), .B(n32329), .Z(n32432) );
  XNOR U32341 ( .A(n32429), .B(n32283), .Z(n32431) );
  XOR U32342 ( .A(n32433), .B(n32434), .Z(n32429) );
  AND U32343 ( .A(n32435), .B(n32436), .Z(n32434) );
  XOR U32344 ( .A(n32433), .B(n32293), .Z(n32435) );
  XOR U32345 ( .A(n32437), .B(n32438), .Z(n32272) );
  AND U32346 ( .A(n1099), .B(n32428), .Z(n32438) );
  XNOR U32347 ( .A(n32426), .B(n32437), .Z(n32428) );
  XNOR U32348 ( .A(n32439), .B(n32440), .Z(n1099) );
  AND U32349 ( .A(n32441), .B(n32442), .Z(n32440) );
  XNOR U32350 ( .A(n32443), .B(n32439), .Z(n32442) );
  IV U32351 ( .A(n32329), .Z(n32443) );
  XNOR U32352 ( .A(n32444), .B(n32445), .Z(n32329) );
  AND U32353 ( .A(n1102), .B(n32446), .Z(n32445) );
  XNOR U32354 ( .A(n32444), .B(n32447), .Z(n32446) );
  XNOR U32355 ( .A(n32283), .B(n32439), .Z(n32441) );
  XOR U32356 ( .A(n32448), .B(n32449), .Z(n32283) );
  AND U32357 ( .A(n1110), .B(n32450), .Z(n32449) );
  XOR U32358 ( .A(n32433), .B(n32451), .Z(n32439) );
  AND U32359 ( .A(n32452), .B(n32436), .Z(n32451) );
  XNOR U32360 ( .A(n32342), .B(n32433), .Z(n32436) );
  XNOR U32361 ( .A(n32453), .B(n32454), .Z(n32342) );
  AND U32362 ( .A(n1102), .B(n32455), .Z(n32454) );
  XOR U32363 ( .A(n32456), .B(n32453), .Z(n32455) );
  XNOR U32364 ( .A(n32457), .B(n32433), .Z(n32452) );
  IV U32365 ( .A(n32293), .Z(n32457) );
  XOR U32366 ( .A(n32458), .B(n32459), .Z(n32293) );
  AND U32367 ( .A(n1110), .B(n32460), .Z(n32459) );
  XOR U32368 ( .A(n32461), .B(n32462), .Z(n32433) );
  AND U32369 ( .A(n32463), .B(n32464), .Z(n32462) );
  XNOR U32370 ( .A(n32367), .B(n32461), .Z(n32464) );
  XNOR U32371 ( .A(n32465), .B(n32466), .Z(n32367) );
  AND U32372 ( .A(n1102), .B(n32467), .Z(n32466) );
  XNOR U32373 ( .A(n32468), .B(n32465), .Z(n32467) );
  XOR U32374 ( .A(n32461), .B(n32304), .Z(n32463) );
  XOR U32375 ( .A(n32469), .B(n32470), .Z(n32304) );
  AND U32376 ( .A(n1110), .B(n32471), .Z(n32470) );
  XOR U32377 ( .A(n32472), .B(n32473), .Z(n32461) );
  AND U32378 ( .A(n32474), .B(n32475), .Z(n32473) );
  XNOR U32379 ( .A(n32472), .B(n32415), .Z(n32475) );
  XNOR U32380 ( .A(n32476), .B(n32477), .Z(n32415) );
  AND U32381 ( .A(n1102), .B(n32478), .Z(n32477) );
  XOR U32382 ( .A(n32479), .B(n32476), .Z(n32478) );
  XNOR U32383 ( .A(n32480), .B(n32472), .Z(n32474) );
  IV U32384 ( .A(n32316), .Z(n32480) );
  XOR U32385 ( .A(n32481), .B(n32482), .Z(n32316) );
  AND U32386 ( .A(n1110), .B(n32483), .Z(n32482) );
  AND U32387 ( .A(n32437), .B(n32426), .Z(n32472) );
  XNOR U32388 ( .A(n32484), .B(n32485), .Z(n32426) );
  AND U32389 ( .A(n1102), .B(n32486), .Z(n32485) );
  XNOR U32390 ( .A(n32487), .B(n32484), .Z(n32486) );
  XNOR U32391 ( .A(n32488), .B(n32489), .Z(n1102) );
  AND U32392 ( .A(n32490), .B(n32491), .Z(n32489) );
  XOR U32393 ( .A(n32447), .B(n32488), .Z(n32491) );
  AND U32394 ( .A(n32492), .B(n32493), .Z(n32447) );
  XOR U32395 ( .A(n32488), .B(n32444), .Z(n32490) );
  XNOR U32396 ( .A(n32494), .B(n32495), .Z(n32444) );
  AND U32397 ( .A(n1106), .B(n32450), .Z(n32495) );
  XOR U32398 ( .A(n32448), .B(n32494), .Z(n32450) );
  XOR U32399 ( .A(n32496), .B(n32497), .Z(n32488) );
  AND U32400 ( .A(n32498), .B(n32499), .Z(n32497) );
  XNOR U32401 ( .A(n32496), .B(n32492), .Z(n32499) );
  IV U32402 ( .A(n32456), .Z(n32492) );
  XOR U32403 ( .A(n32500), .B(n32501), .Z(n32456) );
  XOR U32404 ( .A(n32502), .B(n32493), .Z(n32501) );
  AND U32405 ( .A(n32468), .B(n32503), .Z(n32493) );
  AND U32406 ( .A(n32504), .B(n32505), .Z(n32502) );
  XOR U32407 ( .A(n32506), .B(n32500), .Z(n32504) );
  XNOR U32408 ( .A(n32453), .B(n32496), .Z(n32498) );
  XNOR U32409 ( .A(n32507), .B(n32508), .Z(n32453) );
  AND U32410 ( .A(n1106), .B(n32460), .Z(n32508) );
  XOR U32411 ( .A(n32507), .B(n32458), .Z(n32460) );
  XOR U32412 ( .A(n32509), .B(n32510), .Z(n32496) );
  AND U32413 ( .A(n32511), .B(n32512), .Z(n32510) );
  XNOR U32414 ( .A(n32509), .B(n32468), .Z(n32512) );
  XOR U32415 ( .A(n32513), .B(n32505), .Z(n32468) );
  XNOR U32416 ( .A(n32514), .B(n32500), .Z(n32505) );
  XOR U32417 ( .A(n32515), .B(n32516), .Z(n32500) );
  AND U32418 ( .A(n32517), .B(n32518), .Z(n32516) );
  XOR U32419 ( .A(n32519), .B(n32515), .Z(n32517) );
  XNOR U32420 ( .A(n32520), .B(n32521), .Z(n32514) );
  AND U32421 ( .A(n32522), .B(n32523), .Z(n32521) );
  XOR U32422 ( .A(n32520), .B(n32524), .Z(n32522) );
  XNOR U32423 ( .A(n32506), .B(n32503), .Z(n32513) );
  AND U32424 ( .A(n32525), .B(n32526), .Z(n32503) );
  XOR U32425 ( .A(n32527), .B(n32528), .Z(n32506) );
  AND U32426 ( .A(n32529), .B(n32530), .Z(n32528) );
  XOR U32427 ( .A(n32527), .B(n32531), .Z(n32529) );
  XNOR U32428 ( .A(n32465), .B(n32509), .Z(n32511) );
  XNOR U32429 ( .A(n32532), .B(n32533), .Z(n32465) );
  AND U32430 ( .A(n1106), .B(n32471), .Z(n32533) );
  XOR U32431 ( .A(n32532), .B(n32469), .Z(n32471) );
  XOR U32432 ( .A(n32534), .B(n32535), .Z(n32509) );
  AND U32433 ( .A(n32536), .B(n32537), .Z(n32535) );
  XNOR U32434 ( .A(n32534), .B(n32525), .Z(n32537) );
  IV U32435 ( .A(n32479), .Z(n32525) );
  XNOR U32436 ( .A(n32538), .B(n32518), .Z(n32479) );
  XNOR U32437 ( .A(n32539), .B(n32524), .Z(n32518) );
  XNOR U32438 ( .A(n32540), .B(n32541), .Z(n32524) );
  NOR U32439 ( .A(n32542), .B(n32543), .Z(n32541) );
  XOR U32440 ( .A(n32540), .B(n32544), .Z(n32542) );
  XNOR U32441 ( .A(n32523), .B(n32515), .Z(n32539) );
  XOR U32442 ( .A(n32545), .B(n32546), .Z(n32515) );
  AND U32443 ( .A(n32547), .B(n32548), .Z(n32546) );
  XOR U32444 ( .A(n32545), .B(n32549), .Z(n32547) );
  XNOR U32445 ( .A(n32550), .B(n32520), .Z(n32523) );
  XOR U32446 ( .A(n32551), .B(n32552), .Z(n32520) );
  AND U32447 ( .A(n32553), .B(n32554), .Z(n32552) );
  XNOR U32448 ( .A(n32555), .B(n32556), .Z(n32553) );
  IV U32449 ( .A(n32551), .Z(n32555) );
  XNOR U32450 ( .A(n32557), .B(n32558), .Z(n32550) );
  NOR U32451 ( .A(n32559), .B(n32560), .Z(n32558) );
  XNOR U32452 ( .A(n32557), .B(n32561), .Z(n32559) );
  XNOR U32453 ( .A(n32519), .B(n32526), .Z(n32538) );
  NOR U32454 ( .A(n32487), .B(n32562), .Z(n32526) );
  XOR U32455 ( .A(n32531), .B(n32530), .Z(n32519) );
  XNOR U32456 ( .A(n32563), .B(n32527), .Z(n32530) );
  XOR U32457 ( .A(n32564), .B(n32565), .Z(n32527) );
  AND U32458 ( .A(n32566), .B(n32567), .Z(n32565) );
  XNOR U32459 ( .A(n32568), .B(n32569), .Z(n32566) );
  IV U32460 ( .A(n32564), .Z(n32568) );
  XNOR U32461 ( .A(n32570), .B(n32571), .Z(n32563) );
  NOR U32462 ( .A(n32572), .B(n32573), .Z(n32571) );
  XNOR U32463 ( .A(n32570), .B(n32574), .Z(n32572) );
  XOR U32464 ( .A(n32575), .B(n32576), .Z(n32531) );
  NOR U32465 ( .A(n32577), .B(n32578), .Z(n32576) );
  XNOR U32466 ( .A(n32575), .B(n32579), .Z(n32577) );
  XNOR U32467 ( .A(n32476), .B(n32534), .Z(n32536) );
  XNOR U32468 ( .A(n32580), .B(n32581), .Z(n32476) );
  AND U32469 ( .A(n1106), .B(n32483), .Z(n32581) );
  XOR U32470 ( .A(n32580), .B(n32481), .Z(n32483) );
  AND U32471 ( .A(n32484), .B(n32487), .Z(n32534) );
  XOR U32472 ( .A(n32582), .B(n32562), .Z(n32487) );
  XNOR U32473 ( .A(p_input[1552]), .B(p_input[2048]), .Z(n32562) );
  XNOR U32474 ( .A(n32549), .B(n32548), .Z(n32582) );
  XNOR U32475 ( .A(n32583), .B(n32556), .Z(n32548) );
  XNOR U32476 ( .A(n32544), .B(n32543), .Z(n32556) );
  XNOR U32477 ( .A(n32584), .B(n32540), .Z(n32543) );
  XNOR U32478 ( .A(p_input[1562]), .B(p_input[2058]), .Z(n32540) );
  XOR U32479 ( .A(p_input[1563]), .B(n16732), .Z(n32584) );
  XOR U32480 ( .A(p_input[1564]), .B(p_input[2060]), .Z(n32544) );
  XOR U32481 ( .A(n32554), .B(n32585), .Z(n32583) );
  IV U32482 ( .A(n32545), .Z(n32585) );
  XOR U32483 ( .A(p_input[1553]), .B(p_input[2049]), .Z(n32545) );
  XNOR U32484 ( .A(n32586), .B(n32561), .Z(n32554) );
  XNOR U32485 ( .A(p_input[1567]), .B(n16735), .Z(n32561) );
  XOR U32486 ( .A(n32551), .B(n32560), .Z(n32586) );
  XOR U32487 ( .A(n32587), .B(n32557), .Z(n32560) );
  XOR U32488 ( .A(p_input[1565]), .B(p_input[2061]), .Z(n32557) );
  XOR U32489 ( .A(p_input[1566]), .B(n16737), .Z(n32587) );
  XOR U32490 ( .A(p_input[1561]), .B(p_input[2057]), .Z(n32551) );
  XOR U32491 ( .A(n32569), .B(n32567), .Z(n32549) );
  XNOR U32492 ( .A(n32588), .B(n32574), .Z(n32567) );
  XOR U32493 ( .A(p_input[1560]), .B(p_input[2056]), .Z(n32574) );
  XOR U32494 ( .A(n32564), .B(n32573), .Z(n32588) );
  XOR U32495 ( .A(n32589), .B(n32570), .Z(n32573) );
  XOR U32496 ( .A(p_input[1558]), .B(p_input[2054]), .Z(n32570) );
  XOR U32497 ( .A(p_input[1559]), .B(n17722), .Z(n32589) );
  XOR U32498 ( .A(p_input[1554]), .B(p_input[2050]), .Z(n32564) );
  XNOR U32499 ( .A(n32579), .B(n32578), .Z(n32569) );
  XOR U32500 ( .A(n32590), .B(n32575), .Z(n32578) );
  XOR U32501 ( .A(p_input[1555]), .B(p_input[2051]), .Z(n32575) );
  XOR U32502 ( .A(p_input[1556]), .B(n17724), .Z(n32590) );
  XOR U32503 ( .A(p_input[1557]), .B(p_input[2053]), .Z(n32579) );
  XNOR U32504 ( .A(n32591), .B(n32592), .Z(n32484) );
  AND U32505 ( .A(n1106), .B(n32593), .Z(n32592) );
  XNOR U32506 ( .A(n32594), .B(n32595), .Z(n1106) );
  AND U32507 ( .A(n32596), .B(n32597), .Z(n32595) );
  XOR U32508 ( .A(n32594), .B(n32494), .Z(n32597) );
  XNOR U32509 ( .A(n32594), .B(n32448), .Z(n32596) );
  XOR U32510 ( .A(n32598), .B(n32599), .Z(n32594) );
  AND U32511 ( .A(n32600), .B(n32601), .Z(n32599) );
  XOR U32512 ( .A(n32598), .B(n32458), .Z(n32600) );
  XOR U32513 ( .A(n32602), .B(n32603), .Z(n32437) );
  AND U32514 ( .A(n1110), .B(n32593), .Z(n32603) );
  XNOR U32515 ( .A(n32591), .B(n32602), .Z(n32593) );
  XNOR U32516 ( .A(n32604), .B(n32605), .Z(n1110) );
  AND U32517 ( .A(n32606), .B(n32607), .Z(n32605) );
  XNOR U32518 ( .A(n32608), .B(n32604), .Z(n32607) );
  IV U32519 ( .A(n32494), .Z(n32608) );
  XNOR U32520 ( .A(n32609), .B(n32610), .Z(n32494) );
  AND U32521 ( .A(n1113), .B(n32611), .Z(n32610) );
  XNOR U32522 ( .A(n32609), .B(n32612), .Z(n32611) );
  XNOR U32523 ( .A(n32448), .B(n32604), .Z(n32606) );
  XOR U32524 ( .A(n32613), .B(n32614), .Z(n32448) );
  AND U32525 ( .A(n1121), .B(n32615), .Z(n32614) );
  XOR U32526 ( .A(n32598), .B(n32616), .Z(n32604) );
  AND U32527 ( .A(n32617), .B(n32601), .Z(n32616) );
  XNOR U32528 ( .A(n32507), .B(n32598), .Z(n32601) );
  XNOR U32529 ( .A(n32618), .B(n32619), .Z(n32507) );
  AND U32530 ( .A(n1113), .B(n32620), .Z(n32619) );
  XOR U32531 ( .A(n32621), .B(n32618), .Z(n32620) );
  XNOR U32532 ( .A(n32622), .B(n32598), .Z(n32617) );
  IV U32533 ( .A(n32458), .Z(n32622) );
  XOR U32534 ( .A(n32623), .B(n32624), .Z(n32458) );
  AND U32535 ( .A(n1121), .B(n32625), .Z(n32624) );
  XOR U32536 ( .A(n32626), .B(n32627), .Z(n32598) );
  AND U32537 ( .A(n32628), .B(n32629), .Z(n32627) );
  XNOR U32538 ( .A(n32532), .B(n32626), .Z(n32629) );
  XNOR U32539 ( .A(n32630), .B(n32631), .Z(n32532) );
  AND U32540 ( .A(n1113), .B(n32632), .Z(n32631) );
  XNOR U32541 ( .A(n32633), .B(n32630), .Z(n32632) );
  XOR U32542 ( .A(n32626), .B(n32469), .Z(n32628) );
  XOR U32543 ( .A(n32634), .B(n32635), .Z(n32469) );
  AND U32544 ( .A(n1121), .B(n32636), .Z(n32635) );
  XOR U32545 ( .A(n32637), .B(n32638), .Z(n32626) );
  AND U32546 ( .A(n32639), .B(n32640), .Z(n32638) );
  XNOR U32547 ( .A(n32637), .B(n32580), .Z(n32640) );
  XNOR U32548 ( .A(n32641), .B(n32642), .Z(n32580) );
  AND U32549 ( .A(n1113), .B(n32643), .Z(n32642) );
  XOR U32550 ( .A(n32644), .B(n32641), .Z(n32643) );
  XNOR U32551 ( .A(n32645), .B(n32637), .Z(n32639) );
  IV U32552 ( .A(n32481), .Z(n32645) );
  XOR U32553 ( .A(n32646), .B(n32647), .Z(n32481) );
  AND U32554 ( .A(n1121), .B(n32648), .Z(n32647) );
  AND U32555 ( .A(n32602), .B(n32591), .Z(n32637) );
  XNOR U32556 ( .A(n32649), .B(n32650), .Z(n32591) );
  AND U32557 ( .A(n1113), .B(n32651), .Z(n32650) );
  XNOR U32558 ( .A(n32652), .B(n32649), .Z(n32651) );
  XNOR U32559 ( .A(n32653), .B(n32654), .Z(n1113) );
  AND U32560 ( .A(n32655), .B(n32656), .Z(n32654) );
  XOR U32561 ( .A(n32612), .B(n32653), .Z(n32656) );
  AND U32562 ( .A(n32657), .B(n32658), .Z(n32612) );
  XOR U32563 ( .A(n32653), .B(n32609), .Z(n32655) );
  XNOR U32564 ( .A(n32659), .B(n32660), .Z(n32609) );
  AND U32565 ( .A(n1117), .B(n32615), .Z(n32660) );
  XOR U32566 ( .A(n32613), .B(n32659), .Z(n32615) );
  XOR U32567 ( .A(n32661), .B(n32662), .Z(n32653) );
  AND U32568 ( .A(n32663), .B(n32664), .Z(n32662) );
  XNOR U32569 ( .A(n32661), .B(n32657), .Z(n32664) );
  IV U32570 ( .A(n32621), .Z(n32657) );
  XOR U32571 ( .A(n32665), .B(n32666), .Z(n32621) );
  XOR U32572 ( .A(n32667), .B(n32658), .Z(n32666) );
  AND U32573 ( .A(n32633), .B(n32668), .Z(n32658) );
  AND U32574 ( .A(n32669), .B(n32670), .Z(n32667) );
  XOR U32575 ( .A(n32671), .B(n32665), .Z(n32669) );
  XNOR U32576 ( .A(n32618), .B(n32661), .Z(n32663) );
  XNOR U32577 ( .A(n32672), .B(n32673), .Z(n32618) );
  AND U32578 ( .A(n1117), .B(n32625), .Z(n32673) );
  XOR U32579 ( .A(n32672), .B(n32623), .Z(n32625) );
  XOR U32580 ( .A(n32674), .B(n32675), .Z(n32661) );
  AND U32581 ( .A(n32676), .B(n32677), .Z(n32675) );
  XNOR U32582 ( .A(n32674), .B(n32633), .Z(n32677) );
  XOR U32583 ( .A(n32678), .B(n32670), .Z(n32633) );
  XNOR U32584 ( .A(n32679), .B(n32665), .Z(n32670) );
  XOR U32585 ( .A(n32680), .B(n32681), .Z(n32665) );
  AND U32586 ( .A(n32682), .B(n32683), .Z(n32681) );
  XOR U32587 ( .A(n32684), .B(n32680), .Z(n32682) );
  XNOR U32588 ( .A(n32685), .B(n32686), .Z(n32679) );
  AND U32589 ( .A(n32687), .B(n32688), .Z(n32686) );
  XOR U32590 ( .A(n32685), .B(n32689), .Z(n32687) );
  XNOR U32591 ( .A(n32671), .B(n32668), .Z(n32678) );
  AND U32592 ( .A(n32690), .B(n32691), .Z(n32668) );
  XOR U32593 ( .A(n32692), .B(n32693), .Z(n32671) );
  AND U32594 ( .A(n32694), .B(n32695), .Z(n32693) );
  XOR U32595 ( .A(n32692), .B(n32696), .Z(n32694) );
  XNOR U32596 ( .A(n32630), .B(n32674), .Z(n32676) );
  XNOR U32597 ( .A(n32697), .B(n32698), .Z(n32630) );
  AND U32598 ( .A(n1117), .B(n32636), .Z(n32698) );
  XOR U32599 ( .A(n32697), .B(n32634), .Z(n32636) );
  XOR U32600 ( .A(n32699), .B(n32700), .Z(n32674) );
  AND U32601 ( .A(n32701), .B(n32702), .Z(n32700) );
  XNOR U32602 ( .A(n32699), .B(n32690), .Z(n32702) );
  IV U32603 ( .A(n32644), .Z(n32690) );
  XNOR U32604 ( .A(n32703), .B(n32683), .Z(n32644) );
  XNOR U32605 ( .A(n32704), .B(n32689), .Z(n32683) );
  XNOR U32606 ( .A(n32705), .B(n32706), .Z(n32689) );
  NOR U32607 ( .A(n32707), .B(n32708), .Z(n32706) );
  XOR U32608 ( .A(n32705), .B(n32709), .Z(n32707) );
  XNOR U32609 ( .A(n32688), .B(n32680), .Z(n32704) );
  XOR U32610 ( .A(n32710), .B(n32711), .Z(n32680) );
  AND U32611 ( .A(n32712), .B(n32713), .Z(n32711) );
  XOR U32612 ( .A(n32710), .B(n32714), .Z(n32712) );
  XNOR U32613 ( .A(n32715), .B(n32685), .Z(n32688) );
  XOR U32614 ( .A(n32716), .B(n32717), .Z(n32685) );
  AND U32615 ( .A(n32718), .B(n32719), .Z(n32717) );
  XNOR U32616 ( .A(n32720), .B(n32721), .Z(n32718) );
  IV U32617 ( .A(n32716), .Z(n32720) );
  XNOR U32618 ( .A(n32722), .B(n32723), .Z(n32715) );
  NOR U32619 ( .A(n32724), .B(n32725), .Z(n32723) );
  XNOR U32620 ( .A(n32722), .B(n32726), .Z(n32724) );
  XNOR U32621 ( .A(n32684), .B(n32691), .Z(n32703) );
  NOR U32622 ( .A(n32652), .B(n32727), .Z(n32691) );
  XOR U32623 ( .A(n32696), .B(n32695), .Z(n32684) );
  XNOR U32624 ( .A(n32728), .B(n32692), .Z(n32695) );
  XOR U32625 ( .A(n32729), .B(n32730), .Z(n32692) );
  AND U32626 ( .A(n32731), .B(n32732), .Z(n32730) );
  XNOR U32627 ( .A(n32733), .B(n32734), .Z(n32731) );
  IV U32628 ( .A(n32729), .Z(n32733) );
  XNOR U32629 ( .A(n32735), .B(n32736), .Z(n32728) );
  NOR U32630 ( .A(n32737), .B(n32738), .Z(n32736) );
  XNOR U32631 ( .A(n32735), .B(n32739), .Z(n32737) );
  XOR U32632 ( .A(n32740), .B(n32741), .Z(n32696) );
  NOR U32633 ( .A(n32742), .B(n32743), .Z(n32741) );
  XNOR U32634 ( .A(n32740), .B(n32744), .Z(n32742) );
  XNOR U32635 ( .A(n32641), .B(n32699), .Z(n32701) );
  XNOR U32636 ( .A(n32745), .B(n32746), .Z(n32641) );
  AND U32637 ( .A(n1117), .B(n32648), .Z(n32746) );
  XOR U32638 ( .A(n32745), .B(n32646), .Z(n32648) );
  AND U32639 ( .A(n32649), .B(n32652), .Z(n32699) );
  XOR U32640 ( .A(n32747), .B(n32727), .Z(n32652) );
  XNOR U32641 ( .A(p_input[1568]), .B(p_input[2048]), .Z(n32727) );
  XNOR U32642 ( .A(n32714), .B(n32713), .Z(n32747) );
  XNOR U32643 ( .A(n32748), .B(n32721), .Z(n32713) );
  XNOR U32644 ( .A(n32709), .B(n32708), .Z(n32721) );
  XNOR U32645 ( .A(n32749), .B(n32705), .Z(n32708) );
  XNOR U32646 ( .A(p_input[1578]), .B(p_input[2058]), .Z(n32705) );
  XOR U32647 ( .A(p_input[1579]), .B(n16732), .Z(n32749) );
  XOR U32648 ( .A(p_input[1580]), .B(p_input[2060]), .Z(n32709) );
  XOR U32649 ( .A(n32719), .B(n32750), .Z(n32748) );
  IV U32650 ( .A(n32710), .Z(n32750) );
  XOR U32651 ( .A(p_input[1569]), .B(p_input[2049]), .Z(n32710) );
  XNOR U32652 ( .A(n32751), .B(n32726), .Z(n32719) );
  XNOR U32653 ( .A(p_input[1583]), .B(n16735), .Z(n32726) );
  XOR U32654 ( .A(n32716), .B(n32725), .Z(n32751) );
  XOR U32655 ( .A(n32752), .B(n32722), .Z(n32725) );
  XOR U32656 ( .A(p_input[1581]), .B(p_input[2061]), .Z(n32722) );
  XOR U32657 ( .A(p_input[1582]), .B(n16737), .Z(n32752) );
  XOR U32658 ( .A(p_input[1577]), .B(p_input[2057]), .Z(n32716) );
  XOR U32659 ( .A(n32734), .B(n32732), .Z(n32714) );
  XNOR U32660 ( .A(n32753), .B(n32739), .Z(n32732) );
  XOR U32661 ( .A(p_input[1576]), .B(p_input[2056]), .Z(n32739) );
  XOR U32662 ( .A(n32729), .B(n32738), .Z(n32753) );
  XOR U32663 ( .A(n32754), .B(n32735), .Z(n32738) );
  XOR U32664 ( .A(p_input[1574]), .B(p_input[2054]), .Z(n32735) );
  XOR U32665 ( .A(p_input[1575]), .B(n17722), .Z(n32754) );
  XOR U32666 ( .A(p_input[1570]), .B(p_input[2050]), .Z(n32729) );
  XNOR U32667 ( .A(n32744), .B(n32743), .Z(n32734) );
  XOR U32668 ( .A(n32755), .B(n32740), .Z(n32743) );
  XOR U32669 ( .A(p_input[1571]), .B(p_input[2051]), .Z(n32740) );
  XOR U32670 ( .A(p_input[1572]), .B(n17724), .Z(n32755) );
  XOR U32671 ( .A(p_input[1573]), .B(p_input[2053]), .Z(n32744) );
  XNOR U32672 ( .A(n32756), .B(n32757), .Z(n32649) );
  AND U32673 ( .A(n1117), .B(n32758), .Z(n32757) );
  XNOR U32674 ( .A(n32759), .B(n32760), .Z(n1117) );
  AND U32675 ( .A(n32761), .B(n32762), .Z(n32760) );
  XOR U32676 ( .A(n32759), .B(n32659), .Z(n32762) );
  XNOR U32677 ( .A(n32759), .B(n32613), .Z(n32761) );
  XOR U32678 ( .A(n32763), .B(n32764), .Z(n32759) );
  AND U32679 ( .A(n32765), .B(n32766), .Z(n32764) );
  XOR U32680 ( .A(n32763), .B(n32623), .Z(n32765) );
  XOR U32681 ( .A(n32767), .B(n32768), .Z(n32602) );
  AND U32682 ( .A(n1121), .B(n32758), .Z(n32768) );
  XNOR U32683 ( .A(n32756), .B(n32767), .Z(n32758) );
  XNOR U32684 ( .A(n32769), .B(n32770), .Z(n1121) );
  AND U32685 ( .A(n32771), .B(n32772), .Z(n32770) );
  XNOR U32686 ( .A(n32773), .B(n32769), .Z(n32772) );
  IV U32687 ( .A(n32659), .Z(n32773) );
  XNOR U32688 ( .A(n32774), .B(n32775), .Z(n32659) );
  AND U32689 ( .A(n1124), .B(n32776), .Z(n32775) );
  XNOR U32690 ( .A(n32774), .B(n32777), .Z(n32776) );
  XNOR U32691 ( .A(n32613), .B(n32769), .Z(n32771) );
  XOR U32692 ( .A(n32778), .B(n32779), .Z(n32613) );
  AND U32693 ( .A(n1132), .B(n32780), .Z(n32779) );
  XOR U32694 ( .A(n32763), .B(n32781), .Z(n32769) );
  AND U32695 ( .A(n32782), .B(n32766), .Z(n32781) );
  XNOR U32696 ( .A(n32672), .B(n32763), .Z(n32766) );
  XNOR U32697 ( .A(n32783), .B(n32784), .Z(n32672) );
  AND U32698 ( .A(n1124), .B(n32785), .Z(n32784) );
  XOR U32699 ( .A(n32786), .B(n32783), .Z(n32785) );
  XNOR U32700 ( .A(n32787), .B(n32763), .Z(n32782) );
  IV U32701 ( .A(n32623), .Z(n32787) );
  XOR U32702 ( .A(n32788), .B(n32789), .Z(n32623) );
  AND U32703 ( .A(n1132), .B(n32790), .Z(n32789) );
  XOR U32704 ( .A(n32791), .B(n32792), .Z(n32763) );
  AND U32705 ( .A(n32793), .B(n32794), .Z(n32792) );
  XNOR U32706 ( .A(n32697), .B(n32791), .Z(n32794) );
  XNOR U32707 ( .A(n32795), .B(n32796), .Z(n32697) );
  AND U32708 ( .A(n1124), .B(n32797), .Z(n32796) );
  XNOR U32709 ( .A(n32798), .B(n32795), .Z(n32797) );
  XOR U32710 ( .A(n32791), .B(n32634), .Z(n32793) );
  XOR U32711 ( .A(n32799), .B(n32800), .Z(n32634) );
  AND U32712 ( .A(n1132), .B(n32801), .Z(n32800) );
  XOR U32713 ( .A(n32802), .B(n32803), .Z(n32791) );
  AND U32714 ( .A(n32804), .B(n32805), .Z(n32803) );
  XNOR U32715 ( .A(n32802), .B(n32745), .Z(n32805) );
  XNOR U32716 ( .A(n32806), .B(n32807), .Z(n32745) );
  AND U32717 ( .A(n1124), .B(n32808), .Z(n32807) );
  XOR U32718 ( .A(n32809), .B(n32806), .Z(n32808) );
  XNOR U32719 ( .A(n32810), .B(n32802), .Z(n32804) );
  IV U32720 ( .A(n32646), .Z(n32810) );
  XOR U32721 ( .A(n32811), .B(n32812), .Z(n32646) );
  AND U32722 ( .A(n1132), .B(n32813), .Z(n32812) );
  AND U32723 ( .A(n32767), .B(n32756), .Z(n32802) );
  XNOR U32724 ( .A(n32814), .B(n32815), .Z(n32756) );
  AND U32725 ( .A(n1124), .B(n32816), .Z(n32815) );
  XNOR U32726 ( .A(n32817), .B(n32814), .Z(n32816) );
  XNOR U32727 ( .A(n32818), .B(n32819), .Z(n1124) );
  AND U32728 ( .A(n32820), .B(n32821), .Z(n32819) );
  XOR U32729 ( .A(n32777), .B(n32818), .Z(n32821) );
  AND U32730 ( .A(n32822), .B(n32823), .Z(n32777) );
  XOR U32731 ( .A(n32818), .B(n32774), .Z(n32820) );
  XNOR U32732 ( .A(n32824), .B(n32825), .Z(n32774) );
  AND U32733 ( .A(n1128), .B(n32780), .Z(n32825) );
  XOR U32734 ( .A(n32778), .B(n32824), .Z(n32780) );
  XOR U32735 ( .A(n32826), .B(n32827), .Z(n32818) );
  AND U32736 ( .A(n32828), .B(n32829), .Z(n32827) );
  XNOR U32737 ( .A(n32826), .B(n32822), .Z(n32829) );
  IV U32738 ( .A(n32786), .Z(n32822) );
  XOR U32739 ( .A(n32830), .B(n32831), .Z(n32786) );
  XOR U32740 ( .A(n32832), .B(n32823), .Z(n32831) );
  AND U32741 ( .A(n32798), .B(n32833), .Z(n32823) );
  AND U32742 ( .A(n32834), .B(n32835), .Z(n32832) );
  XOR U32743 ( .A(n32836), .B(n32830), .Z(n32834) );
  XNOR U32744 ( .A(n32783), .B(n32826), .Z(n32828) );
  XNOR U32745 ( .A(n32837), .B(n32838), .Z(n32783) );
  AND U32746 ( .A(n1128), .B(n32790), .Z(n32838) );
  XOR U32747 ( .A(n32837), .B(n32788), .Z(n32790) );
  XOR U32748 ( .A(n32839), .B(n32840), .Z(n32826) );
  AND U32749 ( .A(n32841), .B(n32842), .Z(n32840) );
  XNOR U32750 ( .A(n32839), .B(n32798), .Z(n32842) );
  XOR U32751 ( .A(n32843), .B(n32835), .Z(n32798) );
  XNOR U32752 ( .A(n32844), .B(n32830), .Z(n32835) );
  XOR U32753 ( .A(n32845), .B(n32846), .Z(n32830) );
  AND U32754 ( .A(n32847), .B(n32848), .Z(n32846) );
  XOR U32755 ( .A(n32849), .B(n32845), .Z(n32847) );
  XNOR U32756 ( .A(n32850), .B(n32851), .Z(n32844) );
  AND U32757 ( .A(n32852), .B(n32853), .Z(n32851) );
  XOR U32758 ( .A(n32850), .B(n32854), .Z(n32852) );
  XNOR U32759 ( .A(n32836), .B(n32833), .Z(n32843) );
  AND U32760 ( .A(n32855), .B(n32856), .Z(n32833) );
  XOR U32761 ( .A(n32857), .B(n32858), .Z(n32836) );
  AND U32762 ( .A(n32859), .B(n32860), .Z(n32858) );
  XOR U32763 ( .A(n32857), .B(n32861), .Z(n32859) );
  XNOR U32764 ( .A(n32795), .B(n32839), .Z(n32841) );
  XNOR U32765 ( .A(n32862), .B(n32863), .Z(n32795) );
  AND U32766 ( .A(n1128), .B(n32801), .Z(n32863) );
  XOR U32767 ( .A(n32862), .B(n32799), .Z(n32801) );
  XOR U32768 ( .A(n32864), .B(n32865), .Z(n32839) );
  AND U32769 ( .A(n32866), .B(n32867), .Z(n32865) );
  XNOR U32770 ( .A(n32864), .B(n32855), .Z(n32867) );
  IV U32771 ( .A(n32809), .Z(n32855) );
  XNOR U32772 ( .A(n32868), .B(n32848), .Z(n32809) );
  XNOR U32773 ( .A(n32869), .B(n32854), .Z(n32848) );
  XNOR U32774 ( .A(n32870), .B(n32871), .Z(n32854) );
  NOR U32775 ( .A(n32872), .B(n32873), .Z(n32871) );
  XOR U32776 ( .A(n32870), .B(n32874), .Z(n32872) );
  XNOR U32777 ( .A(n32853), .B(n32845), .Z(n32869) );
  XOR U32778 ( .A(n32875), .B(n32876), .Z(n32845) );
  AND U32779 ( .A(n32877), .B(n32878), .Z(n32876) );
  XOR U32780 ( .A(n32875), .B(n32879), .Z(n32877) );
  XNOR U32781 ( .A(n32880), .B(n32850), .Z(n32853) );
  XOR U32782 ( .A(n32881), .B(n32882), .Z(n32850) );
  AND U32783 ( .A(n32883), .B(n32884), .Z(n32882) );
  XNOR U32784 ( .A(n32885), .B(n32886), .Z(n32883) );
  IV U32785 ( .A(n32881), .Z(n32885) );
  XNOR U32786 ( .A(n32887), .B(n32888), .Z(n32880) );
  NOR U32787 ( .A(n32889), .B(n32890), .Z(n32888) );
  XNOR U32788 ( .A(n32887), .B(n32891), .Z(n32889) );
  XNOR U32789 ( .A(n32849), .B(n32856), .Z(n32868) );
  NOR U32790 ( .A(n32817), .B(n32892), .Z(n32856) );
  XOR U32791 ( .A(n32861), .B(n32860), .Z(n32849) );
  XNOR U32792 ( .A(n32893), .B(n32857), .Z(n32860) );
  XOR U32793 ( .A(n32894), .B(n32895), .Z(n32857) );
  AND U32794 ( .A(n32896), .B(n32897), .Z(n32895) );
  XNOR U32795 ( .A(n32898), .B(n32899), .Z(n32896) );
  IV U32796 ( .A(n32894), .Z(n32898) );
  XNOR U32797 ( .A(n32900), .B(n32901), .Z(n32893) );
  NOR U32798 ( .A(n32902), .B(n32903), .Z(n32901) );
  XNOR U32799 ( .A(n32900), .B(n32904), .Z(n32902) );
  XOR U32800 ( .A(n32905), .B(n32906), .Z(n32861) );
  NOR U32801 ( .A(n32907), .B(n32908), .Z(n32906) );
  XNOR U32802 ( .A(n32905), .B(n32909), .Z(n32907) );
  XNOR U32803 ( .A(n32806), .B(n32864), .Z(n32866) );
  XNOR U32804 ( .A(n32910), .B(n32911), .Z(n32806) );
  AND U32805 ( .A(n1128), .B(n32813), .Z(n32911) );
  XOR U32806 ( .A(n32910), .B(n32811), .Z(n32813) );
  AND U32807 ( .A(n32814), .B(n32817), .Z(n32864) );
  XOR U32808 ( .A(n32912), .B(n32892), .Z(n32817) );
  XNOR U32809 ( .A(p_input[1584]), .B(p_input[2048]), .Z(n32892) );
  XNOR U32810 ( .A(n32879), .B(n32878), .Z(n32912) );
  XNOR U32811 ( .A(n32913), .B(n32886), .Z(n32878) );
  XNOR U32812 ( .A(n32874), .B(n32873), .Z(n32886) );
  XNOR U32813 ( .A(n32914), .B(n32870), .Z(n32873) );
  XNOR U32814 ( .A(p_input[1594]), .B(p_input[2058]), .Z(n32870) );
  XOR U32815 ( .A(p_input[1595]), .B(n16732), .Z(n32914) );
  XOR U32816 ( .A(p_input[1596]), .B(p_input[2060]), .Z(n32874) );
  XOR U32817 ( .A(n32884), .B(n32915), .Z(n32913) );
  IV U32818 ( .A(n32875), .Z(n32915) );
  XOR U32819 ( .A(p_input[1585]), .B(p_input[2049]), .Z(n32875) );
  XNOR U32820 ( .A(n32916), .B(n32891), .Z(n32884) );
  XNOR U32821 ( .A(p_input[1599]), .B(n16735), .Z(n32891) );
  XOR U32822 ( .A(n32881), .B(n32890), .Z(n32916) );
  XOR U32823 ( .A(n32917), .B(n32887), .Z(n32890) );
  XOR U32824 ( .A(p_input[1597]), .B(p_input[2061]), .Z(n32887) );
  XOR U32825 ( .A(p_input[1598]), .B(n16737), .Z(n32917) );
  XOR U32826 ( .A(p_input[1593]), .B(p_input[2057]), .Z(n32881) );
  XOR U32827 ( .A(n32899), .B(n32897), .Z(n32879) );
  XNOR U32828 ( .A(n32918), .B(n32904), .Z(n32897) );
  XOR U32829 ( .A(p_input[1592]), .B(p_input[2056]), .Z(n32904) );
  XOR U32830 ( .A(n32894), .B(n32903), .Z(n32918) );
  XOR U32831 ( .A(n32919), .B(n32900), .Z(n32903) );
  XOR U32832 ( .A(p_input[1590]), .B(p_input[2054]), .Z(n32900) );
  XOR U32833 ( .A(p_input[1591]), .B(n17722), .Z(n32919) );
  XOR U32834 ( .A(p_input[1586]), .B(p_input[2050]), .Z(n32894) );
  XNOR U32835 ( .A(n32909), .B(n32908), .Z(n32899) );
  XOR U32836 ( .A(n32920), .B(n32905), .Z(n32908) );
  XOR U32837 ( .A(p_input[1587]), .B(p_input[2051]), .Z(n32905) );
  XOR U32838 ( .A(p_input[1588]), .B(n17724), .Z(n32920) );
  XOR U32839 ( .A(p_input[1589]), .B(p_input[2053]), .Z(n32909) );
  XNOR U32840 ( .A(n32921), .B(n32922), .Z(n32814) );
  AND U32841 ( .A(n1128), .B(n32923), .Z(n32922) );
  XNOR U32842 ( .A(n32924), .B(n32925), .Z(n1128) );
  AND U32843 ( .A(n32926), .B(n32927), .Z(n32925) );
  XOR U32844 ( .A(n32924), .B(n32824), .Z(n32927) );
  XNOR U32845 ( .A(n32924), .B(n32778), .Z(n32926) );
  XOR U32846 ( .A(n32928), .B(n32929), .Z(n32924) );
  AND U32847 ( .A(n32930), .B(n32931), .Z(n32929) );
  XOR U32848 ( .A(n32928), .B(n32788), .Z(n32930) );
  XOR U32849 ( .A(n32932), .B(n32933), .Z(n32767) );
  AND U32850 ( .A(n1132), .B(n32923), .Z(n32933) );
  XNOR U32851 ( .A(n32921), .B(n32932), .Z(n32923) );
  XNOR U32852 ( .A(n32934), .B(n32935), .Z(n1132) );
  AND U32853 ( .A(n32936), .B(n32937), .Z(n32935) );
  XNOR U32854 ( .A(n32938), .B(n32934), .Z(n32937) );
  IV U32855 ( .A(n32824), .Z(n32938) );
  XNOR U32856 ( .A(n32939), .B(n32940), .Z(n32824) );
  AND U32857 ( .A(n1135), .B(n32941), .Z(n32940) );
  XNOR U32858 ( .A(n32939), .B(n32942), .Z(n32941) );
  XNOR U32859 ( .A(n32778), .B(n32934), .Z(n32936) );
  XOR U32860 ( .A(n32943), .B(n32944), .Z(n32778) );
  AND U32861 ( .A(n1143), .B(n32945), .Z(n32944) );
  XOR U32862 ( .A(n32928), .B(n32946), .Z(n32934) );
  AND U32863 ( .A(n32947), .B(n32931), .Z(n32946) );
  XNOR U32864 ( .A(n32837), .B(n32928), .Z(n32931) );
  XNOR U32865 ( .A(n32948), .B(n32949), .Z(n32837) );
  AND U32866 ( .A(n1135), .B(n32950), .Z(n32949) );
  XOR U32867 ( .A(n32951), .B(n32948), .Z(n32950) );
  XNOR U32868 ( .A(n32952), .B(n32928), .Z(n32947) );
  IV U32869 ( .A(n32788), .Z(n32952) );
  XOR U32870 ( .A(n32953), .B(n32954), .Z(n32788) );
  AND U32871 ( .A(n1143), .B(n32955), .Z(n32954) );
  XOR U32872 ( .A(n32956), .B(n32957), .Z(n32928) );
  AND U32873 ( .A(n32958), .B(n32959), .Z(n32957) );
  XNOR U32874 ( .A(n32862), .B(n32956), .Z(n32959) );
  XNOR U32875 ( .A(n32960), .B(n32961), .Z(n32862) );
  AND U32876 ( .A(n1135), .B(n32962), .Z(n32961) );
  XNOR U32877 ( .A(n32963), .B(n32960), .Z(n32962) );
  XOR U32878 ( .A(n32956), .B(n32799), .Z(n32958) );
  XOR U32879 ( .A(n32964), .B(n32965), .Z(n32799) );
  AND U32880 ( .A(n1143), .B(n32966), .Z(n32965) );
  XOR U32881 ( .A(n32967), .B(n32968), .Z(n32956) );
  AND U32882 ( .A(n32969), .B(n32970), .Z(n32968) );
  XNOR U32883 ( .A(n32967), .B(n32910), .Z(n32970) );
  XNOR U32884 ( .A(n32971), .B(n32972), .Z(n32910) );
  AND U32885 ( .A(n1135), .B(n32973), .Z(n32972) );
  XOR U32886 ( .A(n32974), .B(n32971), .Z(n32973) );
  XNOR U32887 ( .A(n32975), .B(n32967), .Z(n32969) );
  IV U32888 ( .A(n32811), .Z(n32975) );
  XOR U32889 ( .A(n32976), .B(n32977), .Z(n32811) );
  AND U32890 ( .A(n1143), .B(n32978), .Z(n32977) );
  AND U32891 ( .A(n32932), .B(n32921), .Z(n32967) );
  XNOR U32892 ( .A(n32979), .B(n32980), .Z(n32921) );
  AND U32893 ( .A(n1135), .B(n32981), .Z(n32980) );
  XNOR U32894 ( .A(n32982), .B(n32979), .Z(n32981) );
  XNOR U32895 ( .A(n32983), .B(n32984), .Z(n1135) );
  AND U32896 ( .A(n32985), .B(n32986), .Z(n32984) );
  XOR U32897 ( .A(n32942), .B(n32983), .Z(n32986) );
  AND U32898 ( .A(n32987), .B(n32988), .Z(n32942) );
  XOR U32899 ( .A(n32983), .B(n32939), .Z(n32985) );
  XNOR U32900 ( .A(n32989), .B(n32990), .Z(n32939) );
  AND U32901 ( .A(n1139), .B(n32945), .Z(n32990) );
  XOR U32902 ( .A(n32943), .B(n32989), .Z(n32945) );
  XOR U32903 ( .A(n32991), .B(n32992), .Z(n32983) );
  AND U32904 ( .A(n32993), .B(n32994), .Z(n32992) );
  XNOR U32905 ( .A(n32991), .B(n32987), .Z(n32994) );
  IV U32906 ( .A(n32951), .Z(n32987) );
  XOR U32907 ( .A(n32995), .B(n32996), .Z(n32951) );
  XOR U32908 ( .A(n32997), .B(n32988), .Z(n32996) );
  AND U32909 ( .A(n32963), .B(n32998), .Z(n32988) );
  AND U32910 ( .A(n32999), .B(n33000), .Z(n32997) );
  XOR U32911 ( .A(n33001), .B(n32995), .Z(n32999) );
  XNOR U32912 ( .A(n32948), .B(n32991), .Z(n32993) );
  XNOR U32913 ( .A(n33002), .B(n33003), .Z(n32948) );
  AND U32914 ( .A(n1139), .B(n32955), .Z(n33003) );
  XOR U32915 ( .A(n33002), .B(n32953), .Z(n32955) );
  XOR U32916 ( .A(n33004), .B(n33005), .Z(n32991) );
  AND U32917 ( .A(n33006), .B(n33007), .Z(n33005) );
  XNOR U32918 ( .A(n33004), .B(n32963), .Z(n33007) );
  XOR U32919 ( .A(n33008), .B(n33000), .Z(n32963) );
  XNOR U32920 ( .A(n33009), .B(n32995), .Z(n33000) );
  XOR U32921 ( .A(n33010), .B(n33011), .Z(n32995) );
  AND U32922 ( .A(n33012), .B(n33013), .Z(n33011) );
  XOR U32923 ( .A(n33014), .B(n33010), .Z(n33012) );
  XNOR U32924 ( .A(n33015), .B(n33016), .Z(n33009) );
  AND U32925 ( .A(n33017), .B(n33018), .Z(n33016) );
  XOR U32926 ( .A(n33015), .B(n33019), .Z(n33017) );
  XNOR U32927 ( .A(n33001), .B(n32998), .Z(n33008) );
  AND U32928 ( .A(n33020), .B(n33021), .Z(n32998) );
  XOR U32929 ( .A(n33022), .B(n33023), .Z(n33001) );
  AND U32930 ( .A(n33024), .B(n33025), .Z(n33023) );
  XOR U32931 ( .A(n33022), .B(n33026), .Z(n33024) );
  XNOR U32932 ( .A(n32960), .B(n33004), .Z(n33006) );
  XNOR U32933 ( .A(n33027), .B(n33028), .Z(n32960) );
  AND U32934 ( .A(n1139), .B(n32966), .Z(n33028) );
  XOR U32935 ( .A(n33027), .B(n32964), .Z(n32966) );
  XOR U32936 ( .A(n33029), .B(n33030), .Z(n33004) );
  AND U32937 ( .A(n33031), .B(n33032), .Z(n33030) );
  XNOR U32938 ( .A(n33029), .B(n33020), .Z(n33032) );
  IV U32939 ( .A(n32974), .Z(n33020) );
  XNOR U32940 ( .A(n33033), .B(n33013), .Z(n32974) );
  XNOR U32941 ( .A(n33034), .B(n33019), .Z(n33013) );
  XNOR U32942 ( .A(n33035), .B(n33036), .Z(n33019) );
  NOR U32943 ( .A(n33037), .B(n33038), .Z(n33036) );
  XOR U32944 ( .A(n33035), .B(n33039), .Z(n33037) );
  XNOR U32945 ( .A(n33018), .B(n33010), .Z(n33034) );
  XOR U32946 ( .A(n33040), .B(n33041), .Z(n33010) );
  AND U32947 ( .A(n33042), .B(n33043), .Z(n33041) );
  XOR U32948 ( .A(n33040), .B(n33044), .Z(n33042) );
  XNOR U32949 ( .A(n33045), .B(n33015), .Z(n33018) );
  XOR U32950 ( .A(n33046), .B(n33047), .Z(n33015) );
  AND U32951 ( .A(n33048), .B(n33049), .Z(n33047) );
  XNOR U32952 ( .A(n33050), .B(n33051), .Z(n33048) );
  IV U32953 ( .A(n33046), .Z(n33050) );
  XNOR U32954 ( .A(n33052), .B(n33053), .Z(n33045) );
  NOR U32955 ( .A(n33054), .B(n33055), .Z(n33053) );
  XNOR U32956 ( .A(n33052), .B(n33056), .Z(n33054) );
  XNOR U32957 ( .A(n33014), .B(n33021), .Z(n33033) );
  NOR U32958 ( .A(n32982), .B(n33057), .Z(n33021) );
  XOR U32959 ( .A(n33026), .B(n33025), .Z(n33014) );
  XNOR U32960 ( .A(n33058), .B(n33022), .Z(n33025) );
  XOR U32961 ( .A(n33059), .B(n33060), .Z(n33022) );
  AND U32962 ( .A(n33061), .B(n33062), .Z(n33060) );
  XNOR U32963 ( .A(n33063), .B(n33064), .Z(n33061) );
  IV U32964 ( .A(n33059), .Z(n33063) );
  XNOR U32965 ( .A(n33065), .B(n33066), .Z(n33058) );
  NOR U32966 ( .A(n33067), .B(n33068), .Z(n33066) );
  XNOR U32967 ( .A(n33065), .B(n33069), .Z(n33067) );
  XOR U32968 ( .A(n33070), .B(n33071), .Z(n33026) );
  NOR U32969 ( .A(n33072), .B(n33073), .Z(n33071) );
  XNOR U32970 ( .A(n33070), .B(n33074), .Z(n33072) );
  XNOR U32971 ( .A(n32971), .B(n33029), .Z(n33031) );
  XNOR U32972 ( .A(n33075), .B(n33076), .Z(n32971) );
  AND U32973 ( .A(n1139), .B(n32978), .Z(n33076) );
  XOR U32974 ( .A(n33075), .B(n32976), .Z(n32978) );
  AND U32975 ( .A(n32979), .B(n32982), .Z(n33029) );
  XOR U32976 ( .A(n33077), .B(n33057), .Z(n32982) );
  XNOR U32977 ( .A(p_input[1600]), .B(p_input[2048]), .Z(n33057) );
  XNOR U32978 ( .A(n33044), .B(n33043), .Z(n33077) );
  XNOR U32979 ( .A(n33078), .B(n33051), .Z(n33043) );
  XNOR U32980 ( .A(n33039), .B(n33038), .Z(n33051) );
  XNOR U32981 ( .A(n33079), .B(n33035), .Z(n33038) );
  XNOR U32982 ( .A(p_input[1610]), .B(p_input[2058]), .Z(n33035) );
  XOR U32983 ( .A(p_input[1611]), .B(n16732), .Z(n33079) );
  XOR U32984 ( .A(p_input[1612]), .B(p_input[2060]), .Z(n33039) );
  XOR U32985 ( .A(n33049), .B(n33080), .Z(n33078) );
  IV U32986 ( .A(n33040), .Z(n33080) );
  XOR U32987 ( .A(p_input[1601]), .B(p_input[2049]), .Z(n33040) );
  XNOR U32988 ( .A(n33081), .B(n33056), .Z(n33049) );
  XNOR U32989 ( .A(p_input[1615]), .B(n16735), .Z(n33056) );
  XOR U32990 ( .A(n33046), .B(n33055), .Z(n33081) );
  XOR U32991 ( .A(n33082), .B(n33052), .Z(n33055) );
  XOR U32992 ( .A(p_input[1613]), .B(p_input[2061]), .Z(n33052) );
  XOR U32993 ( .A(p_input[1614]), .B(n16737), .Z(n33082) );
  XOR U32994 ( .A(p_input[1609]), .B(p_input[2057]), .Z(n33046) );
  XOR U32995 ( .A(n33064), .B(n33062), .Z(n33044) );
  XNOR U32996 ( .A(n33083), .B(n33069), .Z(n33062) );
  XOR U32997 ( .A(p_input[1608]), .B(p_input[2056]), .Z(n33069) );
  XOR U32998 ( .A(n33059), .B(n33068), .Z(n33083) );
  XOR U32999 ( .A(n33084), .B(n33065), .Z(n33068) );
  XOR U33000 ( .A(p_input[1606]), .B(p_input[2054]), .Z(n33065) );
  XOR U33001 ( .A(p_input[1607]), .B(n17722), .Z(n33084) );
  XOR U33002 ( .A(p_input[1602]), .B(p_input[2050]), .Z(n33059) );
  XNOR U33003 ( .A(n33074), .B(n33073), .Z(n33064) );
  XOR U33004 ( .A(n33085), .B(n33070), .Z(n33073) );
  XOR U33005 ( .A(p_input[1603]), .B(p_input[2051]), .Z(n33070) );
  XOR U33006 ( .A(p_input[1604]), .B(n17724), .Z(n33085) );
  XOR U33007 ( .A(p_input[1605]), .B(p_input[2053]), .Z(n33074) );
  XNOR U33008 ( .A(n33086), .B(n33087), .Z(n32979) );
  AND U33009 ( .A(n1139), .B(n33088), .Z(n33087) );
  XNOR U33010 ( .A(n33089), .B(n33090), .Z(n1139) );
  AND U33011 ( .A(n33091), .B(n33092), .Z(n33090) );
  XOR U33012 ( .A(n33089), .B(n32989), .Z(n33092) );
  XNOR U33013 ( .A(n33089), .B(n32943), .Z(n33091) );
  XOR U33014 ( .A(n33093), .B(n33094), .Z(n33089) );
  AND U33015 ( .A(n33095), .B(n33096), .Z(n33094) );
  XOR U33016 ( .A(n33093), .B(n32953), .Z(n33095) );
  XOR U33017 ( .A(n33097), .B(n33098), .Z(n32932) );
  AND U33018 ( .A(n1143), .B(n33088), .Z(n33098) );
  XNOR U33019 ( .A(n33086), .B(n33097), .Z(n33088) );
  XNOR U33020 ( .A(n33099), .B(n33100), .Z(n1143) );
  AND U33021 ( .A(n33101), .B(n33102), .Z(n33100) );
  XNOR U33022 ( .A(n33103), .B(n33099), .Z(n33102) );
  IV U33023 ( .A(n32989), .Z(n33103) );
  XNOR U33024 ( .A(n33104), .B(n33105), .Z(n32989) );
  AND U33025 ( .A(n1146), .B(n33106), .Z(n33105) );
  XNOR U33026 ( .A(n33104), .B(n33107), .Z(n33106) );
  XNOR U33027 ( .A(n32943), .B(n33099), .Z(n33101) );
  XOR U33028 ( .A(n33108), .B(n33109), .Z(n32943) );
  AND U33029 ( .A(n1154), .B(n33110), .Z(n33109) );
  XOR U33030 ( .A(n33093), .B(n33111), .Z(n33099) );
  AND U33031 ( .A(n33112), .B(n33096), .Z(n33111) );
  XNOR U33032 ( .A(n33002), .B(n33093), .Z(n33096) );
  XNOR U33033 ( .A(n33113), .B(n33114), .Z(n33002) );
  AND U33034 ( .A(n1146), .B(n33115), .Z(n33114) );
  XOR U33035 ( .A(n33116), .B(n33113), .Z(n33115) );
  XNOR U33036 ( .A(n33117), .B(n33093), .Z(n33112) );
  IV U33037 ( .A(n32953), .Z(n33117) );
  XOR U33038 ( .A(n33118), .B(n33119), .Z(n32953) );
  AND U33039 ( .A(n1154), .B(n33120), .Z(n33119) );
  XOR U33040 ( .A(n33121), .B(n33122), .Z(n33093) );
  AND U33041 ( .A(n33123), .B(n33124), .Z(n33122) );
  XNOR U33042 ( .A(n33027), .B(n33121), .Z(n33124) );
  XNOR U33043 ( .A(n33125), .B(n33126), .Z(n33027) );
  AND U33044 ( .A(n1146), .B(n33127), .Z(n33126) );
  XNOR U33045 ( .A(n33128), .B(n33125), .Z(n33127) );
  XOR U33046 ( .A(n33121), .B(n32964), .Z(n33123) );
  XOR U33047 ( .A(n33129), .B(n33130), .Z(n32964) );
  AND U33048 ( .A(n1154), .B(n33131), .Z(n33130) );
  XOR U33049 ( .A(n33132), .B(n33133), .Z(n33121) );
  AND U33050 ( .A(n33134), .B(n33135), .Z(n33133) );
  XNOR U33051 ( .A(n33132), .B(n33075), .Z(n33135) );
  XNOR U33052 ( .A(n33136), .B(n33137), .Z(n33075) );
  AND U33053 ( .A(n1146), .B(n33138), .Z(n33137) );
  XOR U33054 ( .A(n33139), .B(n33136), .Z(n33138) );
  XNOR U33055 ( .A(n33140), .B(n33132), .Z(n33134) );
  IV U33056 ( .A(n32976), .Z(n33140) );
  XOR U33057 ( .A(n33141), .B(n33142), .Z(n32976) );
  AND U33058 ( .A(n1154), .B(n33143), .Z(n33142) );
  AND U33059 ( .A(n33097), .B(n33086), .Z(n33132) );
  XNOR U33060 ( .A(n33144), .B(n33145), .Z(n33086) );
  AND U33061 ( .A(n1146), .B(n33146), .Z(n33145) );
  XNOR U33062 ( .A(n33147), .B(n33144), .Z(n33146) );
  XNOR U33063 ( .A(n33148), .B(n33149), .Z(n1146) );
  AND U33064 ( .A(n33150), .B(n33151), .Z(n33149) );
  XOR U33065 ( .A(n33107), .B(n33148), .Z(n33151) );
  AND U33066 ( .A(n33152), .B(n33153), .Z(n33107) );
  XOR U33067 ( .A(n33148), .B(n33104), .Z(n33150) );
  XNOR U33068 ( .A(n33154), .B(n33155), .Z(n33104) );
  AND U33069 ( .A(n1150), .B(n33110), .Z(n33155) );
  XOR U33070 ( .A(n33108), .B(n33154), .Z(n33110) );
  XOR U33071 ( .A(n33156), .B(n33157), .Z(n33148) );
  AND U33072 ( .A(n33158), .B(n33159), .Z(n33157) );
  XNOR U33073 ( .A(n33156), .B(n33152), .Z(n33159) );
  IV U33074 ( .A(n33116), .Z(n33152) );
  XOR U33075 ( .A(n33160), .B(n33161), .Z(n33116) );
  XOR U33076 ( .A(n33162), .B(n33153), .Z(n33161) );
  AND U33077 ( .A(n33128), .B(n33163), .Z(n33153) );
  AND U33078 ( .A(n33164), .B(n33165), .Z(n33162) );
  XOR U33079 ( .A(n33166), .B(n33160), .Z(n33164) );
  XNOR U33080 ( .A(n33113), .B(n33156), .Z(n33158) );
  XNOR U33081 ( .A(n33167), .B(n33168), .Z(n33113) );
  AND U33082 ( .A(n1150), .B(n33120), .Z(n33168) );
  XOR U33083 ( .A(n33167), .B(n33118), .Z(n33120) );
  XOR U33084 ( .A(n33169), .B(n33170), .Z(n33156) );
  AND U33085 ( .A(n33171), .B(n33172), .Z(n33170) );
  XNOR U33086 ( .A(n33169), .B(n33128), .Z(n33172) );
  XOR U33087 ( .A(n33173), .B(n33165), .Z(n33128) );
  XNOR U33088 ( .A(n33174), .B(n33160), .Z(n33165) );
  XOR U33089 ( .A(n33175), .B(n33176), .Z(n33160) );
  AND U33090 ( .A(n33177), .B(n33178), .Z(n33176) );
  XOR U33091 ( .A(n33179), .B(n33175), .Z(n33177) );
  XNOR U33092 ( .A(n33180), .B(n33181), .Z(n33174) );
  AND U33093 ( .A(n33182), .B(n33183), .Z(n33181) );
  XOR U33094 ( .A(n33180), .B(n33184), .Z(n33182) );
  XNOR U33095 ( .A(n33166), .B(n33163), .Z(n33173) );
  AND U33096 ( .A(n33185), .B(n33186), .Z(n33163) );
  XOR U33097 ( .A(n33187), .B(n33188), .Z(n33166) );
  AND U33098 ( .A(n33189), .B(n33190), .Z(n33188) );
  XOR U33099 ( .A(n33187), .B(n33191), .Z(n33189) );
  XNOR U33100 ( .A(n33125), .B(n33169), .Z(n33171) );
  XNOR U33101 ( .A(n33192), .B(n33193), .Z(n33125) );
  AND U33102 ( .A(n1150), .B(n33131), .Z(n33193) );
  XOR U33103 ( .A(n33192), .B(n33129), .Z(n33131) );
  XOR U33104 ( .A(n33194), .B(n33195), .Z(n33169) );
  AND U33105 ( .A(n33196), .B(n33197), .Z(n33195) );
  XNOR U33106 ( .A(n33194), .B(n33185), .Z(n33197) );
  IV U33107 ( .A(n33139), .Z(n33185) );
  XNOR U33108 ( .A(n33198), .B(n33178), .Z(n33139) );
  XNOR U33109 ( .A(n33199), .B(n33184), .Z(n33178) );
  XNOR U33110 ( .A(n33200), .B(n33201), .Z(n33184) );
  NOR U33111 ( .A(n33202), .B(n33203), .Z(n33201) );
  XOR U33112 ( .A(n33200), .B(n33204), .Z(n33202) );
  XNOR U33113 ( .A(n33183), .B(n33175), .Z(n33199) );
  XOR U33114 ( .A(n33205), .B(n33206), .Z(n33175) );
  AND U33115 ( .A(n33207), .B(n33208), .Z(n33206) );
  XOR U33116 ( .A(n33205), .B(n33209), .Z(n33207) );
  XNOR U33117 ( .A(n33210), .B(n33180), .Z(n33183) );
  XOR U33118 ( .A(n33211), .B(n33212), .Z(n33180) );
  AND U33119 ( .A(n33213), .B(n33214), .Z(n33212) );
  XNOR U33120 ( .A(n33215), .B(n33216), .Z(n33213) );
  IV U33121 ( .A(n33211), .Z(n33215) );
  XNOR U33122 ( .A(n33217), .B(n33218), .Z(n33210) );
  NOR U33123 ( .A(n33219), .B(n33220), .Z(n33218) );
  XNOR U33124 ( .A(n33217), .B(n33221), .Z(n33219) );
  XNOR U33125 ( .A(n33179), .B(n33186), .Z(n33198) );
  NOR U33126 ( .A(n33147), .B(n33222), .Z(n33186) );
  XOR U33127 ( .A(n33191), .B(n33190), .Z(n33179) );
  XNOR U33128 ( .A(n33223), .B(n33187), .Z(n33190) );
  XOR U33129 ( .A(n33224), .B(n33225), .Z(n33187) );
  AND U33130 ( .A(n33226), .B(n33227), .Z(n33225) );
  XNOR U33131 ( .A(n33228), .B(n33229), .Z(n33226) );
  IV U33132 ( .A(n33224), .Z(n33228) );
  XNOR U33133 ( .A(n33230), .B(n33231), .Z(n33223) );
  NOR U33134 ( .A(n33232), .B(n33233), .Z(n33231) );
  XNOR U33135 ( .A(n33230), .B(n33234), .Z(n33232) );
  XOR U33136 ( .A(n33235), .B(n33236), .Z(n33191) );
  NOR U33137 ( .A(n33237), .B(n33238), .Z(n33236) );
  XNOR U33138 ( .A(n33235), .B(n33239), .Z(n33237) );
  XNOR U33139 ( .A(n33136), .B(n33194), .Z(n33196) );
  XNOR U33140 ( .A(n33240), .B(n33241), .Z(n33136) );
  AND U33141 ( .A(n1150), .B(n33143), .Z(n33241) );
  XOR U33142 ( .A(n33240), .B(n33141), .Z(n33143) );
  AND U33143 ( .A(n33144), .B(n33147), .Z(n33194) );
  XOR U33144 ( .A(n33242), .B(n33222), .Z(n33147) );
  XNOR U33145 ( .A(p_input[1616]), .B(p_input[2048]), .Z(n33222) );
  XNOR U33146 ( .A(n33209), .B(n33208), .Z(n33242) );
  XNOR U33147 ( .A(n33243), .B(n33216), .Z(n33208) );
  XNOR U33148 ( .A(n33204), .B(n33203), .Z(n33216) );
  XNOR U33149 ( .A(n33244), .B(n33200), .Z(n33203) );
  XNOR U33150 ( .A(p_input[1626]), .B(p_input[2058]), .Z(n33200) );
  XOR U33151 ( .A(p_input[1627]), .B(n16732), .Z(n33244) );
  XOR U33152 ( .A(p_input[1628]), .B(p_input[2060]), .Z(n33204) );
  XOR U33153 ( .A(n33214), .B(n33245), .Z(n33243) );
  IV U33154 ( .A(n33205), .Z(n33245) );
  XOR U33155 ( .A(p_input[1617]), .B(p_input[2049]), .Z(n33205) );
  XNOR U33156 ( .A(n33246), .B(n33221), .Z(n33214) );
  XNOR U33157 ( .A(p_input[1631]), .B(n16735), .Z(n33221) );
  XOR U33158 ( .A(n33211), .B(n33220), .Z(n33246) );
  XOR U33159 ( .A(n33247), .B(n33217), .Z(n33220) );
  XOR U33160 ( .A(p_input[1629]), .B(p_input[2061]), .Z(n33217) );
  XOR U33161 ( .A(p_input[1630]), .B(n16737), .Z(n33247) );
  XOR U33162 ( .A(p_input[1625]), .B(p_input[2057]), .Z(n33211) );
  XOR U33163 ( .A(n33229), .B(n33227), .Z(n33209) );
  XNOR U33164 ( .A(n33248), .B(n33234), .Z(n33227) );
  XOR U33165 ( .A(p_input[1624]), .B(p_input[2056]), .Z(n33234) );
  XOR U33166 ( .A(n33224), .B(n33233), .Z(n33248) );
  XOR U33167 ( .A(n33249), .B(n33230), .Z(n33233) );
  XOR U33168 ( .A(p_input[1622]), .B(p_input[2054]), .Z(n33230) );
  XOR U33169 ( .A(p_input[1623]), .B(n17722), .Z(n33249) );
  XOR U33170 ( .A(p_input[1618]), .B(p_input[2050]), .Z(n33224) );
  XNOR U33171 ( .A(n33239), .B(n33238), .Z(n33229) );
  XOR U33172 ( .A(n33250), .B(n33235), .Z(n33238) );
  XOR U33173 ( .A(p_input[1619]), .B(p_input[2051]), .Z(n33235) );
  XOR U33174 ( .A(p_input[1620]), .B(n17724), .Z(n33250) );
  XOR U33175 ( .A(p_input[1621]), .B(p_input[2053]), .Z(n33239) );
  XNOR U33176 ( .A(n33251), .B(n33252), .Z(n33144) );
  AND U33177 ( .A(n1150), .B(n33253), .Z(n33252) );
  XNOR U33178 ( .A(n33254), .B(n33255), .Z(n1150) );
  AND U33179 ( .A(n33256), .B(n33257), .Z(n33255) );
  XOR U33180 ( .A(n33254), .B(n33154), .Z(n33257) );
  XNOR U33181 ( .A(n33254), .B(n33108), .Z(n33256) );
  XOR U33182 ( .A(n33258), .B(n33259), .Z(n33254) );
  AND U33183 ( .A(n33260), .B(n33261), .Z(n33259) );
  XOR U33184 ( .A(n33258), .B(n33118), .Z(n33260) );
  XOR U33185 ( .A(n33262), .B(n33263), .Z(n33097) );
  AND U33186 ( .A(n1154), .B(n33253), .Z(n33263) );
  XNOR U33187 ( .A(n33251), .B(n33262), .Z(n33253) );
  XNOR U33188 ( .A(n33264), .B(n33265), .Z(n1154) );
  AND U33189 ( .A(n33266), .B(n33267), .Z(n33265) );
  XNOR U33190 ( .A(n33268), .B(n33264), .Z(n33267) );
  IV U33191 ( .A(n33154), .Z(n33268) );
  XNOR U33192 ( .A(n33269), .B(n33270), .Z(n33154) );
  AND U33193 ( .A(n1157), .B(n33271), .Z(n33270) );
  XNOR U33194 ( .A(n33269), .B(n33272), .Z(n33271) );
  XNOR U33195 ( .A(n33108), .B(n33264), .Z(n33266) );
  XOR U33196 ( .A(n33273), .B(n33274), .Z(n33108) );
  AND U33197 ( .A(n1165), .B(n33275), .Z(n33274) );
  XOR U33198 ( .A(n33258), .B(n33276), .Z(n33264) );
  AND U33199 ( .A(n33277), .B(n33261), .Z(n33276) );
  XNOR U33200 ( .A(n33167), .B(n33258), .Z(n33261) );
  XNOR U33201 ( .A(n33278), .B(n33279), .Z(n33167) );
  AND U33202 ( .A(n1157), .B(n33280), .Z(n33279) );
  XOR U33203 ( .A(n33281), .B(n33278), .Z(n33280) );
  XNOR U33204 ( .A(n33282), .B(n33258), .Z(n33277) );
  IV U33205 ( .A(n33118), .Z(n33282) );
  XOR U33206 ( .A(n33283), .B(n33284), .Z(n33118) );
  AND U33207 ( .A(n1165), .B(n33285), .Z(n33284) );
  XOR U33208 ( .A(n33286), .B(n33287), .Z(n33258) );
  AND U33209 ( .A(n33288), .B(n33289), .Z(n33287) );
  XNOR U33210 ( .A(n33192), .B(n33286), .Z(n33289) );
  XNOR U33211 ( .A(n33290), .B(n33291), .Z(n33192) );
  AND U33212 ( .A(n1157), .B(n33292), .Z(n33291) );
  XNOR U33213 ( .A(n33293), .B(n33290), .Z(n33292) );
  XOR U33214 ( .A(n33286), .B(n33129), .Z(n33288) );
  XOR U33215 ( .A(n33294), .B(n33295), .Z(n33129) );
  AND U33216 ( .A(n1165), .B(n33296), .Z(n33295) );
  XOR U33217 ( .A(n33297), .B(n33298), .Z(n33286) );
  AND U33218 ( .A(n33299), .B(n33300), .Z(n33298) );
  XNOR U33219 ( .A(n33297), .B(n33240), .Z(n33300) );
  XNOR U33220 ( .A(n33301), .B(n33302), .Z(n33240) );
  AND U33221 ( .A(n1157), .B(n33303), .Z(n33302) );
  XOR U33222 ( .A(n33304), .B(n33301), .Z(n33303) );
  XNOR U33223 ( .A(n33305), .B(n33297), .Z(n33299) );
  IV U33224 ( .A(n33141), .Z(n33305) );
  XOR U33225 ( .A(n33306), .B(n33307), .Z(n33141) );
  AND U33226 ( .A(n1165), .B(n33308), .Z(n33307) );
  AND U33227 ( .A(n33262), .B(n33251), .Z(n33297) );
  XNOR U33228 ( .A(n33309), .B(n33310), .Z(n33251) );
  AND U33229 ( .A(n1157), .B(n33311), .Z(n33310) );
  XNOR U33230 ( .A(n33312), .B(n33309), .Z(n33311) );
  XNOR U33231 ( .A(n33313), .B(n33314), .Z(n1157) );
  AND U33232 ( .A(n33315), .B(n33316), .Z(n33314) );
  XOR U33233 ( .A(n33272), .B(n33313), .Z(n33316) );
  AND U33234 ( .A(n33317), .B(n33318), .Z(n33272) );
  XOR U33235 ( .A(n33313), .B(n33269), .Z(n33315) );
  XNOR U33236 ( .A(n33319), .B(n33320), .Z(n33269) );
  AND U33237 ( .A(n1161), .B(n33275), .Z(n33320) );
  XOR U33238 ( .A(n33273), .B(n33319), .Z(n33275) );
  XOR U33239 ( .A(n33321), .B(n33322), .Z(n33313) );
  AND U33240 ( .A(n33323), .B(n33324), .Z(n33322) );
  XNOR U33241 ( .A(n33321), .B(n33317), .Z(n33324) );
  IV U33242 ( .A(n33281), .Z(n33317) );
  XOR U33243 ( .A(n33325), .B(n33326), .Z(n33281) );
  XOR U33244 ( .A(n33327), .B(n33318), .Z(n33326) );
  AND U33245 ( .A(n33293), .B(n33328), .Z(n33318) );
  AND U33246 ( .A(n33329), .B(n33330), .Z(n33327) );
  XOR U33247 ( .A(n33331), .B(n33325), .Z(n33329) );
  XNOR U33248 ( .A(n33278), .B(n33321), .Z(n33323) );
  XNOR U33249 ( .A(n33332), .B(n33333), .Z(n33278) );
  AND U33250 ( .A(n1161), .B(n33285), .Z(n33333) );
  XOR U33251 ( .A(n33332), .B(n33283), .Z(n33285) );
  XOR U33252 ( .A(n33334), .B(n33335), .Z(n33321) );
  AND U33253 ( .A(n33336), .B(n33337), .Z(n33335) );
  XNOR U33254 ( .A(n33334), .B(n33293), .Z(n33337) );
  XOR U33255 ( .A(n33338), .B(n33330), .Z(n33293) );
  XNOR U33256 ( .A(n33339), .B(n33325), .Z(n33330) );
  XOR U33257 ( .A(n33340), .B(n33341), .Z(n33325) );
  AND U33258 ( .A(n33342), .B(n33343), .Z(n33341) );
  XOR U33259 ( .A(n33344), .B(n33340), .Z(n33342) );
  XNOR U33260 ( .A(n33345), .B(n33346), .Z(n33339) );
  AND U33261 ( .A(n33347), .B(n33348), .Z(n33346) );
  XOR U33262 ( .A(n33345), .B(n33349), .Z(n33347) );
  XNOR U33263 ( .A(n33331), .B(n33328), .Z(n33338) );
  AND U33264 ( .A(n33350), .B(n33351), .Z(n33328) );
  XOR U33265 ( .A(n33352), .B(n33353), .Z(n33331) );
  AND U33266 ( .A(n33354), .B(n33355), .Z(n33353) );
  XOR U33267 ( .A(n33352), .B(n33356), .Z(n33354) );
  XNOR U33268 ( .A(n33290), .B(n33334), .Z(n33336) );
  XNOR U33269 ( .A(n33357), .B(n33358), .Z(n33290) );
  AND U33270 ( .A(n1161), .B(n33296), .Z(n33358) );
  XOR U33271 ( .A(n33357), .B(n33294), .Z(n33296) );
  XOR U33272 ( .A(n33359), .B(n33360), .Z(n33334) );
  AND U33273 ( .A(n33361), .B(n33362), .Z(n33360) );
  XNOR U33274 ( .A(n33359), .B(n33350), .Z(n33362) );
  IV U33275 ( .A(n33304), .Z(n33350) );
  XNOR U33276 ( .A(n33363), .B(n33343), .Z(n33304) );
  XNOR U33277 ( .A(n33364), .B(n33349), .Z(n33343) );
  XNOR U33278 ( .A(n33365), .B(n33366), .Z(n33349) );
  NOR U33279 ( .A(n33367), .B(n33368), .Z(n33366) );
  XOR U33280 ( .A(n33365), .B(n33369), .Z(n33367) );
  XNOR U33281 ( .A(n33348), .B(n33340), .Z(n33364) );
  XOR U33282 ( .A(n33370), .B(n33371), .Z(n33340) );
  AND U33283 ( .A(n33372), .B(n33373), .Z(n33371) );
  XOR U33284 ( .A(n33370), .B(n33374), .Z(n33372) );
  XNOR U33285 ( .A(n33375), .B(n33345), .Z(n33348) );
  XOR U33286 ( .A(n33376), .B(n33377), .Z(n33345) );
  AND U33287 ( .A(n33378), .B(n33379), .Z(n33377) );
  XNOR U33288 ( .A(n33380), .B(n33381), .Z(n33378) );
  IV U33289 ( .A(n33376), .Z(n33380) );
  XNOR U33290 ( .A(n33382), .B(n33383), .Z(n33375) );
  NOR U33291 ( .A(n33384), .B(n33385), .Z(n33383) );
  XNOR U33292 ( .A(n33382), .B(n33386), .Z(n33384) );
  XNOR U33293 ( .A(n33344), .B(n33351), .Z(n33363) );
  NOR U33294 ( .A(n33312), .B(n33387), .Z(n33351) );
  XOR U33295 ( .A(n33356), .B(n33355), .Z(n33344) );
  XNOR U33296 ( .A(n33388), .B(n33352), .Z(n33355) );
  XOR U33297 ( .A(n33389), .B(n33390), .Z(n33352) );
  AND U33298 ( .A(n33391), .B(n33392), .Z(n33390) );
  XNOR U33299 ( .A(n33393), .B(n33394), .Z(n33391) );
  IV U33300 ( .A(n33389), .Z(n33393) );
  XNOR U33301 ( .A(n33395), .B(n33396), .Z(n33388) );
  NOR U33302 ( .A(n33397), .B(n33398), .Z(n33396) );
  XNOR U33303 ( .A(n33395), .B(n33399), .Z(n33397) );
  XOR U33304 ( .A(n33400), .B(n33401), .Z(n33356) );
  NOR U33305 ( .A(n33402), .B(n33403), .Z(n33401) );
  XNOR U33306 ( .A(n33400), .B(n33404), .Z(n33402) );
  XNOR U33307 ( .A(n33301), .B(n33359), .Z(n33361) );
  XNOR U33308 ( .A(n33405), .B(n33406), .Z(n33301) );
  AND U33309 ( .A(n1161), .B(n33308), .Z(n33406) );
  XOR U33310 ( .A(n33405), .B(n33306), .Z(n33308) );
  AND U33311 ( .A(n33309), .B(n33312), .Z(n33359) );
  XOR U33312 ( .A(n33407), .B(n33387), .Z(n33312) );
  XNOR U33313 ( .A(p_input[1632]), .B(p_input[2048]), .Z(n33387) );
  XNOR U33314 ( .A(n33374), .B(n33373), .Z(n33407) );
  XNOR U33315 ( .A(n33408), .B(n33381), .Z(n33373) );
  XNOR U33316 ( .A(n33369), .B(n33368), .Z(n33381) );
  XNOR U33317 ( .A(n33409), .B(n33365), .Z(n33368) );
  XNOR U33318 ( .A(p_input[1642]), .B(p_input[2058]), .Z(n33365) );
  XOR U33319 ( .A(p_input[1643]), .B(n16732), .Z(n33409) );
  XOR U33320 ( .A(p_input[1644]), .B(p_input[2060]), .Z(n33369) );
  XOR U33321 ( .A(n33379), .B(n33410), .Z(n33408) );
  IV U33322 ( .A(n33370), .Z(n33410) );
  XOR U33323 ( .A(p_input[1633]), .B(p_input[2049]), .Z(n33370) );
  XNOR U33324 ( .A(n33411), .B(n33386), .Z(n33379) );
  XNOR U33325 ( .A(p_input[1647]), .B(n16735), .Z(n33386) );
  XOR U33326 ( .A(n33376), .B(n33385), .Z(n33411) );
  XOR U33327 ( .A(n33412), .B(n33382), .Z(n33385) );
  XOR U33328 ( .A(p_input[1645]), .B(p_input[2061]), .Z(n33382) );
  XOR U33329 ( .A(p_input[1646]), .B(n16737), .Z(n33412) );
  XOR U33330 ( .A(p_input[1641]), .B(p_input[2057]), .Z(n33376) );
  XOR U33331 ( .A(n33394), .B(n33392), .Z(n33374) );
  XNOR U33332 ( .A(n33413), .B(n33399), .Z(n33392) );
  XOR U33333 ( .A(p_input[1640]), .B(p_input[2056]), .Z(n33399) );
  XOR U33334 ( .A(n33389), .B(n33398), .Z(n33413) );
  XOR U33335 ( .A(n33414), .B(n33395), .Z(n33398) );
  XOR U33336 ( .A(p_input[1638]), .B(p_input[2054]), .Z(n33395) );
  XOR U33337 ( .A(p_input[1639]), .B(n17722), .Z(n33414) );
  XOR U33338 ( .A(p_input[1634]), .B(p_input[2050]), .Z(n33389) );
  XNOR U33339 ( .A(n33404), .B(n33403), .Z(n33394) );
  XOR U33340 ( .A(n33415), .B(n33400), .Z(n33403) );
  XOR U33341 ( .A(p_input[1635]), .B(p_input[2051]), .Z(n33400) );
  XOR U33342 ( .A(p_input[1636]), .B(n17724), .Z(n33415) );
  XOR U33343 ( .A(p_input[1637]), .B(p_input[2053]), .Z(n33404) );
  XNOR U33344 ( .A(n33416), .B(n33417), .Z(n33309) );
  AND U33345 ( .A(n1161), .B(n33418), .Z(n33417) );
  XNOR U33346 ( .A(n33419), .B(n33420), .Z(n1161) );
  AND U33347 ( .A(n33421), .B(n33422), .Z(n33420) );
  XOR U33348 ( .A(n33419), .B(n33319), .Z(n33422) );
  XNOR U33349 ( .A(n33419), .B(n33273), .Z(n33421) );
  XOR U33350 ( .A(n33423), .B(n33424), .Z(n33419) );
  AND U33351 ( .A(n33425), .B(n33426), .Z(n33424) );
  XOR U33352 ( .A(n33423), .B(n33283), .Z(n33425) );
  XOR U33353 ( .A(n33427), .B(n33428), .Z(n33262) );
  AND U33354 ( .A(n1165), .B(n33418), .Z(n33428) );
  XNOR U33355 ( .A(n33416), .B(n33427), .Z(n33418) );
  XNOR U33356 ( .A(n33429), .B(n33430), .Z(n1165) );
  AND U33357 ( .A(n33431), .B(n33432), .Z(n33430) );
  XNOR U33358 ( .A(n33433), .B(n33429), .Z(n33432) );
  IV U33359 ( .A(n33319), .Z(n33433) );
  XNOR U33360 ( .A(n33434), .B(n33435), .Z(n33319) );
  AND U33361 ( .A(n1168), .B(n33436), .Z(n33435) );
  XNOR U33362 ( .A(n33434), .B(n33437), .Z(n33436) );
  XNOR U33363 ( .A(n33273), .B(n33429), .Z(n33431) );
  XOR U33364 ( .A(n33438), .B(n33439), .Z(n33273) );
  AND U33365 ( .A(n1176), .B(n33440), .Z(n33439) );
  XOR U33366 ( .A(n33423), .B(n33441), .Z(n33429) );
  AND U33367 ( .A(n33442), .B(n33426), .Z(n33441) );
  XNOR U33368 ( .A(n33332), .B(n33423), .Z(n33426) );
  XNOR U33369 ( .A(n33443), .B(n33444), .Z(n33332) );
  AND U33370 ( .A(n1168), .B(n33445), .Z(n33444) );
  XOR U33371 ( .A(n33446), .B(n33443), .Z(n33445) );
  XNOR U33372 ( .A(n33447), .B(n33423), .Z(n33442) );
  IV U33373 ( .A(n33283), .Z(n33447) );
  XOR U33374 ( .A(n33448), .B(n33449), .Z(n33283) );
  AND U33375 ( .A(n1176), .B(n33450), .Z(n33449) );
  XOR U33376 ( .A(n33451), .B(n33452), .Z(n33423) );
  AND U33377 ( .A(n33453), .B(n33454), .Z(n33452) );
  XNOR U33378 ( .A(n33357), .B(n33451), .Z(n33454) );
  XNOR U33379 ( .A(n33455), .B(n33456), .Z(n33357) );
  AND U33380 ( .A(n1168), .B(n33457), .Z(n33456) );
  XNOR U33381 ( .A(n33458), .B(n33455), .Z(n33457) );
  XOR U33382 ( .A(n33451), .B(n33294), .Z(n33453) );
  XOR U33383 ( .A(n33459), .B(n33460), .Z(n33294) );
  AND U33384 ( .A(n1176), .B(n33461), .Z(n33460) );
  XOR U33385 ( .A(n33462), .B(n33463), .Z(n33451) );
  AND U33386 ( .A(n33464), .B(n33465), .Z(n33463) );
  XNOR U33387 ( .A(n33462), .B(n33405), .Z(n33465) );
  XNOR U33388 ( .A(n33466), .B(n33467), .Z(n33405) );
  AND U33389 ( .A(n1168), .B(n33468), .Z(n33467) );
  XOR U33390 ( .A(n33469), .B(n33466), .Z(n33468) );
  XNOR U33391 ( .A(n33470), .B(n33462), .Z(n33464) );
  IV U33392 ( .A(n33306), .Z(n33470) );
  XOR U33393 ( .A(n33471), .B(n33472), .Z(n33306) );
  AND U33394 ( .A(n1176), .B(n33473), .Z(n33472) );
  AND U33395 ( .A(n33427), .B(n33416), .Z(n33462) );
  XNOR U33396 ( .A(n33474), .B(n33475), .Z(n33416) );
  AND U33397 ( .A(n1168), .B(n33476), .Z(n33475) );
  XNOR U33398 ( .A(n33477), .B(n33474), .Z(n33476) );
  XNOR U33399 ( .A(n33478), .B(n33479), .Z(n1168) );
  AND U33400 ( .A(n33480), .B(n33481), .Z(n33479) );
  XOR U33401 ( .A(n33437), .B(n33478), .Z(n33481) );
  AND U33402 ( .A(n33482), .B(n33483), .Z(n33437) );
  XOR U33403 ( .A(n33478), .B(n33434), .Z(n33480) );
  XNOR U33404 ( .A(n33484), .B(n33485), .Z(n33434) );
  AND U33405 ( .A(n1172), .B(n33440), .Z(n33485) );
  XOR U33406 ( .A(n33438), .B(n33484), .Z(n33440) );
  XOR U33407 ( .A(n33486), .B(n33487), .Z(n33478) );
  AND U33408 ( .A(n33488), .B(n33489), .Z(n33487) );
  XNOR U33409 ( .A(n33486), .B(n33482), .Z(n33489) );
  IV U33410 ( .A(n33446), .Z(n33482) );
  XOR U33411 ( .A(n33490), .B(n33491), .Z(n33446) );
  XOR U33412 ( .A(n33492), .B(n33483), .Z(n33491) );
  AND U33413 ( .A(n33458), .B(n33493), .Z(n33483) );
  AND U33414 ( .A(n33494), .B(n33495), .Z(n33492) );
  XOR U33415 ( .A(n33496), .B(n33490), .Z(n33494) );
  XNOR U33416 ( .A(n33443), .B(n33486), .Z(n33488) );
  XNOR U33417 ( .A(n33497), .B(n33498), .Z(n33443) );
  AND U33418 ( .A(n1172), .B(n33450), .Z(n33498) );
  XOR U33419 ( .A(n33497), .B(n33448), .Z(n33450) );
  XOR U33420 ( .A(n33499), .B(n33500), .Z(n33486) );
  AND U33421 ( .A(n33501), .B(n33502), .Z(n33500) );
  XNOR U33422 ( .A(n33499), .B(n33458), .Z(n33502) );
  XOR U33423 ( .A(n33503), .B(n33495), .Z(n33458) );
  XNOR U33424 ( .A(n33504), .B(n33490), .Z(n33495) );
  XOR U33425 ( .A(n33505), .B(n33506), .Z(n33490) );
  AND U33426 ( .A(n33507), .B(n33508), .Z(n33506) );
  XOR U33427 ( .A(n33509), .B(n33505), .Z(n33507) );
  XNOR U33428 ( .A(n33510), .B(n33511), .Z(n33504) );
  AND U33429 ( .A(n33512), .B(n33513), .Z(n33511) );
  XOR U33430 ( .A(n33510), .B(n33514), .Z(n33512) );
  XNOR U33431 ( .A(n33496), .B(n33493), .Z(n33503) );
  AND U33432 ( .A(n33515), .B(n33516), .Z(n33493) );
  XOR U33433 ( .A(n33517), .B(n33518), .Z(n33496) );
  AND U33434 ( .A(n33519), .B(n33520), .Z(n33518) );
  XOR U33435 ( .A(n33517), .B(n33521), .Z(n33519) );
  XNOR U33436 ( .A(n33455), .B(n33499), .Z(n33501) );
  XNOR U33437 ( .A(n33522), .B(n33523), .Z(n33455) );
  AND U33438 ( .A(n1172), .B(n33461), .Z(n33523) );
  XOR U33439 ( .A(n33522), .B(n33459), .Z(n33461) );
  XOR U33440 ( .A(n33524), .B(n33525), .Z(n33499) );
  AND U33441 ( .A(n33526), .B(n33527), .Z(n33525) );
  XNOR U33442 ( .A(n33524), .B(n33515), .Z(n33527) );
  IV U33443 ( .A(n33469), .Z(n33515) );
  XNOR U33444 ( .A(n33528), .B(n33508), .Z(n33469) );
  XNOR U33445 ( .A(n33529), .B(n33514), .Z(n33508) );
  XNOR U33446 ( .A(n33530), .B(n33531), .Z(n33514) );
  NOR U33447 ( .A(n33532), .B(n33533), .Z(n33531) );
  XOR U33448 ( .A(n33530), .B(n33534), .Z(n33532) );
  XNOR U33449 ( .A(n33513), .B(n33505), .Z(n33529) );
  XOR U33450 ( .A(n33535), .B(n33536), .Z(n33505) );
  AND U33451 ( .A(n33537), .B(n33538), .Z(n33536) );
  XOR U33452 ( .A(n33535), .B(n33539), .Z(n33537) );
  XNOR U33453 ( .A(n33540), .B(n33510), .Z(n33513) );
  XOR U33454 ( .A(n33541), .B(n33542), .Z(n33510) );
  AND U33455 ( .A(n33543), .B(n33544), .Z(n33542) );
  XNOR U33456 ( .A(n33545), .B(n33546), .Z(n33543) );
  IV U33457 ( .A(n33541), .Z(n33545) );
  XNOR U33458 ( .A(n33547), .B(n33548), .Z(n33540) );
  NOR U33459 ( .A(n33549), .B(n33550), .Z(n33548) );
  XNOR U33460 ( .A(n33547), .B(n33551), .Z(n33549) );
  XNOR U33461 ( .A(n33509), .B(n33516), .Z(n33528) );
  NOR U33462 ( .A(n33477), .B(n33552), .Z(n33516) );
  XOR U33463 ( .A(n33521), .B(n33520), .Z(n33509) );
  XNOR U33464 ( .A(n33553), .B(n33517), .Z(n33520) );
  XOR U33465 ( .A(n33554), .B(n33555), .Z(n33517) );
  AND U33466 ( .A(n33556), .B(n33557), .Z(n33555) );
  XNOR U33467 ( .A(n33558), .B(n33559), .Z(n33556) );
  IV U33468 ( .A(n33554), .Z(n33558) );
  XNOR U33469 ( .A(n33560), .B(n33561), .Z(n33553) );
  NOR U33470 ( .A(n33562), .B(n33563), .Z(n33561) );
  XNOR U33471 ( .A(n33560), .B(n33564), .Z(n33562) );
  XOR U33472 ( .A(n33565), .B(n33566), .Z(n33521) );
  NOR U33473 ( .A(n33567), .B(n33568), .Z(n33566) );
  XNOR U33474 ( .A(n33565), .B(n33569), .Z(n33567) );
  XNOR U33475 ( .A(n33466), .B(n33524), .Z(n33526) );
  XNOR U33476 ( .A(n33570), .B(n33571), .Z(n33466) );
  AND U33477 ( .A(n1172), .B(n33473), .Z(n33571) );
  XOR U33478 ( .A(n33570), .B(n33471), .Z(n33473) );
  AND U33479 ( .A(n33474), .B(n33477), .Z(n33524) );
  XOR U33480 ( .A(n33572), .B(n33552), .Z(n33477) );
  XNOR U33481 ( .A(p_input[1648]), .B(p_input[2048]), .Z(n33552) );
  XNOR U33482 ( .A(n33539), .B(n33538), .Z(n33572) );
  XNOR U33483 ( .A(n33573), .B(n33546), .Z(n33538) );
  XNOR U33484 ( .A(n33534), .B(n33533), .Z(n33546) );
  XNOR U33485 ( .A(n33574), .B(n33530), .Z(n33533) );
  XNOR U33486 ( .A(p_input[1658]), .B(p_input[2058]), .Z(n33530) );
  XOR U33487 ( .A(p_input[1659]), .B(n16732), .Z(n33574) );
  XOR U33488 ( .A(p_input[1660]), .B(p_input[2060]), .Z(n33534) );
  XOR U33489 ( .A(n33544), .B(n33575), .Z(n33573) );
  IV U33490 ( .A(n33535), .Z(n33575) );
  XOR U33491 ( .A(p_input[1649]), .B(p_input[2049]), .Z(n33535) );
  XNOR U33492 ( .A(n33576), .B(n33551), .Z(n33544) );
  XNOR U33493 ( .A(p_input[1663]), .B(n16735), .Z(n33551) );
  XOR U33494 ( .A(n33541), .B(n33550), .Z(n33576) );
  XOR U33495 ( .A(n33577), .B(n33547), .Z(n33550) );
  XOR U33496 ( .A(p_input[1661]), .B(p_input[2061]), .Z(n33547) );
  XOR U33497 ( .A(p_input[1662]), .B(n16737), .Z(n33577) );
  XOR U33498 ( .A(p_input[1657]), .B(p_input[2057]), .Z(n33541) );
  XOR U33499 ( .A(n33559), .B(n33557), .Z(n33539) );
  XNOR U33500 ( .A(n33578), .B(n33564), .Z(n33557) );
  XOR U33501 ( .A(p_input[1656]), .B(p_input[2056]), .Z(n33564) );
  XOR U33502 ( .A(n33554), .B(n33563), .Z(n33578) );
  XOR U33503 ( .A(n33579), .B(n33560), .Z(n33563) );
  XOR U33504 ( .A(p_input[1654]), .B(p_input[2054]), .Z(n33560) );
  XOR U33505 ( .A(p_input[1655]), .B(n17722), .Z(n33579) );
  XOR U33506 ( .A(p_input[1650]), .B(p_input[2050]), .Z(n33554) );
  XNOR U33507 ( .A(n33569), .B(n33568), .Z(n33559) );
  XOR U33508 ( .A(n33580), .B(n33565), .Z(n33568) );
  XOR U33509 ( .A(p_input[1651]), .B(p_input[2051]), .Z(n33565) );
  XOR U33510 ( .A(p_input[1652]), .B(n17724), .Z(n33580) );
  XOR U33511 ( .A(p_input[1653]), .B(p_input[2053]), .Z(n33569) );
  XNOR U33512 ( .A(n33581), .B(n33582), .Z(n33474) );
  AND U33513 ( .A(n1172), .B(n33583), .Z(n33582) );
  XNOR U33514 ( .A(n33584), .B(n33585), .Z(n1172) );
  AND U33515 ( .A(n33586), .B(n33587), .Z(n33585) );
  XOR U33516 ( .A(n33584), .B(n33484), .Z(n33587) );
  XNOR U33517 ( .A(n33584), .B(n33438), .Z(n33586) );
  XOR U33518 ( .A(n33588), .B(n33589), .Z(n33584) );
  AND U33519 ( .A(n33590), .B(n33591), .Z(n33589) );
  XOR U33520 ( .A(n33588), .B(n33448), .Z(n33590) );
  XOR U33521 ( .A(n33592), .B(n33593), .Z(n33427) );
  AND U33522 ( .A(n1176), .B(n33583), .Z(n33593) );
  XNOR U33523 ( .A(n33581), .B(n33592), .Z(n33583) );
  XNOR U33524 ( .A(n33594), .B(n33595), .Z(n1176) );
  AND U33525 ( .A(n33596), .B(n33597), .Z(n33595) );
  XNOR U33526 ( .A(n33598), .B(n33594), .Z(n33597) );
  IV U33527 ( .A(n33484), .Z(n33598) );
  XNOR U33528 ( .A(n33599), .B(n33600), .Z(n33484) );
  AND U33529 ( .A(n1179), .B(n33601), .Z(n33600) );
  XNOR U33530 ( .A(n33599), .B(n33602), .Z(n33601) );
  XNOR U33531 ( .A(n33438), .B(n33594), .Z(n33596) );
  XOR U33532 ( .A(n33603), .B(n33604), .Z(n33438) );
  AND U33533 ( .A(n1187), .B(n33605), .Z(n33604) );
  XOR U33534 ( .A(n33588), .B(n33606), .Z(n33594) );
  AND U33535 ( .A(n33607), .B(n33591), .Z(n33606) );
  XNOR U33536 ( .A(n33497), .B(n33588), .Z(n33591) );
  XNOR U33537 ( .A(n33608), .B(n33609), .Z(n33497) );
  AND U33538 ( .A(n1179), .B(n33610), .Z(n33609) );
  XOR U33539 ( .A(n33611), .B(n33608), .Z(n33610) );
  XNOR U33540 ( .A(n33612), .B(n33588), .Z(n33607) );
  IV U33541 ( .A(n33448), .Z(n33612) );
  XOR U33542 ( .A(n33613), .B(n33614), .Z(n33448) );
  AND U33543 ( .A(n1187), .B(n33615), .Z(n33614) );
  XOR U33544 ( .A(n33616), .B(n33617), .Z(n33588) );
  AND U33545 ( .A(n33618), .B(n33619), .Z(n33617) );
  XNOR U33546 ( .A(n33522), .B(n33616), .Z(n33619) );
  XNOR U33547 ( .A(n33620), .B(n33621), .Z(n33522) );
  AND U33548 ( .A(n1179), .B(n33622), .Z(n33621) );
  XNOR U33549 ( .A(n33623), .B(n33620), .Z(n33622) );
  XOR U33550 ( .A(n33616), .B(n33459), .Z(n33618) );
  XOR U33551 ( .A(n33624), .B(n33625), .Z(n33459) );
  AND U33552 ( .A(n1187), .B(n33626), .Z(n33625) );
  XOR U33553 ( .A(n33627), .B(n33628), .Z(n33616) );
  AND U33554 ( .A(n33629), .B(n33630), .Z(n33628) );
  XNOR U33555 ( .A(n33627), .B(n33570), .Z(n33630) );
  XNOR U33556 ( .A(n33631), .B(n33632), .Z(n33570) );
  AND U33557 ( .A(n1179), .B(n33633), .Z(n33632) );
  XOR U33558 ( .A(n33634), .B(n33631), .Z(n33633) );
  XNOR U33559 ( .A(n33635), .B(n33627), .Z(n33629) );
  IV U33560 ( .A(n33471), .Z(n33635) );
  XOR U33561 ( .A(n33636), .B(n33637), .Z(n33471) );
  AND U33562 ( .A(n1187), .B(n33638), .Z(n33637) );
  AND U33563 ( .A(n33592), .B(n33581), .Z(n33627) );
  XNOR U33564 ( .A(n33639), .B(n33640), .Z(n33581) );
  AND U33565 ( .A(n1179), .B(n33641), .Z(n33640) );
  XNOR U33566 ( .A(n33642), .B(n33639), .Z(n33641) );
  XNOR U33567 ( .A(n33643), .B(n33644), .Z(n1179) );
  AND U33568 ( .A(n33645), .B(n33646), .Z(n33644) );
  XOR U33569 ( .A(n33602), .B(n33643), .Z(n33646) );
  AND U33570 ( .A(n33647), .B(n33648), .Z(n33602) );
  XOR U33571 ( .A(n33643), .B(n33599), .Z(n33645) );
  XNOR U33572 ( .A(n33649), .B(n33650), .Z(n33599) );
  AND U33573 ( .A(n1183), .B(n33605), .Z(n33650) );
  XOR U33574 ( .A(n33603), .B(n33649), .Z(n33605) );
  XOR U33575 ( .A(n33651), .B(n33652), .Z(n33643) );
  AND U33576 ( .A(n33653), .B(n33654), .Z(n33652) );
  XNOR U33577 ( .A(n33651), .B(n33647), .Z(n33654) );
  IV U33578 ( .A(n33611), .Z(n33647) );
  XOR U33579 ( .A(n33655), .B(n33656), .Z(n33611) );
  XOR U33580 ( .A(n33657), .B(n33648), .Z(n33656) );
  AND U33581 ( .A(n33623), .B(n33658), .Z(n33648) );
  AND U33582 ( .A(n33659), .B(n33660), .Z(n33657) );
  XOR U33583 ( .A(n33661), .B(n33655), .Z(n33659) );
  XNOR U33584 ( .A(n33608), .B(n33651), .Z(n33653) );
  XNOR U33585 ( .A(n33662), .B(n33663), .Z(n33608) );
  AND U33586 ( .A(n1183), .B(n33615), .Z(n33663) );
  XOR U33587 ( .A(n33662), .B(n33613), .Z(n33615) );
  XOR U33588 ( .A(n33664), .B(n33665), .Z(n33651) );
  AND U33589 ( .A(n33666), .B(n33667), .Z(n33665) );
  XNOR U33590 ( .A(n33664), .B(n33623), .Z(n33667) );
  XOR U33591 ( .A(n33668), .B(n33660), .Z(n33623) );
  XNOR U33592 ( .A(n33669), .B(n33655), .Z(n33660) );
  XOR U33593 ( .A(n33670), .B(n33671), .Z(n33655) );
  AND U33594 ( .A(n33672), .B(n33673), .Z(n33671) );
  XOR U33595 ( .A(n33674), .B(n33670), .Z(n33672) );
  XNOR U33596 ( .A(n33675), .B(n33676), .Z(n33669) );
  AND U33597 ( .A(n33677), .B(n33678), .Z(n33676) );
  XOR U33598 ( .A(n33675), .B(n33679), .Z(n33677) );
  XNOR U33599 ( .A(n33661), .B(n33658), .Z(n33668) );
  AND U33600 ( .A(n33680), .B(n33681), .Z(n33658) );
  XOR U33601 ( .A(n33682), .B(n33683), .Z(n33661) );
  AND U33602 ( .A(n33684), .B(n33685), .Z(n33683) );
  XOR U33603 ( .A(n33682), .B(n33686), .Z(n33684) );
  XNOR U33604 ( .A(n33620), .B(n33664), .Z(n33666) );
  XNOR U33605 ( .A(n33687), .B(n33688), .Z(n33620) );
  AND U33606 ( .A(n1183), .B(n33626), .Z(n33688) );
  XOR U33607 ( .A(n33687), .B(n33624), .Z(n33626) );
  XOR U33608 ( .A(n33689), .B(n33690), .Z(n33664) );
  AND U33609 ( .A(n33691), .B(n33692), .Z(n33690) );
  XNOR U33610 ( .A(n33689), .B(n33680), .Z(n33692) );
  IV U33611 ( .A(n33634), .Z(n33680) );
  XNOR U33612 ( .A(n33693), .B(n33673), .Z(n33634) );
  XNOR U33613 ( .A(n33694), .B(n33679), .Z(n33673) );
  XNOR U33614 ( .A(n33695), .B(n33696), .Z(n33679) );
  NOR U33615 ( .A(n33697), .B(n33698), .Z(n33696) );
  XOR U33616 ( .A(n33695), .B(n33699), .Z(n33697) );
  XNOR U33617 ( .A(n33678), .B(n33670), .Z(n33694) );
  XOR U33618 ( .A(n33700), .B(n33701), .Z(n33670) );
  AND U33619 ( .A(n33702), .B(n33703), .Z(n33701) );
  XOR U33620 ( .A(n33700), .B(n33704), .Z(n33702) );
  XNOR U33621 ( .A(n33705), .B(n33675), .Z(n33678) );
  XOR U33622 ( .A(n33706), .B(n33707), .Z(n33675) );
  AND U33623 ( .A(n33708), .B(n33709), .Z(n33707) );
  XNOR U33624 ( .A(n33710), .B(n33711), .Z(n33708) );
  IV U33625 ( .A(n33706), .Z(n33710) );
  XNOR U33626 ( .A(n33712), .B(n33713), .Z(n33705) );
  NOR U33627 ( .A(n33714), .B(n33715), .Z(n33713) );
  XNOR U33628 ( .A(n33712), .B(n33716), .Z(n33714) );
  XNOR U33629 ( .A(n33674), .B(n33681), .Z(n33693) );
  NOR U33630 ( .A(n33642), .B(n33717), .Z(n33681) );
  XOR U33631 ( .A(n33686), .B(n33685), .Z(n33674) );
  XNOR U33632 ( .A(n33718), .B(n33682), .Z(n33685) );
  XOR U33633 ( .A(n33719), .B(n33720), .Z(n33682) );
  AND U33634 ( .A(n33721), .B(n33722), .Z(n33720) );
  XNOR U33635 ( .A(n33723), .B(n33724), .Z(n33721) );
  IV U33636 ( .A(n33719), .Z(n33723) );
  XNOR U33637 ( .A(n33725), .B(n33726), .Z(n33718) );
  NOR U33638 ( .A(n33727), .B(n33728), .Z(n33726) );
  XNOR U33639 ( .A(n33725), .B(n33729), .Z(n33727) );
  XOR U33640 ( .A(n33730), .B(n33731), .Z(n33686) );
  NOR U33641 ( .A(n33732), .B(n33733), .Z(n33731) );
  XNOR U33642 ( .A(n33730), .B(n33734), .Z(n33732) );
  XNOR U33643 ( .A(n33631), .B(n33689), .Z(n33691) );
  XNOR U33644 ( .A(n33735), .B(n33736), .Z(n33631) );
  AND U33645 ( .A(n1183), .B(n33638), .Z(n33736) );
  XOR U33646 ( .A(n33735), .B(n33636), .Z(n33638) );
  AND U33647 ( .A(n33639), .B(n33642), .Z(n33689) );
  XOR U33648 ( .A(n33737), .B(n33717), .Z(n33642) );
  XNOR U33649 ( .A(p_input[1664]), .B(p_input[2048]), .Z(n33717) );
  XNOR U33650 ( .A(n33704), .B(n33703), .Z(n33737) );
  XNOR U33651 ( .A(n33738), .B(n33711), .Z(n33703) );
  XNOR U33652 ( .A(n33699), .B(n33698), .Z(n33711) );
  XNOR U33653 ( .A(n33739), .B(n33695), .Z(n33698) );
  XNOR U33654 ( .A(p_input[1674]), .B(p_input[2058]), .Z(n33695) );
  XOR U33655 ( .A(p_input[1675]), .B(n16732), .Z(n33739) );
  XOR U33656 ( .A(p_input[1676]), .B(p_input[2060]), .Z(n33699) );
  XOR U33657 ( .A(n33709), .B(n33740), .Z(n33738) );
  IV U33658 ( .A(n33700), .Z(n33740) );
  XOR U33659 ( .A(p_input[1665]), .B(p_input[2049]), .Z(n33700) );
  XNOR U33660 ( .A(n33741), .B(n33716), .Z(n33709) );
  XNOR U33661 ( .A(p_input[1679]), .B(n16735), .Z(n33716) );
  XOR U33662 ( .A(n33706), .B(n33715), .Z(n33741) );
  XOR U33663 ( .A(n33742), .B(n33712), .Z(n33715) );
  XOR U33664 ( .A(p_input[1677]), .B(p_input[2061]), .Z(n33712) );
  XOR U33665 ( .A(p_input[1678]), .B(n16737), .Z(n33742) );
  XOR U33666 ( .A(p_input[1673]), .B(p_input[2057]), .Z(n33706) );
  XOR U33667 ( .A(n33724), .B(n33722), .Z(n33704) );
  XNOR U33668 ( .A(n33743), .B(n33729), .Z(n33722) );
  XOR U33669 ( .A(p_input[1672]), .B(p_input[2056]), .Z(n33729) );
  XOR U33670 ( .A(n33719), .B(n33728), .Z(n33743) );
  XOR U33671 ( .A(n33744), .B(n33725), .Z(n33728) );
  XOR U33672 ( .A(p_input[1670]), .B(p_input[2054]), .Z(n33725) );
  XOR U33673 ( .A(p_input[1671]), .B(n17722), .Z(n33744) );
  XOR U33674 ( .A(p_input[1666]), .B(p_input[2050]), .Z(n33719) );
  XNOR U33675 ( .A(n33734), .B(n33733), .Z(n33724) );
  XOR U33676 ( .A(n33745), .B(n33730), .Z(n33733) );
  XOR U33677 ( .A(p_input[1667]), .B(p_input[2051]), .Z(n33730) );
  XOR U33678 ( .A(p_input[1668]), .B(n17724), .Z(n33745) );
  XOR U33679 ( .A(p_input[1669]), .B(p_input[2053]), .Z(n33734) );
  XNOR U33680 ( .A(n33746), .B(n33747), .Z(n33639) );
  AND U33681 ( .A(n1183), .B(n33748), .Z(n33747) );
  XNOR U33682 ( .A(n33749), .B(n33750), .Z(n1183) );
  AND U33683 ( .A(n33751), .B(n33752), .Z(n33750) );
  XOR U33684 ( .A(n33749), .B(n33649), .Z(n33752) );
  XNOR U33685 ( .A(n33749), .B(n33603), .Z(n33751) );
  XOR U33686 ( .A(n33753), .B(n33754), .Z(n33749) );
  AND U33687 ( .A(n33755), .B(n33756), .Z(n33754) );
  XOR U33688 ( .A(n33753), .B(n33613), .Z(n33755) );
  XOR U33689 ( .A(n33757), .B(n33758), .Z(n33592) );
  AND U33690 ( .A(n1187), .B(n33748), .Z(n33758) );
  XNOR U33691 ( .A(n33746), .B(n33757), .Z(n33748) );
  XNOR U33692 ( .A(n33759), .B(n33760), .Z(n1187) );
  AND U33693 ( .A(n33761), .B(n33762), .Z(n33760) );
  XNOR U33694 ( .A(n33763), .B(n33759), .Z(n33762) );
  IV U33695 ( .A(n33649), .Z(n33763) );
  XNOR U33696 ( .A(n33764), .B(n33765), .Z(n33649) );
  AND U33697 ( .A(n1190), .B(n33766), .Z(n33765) );
  XNOR U33698 ( .A(n33764), .B(n33767), .Z(n33766) );
  XNOR U33699 ( .A(n33603), .B(n33759), .Z(n33761) );
  XOR U33700 ( .A(n33768), .B(n33769), .Z(n33603) );
  AND U33701 ( .A(n1198), .B(n33770), .Z(n33769) );
  XOR U33702 ( .A(n33753), .B(n33771), .Z(n33759) );
  AND U33703 ( .A(n33772), .B(n33756), .Z(n33771) );
  XNOR U33704 ( .A(n33662), .B(n33753), .Z(n33756) );
  XNOR U33705 ( .A(n33773), .B(n33774), .Z(n33662) );
  AND U33706 ( .A(n1190), .B(n33775), .Z(n33774) );
  XOR U33707 ( .A(n33776), .B(n33773), .Z(n33775) );
  XNOR U33708 ( .A(n33777), .B(n33753), .Z(n33772) );
  IV U33709 ( .A(n33613), .Z(n33777) );
  XOR U33710 ( .A(n33778), .B(n33779), .Z(n33613) );
  AND U33711 ( .A(n1198), .B(n33780), .Z(n33779) );
  XOR U33712 ( .A(n33781), .B(n33782), .Z(n33753) );
  AND U33713 ( .A(n33783), .B(n33784), .Z(n33782) );
  XNOR U33714 ( .A(n33687), .B(n33781), .Z(n33784) );
  XNOR U33715 ( .A(n33785), .B(n33786), .Z(n33687) );
  AND U33716 ( .A(n1190), .B(n33787), .Z(n33786) );
  XNOR U33717 ( .A(n33788), .B(n33785), .Z(n33787) );
  XOR U33718 ( .A(n33781), .B(n33624), .Z(n33783) );
  XOR U33719 ( .A(n33789), .B(n33790), .Z(n33624) );
  AND U33720 ( .A(n1198), .B(n33791), .Z(n33790) );
  XOR U33721 ( .A(n33792), .B(n33793), .Z(n33781) );
  AND U33722 ( .A(n33794), .B(n33795), .Z(n33793) );
  XNOR U33723 ( .A(n33792), .B(n33735), .Z(n33795) );
  XNOR U33724 ( .A(n33796), .B(n33797), .Z(n33735) );
  AND U33725 ( .A(n1190), .B(n33798), .Z(n33797) );
  XOR U33726 ( .A(n33799), .B(n33796), .Z(n33798) );
  XNOR U33727 ( .A(n33800), .B(n33792), .Z(n33794) );
  IV U33728 ( .A(n33636), .Z(n33800) );
  XOR U33729 ( .A(n33801), .B(n33802), .Z(n33636) );
  AND U33730 ( .A(n1198), .B(n33803), .Z(n33802) );
  AND U33731 ( .A(n33757), .B(n33746), .Z(n33792) );
  XNOR U33732 ( .A(n33804), .B(n33805), .Z(n33746) );
  AND U33733 ( .A(n1190), .B(n33806), .Z(n33805) );
  XNOR U33734 ( .A(n33807), .B(n33804), .Z(n33806) );
  XNOR U33735 ( .A(n33808), .B(n33809), .Z(n1190) );
  AND U33736 ( .A(n33810), .B(n33811), .Z(n33809) );
  XOR U33737 ( .A(n33767), .B(n33808), .Z(n33811) );
  AND U33738 ( .A(n33812), .B(n33813), .Z(n33767) );
  XOR U33739 ( .A(n33808), .B(n33764), .Z(n33810) );
  XNOR U33740 ( .A(n33814), .B(n33815), .Z(n33764) );
  AND U33741 ( .A(n1194), .B(n33770), .Z(n33815) );
  XOR U33742 ( .A(n33768), .B(n33814), .Z(n33770) );
  XOR U33743 ( .A(n33816), .B(n33817), .Z(n33808) );
  AND U33744 ( .A(n33818), .B(n33819), .Z(n33817) );
  XNOR U33745 ( .A(n33816), .B(n33812), .Z(n33819) );
  IV U33746 ( .A(n33776), .Z(n33812) );
  XOR U33747 ( .A(n33820), .B(n33821), .Z(n33776) );
  XOR U33748 ( .A(n33822), .B(n33813), .Z(n33821) );
  AND U33749 ( .A(n33788), .B(n33823), .Z(n33813) );
  AND U33750 ( .A(n33824), .B(n33825), .Z(n33822) );
  XOR U33751 ( .A(n33826), .B(n33820), .Z(n33824) );
  XNOR U33752 ( .A(n33773), .B(n33816), .Z(n33818) );
  XNOR U33753 ( .A(n33827), .B(n33828), .Z(n33773) );
  AND U33754 ( .A(n1194), .B(n33780), .Z(n33828) );
  XOR U33755 ( .A(n33827), .B(n33778), .Z(n33780) );
  XOR U33756 ( .A(n33829), .B(n33830), .Z(n33816) );
  AND U33757 ( .A(n33831), .B(n33832), .Z(n33830) );
  XNOR U33758 ( .A(n33829), .B(n33788), .Z(n33832) );
  XOR U33759 ( .A(n33833), .B(n33825), .Z(n33788) );
  XNOR U33760 ( .A(n33834), .B(n33820), .Z(n33825) );
  XOR U33761 ( .A(n33835), .B(n33836), .Z(n33820) );
  AND U33762 ( .A(n33837), .B(n33838), .Z(n33836) );
  XOR U33763 ( .A(n33839), .B(n33835), .Z(n33837) );
  XNOR U33764 ( .A(n33840), .B(n33841), .Z(n33834) );
  AND U33765 ( .A(n33842), .B(n33843), .Z(n33841) );
  XOR U33766 ( .A(n33840), .B(n33844), .Z(n33842) );
  XNOR U33767 ( .A(n33826), .B(n33823), .Z(n33833) );
  AND U33768 ( .A(n33845), .B(n33846), .Z(n33823) );
  XOR U33769 ( .A(n33847), .B(n33848), .Z(n33826) );
  AND U33770 ( .A(n33849), .B(n33850), .Z(n33848) );
  XOR U33771 ( .A(n33847), .B(n33851), .Z(n33849) );
  XNOR U33772 ( .A(n33785), .B(n33829), .Z(n33831) );
  XNOR U33773 ( .A(n33852), .B(n33853), .Z(n33785) );
  AND U33774 ( .A(n1194), .B(n33791), .Z(n33853) );
  XOR U33775 ( .A(n33852), .B(n33789), .Z(n33791) );
  XOR U33776 ( .A(n33854), .B(n33855), .Z(n33829) );
  AND U33777 ( .A(n33856), .B(n33857), .Z(n33855) );
  XNOR U33778 ( .A(n33854), .B(n33845), .Z(n33857) );
  IV U33779 ( .A(n33799), .Z(n33845) );
  XNOR U33780 ( .A(n33858), .B(n33838), .Z(n33799) );
  XNOR U33781 ( .A(n33859), .B(n33844), .Z(n33838) );
  XNOR U33782 ( .A(n33860), .B(n33861), .Z(n33844) );
  NOR U33783 ( .A(n33862), .B(n33863), .Z(n33861) );
  XOR U33784 ( .A(n33860), .B(n33864), .Z(n33862) );
  XNOR U33785 ( .A(n33843), .B(n33835), .Z(n33859) );
  XOR U33786 ( .A(n33865), .B(n33866), .Z(n33835) );
  AND U33787 ( .A(n33867), .B(n33868), .Z(n33866) );
  XOR U33788 ( .A(n33865), .B(n33869), .Z(n33867) );
  XNOR U33789 ( .A(n33870), .B(n33840), .Z(n33843) );
  XOR U33790 ( .A(n33871), .B(n33872), .Z(n33840) );
  AND U33791 ( .A(n33873), .B(n33874), .Z(n33872) );
  XNOR U33792 ( .A(n33875), .B(n33876), .Z(n33873) );
  IV U33793 ( .A(n33871), .Z(n33875) );
  XNOR U33794 ( .A(n33877), .B(n33878), .Z(n33870) );
  NOR U33795 ( .A(n33879), .B(n33880), .Z(n33878) );
  XNOR U33796 ( .A(n33877), .B(n33881), .Z(n33879) );
  XNOR U33797 ( .A(n33839), .B(n33846), .Z(n33858) );
  NOR U33798 ( .A(n33807), .B(n33882), .Z(n33846) );
  XOR U33799 ( .A(n33851), .B(n33850), .Z(n33839) );
  XNOR U33800 ( .A(n33883), .B(n33847), .Z(n33850) );
  XOR U33801 ( .A(n33884), .B(n33885), .Z(n33847) );
  AND U33802 ( .A(n33886), .B(n33887), .Z(n33885) );
  XNOR U33803 ( .A(n33888), .B(n33889), .Z(n33886) );
  IV U33804 ( .A(n33884), .Z(n33888) );
  XNOR U33805 ( .A(n33890), .B(n33891), .Z(n33883) );
  NOR U33806 ( .A(n33892), .B(n33893), .Z(n33891) );
  XNOR U33807 ( .A(n33890), .B(n33894), .Z(n33892) );
  XOR U33808 ( .A(n33895), .B(n33896), .Z(n33851) );
  NOR U33809 ( .A(n33897), .B(n33898), .Z(n33896) );
  XNOR U33810 ( .A(n33895), .B(n33899), .Z(n33897) );
  XNOR U33811 ( .A(n33796), .B(n33854), .Z(n33856) );
  XNOR U33812 ( .A(n33900), .B(n33901), .Z(n33796) );
  AND U33813 ( .A(n1194), .B(n33803), .Z(n33901) );
  XOR U33814 ( .A(n33900), .B(n33801), .Z(n33803) );
  AND U33815 ( .A(n33804), .B(n33807), .Z(n33854) );
  XOR U33816 ( .A(n33902), .B(n33882), .Z(n33807) );
  XNOR U33817 ( .A(p_input[1680]), .B(p_input[2048]), .Z(n33882) );
  XNOR U33818 ( .A(n33869), .B(n33868), .Z(n33902) );
  XNOR U33819 ( .A(n33903), .B(n33876), .Z(n33868) );
  XNOR U33820 ( .A(n33864), .B(n33863), .Z(n33876) );
  XNOR U33821 ( .A(n33904), .B(n33860), .Z(n33863) );
  XNOR U33822 ( .A(p_input[1690]), .B(p_input[2058]), .Z(n33860) );
  XOR U33823 ( .A(p_input[1691]), .B(n16732), .Z(n33904) );
  XOR U33824 ( .A(p_input[1692]), .B(p_input[2060]), .Z(n33864) );
  XOR U33825 ( .A(n33874), .B(n33905), .Z(n33903) );
  IV U33826 ( .A(n33865), .Z(n33905) );
  XOR U33827 ( .A(p_input[1681]), .B(p_input[2049]), .Z(n33865) );
  XNOR U33828 ( .A(n33906), .B(n33881), .Z(n33874) );
  XNOR U33829 ( .A(p_input[1695]), .B(n16735), .Z(n33881) );
  XOR U33830 ( .A(n33871), .B(n33880), .Z(n33906) );
  XOR U33831 ( .A(n33907), .B(n33877), .Z(n33880) );
  XOR U33832 ( .A(p_input[1693]), .B(p_input[2061]), .Z(n33877) );
  XOR U33833 ( .A(p_input[1694]), .B(n16737), .Z(n33907) );
  XOR U33834 ( .A(p_input[1689]), .B(p_input[2057]), .Z(n33871) );
  XOR U33835 ( .A(n33889), .B(n33887), .Z(n33869) );
  XNOR U33836 ( .A(n33908), .B(n33894), .Z(n33887) );
  XOR U33837 ( .A(p_input[1688]), .B(p_input[2056]), .Z(n33894) );
  XOR U33838 ( .A(n33884), .B(n33893), .Z(n33908) );
  XOR U33839 ( .A(n33909), .B(n33890), .Z(n33893) );
  XOR U33840 ( .A(p_input[1686]), .B(p_input[2054]), .Z(n33890) );
  XOR U33841 ( .A(p_input[1687]), .B(n17722), .Z(n33909) );
  XOR U33842 ( .A(p_input[1682]), .B(p_input[2050]), .Z(n33884) );
  XNOR U33843 ( .A(n33899), .B(n33898), .Z(n33889) );
  XOR U33844 ( .A(n33910), .B(n33895), .Z(n33898) );
  XOR U33845 ( .A(p_input[1683]), .B(p_input[2051]), .Z(n33895) );
  XOR U33846 ( .A(p_input[1684]), .B(n17724), .Z(n33910) );
  XOR U33847 ( .A(p_input[1685]), .B(p_input[2053]), .Z(n33899) );
  XNOR U33848 ( .A(n33911), .B(n33912), .Z(n33804) );
  AND U33849 ( .A(n1194), .B(n33913), .Z(n33912) );
  XNOR U33850 ( .A(n33914), .B(n33915), .Z(n1194) );
  AND U33851 ( .A(n33916), .B(n33917), .Z(n33915) );
  XOR U33852 ( .A(n33914), .B(n33814), .Z(n33917) );
  XNOR U33853 ( .A(n33914), .B(n33768), .Z(n33916) );
  XOR U33854 ( .A(n33918), .B(n33919), .Z(n33914) );
  AND U33855 ( .A(n33920), .B(n33921), .Z(n33919) );
  XOR U33856 ( .A(n33918), .B(n33778), .Z(n33920) );
  XOR U33857 ( .A(n33922), .B(n33923), .Z(n33757) );
  AND U33858 ( .A(n1198), .B(n33913), .Z(n33923) );
  XNOR U33859 ( .A(n33911), .B(n33922), .Z(n33913) );
  XNOR U33860 ( .A(n33924), .B(n33925), .Z(n1198) );
  AND U33861 ( .A(n33926), .B(n33927), .Z(n33925) );
  XNOR U33862 ( .A(n33928), .B(n33924), .Z(n33927) );
  IV U33863 ( .A(n33814), .Z(n33928) );
  XNOR U33864 ( .A(n33929), .B(n33930), .Z(n33814) );
  AND U33865 ( .A(n1201), .B(n33931), .Z(n33930) );
  XNOR U33866 ( .A(n33929), .B(n33932), .Z(n33931) );
  XNOR U33867 ( .A(n33768), .B(n33924), .Z(n33926) );
  XOR U33868 ( .A(n33933), .B(n33934), .Z(n33768) );
  AND U33869 ( .A(n1209), .B(n33935), .Z(n33934) );
  XOR U33870 ( .A(n33918), .B(n33936), .Z(n33924) );
  AND U33871 ( .A(n33937), .B(n33921), .Z(n33936) );
  XNOR U33872 ( .A(n33827), .B(n33918), .Z(n33921) );
  XNOR U33873 ( .A(n33938), .B(n33939), .Z(n33827) );
  AND U33874 ( .A(n1201), .B(n33940), .Z(n33939) );
  XOR U33875 ( .A(n33941), .B(n33938), .Z(n33940) );
  XNOR U33876 ( .A(n33942), .B(n33918), .Z(n33937) );
  IV U33877 ( .A(n33778), .Z(n33942) );
  XOR U33878 ( .A(n33943), .B(n33944), .Z(n33778) );
  AND U33879 ( .A(n1209), .B(n33945), .Z(n33944) );
  XOR U33880 ( .A(n33946), .B(n33947), .Z(n33918) );
  AND U33881 ( .A(n33948), .B(n33949), .Z(n33947) );
  XNOR U33882 ( .A(n33852), .B(n33946), .Z(n33949) );
  XNOR U33883 ( .A(n33950), .B(n33951), .Z(n33852) );
  AND U33884 ( .A(n1201), .B(n33952), .Z(n33951) );
  XNOR U33885 ( .A(n33953), .B(n33950), .Z(n33952) );
  XOR U33886 ( .A(n33946), .B(n33789), .Z(n33948) );
  XOR U33887 ( .A(n33954), .B(n33955), .Z(n33789) );
  AND U33888 ( .A(n1209), .B(n33956), .Z(n33955) );
  XOR U33889 ( .A(n33957), .B(n33958), .Z(n33946) );
  AND U33890 ( .A(n33959), .B(n33960), .Z(n33958) );
  XNOR U33891 ( .A(n33957), .B(n33900), .Z(n33960) );
  XNOR U33892 ( .A(n33961), .B(n33962), .Z(n33900) );
  AND U33893 ( .A(n1201), .B(n33963), .Z(n33962) );
  XOR U33894 ( .A(n33964), .B(n33961), .Z(n33963) );
  XNOR U33895 ( .A(n33965), .B(n33957), .Z(n33959) );
  IV U33896 ( .A(n33801), .Z(n33965) );
  XOR U33897 ( .A(n33966), .B(n33967), .Z(n33801) );
  AND U33898 ( .A(n1209), .B(n33968), .Z(n33967) );
  AND U33899 ( .A(n33922), .B(n33911), .Z(n33957) );
  XNOR U33900 ( .A(n33969), .B(n33970), .Z(n33911) );
  AND U33901 ( .A(n1201), .B(n33971), .Z(n33970) );
  XNOR U33902 ( .A(n33972), .B(n33969), .Z(n33971) );
  XNOR U33903 ( .A(n33973), .B(n33974), .Z(n1201) );
  AND U33904 ( .A(n33975), .B(n33976), .Z(n33974) );
  XOR U33905 ( .A(n33932), .B(n33973), .Z(n33976) );
  AND U33906 ( .A(n33977), .B(n33978), .Z(n33932) );
  XOR U33907 ( .A(n33973), .B(n33929), .Z(n33975) );
  XNOR U33908 ( .A(n33979), .B(n33980), .Z(n33929) );
  AND U33909 ( .A(n1205), .B(n33935), .Z(n33980) );
  XOR U33910 ( .A(n33933), .B(n33979), .Z(n33935) );
  XOR U33911 ( .A(n33981), .B(n33982), .Z(n33973) );
  AND U33912 ( .A(n33983), .B(n33984), .Z(n33982) );
  XNOR U33913 ( .A(n33981), .B(n33977), .Z(n33984) );
  IV U33914 ( .A(n33941), .Z(n33977) );
  XOR U33915 ( .A(n33985), .B(n33986), .Z(n33941) );
  XOR U33916 ( .A(n33987), .B(n33978), .Z(n33986) );
  AND U33917 ( .A(n33953), .B(n33988), .Z(n33978) );
  AND U33918 ( .A(n33989), .B(n33990), .Z(n33987) );
  XOR U33919 ( .A(n33991), .B(n33985), .Z(n33989) );
  XNOR U33920 ( .A(n33938), .B(n33981), .Z(n33983) );
  XNOR U33921 ( .A(n33992), .B(n33993), .Z(n33938) );
  AND U33922 ( .A(n1205), .B(n33945), .Z(n33993) );
  XOR U33923 ( .A(n33992), .B(n33943), .Z(n33945) );
  XOR U33924 ( .A(n33994), .B(n33995), .Z(n33981) );
  AND U33925 ( .A(n33996), .B(n33997), .Z(n33995) );
  XNOR U33926 ( .A(n33994), .B(n33953), .Z(n33997) );
  XOR U33927 ( .A(n33998), .B(n33990), .Z(n33953) );
  XNOR U33928 ( .A(n33999), .B(n33985), .Z(n33990) );
  XOR U33929 ( .A(n34000), .B(n34001), .Z(n33985) );
  AND U33930 ( .A(n34002), .B(n34003), .Z(n34001) );
  XOR U33931 ( .A(n34004), .B(n34000), .Z(n34002) );
  XNOR U33932 ( .A(n34005), .B(n34006), .Z(n33999) );
  AND U33933 ( .A(n34007), .B(n34008), .Z(n34006) );
  XOR U33934 ( .A(n34005), .B(n34009), .Z(n34007) );
  XNOR U33935 ( .A(n33991), .B(n33988), .Z(n33998) );
  AND U33936 ( .A(n34010), .B(n34011), .Z(n33988) );
  XOR U33937 ( .A(n34012), .B(n34013), .Z(n33991) );
  AND U33938 ( .A(n34014), .B(n34015), .Z(n34013) );
  XOR U33939 ( .A(n34012), .B(n34016), .Z(n34014) );
  XNOR U33940 ( .A(n33950), .B(n33994), .Z(n33996) );
  XNOR U33941 ( .A(n34017), .B(n34018), .Z(n33950) );
  AND U33942 ( .A(n1205), .B(n33956), .Z(n34018) );
  XOR U33943 ( .A(n34017), .B(n33954), .Z(n33956) );
  XOR U33944 ( .A(n34019), .B(n34020), .Z(n33994) );
  AND U33945 ( .A(n34021), .B(n34022), .Z(n34020) );
  XNOR U33946 ( .A(n34019), .B(n34010), .Z(n34022) );
  IV U33947 ( .A(n33964), .Z(n34010) );
  XNOR U33948 ( .A(n34023), .B(n34003), .Z(n33964) );
  XNOR U33949 ( .A(n34024), .B(n34009), .Z(n34003) );
  XNOR U33950 ( .A(n34025), .B(n34026), .Z(n34009) );
  NOR U33951 ( .A(n34027), .B(n34028), .Z(n34026) );
  XOR U33952 ( .A(n34025), .B(n34029), .Z(n34027) );
  XNOR U33953 ( .A(n34008), .B(n34000), .Z(n34024) );
  XOR U33954 ( .A(n34030), .B(n34031), .Z(n34000) );
  AND U33955 ( .A(n34032), .B(n34033), .Z(n34031) );
  XOR U33956 ( .A(n34030), .B(n34034), .Z(n34032) );
  XNOR U33957 ( .A(n34035), .B(n34005), .Z(n34008) );
  XOR U33958 ( .A(n34036), .B(n34037), .Z(n34005) );
  AND U33959 ( .A(n34038), .B(n34039), .Z(n34037) );
  XNOR U33960 ( .A(n34040), .B(n34041), .Z(n34038) );
  IV U33961 ( .A(n34036), .Z(n34040) );
  XNOR U33962 ( .A(n34042), .B(n34043), .Z(n34035) );
  NOR U33963 ( .A(n34044), .B(n34045), .Z(n34043) );
  XNOR U33964 ( .A(n34042), .B(n34046), .Z(n34044) );
  XNOR U33965 ( .A(n34004), .B(n34011), .Z(n34023) );
  NOR U33966 ( .A(n33972), .B(n34047), .Z(n34011) );
  XOR U33967 ( .A(n34016), .B(n34015), .Z(n34004) );
  XNOR U33968 ( .A(n34048), .B(n34012), .Z(n34015) );
  XOR U33969 ( .A(n34049), .B(n34050), .Z(n34012) );
  AND U33970 ( .A(n34051), .B(n34052), .Z(n34050) );
  XNOR U33971 ( .A(n34053), .B(n34054), .Z(n34051) );
  IV U33972 ( .A(n34049), .Z(n34053) );
  XNOR U33973 ( .A(n34055), .B(n34056), .Z(n34048) );
  NOR U33974 ( .A(n34057), .B(n34058), .Z(n34056) );
  XNOR U33975 ( .A(n34055), .B(n34059), .Z(n34057) );
  XOR U33976 ( .A(n34060), .B(n34061), .Z(n34016) );
  NOR U33977 ( .A(n34062), .B(n34063), .Z(n34061) );
  XNOR U33978 ( .A(n34060), .B(n34064), .Z(n34062) );
  XNOR U33979 ( .A(n33961), .B(n34019), .Z(n34021) );
  XNOR U33980 ( .A(n34065), .B(n34066), .Z(n33961) );
  AND U33981 ( .A(n1205), .B(n33968), .Z(n34066) );
  XOR U33982 ( .A(n34065), .B(n33966), .Z(n33968) );
  AND U33983 ( .A(n33969), .B(n33972), .Z(n34019) );
  XOR U33984 ( .A(n34067), .B(n34047), .Z(n33972) );
  XNOR U33985 ( .A(p_input[1696]), .B(p_input[2048]), .Z(n34047) );
  XNOR U33986 ( .A(n34034), .B(n34033), .Z(n34067) );
  XNOR U33987 ( .A(n34068), .B(n34041), .Z(n34033) );
  XNOR U33988 ( .A(n34029), .B(n34028), .Z(n34041) );
  XNOR U33989 ( .A(n34069), .B(n34025), .Z(n34028) );
  XNOR U33990 ( .A(p_input[1706]), .B(p_input[2058]), .Z(n34025) );
  XOR U33991 ( .A(p_input[1707]), .B(n16732), .Z(n34069) );
  XOR U33992 ( .A(p_input[1708]), .B(p_input[2060]), .Z(n34029) );
  XOR U33993 ( .A(n34039), .B(n34070), .Z(n34068) );
  IV U33994 ( .A(n34030), .Z(n34070) );
  XOR U33995 ( .A(p_input[1697]), .B(p_input[2049]), .Z(n34030) );
  XNOR U33996 ( .A(n34071), .B(n34046), .Z(n34039) );
  XNOR U33997 ( .A(p_input[1711]), .B(n16735), .Z(n34046) );
  XOR U33998 ( .A(n34036), .B(n34045), .Z(n34071) );
  XOR U33999 ( .A(n34072), .B(n34042), .Z(n34045) );
  XOR U34000 ( .A(p_input[1709]), .B(p_input[2061]), .Z(n34042) );
  XOR U34001 ( .A(p_input[1710]), .B(n16737), .Z(n34072) );
  XOR U34002 ( .A(p_input[1705]), .B(p_input[2057]), .Z(n34036) );
  XOR U34003 ( .A(n34054), .B(n34052), .Z(n34034) );
  XNOR U34004 ( .A(n34073), .B(n34059), .Z(n34052) );
  XOR U34005 ( .A(p_input[1704]), .B(p_input[2056]), .Z(n34059) );
  XOR U34006 ( .A(n34049), .B(n34058), .Z(n34073) );
  XOR U34007 ( .A(n34074), .B(n34055), .Z(n34058) );
  XOR U34008 ( .A(p_input[1702]), .B(p_input[2054]), .Z(n34055) );
  XOR U34009 ( .A(p_input[1703]), .B(n17722), .Z(n34074) );
  XOR U34010 ( .A(p_input[1698]), .B(p_input[2050]), .Z(n34049) );
  XNOR U34011 ( .A(n34064), .B(n34063), .Z(n34054) );
  XOR U34012 ( .A(n34075), .B(n34060), .Z(n34063) );
  XOR U34013 ( .A(p_input[1699]), .B(p_input[2051]), .Z(n34060) );
  XOR U34014 ( .A(p_input[1700]), .B(n17724), .Z(n34075) );
  XOR U34015 ( .A(p_input[1701]), .B(p_input[2053]), .Z(n34064) );
  XNOR U34016 ( .A(n34076), .B(n34077), .Z(n33969) );
  AND U34017 ( .A(n1205), .B(n34078), .Z(n34077) );
  XNOR U34018 ( .A(n34079), .B(n34080), .Z(n1205) );
  AND U34019 ( .A(n34081), .B(n34082), .Z(n34080) );
  XOR U34020 ( .A(n34079), .B(n33979), .Z(n34082) );
  XNOR U34021 ( .A(n34079), .B(n33933), .Z(n34081) );
  XOR U34022 ( .A(n34083), .B(n34084), .Z(n34079) );
  AND U34023 ( .A(n34085), .B(n34086), .Z(n34084) );
  XOR U34024 ( .A(n34083), .B(n33943), .Z(n34085) );
  XOR U34025 ( .A(n34087), .B(n34088), .Z(n33922) );
  AND U34026 ( .A(n1209), .B(n34078), .Z(n34088) );
  XNOR U34027 ( .A(n34076), .B(n34087), .Z(n34078) );
  XNOR U34028 ( .A(n34089), .B(n34090), .Z(n1209) );
  AND U34029 ( .A(n34091), .B(n34092), .Z(n34090) );
  XNOR U34030 ( .A(n34093), .B(n34089), .Z(n34092) );
  IV U34031 ( .A(n33979), .Z(n34093) );
  XNOR U34032 ( .A(n34094), .B(n34095), .Z(n33979) );
  AND U34033 ( .A(n1212), .B(n34096), .Z(n34095) );
  XNOR U34034 ( .A(n34094), .B(n34097), .Z(n34096) );
  XNOR U34035 ( .A(n33933), .B(n34089), .Z(n34091) );
  XOR U34036 ( .A(n34098), .B(n34099), .Z(n33933) );
  AND U34037 ( .A(n1220), .B(n34100), .Z(n34099) );
  XOR U34038 ( .A(n34083), .B(n34101), .Z(n34089) );
  AND U34039 ( .A(n34102), .B(n34086), .Z(n34101) );
  XNOR U34040 ( .A(n33992), .B(n34083), .Z(n34086) );
  XNOR U34041 ( .A(n34103), .B(n34104), .Z(n33992) );
  AND U34042 ( .A(n1212), .B(n34105), .Z(n34104) );
  XOR U34043 ( .A(n34106), .B(n34103), .Z(n34105) );
  XNOR U34044 ( .A(n34107), .B(n34083), .Z(n34102) );
  IV U34045 ( .A(n33943), .Z(n34107) );
  XOR U34046 ( .A(n34108), .B(n34109), .Z(n33943) );
  AND U34047 ( .A(n1220), .B(n34110), .Z(n34109) );
  XOR U34048 ( .A(n34111), .B(n34112), .Z(n34083) );
  AND U34049 ( .A(n34113), .B(n34114), .Z(n34112) );
  XNOR U34050 ( .A(n34017), .B(n34111), .Z(n34114) );
  XNOR U34051 ( .A(n34115), .B(n34116), .Z(n34017) );
  AND U34052 ( .A(n1212), .B(n34117), .Z(n34116) );
  XNOR U34053 ( .A(n34118), .B(n34115), .Z(n34117) );
  XOR U34054 ( .A(n34111), .B(n33954), .Z(n34113) );
  XOR U34055 ( .A(n34119), .B(n34120), .Z(n33954) );
  AND U34056 ( .A(n1220), .B(n34121), .Z(n34120) );
  XOR U34057 ( .A(n34122), .B(n34123), .Z(n34111) );
  AND U34058 ( .A(n34124), .B(n34125), .Z(n34123) );
  XNOR U34059 ( .A(n34122), .B(n34065), .Z(n34125) );
  XNOR U34060 ( .A(n34126), .B(n34127), .Z(n34065) );
  AND U34061 ( .A(n1212), .B(n34128), .Z(n34127) );
  XOR U34062 ( .A(n34129), .B(n34126), .Z(n34128) );
  XNOR U34063 ( .A(n34130), .B(n34122), .Z(n34124) );
  IV U34064 ( .A(n33966), .Z(n34130) );
  XOR U34065 ( .A(n34131), .B(n34132), .Z(n33966) );
  AND U34066 ( .A(n1220), .B(n34133), .Z(n34132) );
  AND U34067 ( .A(n34087), .B(n34076), .Z(n34122) );
  XNOR U34068 ( .A(n34134), .B(n34135), .Z(n34076) );
  AND U34069 ( .A(n1212), .B(n34136), .Z(n34135) );
  XNOR U34070 ( .A(n34137), .B(n34134), .Z(n34136) );
  XNOR U34071 ( .A(n34138), .B(n34139), .Z(n1212) );
  AND U34072 ( .A(n34140), .B(n34141), .Z(n34139) );
  XOR U34073 ( .A(n34097), .B(n34138), .Z(n34141) );
  AND U34074 ( .A(n34142), .B(n34143), .Z(n34097) );
  XOR U34075 ( .A(n34138), .B(n34094), .Z(n34140) );
  XNOR U34076 ( .A(n34144), .B(n34145), .Z(n34094) );
  AND U34077 ( .A(n1216), .B(n34100), .Z(n34145) );
  XOR U34078 ( .A(n34098), .B(n34144), .Z(n34100) );
  XOR U34079 ( .A(n34146), .B(n34147), .Z(n34138) );
  AND U34080 ( .A(n34148), .B(n34149), .Z(n34147) );
  XNOR U34081 ( .A(n34146), .B(n34142), .Z(n34149) );
  IV U34082 ( .A(n34106), .Z(n34142) );
  XOR U34083 ( .A(n34150), .B(n34151), .Z(n34106) );
  XOR U34084 ( .A(n34152), .B(n34143), .Z(n34151) );
  AND U34085 ( .A(n34118), .B(n34153), .Z(n34143) );
  AND U34086 ( .A(n34154), .B(n34155), .Z(n34152) );
  XOR U34087 ( .A(n34156), .B(n34150), .Z(n34154) );
  XNOR U34088 ( .A(n34103), .B(n34146), .Z(n34148) );
  XNOR U34089 ( .A(n34157), .B(n34158), .Z(n34103) );
  AND U34090 ( .A(n1216), .B(n34110), .Z(n34158) );
  XOR U34091 ( .A(n34157), .B(n34108), .Z(n34110) );
  XOR U34092 ( .A(n34159), .B(n34160), .Z(n34146) );
  AND U34093 ( .A(n34161), .B(n34162), .Z(n34160) );
  XNOR U34094 ( .A(n34159), .B(n34118), .Z(n34162) );
  XOR U34095 ( .A(n34163), .B(n34155), .Z(n34118) );
  XNOR U34096 ( .A(n34164), .B(n34150), .Z(n34155) );
  XOR U34097 ( .A(n34165), .B(n34166), .Z(n34150) );
  AND U34098 ( .A(n34167), .B(n34168), .Z(n34166) );
  XOR U34099 ( .A(n34169), .B(n34165), .Z(n34167) );
  XNOR U34100 ( .A(n34170), .B(n34171), .Z(n34164) );
  AND U34101 ( .A(n34172), .B(n34173), .Z(n34171) );
  XOR U34102 ( .A(n34170), .B(n34174), .Z(n34172) );
  XNOR U34103 ( .A(n34156), .B(n34153), .Z(n34163) );
  AND U34104 ( .A(n34175), .B(n34176), .Z(n34153) );
  XOR U34105 ( .A(n34177), .B(n34178), .Z(n34156) );
  AND U34106 ( .A(n34179), .B(n34180), .Z(n34178) );
  XOR U34107 ( .A(n34177), .B(n34181), .Z(n34179) );
  XNOR U34108 ( .A(n34115), .B(n34159), .Z(n34161) );
  XNOR U34109 ( .A(n34182), .B(n34183), .Z(n34115) );
  AND U34110 ( .A(n1216), .B(n34121), .Z(n34183) );
  XOR U34111 ( .A(n34182), .B(n34119), .Z(n34121) );
  XOR U34112 ( .A(n34184), .B(n34185), .Z(n34159) );
  AND U34113 ( .A(n34186), .B(n34187), .Z(n34185) );
  XNOR U34114 ( .A(n34184), .B(n34175), .Z(n34187) );
  IV U34115 ( .A(n34129), .Z(n34175) );
  XNOR U34116 ( .A(n34188), .B(n34168), .Z(n34129) );
  XNOR U34117 ( .A(n34189), .B(n34174), .Z(n34168) );
  XNOR U34118 ( .A(n34190), .B(n34191), .Z(n34174) );
  NOR U34119 ( .A(n34192), .B(n34193), .Z(n34191) );
  XOR U34120 ( .A(n34190), .B(n34194), .Z(n34192) );
  XNOR U34121 ( .A(n34173), .B(n34165), .Z(n34189) );
  XOR U34122 ( .A(n34195), .B(n34196), .Z(n34165) );
  AND U34123 ( .A(n34197), .B(n34198), .Z(n34196) );
  XOR U34124 ( .A(n34195), .B(n34199), .Z(n34197) );
  XNOR U34125 ( .A(n34200), .B(n34170), .Z(n34173) );
  XOR U34126 ( .A(n34201), .B(n34202), .Z(n34170) );
  AND U34127 ( .A(n34203), .B(n34204), .Z(n34202) );
  XNOR U34128 ( .A(n34205), .B(n34206), .Z(n34203) );
  IV U34129 ( .A(n34201), .Z(n34205) );
  XNOR U34130 ( .A(n34207), .B(n34208), .Z(n34200) );
  NOR U34131 ( .A(n34209), .B(n34210), .Z(n34208) );
  XNOR U34132 ( .A(n34207), .B(n34211), .Z(n34209) );
  XNOR U34133 ( .A(n34169), .B(n34176), .Z(n34188) );
  NOR U34134 ( .A(n34137), .B(n34212), .Z(n34176) );
  XOR U34135 ( .A(n34181), .B(n34180), .Z(n34169) );
  XNOR U34136 ( .A(n34213), .B(n34177), .Z(n34180) );
  XOR U34137 ( .A(n34214), .B(n34215), .Z(n34177) );
  AND U34138 ( .A(n34216), .B(n34217), .Z(n34215) );
  XNOR U34139 ( .A(n34218), .B(n34219), .Z(n34216) );
  IV U34140 ( .A(n34214), .Z(n34218) );
  XNOR U34141 ( .A(n34220), .B(n34221), .Z(n34213) );
  NOR U34142 ( .A(n34222), .B(n34223), .Z(n34221) );
  XNOR U34143 ( .A(n34220), .B(n34224), .Z(n34222) );
  XOR U34144 ( .A(n34225), .B(n34226), .Z(n34181) );
  NOR U34145 ( .A(n34227), .B(n34228), .Z(n34226) );
  XNOR U34146 ( .A(n34225), .B(n34229), .Z(n34227) );
  XNOR U34147 ( .A(n34126), .B(n34184), .Z(n34186) );
  XNOR U34148 ( .A(n34230), .B(n34231), .Z(n34126) );
  AND U34149 ( .A(n1216), .B(n34133), .Z(n34231) );
  XOR U34150 ( .A(n34230), .B(n34131), .Z(n34133) );
  AND U34151 ( .A(n34134), .B(n34137), .Z(n34184) );
  XOR U34152 ( .A(n34232), .B(n34212), .Z(n34137) );
  XNOR U34153 ( .A(p_input[1712]), .B(p_input[2048]), .Z(n34212) );
  XNOR U34154 ( .A(n34199), .B(n34198), .Z(n34232) );
  XNOR U34155 ( .A(n34233), .B(n34206), .Z(n34198) );
  XNOR U34156 ( .A(n34194), .B(n34193), .Z(n34206) );
  XNOR U34157 ( .A(n34234), .B(n34190), .Z(n34193) );
  XNOR U34158 ( .A(p_input[1722]), .B(p_input[2058]), .Z(n34190) );
  XOR U34159 ( .A(p_input[1723]), .B(n16732), .Z(n34234) );
  XOR U34160 ( .A(p_input[1724]), .B(p_input[2060]), .Z(n34194) );
  XOR U34161 ( .A(n34204), .B(n34235), .Z(n34233) );
  IV U34162 ( .A(n34195), .Z(n34235) );
  XOR U34163 ( .A(p_input[1713]), .B(p_input[2049]), .Z(n34195) );
  XNOR U34164 ( .A(n34236), .B(n34211), .Z(n34204) );
  XNOR U34165 ( .A(p_input[1727]), .B(n16735), .Z(n34211) );
  XOR U34166 ( .A(n34201), .B(n34210), .Z(n34236) );
  XOR U34167 ( .A(n34237), .B(n34207), .Z(n34210) );
  XOR U34168 ( .A(p_input[1725]), .B(p_input[2061]), .Z(n34207) );
  XOR U34169 ( .A(p_input[1726]), .B(n16737), .Z(n34237) );
  XOR U34170 ( .A(p_input[1721]), .B(p_input[2057]), .Z(n34201) );
  XOR U34171 ( .A(n34219), .B(n34217), .Z(n34199) );
  XNOR U34172 ( .A(n34238), .B(n34224), .Z(n34217) );
  XOR U34173 ( .A(p_input[1720]), .B(p_input[2056]), .Z(n34224) );
  XOR U34174 ( .A(n34214), .B(n34223), .Z(n34238) );
  XOR U34175 ( .A(n34239), .B(n34220), .Z(n34223) );
  XOR U34176 ( .A(p_input[1718]), .B(p_input[2054]), .Z(n34220) );
  XOR U34177 ( .A(p_input[1719]), .B(n17722), .Z(n34239) );
  XOR U34178 ( .A(p_input[1714]), .B(p_input[2050]), .Z(n34214) );
  XNOR U34179 ( .A(n34229), .B(n34228), .Z(n34219) );
  XOR U34180 ( .A(n34240), .B(n34225), .Z(n34228) );
  XOR U34181 ( .A(p_input[1715]), .B(p_input[2051]), .Z(n34225) );
  XOR U34182 ( .A(p_input[1716]), .B(n17724), .Z(n34240) );
  XOR U34183 ( .A(p_input[1717]), .B(p_input[2053]), .Z(n34229) );
  XNOR U34184 ( .A(n34241), .B(n34242), .Z(n34134) );
  AND U34185 ( .A(n1216), .B(n34243), .Z(n34242) );
  XNOR U34186 ( .A(n34244), .B(n34245), .Z(n1216) );
  AND U34187 ( .A(n34246), .B(n34247), .Z(n34245) );
  XOR U34188 ( .A(n34244), .B(n34144), .Z(n34247) );
  XNOR U34189 ( .A(n34244), .B(n34098), .Z(n34246) );
  XOR U34190 ( .A(n34248), .B(n34249), .Z(n34244) );
  AND U34191 ( .A(n34250), .B(n34251), .Z(n34249) );
  XOR U34192 ( .A(n34248), .B(n34108), .Z(n34250) );
  XOR U34193 ( .A(n34252), .B(n34253), .Z(n34087) );
  AND U34194 ( .A(n1220), .B(n34243), .Z(n34253) );
  XNOR U34195 ( .A(n34241), .B(n34252), .Z(n34243) );
  XNOR U34196 ( .A(n34254), .B(n34255), .Z(n1220) );
  AND U34197 ( .A(n34256), .B(n34257), .Z(n34255) );
  XNOR U34198 ( .A(n34258), .B(n34254), .Z(n34257) );
  IV U34199 ( .A(n34144), .Z(n34258) );
  XNOR U34200 ( .A(n34259), .B(n34260), .Z(n34144) );
  AND U34201 ( .A(n1223), .B(n34261), .Z(n34260) );
  XNOR U34202 ( .A(n34259), .B(n34262), .Z(n34261) );
  XNOR U34203 ( .A(n34098), .B(n34254), .Z(n34256) );
  XOR U34204 ( .A(n34263), .B(n34264), .Z(n34098) );
  AND U34205 ( .A(n1231), .B(n34265), .Z(n34264) );
  XOR U34206 ( .A(n34248), .B(n34266), .Z(n34254) );
  AND U34207 ( .A(n34267), .B(n34251), .Z(n34266) );
  XNOR U34208 ( .A(n34157), .B(n34248), .Z(n34251) );
  XNOR U34209 ( .A(n34268), .B(n34269), .Z(n34157) );
  AND U34210 ( .A(n1223), .B(n34270), .Z(n34269) );
  XOR U34211 ( .A(n34271), .B(n34268), .Z(n34270) );
  XNOR U34212 ( .A(n34272), .B(n34248), .Z(n34267) );
  IV U34213 ( .A(n34108), .Z(n34272) );
  XOR U34214 ( .A(n34273), .B(n34274), .Z(n34108) );
  AND U34215 ( .A(n1231), .B(n34275), .Z(n34274) );
  XOR U34216 ( .A(n34276), .B(n34277), .Z(n34248) );
  AND U34217 ( .A(n34278), .B(n34279), .Z(n34277) );
  XNOR U34218 ( .A(n34182), .B(n34276), .Z(n34279) );
  XNOR U34219 ( .A(n34280), .B(n34281), .Z(n34182) );
  AND U34220 ( .A(n1223), .B(n34282), .Z(n34281) );
  XNOR U34221 ( .A(n34283), .B(n34280), .Z(n34282) );
  XOR U34222 ( .A(n34276), .B(n34119), .Z(n34278) );
  XOR U34223 ( .A(n34284), .B(n34285), .Z(n34119) );
  AND U34224 ( .A(n1231), .B(n34286), .Z(n34285) );
  XOR U34225 ( .A(n34287), .B(n34288), .Z(n34276) );
  AND U34226 ( .A(n34289), .B(n34290), .Z(n34288) );
  XNOR U34227 ( .A(n34287), .B(n34230), .Z(n34290) );
  XNOR U34228 ( .A(n34291), .B(n34292), .Z(n34230) );
  AND U34229 ( .A(n1223), .B(n34293), .Z(n34292) );
  XOR U34230 ( .A(n34294), .B(n34291), .Z(n34293) );
  XNOR U34231 ( .A(n34295), .B(n34287), .Z(n34289) );
  IV U34232 ( .A(n34131), .Z(n34295) );
  XOR U34233 ( .A(n34296), .B(n34297), .Z(n34131) );
  AND U34234 ( .A(n1231), .B(n34298), .Z(n34297) );
  AND U34235 ( .A(n34252), .B(n34241), .Z(n34287) );
  XNOR U34236 ( .A(n34299), .B(n34300), .Z(n34241) );
  AND U34237 ( .A(n1223), .B(n34301), .Z(n34300) );
  XNOR U34238 ( .A(n34302), .B(n34299), .Z(n34301) );
  XNOR U34239 ( .A(n34303), .B(n34304), .Z(n1223) );
  AND U34240 ( .A(n34305), .B(n34306), .Z(n34304) );
  XOR U34241 ( .A(n34262), .B(n34303), .Z(n34306) );
  AND U34242 ( .A(n34307), .B(n34308), .Z(n34262) );
  XOR U34243 ( .A(n34303), .B(n34259), .Z(n34305) );
  XNOR U34244 ( .A(n34309), .B(n34310), .Z(n34259) );
  AND U34245 ( .A(n1227), .B(n34265), .Z(n34310) );
  XOR U34246 ( .A(n34263), .B(n34309), .Z(n34265) );
  XOR U34247 ( .A(n34311), .B(n34312), .Z(n34303) );
  AND U34248 ( .A(n34313), .B(n34314), .Z(n34312) );
  XNOR U34249 ( .A(n34311), .B(n34307), .Z(n34314) );
  IV U34250 ( .A(n34271), .Z(n34307) );
  XOR U34251 ( .A(n34315), .B(n34316), .Z(n34271) );
  XOR U34252 ( .A(n34317), .B(n34308), .Z(n34316) );
  AND U34253 ( .A(n34283), .B(n34318), .Z(n34308) );
  AND U34254 ( .A(n34319), .B(n34320), .Z(n34317) );
  XOR U34255 ( .A(n34321), .B(n34315), .Z(n34319) );
  XNOR U34256 ( .A(n34268), .B(n34311), .Z(n34313) );
  XNOR U34257 ( .A(n34322), .B(n34323), .Z(n34268) );
  AND U34258 ( .A(n1227), .B(n34275), .Z(n34323) );
  XOR U34259 ( .A(n34322), .B(n34273), .Z(n34275) );
  XOR U34260 ( .A(n34324), .B(n34325), .Z(n34311) );
  AND U34261 ( .A(n34326), .B(n34327), .Z(n34325) );
  XNOR U34262 ( .A(n34324), .B(n34283), .Z(n34327) );
  XOR U34263 ( .A(n34328), .B(n34320), .Z(n34283) );
  XNOR U34264 ( .A(n34329), .B(n34315), .Z(n34320) );
  XOR U34265 ( .A(n34330), .B(n34331), .Z(n34315) );
  AND U34266 ( .A(n34332), .B(n34333), .Z(n34331) );
  XOR U34267 ( .A(n34334), .B(n34330), .Z(n34332) );
  XNOR U34268 ( .A(n34335), .B(n34336), .Z(n34329) );
  AND U34269 ( .A(n34337), .B(n34338), .Z(n34336) );
  XOR U34270 ( .A(n34335), .B(n34339), .Z(n34337) );
  XNOR U34271 ( .A(n34321), .B(n34318), .Z(n34328) );
  AND U34272 ( .A(n34340), .B(n34341), .Z(n34318) );
  XOR U34273 ( .A(n34342), .B(n34343), .Z(n34321) );
  AND U34274 ( .A(n34344), .B(n34345), .Z(n34343) );
  XOR U34275 ( .A(n34342), .B(n34346), .Z(n34344) );
  XNOR U34276 ( .A(n34280), .B(n34324), .Z(n34326) );
  XNOR U34277 ( .A(n34347), .B(n34348), .Z(n34280) );
  AND U34278 ( .A(n1227), .B(n34286), .Z(n34348) );
  XOR U34279 ( .A(n34347), .B(n34284), .Z(n34286) );
  XOR U34280 ( .A(n34349), .B(n34350), .Z(n34324) );
  AND U34281 ( .A(n34351), .B(n34352), .Z(n34350) );
  XNOR U34282 ( .A(n34349), .B(n34340), .Z(n34352) );
  IV U34283 ( .A(n34294), .Z(n34340) );
  XNOR U34284 ( .A(n34353), .B(n34333), .Z(n34294) );
  XNOR U34285 ( .A(n34354), .B(n34339), .Z(n34333) );
  XNOR U34286 ( .A(n34355), .B(n34356), .Z(n34339) );
  NOR U34287 ( .A(n34357), .B(n34358), .Z(n34356) );
  XOR U34288 ( .A(n34355), .B(n34359), .Z(n34357) );
  XNOR U34289 ( .A(n34338), .B(n34330), .Z(n34354) );
  XOR U34290 ( .A(n34360), .B(n34361), .Z(n34330) );
  AND U34291 ( .A(n34362), .B(n34363), .Z(n34361) );
  XOR U34292 ( .A(n34360), .B(n34364), .Z(n34362) );
  XNOR U34293 ( .A(n34365), .B(n34335), .Z(n34338) );
  XOR U34294 ( .A(n34366), .B(n34367), .Z(n34335) );
  AND U34295 ( .A(n34368), .B(n34369), .Z(n34367) );
  XNOR U34296 ( .A(n34370), .B(n34371), .Z(n34368) );
  IV U34297 ( .A(n34366), .Z(n34370) );
  XNOR U34298 ( .A(n34372), .B(n34373), .Z(n34365) );
  NOR U34299 ( .A(n34374), .B(n34375), .Z(n34373) );
  XNOR U34300 ( .A(n34372), .B(n34376), .Z(n34374) );
  XNOR U34301 ( .A(n34334), .B(n34341), .Z(n34353) );
  NOR U34302 ( .A(n34302), .B(n34377), .Z(n34341) );
  XOR U34303 ( .A(n34346), .B(n34345), .Z(n34334) );
  XNOR U34304 ( .A(n34378), .B(n34342), .Z(n34345) );
  XOR U34305 ( .A(n34379), .B(n34380), .Z(n34342) );
  AND U34306 ( .A(n34381), .B(n34382), .Z(n34380) );
  XNOR U34307 ( .A(n34383), .B(n34384), .Z(n34381) );
  IV U34308 ( .A(n34379), .Z(n34383) );
  XNOR U34309 ( .A(n34385), .B(n34386), .Z(n34378) );
  NOR U34310 ( .A(n34387), .B(n34388), .Z(n34386) );
  XNOR U34311 ( .A(n34385), .B(n34389), .Z(n34387) );
  XOR U34312 ( .A(n34390), .B(n34391), .Z(n34346) );
  NOR U34313 ( .A(n34392), .B(n34393), .Z(n34391) );
  XNOR U34314 ( .A(n34390), .B(n34394), .Z(n34392) );
  XNOR U34315 ( .A(n34291), .B(n34349), .Z(n34351) );
  XNOR U34316 ( .A(n34395), .B(n34396), .Z(n34291) );
  AND U34317 ( .A(n1227), .B(n34298), .Z(n34396) );
  XOR U34318 ( .A(n34395), .B(n34296), .Z(n34298) );
  AND U34319 ( .A(n34299), .B(n34302), .Z(n34349) );
  XOR U34320 ( .A(n34397), .B(n34377), .Z(n34302) );
  XNOR U34321 ( .A(p_input[1728]), .B(p_input[2048]), .Z(n34377) );
  XNOR U34322 ( .A(n34364), .B(n34363), .Z(n34397) );
  XNOR U34323 ( .A(n34398), .B(n34371), .Z(n34363) );
  XNOR U34324 ( .A(n34359), .B(n34358), .Z(n34371) );
  XNOR U34325 ( .A(n34399), .B(n34355), .Z(n34358) );
  XNOR U34326 ( .A(p_input[1738]), .B(p_input[2058]), .Z(n34355) );
  XOR U34327 ( .A(p_input[1739]), .B(n16732), .Z(n34399) );
  XOR U34328 ( .A(p_input[1740]), .B(p_input[2060]), .Z(n34359) );
  XOR U34329 ( .A(n34369), .B(n34400), .Z(n34398) );
  IV U34330 ( .A(n34360), .Z(n34400) );
  XOR U34331 ( .A(p_input[1729]), .B(p_input[2049]), .Z(n34360) );
  XNOR U34332 ( .A(n34401), .B(n34376), .Z(n34369) );
  XNOR U34333 ( .A(p_input[1743]), .B(n16735), .Z(n34376) );
  XOR U34334 ( .A(n34366), .B(n34375), .Z(n34401) );
  XOR U34335 ( .A(n34402), .B(n34372), .Z(n34375) );
  XOR U34336 ( .A(p_input[1741]), .B(p_input[2061]), .Z(n34372) );
  XOR U34337 ( .A(p_input[1742]), .B(n16737), .Z(n34402) );
  XOR U34338 ( .A(p_input[1737]), .B(p_input[2057]), .Z(n34366) );
  XOR U34339 ( .A(n34384), .B(n34382), .Z(n34364) );
  XNOR U34340 ( .A(n34403), .B(n34389), .Z(n34382) );
  XOR U34341 ( .A(p_input[1736]), .B(p_input[2056]), .Z(n34389) );
  XOR U34342 ( .A(n34379), .B(n34388), .Z(n34403) );
  XOR U34343 ( .A(n34404), .B(n34385), .Z(n34388) );
  XOR U34344 ( .A(p_input[1734]), .B(p_input[2054]), .Z(n34385) );
  XOR U34345 ( .A(p_input[1735]), .B(n17722), .Z(n34404) );
  XOR U34346 ( .A(p_input[1730]), .B(p_input[2050]), .Z(n34379) );
  XNOR U34347 ( .A(n34394), .B(n34393), .Z(n34384) );
  XOR U34348 ( .A(n34405), .B(n34390), .Z(n34393) );
  XOR U34349 ( .A(p_input[1731]), .B(p_input[2051]), .Z(n34390) );
  XOR U34350 ( .A(p_input[1732]), .B(n17724), .Z(n34405) );
  XOR U34351 ( .A(p_input[1733]), .B(p_input[2053]), .Z(n34394) );
  XNOR U34352 ( .A(n34406), .B(n34407), .Z(n34299) );
  AND U34353 ( .A(n1227), .B(n34408), .Z(n34407) );
  XNOR U34354 ( .A(n34409), .B(n34410), .Z(n1227) );
  AND U34355 ( .A(n34411), .B(n34412), .Z(n34410) );
  XOR U34356 ( .A(n34409), .B(n34309), .Z(n34412) );
  XNOR U34357 ( .A(n34409), .B(n34263), .Z(n34411) );
  XOR U34358 ( .A(n34413), .B(n34414), .Z(n34409) );
  AND U34359 ( .A(n34415), .B(n34416), .Z(n34414) );
  XOR U34360 ( .A(n34413), .B(n34273), .Z(n34415) );
  XOR U34361 ( .A(n34417), .B(n34418), .Z(n34252) );
  AND U34362 ( .A(n1231), .B(n34408), .Z(n34418) );
  XNOR U34363 ( .A(n34406), .B(n34417), .Z(n34408) );
  XNOR U34364 ( .A(n34419), .B(n34420), .Z(n1231) );
  AND U34365 ( .A(n34421), .B(n34422), .Z(n34420) );
  XNOR U34366 ( .A(n34423), .B(n34419), .Z(n34422) );
  IV U34367 ( .A(n34309), .Z(n34423) );
  XNOR U34368 ( .A(n34424), .B(n34425), .Z(n34309) );
  AND U34369 ( .A(n1234), .B(n34426), .Z(n34425) );
  XNOR U34370 ( .A(n34424), .B(n34427), .Z(n34426) );
  XNOR U34371 ( .A(n34263), .B(n34419), .Z(n34421) );
  XOR U34372 ( .A(n34428), .B(n34429), .Z(n34263) );
  AND U34373 ( .A(n1242), .B(n34430), .Z(n34429) );
  XOR U34374 ( .A(n34413), .B(n34431), .Z(n34419) );
  AND U34375 ( .A(n34432), .B(n34416), .Z(n34431) );
  XNOR U34376 ( .A(n34322), .B(n34413), .Z(n34416) );
  XNOR U34377 ( .A(n34433), .B(n34434), .Z(n34322) );
  AND U34378 ( .A(n1234), .B(n34435), .Z(n34434) );
  XOR U34379 ( .A(n34436), .B(n34433), .Z(n34435) );
  XNOR U34380 ( .A(n34437), .B(n34413), .Z(n34432) );
  IV U34381 ( .A(n34273), .Z(n34437) );
  XOR U34382 ( .A(n34438), .B(n34439), .Z(n34273) );
  AND U34383 ( .A(n1242), .B(n34440), .Z(n34439) );
  XOR U34384 ( .A(n34441), .B(n34442), .Z(n34413) );
  AND U34385 ( .A(n34443), .B(n34444), .Z(n34442) );
  XNOR U34386 ( .A(n34347), .B(n34441), .Z(n34444) );
  XNOR U34387 ( .A(n34445), .B(n34446), .Z(n34347) );
  AND U34388 ( .A(n1234), .B(n34447), .Z(n34446) );
  XNOR U34389 ( .A(n34448), .B(n34445), .Z(n34447) );
  XOR U34390 ( .A(n34441), .B(n34284), .Z(n34443) );
  XOR U34391 ( .A(n34449), .B(n34450), .Z(n34284) );
  AND U34392 ( .A(n1242), .B(n34451), .Z(n34450) );
  XOR U34393 ( .A(n34452), .B(n34453), .Z(n34441) );
  AND U34394 ( .A(n34454), .B(n34455), .Z(n34453) );
  XNOR U34395 ( .A(n34452), .B(n34395), .Z(n34455) );
  XNOR U34396 ( .A(n34456), .B(n34457), .Z(n34395) );
  AND U34397 ( .A(n1234), .B(n34458), .Z(n34457) );
  XOR U34398 ( .A(n34459), .B(n34456), .Z(n34458) );
  XNOR U34399 ( .A(n34460), .B(n34452), .Z(n34454) );
  IV U34400 ( .A(n34296), .Z(n34460) );
  XOR U34401 ( .A(n34461), .B(n34462), .Z(n34296) );
  AND U34402 ( .A(n1242), .B(n34463), .Z(n34462) );
  AND U34403 ( .A(n34417), .B(n34406), .Z(n34452) );
  XNOR U34404 ( .A(n34464), .B(n34465), .Z(n34406) );
  AND U34405 ( .A(n1234), .B(n34466), .Z(n34465) );
  XNOR U34406 ( .A(n34467), .B(n34464), .Z(n34466) );
  XNOR U34407 ( .A(n34468), .B(n34469), .Z(n1234) );
  AND U34408 ( .A(n34470), .B(n34471), .Z(n34469) );
  XOR U34409 ( .A(n34427), .B(n34468), .Z(n34471) );
  AND U34410 ( .A(n34472), .B(n34473), .Z(n34427) );
  XOR U34411 ( .A(n34468), .B(n34424), .Z(n34470) );
  XNOR U34412 ( .A(n34474), .B(n34475), .Z(n34424) );
  AND U34413 ( .A(n1238), .B(n34430), .Z(n34475) );
  XOR U34414 ( .A(n34428), .B(n34474), .Z(n34430) );
  XOR U34415 ( .A(n34476), .B(n34477), .Z(n34468) );
  AND U34416 ( .A(n34478), .B(n34479), .Z(n34477) );
  XNOR U34417 ( .A(n34476), .B(n34472), .Z(n34479) );
  IV U34418 ( .A(n34436), .Z(n34472) );
  XOR U34419 ( .A(n34480), .B(n34481), .Z(n34436) );
  XOR U34420 ( .A(n34482), .B(n34473), .Z(n34481) );
  AND U34421 ( .A(n34448), .B(n34483), .Z(n34473) );
  AND U34422 ( .A(n34484), .B(n34485), .Z(n34482) );
  XOR U34423 ( .A(n34486), .B(n34480), .Z(n34484) );
  XNOR U34424 ( .A(n34433), .B(n34476), .Z(n34478) );
  XNOR U34425 ( .A(n34487), .B(n34488), .Z(n34433) );
  AND U34426 ( .A(n1238), .B(n34440), .Z(n34488) );
  XOR U34427 ( .A(n34487), .B(n34438), .Z(n34440) );
  XOR U34428 ( .A(n34489), .B(n34490), .Z(n34476) );
  AND U34429 ( .A(n34491), .B(n34492), .Z(n34490) );
  XNOR U34430 ( .A(n34489), .B(n34448), .Z(n34492) );
  XOR U34431 ( .A(n34493), .B(n34485), .Z(n34448) );
  XNOR U34432 ( .A(n34494), .B(n34480), .Z(n34485) );
  XOR U34433 ( .A(n34495), .B(n34496), .Z(n34480) );
  AND U34434 ( .A(n34497), .B(n34498), .Z(n34496) );
  XOR U34435 ( .A(n34499), .B(n34495), .Z(n34497) );
  XNOR U34436 ( .A(n34500), .B(n34501), .Z(n34494) );
  AND U34437 ( .A(n34502), .B(n34503), .Z(n34501) );
  XOR U34438 ( .A(n34500), .B(n34504), .Z(n34502) );
  XNOR U34439 ( .A(n34486), .B(n34483), .Z(n34493) );
  AND U34440 ( .A(n34505), .B(n34506), .Z(n34483) );
  XOR U34441 ( .A(n34507), .B(n34508), .Z(n34486) );
  AND U34442 ( .A(n34509), .B(n34510), .Z(n34508) );
  XOR U34443 ( .A(n34507), .B(n34511), .Z(n34509) );
  XNOR U34444 ( .A(n34445), .B(n34489), .Z(n34491) );
  XNOR U34445 ( .A(n34512), .B(n34513), .Z(n34445) );
  AND U34446 ( .A(n1238), .B(n34451), .Z(n34513) );
  XOR U34447 ( .A(n34512), .B(n34449), .Z(n34451) );
  XOR U34448 ( .A(n34514), .B(n34515), .Z(n34489) );
  AND U34449 ( .A(n34516), .B(n34517), .Z(n34515) );
  XNOR U34450 ( .A(n34514), .B(n34505), .Z(n34517) );
  IV U34451 ( .A(n34459), .Z(n34505) );
  XNOR U34452 ( .A(n34518), .B(n34498), .Z(n34459) );
  XNOR U34453 ( .A(n34519), .B(n34504), .Z(n34498) );
  XNOR U34454 ( .A(n34520), .B(n34521), .Z(n34504) );
  NOR U34455 ( .A(n34522), .B(n34523), .Z(n34521) );
  XOR U34456 ( .A(n34520), .B(n34524), .Z(n34522) );
  XNOR U34457 ( .A(n34503), .B(n34495), .Z(n34519) );
  XOR U34458 ( .A(n34525), .B(n34526), .Z(n34495) );
  AND U34459 ( .A(n34527), .B(n34528), .Z(n34526) );
  XOR U34460 ( .A(n34525), .B(n34529), .Z(n34527) );
  XNOR U34461 ( .A(n34530), .B(n34500), .Z(n34503) );
  XOR U34462 ( .A(n34531), .B(n34532), .Z(n34500) );
  AND U34463 ( .A(n34533), .B(n34534), .Z(n34532) );
  XNOR U34464 ( .A(n34535), .B(n34536), .Z(n34533) );
  IV U34465 ( .A(n34531), .Z(n34535) );
  XNOR U34466 ( .A(n34537), .B(n34538), .Z(n34530) );
  NOR U34467 ( .A(n34539), .B(n34540), .Z(n34538) );
  XNOR U34468 ( .A(n34537), .B(n34541), .Z(n34539) );
  XNOR U34469 ( .A(n34499), .B(n34506), .Z(n34518) );
  NOR U34470 ( .A(n34467), .B(n34542), .Z(n34506) );
  XOR U34471 ( .A(n34511), .B(n34510), .Z(n34499) );
  XNOR U34472 ( .A(n34543), .B(n34507), .Z(n34510) );
  XOR U34473 ( .A(n34544), .B(n34545), .Z(n34507) );
  AND U34474 ( .A(n34546), .B(n34547), .Z(n34545) );
  XNOR U34475 ( .A(n34548), .B(n34549), .Z(n34546) );
  IV U34476 ( .A(n34544), .Z(n34548) );
  XNOR U34477 ( .A(n34550), .B(n34551), .Z(n34543) );
  NOR U34478 ( .A(n34552), .B(n34553), .Z(n34551) );
  XNOR U34479 ( .A(n34550), .B(n34554), .Z(n34552) );
  XOR U34480 ( .A(n34555), .B(n34556), .Z(n34511) );
  NOR U34481 ( .A(n34557), .B(n34558), .Z(n34556) );
  XNOR U34482 ( .A(n34555), .B(n34559), .Z(n34557) );
  XNOR U34483 ( .A(n34456), .B(n34514), .Z(n34516) );
  XNOR U34484 ( .A(n34560), .B(n34561), .Z(n34456) );
  AND U34485 ( .A(n1238), .B(n34463), .Z(n34561) );
  XOR U34486 ( .A(n34560), .B(n34461), .Z(n34463) );
  AND U34487 ( .A(n34464), .B(n34467), .Z(n34514) );
  XOR U34488 ( .A(n34562), .B(n34542), .Z(n34467) );
  XNOR U34489 ( .A(p_input[1744]), .B(p_input[2048]), .Z(n34542) );
  XNOR U34490 ( .A(n34529), .B(n34528), .Z(n34562) );
  XNOR U34491 ( .A(n34563), .B(n34536), .Z(n34528) );
  XNOR U34492 ( .A(n34524), .B(n34523), .Z(n34536) );
  XNOR U34493 ( .A(n34564), .B(n34520), .Z(n34523) );
  XNOR U34494 ( .A(p_input[1754]), .B(p_input[2058]), .Z(n34520) );
  XOR U34495 ( .A(p_input[1755]), .B(n16732), .Z(n34564) );
  XOR U34496 ( .A(p_input[1756]), .B(p_input[2060]), .Z(n34524) );
  XOR U34497 ( .A(n34534), .B(n34565), .Z(n34563) );
  IV U34498 ( .A(n34525), .Z(n34565) );
  XOR U34499 ( .A(p_input[1745]), .B(p_input[2049]), .Z(n34525) );
  XNOR U34500 ( .A(n34566), .B(n34541), .Z(n34534) );
  XNOR U34501 ( .A(p_input[1759]), .B(n16735), .Z(n34541) );
  XOR U34502 ( .A(n34531), .B(n34540), .Z(n34566) );
  XOR U34503 ( .A(n34567), .B(n34537), .Z(n34540) );
  XOR U34504 ( .A(p_input[1757]), .B(p_input[2061]), .Z(n34537) );
  XOR U34505 ( .A(p_input[1758]), .B(n16737), .Z(n34567) );
  XOR U34506 ( .A(p_input[1753]), .B(p_input[2057]), .Z(n34531) );
  XOR U34507 ( .A(n34549), .B(n34547), .Z(n34529) );
  XNOR U34508 ( .A(n34568), .B(n34554), .Z(n34547) );
  XOR U34509 ( .A(p_input[1752]), .B(p_input[2056]), .Z(n34554) );
  XOR U34510 ( .A(n34544), .B(n34553), .Z(n34568) );
  XOR U34511 ( .A(n34569), .B(n34550), .Z(n34553) );
  XOR U34512 ( .A(p_input[1750]), .B(p_input[2054]), .Z(n34550) );
  XOR U34513 ( .A(p_input[1751]), .B(n17722), .Z(n34569) );
  XOR U34514 ( .A(p_input[1746]), .B(p_input[2050]), .Z(n34544) );
  XNOR U34515 ( .A(n34559), .B(n34558), .Z(n34549) );
  XOR U34516 ( .A(n34570), .B(n34555), .Z(n34558) );
  XOR U34517 ( .A(p_input[1747]), .B(p_input[2051]), .Z(n34555) );
  XOR U34518 ( .A(p_input[1748]), .B(n17724), .Z(n34570) );
  XOR U34519 ( .A(p_input[1749]), .B(p_input[2053]), .Z(n34559) );
  XNOR U34520 ( .A(n34571), .B(n34572), .Z(n34464) );
  AND U34521 ( .A(n1238), .B(n34573), .Z(n34572) );
  XNOR U34522 ( .A(n34574), .B(n34575), .Z(n1238) );
  AND U34523 ( .A(n34576), .B(n34577), .Z(n34575) );
  XOR U34524 ( .A(n34574), .B(n34474), .Z(n34577) );
  XNOR U34525 ( .A(n34574), .B(n34428), .Z(n34576) );
  XOR U34526 ( .A(n34578), .B(n34579), .Z(n34574) );
  AND U34527 ( .A(n34580), .B(n34581), .Z(n34579) );
  XOR U34528 ( .A(n34578), .B(n34438), .Z(n34580) );
  XOR U34529 ( .A(n34582), .B(n34583), .Z(n34417) );
  AND U34530 ( .A(n1242), .B(n34573), .Z(n34583) );
  XNOR U34531 ( .A(n34571), .B(n34582), .Z(n34573) );
  XNOR U34532 ( .A(n34584), .B(n34585), .Z(n1242) );
  AND U34533 ( .A(n34586), .B(n34587), .Z(n34585) );
  XNOR U34534 ( .A(n34588), .B(n34584), .Z(n34587) );
  IV U34535 ( .A(n34474), .Z(n34588) );
  XNOR U34536 ( .A(n34589), .B(n34590), .Z(n34474) );
  AND U34537 ( .A(n1245), .B(n34591), .Z(n34590) );
  XNOR U34538 ( .A(n34589), .B(n34592), .Z(n34591) );
  XNOR U34539 ( .A(n34428), .B(n34584), .Z(n34586) );
  XOR U34540 ( .A(n34593), .B(n34594), .Z(n34428) );
  AND U34541 ( .A(n1253), .B(n34595), .Z(n34594) );
  XOR U34542 ( .A(n34578), .B(n34596), .Z(n34584) );
  AND U34543 ( .A(n34597), .B(n34581), .Z(n34596) );
  XNOR U34544 ( .A(n34487), .B(n34578), .Z(n34581) );
  XNOR U34545 ( .A(n34598), .B(n34599), .Z(n34487) );
  AND U34546 ( .A(n1245), .B(n34600), .Z(n34599) );
  XOR U34547 ( .A(n34601), .B(n34598), .Z(n34600) );
  XNOR U34548 ( .A(n34602), .B(n34578), .Z(n34597) );
  IV U34549 ( .A(n34438), .Z(n34602) );
  XOR U34550 ( .A(n34603), .B(n34604), .Z(n34438) );
  AND U34551 ( .A(n1253), .B(n34605), .Z(n34604) );
  XOR U34552 ( .A(n34606), .B(n34607), .Z(n34578) );
  AND U34553 ( .A(n34608), .B(n34609), .Z(n34607) );
  XNOR U34554 ( .A(n34512), .B(n34606), .Z(n34609) );
  XNOR U34555 ( .A(n34610), .B(n34611), .Z(n34512) );
  AND U34556 ( .A(n1245), .B(n34612), .Z(n34611) );
  XNOR U34557 ( .A(n34613), .B(n34610), .Z(n34612) );
  XOR U34558 ( .A(n34606), .B(n34449), .Z(n34608) );
  XOR U34559 ( .A(n34614), .B(n34615), .Z(n34449) );
  AND U34560 ( .A(n1253), .B(n34616), .Z(n34615) );
  XOR U34561 ( .A(n34617), .B(n34618), .Z(n34606) );
  AND U34562 ( .A(n34619), .B(n34620), .Z(n34618) );
  XNOR U34563 ( .A(n34617), .B(n34560), .Z(n34620) );
  XNOR U34564 ( .A(n34621), .B(n34622), .Z(n34560) );
  AND U34565 ( .A(n1245), .B(n34623), .Z(n34622) );
  XOR U34566 ( .A(n34624), .B(n34621), .Z(n34623) );
  XNOR U34567 ( .A(n34625), .B(n34617), .Z(n34619) );
  IV U34568 ( .A(n34461), .Z(n34625) );
  XOR U34569 ( .A(n34626), .B(n34627), .Z(n34461) );
  AND U34570 ( .A(n1253), .B(n34628), .Z(n34627) );
  AND U34571 ( .A(n34582), .B(n34571), .Z(n34617) );
  XNOR U34572 ( .A(n34629), .B(n34630), .Z(n34571) );
  AND U34573 ( .A(n1245), .B(n34631), .Z(n34630) );
  XNOR U34574 ( .A(n34632), .B(n34629), .Z(n34631) );
  XNOR U34575 ( .A(n34633), .B(n34634), .Z(n1245) );
  AND U34576 ( .A(n34635), .B(n34636), .Z(n34634) );
  XOR U34577 ( .A(n34592), .B(n34633), .Z(n34636) );
  AND U34578 ( .A(n34637), .B(n34638), .Z(n34592) );
  XOR U34579 ( .A(n34633), .B(n34589), .Z(n34635) );
  XNOR U34580 ( .A(n34639), .B(n34640), .Z(n34589) );
  AND U34581 ( .A(n1249), .B(n34595), .Z(n34640) );
  XOR U34582 ( .A(n34593), .B(n34639), .Z(n34595) );
  XOR U34583 ( .A(n34641), .B(n34642), .Z(n34633) );
  AND U34584 ( .A(n34643), .B(n34644), .Z(n34642) );
  XNOR U34585 ( .A(n34641), .B(n34637), .Z(n34644) );
  IV U34586 ( .A(n34601), .Z(n34637) );
  XOR U34587 ( .A(n34645), .B(n34646), .Z(n34601) );
  XOR U34588 ( .A(n34647), .B(n34638), .Z(n34646) );
  AND U34589 ( .A(n34613), .B(n34648), .Z(n34638) );
  AND U34590 ( .A(n34649), .B(n34650), .Z(n34647) );
  XOR U34591 ( .A(n34651), .B(n34645), .Z(n34649) );
  XNOR U34592 ( .A(n34598), .B(n34641), .Z(n34643) );
  XNOR U34593 ( .A(n34652), .B(n34653), .Z(n34598) );
  AND U34594 ( .A(n1249), .B(n34605), .Z(n34653) );
  XOR U34595 ( .A(n34652), .B(n34603), .Z(n34605) );
  XOR U34596 ( .A(n34654), .B(n34655), .Z(n34641) );
  AND U34597 ( .A(n34656), .B(n34657), .Z(n34655) );
  XNOR U34598 ( .A(n34654), .B(n34613), .Z(n34657) );
  XOR U34599 ( .A(n34658), .B(n34650), .Z(n34613) );
  XNOR U34600 ( .A(n34659), .B(n34645), .Z(n34650) );
  XOR U34601 ( .A(n34660), .B(n34661), .Z(n34645) );
  AND U34602 ( .A(n34662), .B(n34663), .Z(n34661) );
  XOR U34603 ( .A(n34664), .B(n34660), .Z(n34662) );
  XNOR U34604 ( .A(n34665), .B(n34666), .Z(n34659) );
  AND U34605 ( .A(n34667), .B(n34668), .Z(n34666) );
  XOR U34606 ( .A(n34665), .B(n34669), .Z(n34667) );
  XNOR U34607 ( .A(n34651), .B(n34648), .Z(n34658) );
  AND U34608 ( .A(n34670), .B(n34671), .Z(n34648) );
  XOR U34609 ( .A(n34672), .B(n34673), .Z(n34651) );
  AND U34610 ( .A(n34674), .B(n34675), .Z(n34673) );
  XOR U34611 ( .A(n34672), .B(n34676), .Z(n34674) );
  XNOR U34612 ( .A(n34610), .B(n34654), .Z(n34656) );
  XNOR U34613 ( .A(n34677), .B(n34678), .Z(n34610) );
  AND U34614 ( .A(n1249), .B(n34616), .Z(n34678) );
  XOR U34615 ( .A(n34677), .B(n34614), .Z(n34616) );
  XOR U34616 ( .A(n34679), .B(n34680), .Z(n34654) );
  AND U34617 ( .A(n34681), .B(n34682), .Z(n34680) );
  XNOR U34618 ( .A(n34679), .B(n34670), .Z(n34682) );
  IV U34619 ( .A(n34624), .Z(n34670) );
  XNOR U34620 ( .A(n34683), .B(n34663), .Z(n34624) );
  XNOR U34621 ( .A(n34684), .B(n34669), .Z(n34663) );
  XNOR U34622 ( .A(n34685), .B(n34686), .Z(n34669) );
  NOR U34623 ( .A(n34687), .B(n34688), .Z(n34686) );
  XOR U34624 ( .A(n34685), .B(n34689), .Z(n34687) );
  XNOR U34625 ( .A(n34668), .B(n34660), .Z(n34684) );
  XOR U34626 ( .A(n34690), .B(n34691), .Z(n34660) );
  AND U34627 ( .A(n34692), .B(n34693), .Z(n34691) );
  XOR U34628 ( .A(n34690), .B(n34694), .Z(n34692) );
  XNOR U34629 ( .A(n34695), .B(n34665), .Z(n34668) );
  XOR U34630 ( .A(n34696), .B(n34697), .Z(n34665) );
  AND U34631 ( .A(n34698), .B(n34699), .Z(n34697) );
  XNOR U34632 ( .A(n34700), .B(n34701), .Z(n34698) );
  IV U34633 ( .A(n34696), .Z(n34700) );
  XNOR U34634 ( .A(n34702), .B(n34703), .Z(n34695) );
  NOR U34635 ( .A(n34704), .B(n34705), .Z(n34703) );
  XNOR U34636 ( .A(n34702), .B(n34706), .Z(n34704) );
  XNOR U34637 ( .A(n34664), .B(n34671), .Z(n34683) );
  NOR U34638 ( .A(n34632), .B(n34707), .Z(n34671) );
  XOR U34639 ( .A(n34676), .B(n34675), .Z(n34664) );
  XNOR U34640 ( .A(n34708), .B(n34672), .Z(n34675) );
  XOR U34641 ( .A(n34709), .B(n34710), .Z(n34672) );
  AND U34642 ( .A(n34711), .B(n34712), .Z(n34710) );
  XNOR U34643 ( .A(n34713), .B(n34714), .Z(n34711) );
  IV U34644 ( .A(n34709), .Z(n34713) );
  XNOR U34645 ( .A(n34715), .B(n34716), .Z(n34708) );
  NOR U34646 ( .A(n34717), .B(n34718), .Z(n34716) );
  XNOR U34647 ( .A(n34715), .B(n34719), .Z(n34717) );
  XOR U34648 ( .A(n34720), .B(n34721), .Z(n34676) );
  NOR U34649 ( .A(n34722), .B(n34723), .Z(n34721) );
  XNOR U34650 ( .A(n34720), .B(n34724), .Z(n34722) );
  XNOR U34651 ( .A(n34621), .B(n34679), .Z(n34681) );
  XNOR U34652 ( .A(n34725), .B(n34726), .Z(n34621) );
  AND U34653 ( .A(n1249), .B(n34628), .Z(n34726) );
  XOR U34654 ( .A(n34725), .B(n34626), .Z(n34628) );
  AND U34655 ( .A(n34629), .B(n34632), .Z(n34679) );
  XOR U34656 ( .A(n34727), .B(n34707), .Z(n34632) );
  XNOR U34657 ( .A(p_input[1760]), .B(p_input[2048]), .Z(n34707) );
  XNOR U34658 ( .A(n34694), .B(n34693), .Z(n34727) );
  XNOR U34659 ( .A(n34728), .B(n34701), .Z(n34693) );
  XNOR U34660 ( .A(n34689), .B(n34688), .Z(n34701) );
  XNOR U34661 ( .A(n34729), .B(n34685), .Z(n34688) );
  XNOR U34662 ( .A(p_input[1770]), .B(p_input[2058]), .Z(n34685) );
  XOR U34663 ( .A(p_input[1771]), .B(n16732), .Z(n34729) );
  XOR U34664 ( .A(p_input[1772]), .B(p_input[2060]), .Z(n34689) );
  XOR U34665 ( .A(n34699), .B(n34730), .Z(n34728) );
  IV U34666 ( .A(n34690), .Z(n34730) );
  XOR U34667 ( .A(p_input[1761]), .B(p_input[2049]), .Z(n34690) );
  XNOR U34668 ( .A(n34731), .B(n34706), .Z(n34699) );
  XNOR U34669 ( .A(p_input[1775]), .B(n16735), .Z(n34706) );
  XOR U34670 ( .A(n34696), .B(n34705), .Z(n34731) );
  XOR U34671 ( .A(n34732), .B(n34702), .Z(n34705) );
  XOR U34672 ( .A(p_input[1773]), .B(p_input[2061]), .Z(n34702) );
  XOR U34673 ( .A(p_input[1774]), .B(n16737), .Z(n34732) );
  XOR U34674 ( .A(p_input[1769]), .B(p_input[2057]), .Z(n34696) );
  XOR U34675 ( .A(n34714), .B(n34712), .Z(n34694) );
  XNOR U34676 ( .A(n34733), .B(n34719), .Z(n34712) );
  XOR U34677 ( .A(p_input[1768]), .B(p_input[2056]), .Z(n34719) );
  XOR U34678 ( .A(n34709), .B(n34718), .Z(n34733) );
  XOR U34679 ( .A(n34734), .B(n34715), .Z(n34718) );
  XOR U34680 ( .A(p_input[1766]), .B(p_input[2054]), .Z(n34715) );
  XOR U34681 ( .A(p_input[1767]), .B(n17722), .Z(n34734) );
  XOR U34682 ( .A(p_input[1762]), .B(p_input[2050]), .Z(n34709) );
  XNOR U34683 ( .A(n34724), .B(n34723), .Z(n34714) );
  XOR U34684 ( .A(n34735), .B(n34720), .Z(n34723) );
  XOR U34685 ( .A(p_input[1763]), .B(p_input[2051]), .Z(n34720) );
  XOR U34686 ( .A(p_input[1764]), .B(n17724), .Z(n34735) );
  XOR U34687 ( .A(p_input[1765]), .B(p_input[2053]), .Z(n34724) );
  XNOR U34688 ( .A(n34736), .B(n34737), .Z(n34629) );
  AND U34689 ( .A(n1249), .B(n34738), .Z(n34737) );
  XNOR U34690 ( .A(n34739), .B(n34740), .Z(n1249) );
  AND U34691 ( .A(n34741), .B(n34742), .Z(n34740) );
  XOR U34692 ( .A(n34739), .B(n34639), .Z(n34742) );
  XNOR U34693 ( .A(n34739), .B(n34593), .Z(n34741) );
  XOR U34694 ( .A(n34743), .B(n34744), .Z(n34739) );
  AND U34695 ( .A(n34745), .B(n34746), .Z(n34744) );
  XOR U34696 ( .A(n34743), .B(n34603), .Z(n34745) );
  XOR U34697 ( .A(n34747), .B(n34748), .Z(n34582) );
  AND U34698 ( .A(n1253), .B(n34738), .Z(n34748) );
  XNOR U34699 ( .A(n34736), .B(n34747), .Z(n34738) );
  XNOR U34700 ( .A(n34749), .B(n34750), .Z(n1253) );
  AND U34701 ( .A(n34751), .B(n34752), .Z(n34750) );
  XNOR U34702 ( .A(n34753), .B(n34749), .Z(n34752) );
  IV U34703 ( .A(n34639), .Z(n34753) );
  XNOR U34704 ( .A(n34754), .B(n34755), .Z(n34639) );
  AND U34705 ( .A(n1256), .B(n34756), .Z(n34755) );
  XNOR U34706 ( .A(n34754), .B(n34757), .Z(n34756) );
  XNOR U34707 ( .A(n34593), .B(n34749), .Z(n34751) );
  XOR U34708 ( .A(n34758), .B(n34759), .Z(n34593) );
  AND U34709 ( .A(n1264), .B(n34760), .Z(n34759) );
  XOR U34710 ( .A(n34743), .B(n34761), .Z(n34749) );
  AND U34711 ( .A(n34762), .B(n34746), .Z(n34761) );
  XNOR U34712 ( .A(n34652), .B(n34743), .Z(n34746) );
  XNOR U34713 ( .A(n34763), .B(n34764), .Z(n34652) );
  AND U34714 ( .A(n1256), .B(n34765), .Z(n34764) );
  XOR U34715 ( .A(n34766), .B(n34763), .Z(n34765) );
  XNOR U34716 ( .A(n34767), .B(n34743), .Z(n34762) );
  IV U34717 ( .A(n34603), .Z(n34767) );
  XOR U34718 ( .A(n34768), .B(n34769), .Z(n34603) );
  AND U34719 ( .A(n1264), .B(n34770), .Z(n34769) );
  XOR U34720 ( .A(n34771), .B(n34772), .Z(n34743) );
  AND U34721 ( .A(n34773), .B(n34774), .Z(n34772) );
  XNOR U34722 ( .A(n34677), .B(n34771), .Z(n34774) );
  XNOR U34723 ( .A(n34775), .B(n34776), .Z(n34677) );
  AND U34724 ( .A(n1256), .B(n34777), .Z(n34776) );
  XNOR U34725 ( .A(n34778), .B(n34775), .Z(n34777) );
  XOR U34726 ( .A(n34771), .B(n34614), .Z(n34773) );
  XOR U34727 ( .A(n34779), .B(n34780), .Z(n34614) );
  AND U34728 ( .A(n1264), .B(n34781), .Z(n34780) );
  XOR U34729 ( .A(n34782), .B(n34783), .Z(n34771) );
  AND U34730 ( .A(n34784), .B(n34785), .Z(n34783) );
  XNOR U34731 ( .A(n34782), .B(n34725), .Z(n34785) );
  XNOR U34732 ( .A(n34786), .B(n34787), .Z(n34725) );
  AND U34733 ( .A(n1256), .B(n34788), .Z(n34787) );
  XOR U34734 ( .A(n34789), .B(n34786), .Z(n34788) );
  XNOR U34735 ( .A(n34790), .B(n34782), .Z(n34784) );
  IV U34736 ( .A(n34626), .Z(n34790) );
  XOR U34737 ( .A(n34791), .B(n34792), .Z(n34626) );
  AND U34738 ( .A(n1264), .B(n34793), .Z(n34792) );
  AND U34739 ( .A(n34747), .B(n34736), .Z(n34782) );
  XNOR U34740 ( .A(n34794), .B(n34795), .Z(n34736) );
  AND U34741 ( .A(n1256), .B(n34796), .Z(n34795) );
  XNOR U34742 ( .A(n34797), .B(n34794), .Z(n34796) );
  XNOR U34743 ( .A(n34798), .B(n34799), .Z(n1256) );
  AND U34744 ( .A(n34800), .B(n34801), .Z(n34799) );
  XOR U34745 ( .A(n34757), .B(n34798), .Z(n34801) );
  AND U34746 ( .A(n34802), .B(n34803), .Z(n34757) );
  XOR U34747 ( .A(n34798), .B(n34754), .Z(n34800) );
  XNOR U34748 ( .A(n34804), .B(n34805), .Z(n34754) );
  AND U34749 ( .A(n1260), .B(n34760), .Z(n34805) );
  XOR U34750 ( .A(n34758), .B(n34804), .Z(n34760) );
  XOR U34751 ( .A(n34806), .B(n34807), .Z(n34798) );
  AND U34752 ( .A(n34808), .B(n34809), .Z(n34807) );
  XNOR U34753 ( .A(n34806), .B(n34802), .Z(n34809) );
  IV U34754 ( .A(n34766), .Z(n34802) );
  XOR U34755 ( .A(n34810), .B(n34811), .Z(n34766) );
  XOR U34756 ( .A(n34812), .B(n34803), .Z(n34811) );
  AND U34757 ( .A(n34778), .B(n34813), .Z(n34803) );
  AND U34758 ( .A(n34814), .B(n34815), .Z(n34812) );
  XOR U34759 ( .A(n34816), .B(n34810), .Z(n34814) );
  XNOR U34760 ( .A(n34763), .B(n34806), .Z(n34808) );
  XNOR U34761 ( .A(n34817), .B(n34818), .Z(n34763) );
  AND U34762 ( .A(n1260), .B(n34770), .Z(n34818) );
  XOR U34763 ( .A(n34817), .B(n34768), .Z(n34770) );
  XOR U34764 ( .A(n34819), .B(n34820), .Z(n34806) );
  AND U34765 ( .A(n34821), .B(n34822), .Z(n34820) );
  XNOR U34766 ( .A(n34819), .B(n34778), .Z(n34822) );
  XOR U34767 ( .A(n34823), .B(n34815), .Z(n34778) );
  XNOR U34768 ( .A(n34824), .B(n34810), .Z(n34815) );
  XOR U34769 ( .A(n34825), .B(n34826), .Z(n34810) );
  AND U34770 ( .A(n34827), .B(n34828), .Z(n34826) );
  XOR U34771 ( .A(n34829), .B(n34825), .Z(n34827) );
  XNOR U34772 ( .A(n34830), .B(n34831), .Z(n34824) );
  AND U34773 ( .A(n34832), .B(n34833), .Z(n34831) );
  XOR U34774 ( .A(n34830), .B(n34834), .Z(n34832) );
  XNOR U34775 ( .A(n34816), .B(n34813), .Z(n34823) );
  AND U34776 ( .A(n34835), .B(n34836), .Z(n34813) );
  XOR U34777 ( .A(n34837), .B(n34838), .Z(n34816) );
  AND U34778 ( .A(n34839), .B(n34840), .Z(n34838) );
  XOR U34779 ( .A(n34837), .B(n34841), .Z(n34839) );
  XNOR U34780 ( .A(n34775), .B(n34819), .Z(n34821) );
  XNOR U34781 ( .A(n34842), .B(n34843), .Z(n34775) );
  AND U34782 ( .A(n1260), .B(n34781), .Z(n34843) );
  XOR U34783 ( .A(n34842), .B(n34779), .Z(n34781) );
  XOR U34784 ( .A(n34844), .B(n34845), .Z(n34819) );
  AND U34785 ( .A(n34846), .B(n34847), .Z(n34845) );
  XNOR U34786 ( .A(n34844), .B(n34835), .Z(n34847) );
  IV U34787 ( .A(n34789), .Z(n34835) );
  XNOR U34788 ( .A(n34848), .B(n34828), .Z(n34789) );
  XNOR U34789 ( .A(n34849), .B(n34834), .Z(n34828) );
  XNOR U34790 ( .A(n34850), .B(n34851), .Z(n34834) );
  NOR U34791 ( .A(n34852), .B(n34853), .Z(n34851) );
  XOR U34792 ( .A(n34850), .B(n34854), .Z(n34852) );
  XNOR U34793 ( .A(n34833), .B(n34825), .Z(n34849) );
  XOR U34794 ( .A(n34855), .B(n34856), .Z(n34825) );
  AND U34795 ( .A(n34857), .B(n34858), .Z(n34856) );
  XOR U34796 ( .A(n34855), .B(n34859), .Z(n34857) );
  XNOR U34797 ( .A(n34860), .B(n34830), .Z(n34833) );
  XOR U34798 ( .A(n34861), .B(n34862), .Z(n34830) );
  AND U34799 ( .A(n34863), .B(n34864), .Z(n34862) );
  XNOR U34800 ( .A(n34865), .B(n34866), .Z(n34863) );
  IV U34801 ( .A(n34861), .Z(n34865) );
  XNOR U34802 ( .A(n34867), .B(n34868), .Z(n34860) );
  NOR U34803 ( .A(n34869), .B(n34870), .Z(n34868) );
  XNOR U34804 ( .A(n34867), .B(n34871), .Z(n34869) );
  XNOR U34805 ( .A(n34829), .B(n34836), .Z(n34848) );
  NOR U34806 ( .A(n34797), .B(n34872), .Z(n34836) );
  XOR U34807 ( .A(n34841), .B(n34840), .Z(n34829) );
  XNOR U34808 ( .A(n34873), .B(n34837), .Z(n34840) );
  XOR U34809 ( .A(n34874), .B(n34875), .Z(n34837) );
  AND U34810 ( .A(n34876), .B(n34877), .Z(n34875) );
  XNOR U34811 ( .A(n34878), .B(n34879), .Z(n34876) );
  IV U34812 ( .A(n34874), .Z(n34878) );
  XNOR U34813 ( .A(n34880), .B(n34881), .Z(n34873) );
  NOR U34814 ( .A(n34882), .B(n34883), .Z(n34881) );
  XNOR U34815 ( .A(n34880), .B(n34884), .Z(n34882) );
  XOR U34816 ( .A(n34885), .B(n34886), .Z(n34841) );
  NOR U34817 ( .A(n34887), .B(n34888), .Z(n34886) );
  XNOR U34818 ( .A(n34885), .B(n34889), .Z(n34887) );
  XNOR U34819 ( .A(n34786), .B(n34844), .Z(n34846) );
  XNOR U34820 ( .A(n34890), .B(n34891), .Z(n34786) );
  AND U34821 ( .A(n1260), .B(n34793), .Z(n34891) );
  XOR U34822 ( .A(n34890), .B(n34791), .Z(n34793) );
  AND U34823 ( .A(n34794), .B(n34797), .Z(n34844) );
  XOR U34824 ( .A(n34892), .B(n34872), .Z(n34797) );
  XNOR U34825 ( .A(p_input[1776]), .B(p_input[2048]), .Z(n34872) );
  XNOR U34826 ( .A(n34859), .B(n34858), .Z(n34892) );
  XNOR U34827 ( .A(n34893), .B(n34866), .Z(n34858) );
  XNOR U34828 ( .A(n34854), .B(n34853), .Z(n34866) );
  XNOR U34829 ( .A(n34894), .B(n34850), .Z(n34853) );
  XNOR U34830 ( .A(p_input[1786]), .B(p_input[2058]), .Z(n34850) );
  XOR U34831 ( .A(p_input[1787]), .B(n16732), .Z(n34894) );
  XOR U34832 ( .A(p_input[1788]), .B(p_input[2060]), .Z(n34854) );
  XOR U34833 ( .A(n34864), .B(n34895), .Z(n34893) );
  IV U34834 ( .A(n34855), .Z(n34895) );
  XOR U34835 ( .A(p_input[1777]), .B(p_input[2049]), .Z(n34855) );
  XNOR U34836 ( .A(n34896), .B(n34871), .Z(n34864) );
  XNOR U34837 ( .A(p_input[1791]), .B(n16735), .Z(n34871) );
  XOR U34838 ( .A(n34861), .B(n34870), .Z(n34896) );
  XOR U34839 ( .A(n34897), .B(n34867), .Z(n34870) );
  XOR U34840 ( .A(p_input[1789]), .B(p_input[2061]), .Z(n34867) );
  XOR U34841 ( .A(p_input[1790]), .B(n16737), .Z(n34897) );
  XOR U34842 ( .A(p_input[1785]), .B(p_input[2057]), .Z(n34861) );
  XOR U34843 ( .A(n34879), .B(n34877), .Z(n34859) );
  XNOR U34844 ( .A(n34898), .B(n34884), .Z(n34877) );
  XOR U34845 ( .A(p_input[1784]), .B(p_input[2056]), .Z(n34884) );
  XOR U34846 ( .A(n34874), .B(n34883), .Z(n34898) );
  XOR U34847 ( .A(n34899), .B(n34880), .Z(n34883) );
  XOR U34848 ( .A(p_input[1782]), .B(p_input[2054]), .Z(n34880) );
  XOR U34849 ( .A(p_input[1783]), .B(n17722), .Z(n34899) );
  XOR U34850 ( .A(p_input[1778]), .B(p_input[2050]), .Z(n34874) );
  XNOR U34851 ( .A(n34889), .B(n34888), .Z(n34879) );
  XOR U34852 ( .A(n34900), .B(n34885), .Z(n34888) );
  XOR U34853 ( .A(p_input[1779]), .B(p_input[2051]), .Z(n34885) );
  XOR U34854 ( .A(p_input[1780]), .B(n17724), .Z(n34900) );
  XOR U34855 ( .A(p_input[1781]), .B(p_input[2053]), .Z(n34889) );
  XNOR U34856 ( .A(n34901), .B(n34902), .Z(n34794) );
  AND U34857 ( .A(n1260), .B(n34903), .Z(n34902) );
  XNOR U34858 ( .A(n34904), .B(n34905), .Z(n1260) );
  AND U34859 ( .A(n34906), .B(n34907), .Z(n34905) );
  XOR U34860 ( .A(n34904), .B(n34804), .Z(n34907) );
  XNOR U34861 ( .A(n34904), .B(n34758), .Z(n34906) );
  XOR U34862 ( .A(n34908), .B(n34909), .Z(n34904) );
  AND U34863 ( .A(n34910), .B(n34911), .Z(n34909) );
  XOR U34864 ( .A(n34908), .B(n34768), .Z(n34910) );
  XOR U34865 ( .A(n34912), .B(n34913), .Z(n34747) );
  AND U34866 ( .A(n1264), .B(n34903), .Z(n34913) );
  XNOR U34867 ( .A(n34901), .B(n34912), .Z(n34903) );
  XNOR U34868 ( .A(n34914), .B(n34915), .Z(n1264) );
  AND U34869 ( .A(n34916), .B(n34917), .Z(n34915) );
  XNOR U34870 ( .A(n34918), .B(n34914), .Z(n34917) );
  IV U34871 ( .A(n34804), .Z(n34918) );
  XNOR U34872 ( .A(n34919), .B(n34920), .Z(n34804) );
  AND U34873 ( .A(n1267), .B(n34921), .Z(n34920) );
  XNOR U34874 ( .A(n34919), .B(n34922), .Z(n34921) );
  XNOR U34875 ( .A(n34758), .B(n34914), .Z(n34916) );
  XOR U34876 ( .A(n34923), .B(n34924), .Z(n34758) );
  AND U34877 ( .A(n1275), .B(n34925), .Z(n34924) );
  XOR U34878 ( .A(n34908), .B(n34926), .Z(n34914) );
  AND U34879 ( .A(n34927), .B(n34911), .Z(n34926) );
  XNOR U34880 ( .A(n34817), .B(n34908), .Z(n34911) );
  XNOR U34881 ( .A(n34928), .B(n34929), .Z(n34817) );
  AND U34882 ( .A(n1267), .B(n34930), .Z(n34929) );
  XOR U34883 ( .A(n34931), .B(n34928), .Z(n34930) );
  XNOR U34884 ( .A(n34932), .B(n34908), .Z(n34927) );
  IV U34885 ( .A(n34768), .Z(n34932) );
  XOR U34886 ( .A(n34933), .B(n34934), .Z(n34768) );
  AND U34887 ( .A(n1275), .B(n34935), .Z(n34934) );
  XOR U34888 ( .A(n34936), .B(n34937), .Z(n34908) );
  AND U34889 ( .A(n34938), .B(n34939), .Z(n34937) );
  XNOR U34890 ( .A(n34842), .B(n34936), .Z(n34939) );
  XNOR U34891 ( .A(n34940), .B(n34941), .Z(n34842) );
  AND U34892 ( .A(n1267), .B(n34942), .Z(n34941) );
  XNOR U34893 ( .A(n34943), .B(n34940), .Z(n34942) );
  XOR U34894 ( .A(n34936), .B(n34779), .Z(n34938) );
  XOR U34895 ( .A(n34944), .B(n34945), .Z(n34779) );
  AND U34896 ( .A(n1275), .B(n34946), .Z(n34945) );
  XOR U34897 ( .A(n34947), .B(n34948), .Z(n34936) );
  AND U34898 ( .A(n34949), .B(n34950), .Z(n34948) );
  XNOR U34899 ( .A(n34947), .B(n34890), .Z(n34950) );
  XNOR U34900 ( .A(n34951), .B(n34952), .Z(n34890) );
  AND U34901 ( .A(n1267), .B(n34953), .Z(n34952) );
  XOR U34902 ( .A(n34954), .B(n34951), .Z(n34953) );
  XNOR U34903 ( .A(n34955), .B(n34947), .Z(n34949) );
  IV U34904 ( .A(n34791), .Z(n34955) );
  XOR U34905 ( .A(n34956), .B(n34957), .Z(n34791) );
  AND U34906 ( .A(n1275), .B(n34958), .Z(n34957) );
  AND U34907 ( .A(n34912), .B(n34901), .Z(n34947) );
  XNOR U34908 ( .A(n34959), .B(n34960), .Z(n34901) );
  AND U34909 ( .A(n1267), .B(n34961), .Z(n34960) );
  XNOR U34910 ( .A(n34962), .B(n34959), .Z(n34961) );
  XNOR U34911 ( .A(n34963), .B(n34964), .Z(n1267) );
  AND U34912 ( .A(n34965), .B(n34966), .Z(n34964) );
  XOR U34913 ( .A(n34922), .B(n34963), .Z(n34966) );
  AND U34914 ( .A(n34967), .B(n34968), .Z(n34922) );
  XOR U34915 ( .A(n34963), .B(n34919), .Z(n34965) );
  XNOR U34916 ( .A(n34969), .B(n34970), .Z(n34919) );
  AND U34917 ( .A(n1271), .B(n34925), .Z(n34970) );
  XOR U34918 ( .A(n34923), .B(n34969), .Z(n34925) );
  XOR U34919 ( .A(n34971), .B(n34972), .Z(n34963) );
  AND U34920 ( .A(n34973), .B(n34974), .Z(n34972) );
  XNOR U34921 ( .A(n34971), .B(n34967), .Z(n34974) );
  IV U34922 ( .A(n34931), .Z(n34967) );
  XOR U34923 ( .A(n34975), .B(n34976), .Z(n34931) );
  XOR U34924 ( .A(n34977), .B(n34968), .Z(n34976) );
  AND U34925 ( .A(n34943), .B(n34978), .Z(n34968) );
  AND U34926 ( .A(n34979), .B(n34980), .Z(n34977) );
  XOR U34927 ( .A(n34981), .B(n34975), .Z(n34979) );
  XNOR U34928 ( .A(n34928), .B(n34971), .Z(n34973) );
  XNOR U34929 ( .A(n34982), .B(n34983), .Z(n34928) );
  AND U34930 ( .A(n1271), .B(n34935), .Z(n34983) );
  XOR U34931 ( .A(n34982), .B(n34933), .Z(n34935) );
  XOR U34932 ( .A(n34984), .B(n34985), .Z(n34971) );
  AND U34933 ( .A(n34986), .B(n34987), .Z(n34985) );
  XNOR U34934 ( .A(n34984), .B(n34943), .Z(n34987) );
  XOR U34935 ( .A(n34988), .B(n34980), .Z(n34943) );
  XNOR U34936 ( .A(n34989), .B(n34975), .Z(n34980) );
  XOR U34937 ( .A(n34990), .B(n34991), .Z(n34975) );
  AND U34938 ( .A(n34992), .B(n34993), .Z(n34991) );
  XOR U34939 ( .A(n34994), .B(n34990), .Z(n34992) );
  XNOR U34940 ( .A(n34995), .B(n34996), .Z(n34989) );
  AND U34941 ( .A(n34997), .B(n34998), .Z(n34996) );
  XOR U34942 ( .A(n34995), .B(n34999), .Z(n34997) );
  XNOR U34943 ( .A(n34981), .B(n34978), .Z(n34988) );
  AND U34944 ( .A(n35000), .B(n35001), .Z(n34978) );
  XOR U34945 ( .A(n35002), .B(n35003), .Z(n34981) );
  AND U34946 ( .A(n35004), .B(n35005), .Z(n35003) );
  XOR U34947 ( .A(n35002), .B(n35006), .Z(n35004) );
  XNOR U34948 ( .A(n34940), .B(n34984), .Z(n34986) );
  XNOR U34949 ( .A(n35007), .B(n35008), .Z(n34940) );
  AND U34950 ( .A(n1271), .B(n34946), .Z(n35008) );
  XOR U34951 ( .A(n35007), .B(n34944), .Z(n34946) );
  XOR U34952 ( .A(n35009), .B(n35010), .Z(n34984) );
  AND U34953 ( .A(n35011), .B(n35012), .Z(n35010) );
  XNOR U34954 ( .A(n35009), .B(n35000), .Z(n35012) );
  IV U34955 ( .A(n34954), .Z(n35000) );
  XNOR U34956 ( .A(n35013), .B(n34993), .Z(n34954) );
  XNOR U34957 ( .A(n35014), .B(n34999), .Z(n34993) );
  XNOR U34958 ( .A(n35015), .B(n35016), .Z(n34999) );
  NOR U34959 ( .A(n35017), .B(n35018), .Z(n35016) );
  XOR U34960 ( .A(n35015), .B(n35019), .Z(n35017) );
  XNOR U34961 ( .A(n34998), .B(n34990), .Z(n35014) );
  XOR U34962 ( .A(n35020), .B(n35021), .Z(n34990) );
  AND U34963 ( .A(n35022), .B(n35023), .Z(n35021) );
  XOR U34964 ( .A(n35020), .B(n35024), .Z(n35022) );
  XNOR U34965 ( .A(n35025), .B(n34995), .Z(n34998) );
  XOR U34966 ( .A(n35026), .B(n35027), .Z(n34995) );
  AND U34967 ( .A(n35028), .B(n35029), .Z(n35027) );
  XNOR U34968 ( .A(n35030), .B(n35031), .Z(n35028) );
  IV U34969 ( .A(n35026), .Z(n35030) );
  XNOR U34970 ( .A(n35032), .B(n35033), .Z(n35025) );
  NOR U34971 ( .A(n35034), .B(n35035), .Z(n35033) );
  XNOR U34972 ( .A(n35032), .B(n35036), .Z(n35034) );
  XNOR U34973 ( .A(n34994), .B(n35001), .Z(n35013) );
  NOR U34974 ( .A(n34962), .B(n35037), .Z(n35001) );
  XOR U34975 ( .A(n35006), .B(n35005), .Z(n34994) );
  XNOR U34976 ( .A(n35038), .B(n35002), .Z(n35005) );
  XOR U34977 ( .A(n35039), .B(n35040), .Z(n35002) );
  AND U34978 ( .A(n35041), .B(n35042), .Z(n35040) );
  XNOR U34979 ( .A(n35043), .B(n35044), .Z(n35041) );
  IV U34980 ( .A(n35039), .Z(n35043) );
  XNOR U34981 ( .A(n35045), .B(n35046), .Z(n35038) );
  NOR U34982 ( .A(n35047), .B(n35048), .Z(n35046) );
  XNOR U34983 ( .A(n35045), .B(n35049), .Z(n35047) );
  XOR U34984 ( .A(n35050), .B(n35051), .Z(n35006) );
  NOR U34985 ( .A(n35052), .B(n35053), .Z(n35051) );
  XNOR U34986 ( .A(n35050), .B(n35054), .Z(n35052) );
  XNOR U34987 ( .A(n34951), .B(n35009), .Z(n35011) );
  XNOR U34988 ( .A(n35055), .B(n35056), .Z(n34951) );
  AND U34989 ( .A(n1271), .B(n34958), .Z(n35056) );
  XOR U34990 ( .A(n35055), .B(n34956), .Z(n34958) );
  AND U34991 ( .A(n34959), .B(n34962), .Z(n35009) );
  XOR U34992 ( .A(n35057), .B(n35037), .Z(n34962) );
  XNOR U34993 ( .A(p_input[1792]), .B(p_input[2048]), .Z(n35037) );
  XNOR U34994 ( .A(n35024), .B(n35023), .Z(n35057) );
  XNOR U34995 ( .A(n35058), .B(n35031), .Z(n35023) );
  XNOR U34996 ( .A(n35019), .B(n35018), .Z(n35031) );
  XNOR U34997 ( .A(n35059), .B(n35015), .Z(n35018) );
  XNOR U34998 ( .A(p_input[1802]), .B(p_input[2058]), .Z(n35015) );
  XOR U34999 ( .A(p_input[1803]), .B(n16732), .Z(n35059) );
  XOR U35000 ( .A(p_input[1804]), .B(p_input[2060]), .Z(n35019) );
  XOR U35001 ( .A(n35029), .B(n35060), .Z(n35058) );
  IV U35002 ( .A(n35020), .Z(n35060) );
  XOR U35003 ( .A(p_input[1793]), .B(p_input[2049]), .Z(n35020) );
  XNOR U35004 ( .A(n35061), .B(n35036), .Z(n35029) );
  XNOR U35005 ( .A(p_input[1807]), .B(n16735), .Z(n35036) );
  XOR U35006 ( .A(n35026), .B(n35035), .Z(n35061) );
  XOR U35007 ( .A(n35062), .B(n35032), .Z(n35035) );
  XOR U35008 ( .A(p_input[1805]), .B(p_input[2061]), .Z(n35032) );
  XOR U35009 ( .A(p_input[1806]), .B(n16737), .Z(n35062) );
  XOR U35010 ( .A(p_input[1801]), .B(p_input[2057]), .Z(n35026) );
  XOR U35011 ( .A(n35044), .B(n35042), .Z(n35024) );
  XNOR U35012 ( .A(n35063), .B(n35049), .Z(n35042) );
  XOR U35013 ( .A(p_input[1800]), .B(p_input[2056]), .Z(n35049) );
  XOR U35014 ( .A(n35039), .B(n35048), .Z(n35063) );
  XOR U35015 ( .A(n35064), .B(n35045), .Z(n35048) );
  XOR U35016 ( .A(p_input[1798]), .B(p_input[2054]), .Z(n35045) );
  XOR U35017 ( .A(p_input[1799]), .B(n17722), .Z(n35064) );
  XOR U35018 ( .A(p_input[1794]), .B(p_input[2050]), .Z(n35039) );
  XNOR U35019 ( .A(n35054), .B(n35053), .Z(n35044) );
  XOR U35020 ( .A(n35065), .B(n35050), .Z(n35053) );
  XOR U35021 ( .A(p_input[1795]), .B(p_input[2051]), .Z(n35050) );
  XOR U35022 ( .A(p_input[1796]), .B(n17724), .Z(n35065) );
  XOR U35023 ( .A(p_input[1797]), .B(p_input[2053]), .Z(n35054) );
  XNOR U35024 ( .A(n35066), .B(n35067), .Z(n34959) );
  AND U35025 ( .A(n1271), .B(n35068), .Z(n35067) );
  XNOR U35026 ( .A(n35069), .B(n35070), .Z(n1271) );
  AND U35027 ( .A(n35071), .B(n35072), .Z(n35070) );
  XOR U35028 ( .A(n35069), .B(n34969), .Z(n35072) );
  XNOR U35029 ( .A(n35069), .B(n34923), .Z(n35071) );
  XOR U35030 ( .A(n35073), .B(n35074), .Z(n35069) );
  AND U35031 ( .A(n35075), .B(n35076), .Z(n35074) );
  XOR U35032 ( .A(n35073), .B(n34933), .Z(n35075) );
  XOR U35033 ( .A(n35077), .B(n35078), .Z(n34912) );
  AND U35034 ( .A(n1275), .B(n35068), .Z(n35078) );
  XNOR U35035 ( .A(n35066), .B(n35077), .Z(n35068) );
  XNOR U35036 ( .A(n35079), .B(n35080), .Z(n1275) );
  AND U35037 ( .A(n35081), .B(n35082), .Z(n35080) );
  XNOR U35038 ( .A(n35083), .B(n35079), .Z(n35082) );
  IV U35039 ( .A(n34969), .Z(n35083) );
  XNOR U35040 ( .A(n35084), .B(n35085), .Z(n34969) );
  AND U35041 ( .A(n1278), .B(n35086), .Z(n35085) );
  XNOR U35042 ( .A(n35084), .B(n35087), .Z(n35086) );
  XNOR U35043 ( .A(n34923), .B(n35079), .Z(n35081) );
  XOR U35044 ( .A(n35088), .B(n35089), .Z(n34923) );
  AND U35045 ( .A(n1286), .B(n35090), .Z(n35089) );
  XOR U35046 ( .A(n35073), .B(n35091), .Z(n35079) );
  AND U35047 ( .A(n35092), .B(n35076), .Z(n35091) );
  XNOR U35048 ( .A(n34982), .B(n35073), .Z(n35076) );
  XNOR U35049 ( .A(n35093), .B(n35094), .Z(n34982) );
  AND U35050 ( .A(n1278), .B(n35095), .Z(n35094) );
  XOR U35051 ( .A(n35096), .B(n35093), .Z(n35095) );
  XNOR U35052 ( .A(n35097), .B(n35073), .Z(n35092) );
  IV U35053 ( .A(n34933), .Z(n35097) );
  XOR U35054 ( .A(n35098), .B(n35099), .Z(n34933) );
  AND U35055 ( .A(n1286), .B(n35100), .Z(n35099) );
  XOR U35056 ( .A(n35101), .B(n35102), .Z(n35073) );
  AND U35057 ( .A(n35103), .B(n35104), .Z(n35102) );
  XNOR U35058 ( .A(n35007), .B(n35101), .Z(n35104) );
  XNOR U35059 ( .A(n35105), .B(n35106), .Z(n35007) );
  AND U35060 ( .A(n1278), .B(n35107), .Z(n35106) );
  XNOR U35061 ( .A(n35108), .B(n35105), .Z(n35107) );
  XOR U35062 ( .A(n35101), .B(n34944), .Z(n35103) );
  XOR U35063 ( .A(n35109), .B(n35110), .Z(n34944) );
  AND U35064 ( .A(n1286), .B(n35111), .Z(n35110) );
  XOR U35065 ( .A(n35112), .B(n35113), .Z(n35101) );
  AND U35066 ( .A(n35114), .B(n35115), .Z(n35113) );
  XNOR U35067 ( .A(n35112), .B(n35055), .Z(n35115) );
  XNOR U35068 ( .A(n35116), .B(n35117), .Z(n35055) );
  AND U35069 ( .A(n1278), .B(n35118), .Z(n35117) );
  XOR U35070 ( .A(n35119), .B(n35116), .Z(n35118) );
  XNOR U35071 ( .A(n35120), .B(n35112), .Z(n35114) );
  IV U35072 ( .A(n34956), .Z(n35120) );
  XOR U35073 ( .A(n35121), .B(n35122), .Z(n34956) );
  AND U35074 ( .A(n1286), .B(n35123), .Z(n35122) );
  AND U35075 ( .A(n35077), .B(n35066), .Z(n35112) );
  XNOR U35076 ( .A(n35124), .B(n35125), .Z(n35066) );
  AND U35077 ( .A(n1278), .B(n35126), .Z(n35125) );
  XNOR U35078 ( .A(n35127), .B(n35124), .Z(n35126) );
  XNOR U35079 ( .A(n35128), .B(n35129), .Z(n1278) );
  AND U35080 ( .A(n35130), .B(n35131), .Z(n35129) );
  XOR U35081 ( .A(n35087), .B(n35128), .Z(n35131) );
  AND U35082 ( .A(n35132), .B(n35133), .Z(n35087) );
  XOR U35083 ( .A(n35128), .B(n35084), .Z(n35130) );
  XNOR U35084 ( .A(n35134), .B(n35135), .Z(n35084) );
  AND U35085 ( .A(n1282), .B(n35090), .Z(n35135) );
  XOR U35086 ( .A(n35088), .B(n35134), .Z(n35090) );
  XOR U35087 ( .A(n35136), .B(n35137), .Z(n35128) );
  AND U35088 ( .A(n35138), .B(n35139), .Z(n35137) );
  XNOR U35089 ( .A(n35136), .B(n35132), .Z(n35139) );
  IV U35090 ( .A(n35096), .Z(n35132) );
  XOR U35091 ( .A(n35140), .B(n35141), .Z(n35096) );
  XOR U35092 ( .A(n35142), .B(n35133), .Z(n35141) );
  AND U35093 ( .A(n35108), .B(n35143), .Z(n35133) );
  AND U35094 ( .A(n35144), .B(n35145), .Z(n35142) );
  XOR U35095 ( .A(n35146), .B(n35140), .Z(n35144) );
  XNOR U35096 ( .A(n35093), .B(n35136), .Z(n35138) );
  XNOR U35097 ( .A(n35147), .B(n35148), .Z(n35093) );
  AND U35098 ( .A(n1282), .B(n35100), .Z(n35148) );
  XOR U35099 ( .A(n35147), .B(n35098), .Z(n35100) );
  XOR U35100 ( .A(n35149), .B(n35150), .Z(n35136) );
  AND U35101 ( .A(n35151), .B(n35152), .Z(n35150) );
  XNOR U35102 ( .A(n35149), .B(n35108), .Z(n35152) );
  XOR U35103 ( .A(n35153), .B(n35145), .Z(n35108) );
  XNOR U35104 ( .A(n35154), .B(n35140), .Z(n35145) );
  XOR U35105 ( .A(n35155), .B(n35156), .Z(n35140) );
  AND U35106 ( .A(n35157), .B(n35158), .Z(n35156) );
  XOR U35107 ( .A(n35159), .B(n35155), .Z(n35157) );
  XNOR U35108 ( .A(n35160), .B(n35161), .Z(n35154) );
  AND U35109 ( .A(n35162), .B(n35163), .Z(n35161) );
  XOR U35110 ( .A(n35160), .B(n35164), .Z(n35162) );
  XNOR U35111 ( .A(n35146), .B(n35143), .Z(n35153) );
  AND U35112 ( .A(n35165), .B(n35166), .Z(n35143) );
  XOR U35113 ( .A(n35167), .B(n35168), .Z(n35146) );
  AND U35114 ( .A(n35169), .B(n35170), .Z(n35168) );
  XOR U35115 ( .A(n35167), .B(n35171), .Z(n35169) );
  XNOR U35116 ( .A(n35105), .B(n35149), .Z(n35151) );
  XNOR U35117 ( .A(n35172), .B(n35173), .Z(n35105) );
  AND U35118 ( .A(n1282), .B(n35111), .Z(n35173) );
  XOR U35119 ( .A(n35172), .B(n35109), .Z(n35111) );
  XOR U35120 ( .A(n35174), .B(n35175), .Z(n35149) );
  AND U35121 ( .A(n35176), .B(n35177), .Z(n35175) );
  XNOR U35122 ( .A(n35174), .B(n35165), .Z(n35177) );
  IV U35123 ( .A(n35119), .Z(n35165) );
  XNOR U35124 ( .A(n35178), .B(n35158), .Z(n35119) );
  XNOR U35125 ( .A(n35179), .B(n35164), .Z(n35158) );
  XNOR U35126 ( .A(n35180), .B(n35181), .Z(n35164) );
  NOR U35127 ( .A(n35182), .B(n35183), .Z(n35181) );
  XOR U35128 ( .A(n35180), .B(n35184), .Z(n35182) );
  XNOR U35129 ( .A(n35163), .B(n35155), .Z(n35179) );
  XOR U35130 ( .A(n35185), .B(n35186), .Z(n35155) );
  AND U35131 ( .A(n35187), .B(n35188), .Z(n35186) );
  XOR U35132 ( .A(n35185), .B(n35189), .Z(n35187) );
  XNOR U35133 ( .A(n35190), .B(n35160), .Z(n35163) );
  XOR U35134 ( .A(n35191), .B(n35192), .Z(n35160) );
  AND U35135 ( .A(n35193), .B(n35194), .Z(n35192) );
  XNOR U35136 ( .A(n35195), .B(n35196), .Z(n35193) );
  IV U35137 ( .A(n35191), .Z(n35195) );
  XNOR U35138 ( .A(n35197), .B(n35198), .Z(n35190) );
  NOR U35139 ( .A(n35199), .B(n35200), .Z(n35198) );
  XNOR U35140 ( .A(n35197), .B(n35201), .Z(n35199) );
  XNOR U35141 ( .A(n35159), .B(n35166), .Z(n35178) );
  NOR U35142 ( .A(n35127), .B(n35202), .Z(n35166) );
  XOR U35143 ( .A(n35171), .B(n35170), .Z(n35159) );
  XNOR U35144 ( .A(n35203), .B(n35167), .Z(n35170) );
  XOR U35145 ( .A(n35204), .B(n35205), .Z(n35167) );
  AND U35146 ( .A(n35206), .B(n35207), .Z(n35205) );
  XNOR U35147 ( .A(n35208), .B(n35209), .Z(n35206) );
  IV U35148 ( .A(n35204), .Z(n35208) );
  XNOR U35149 ( .A(n35210), .B(n35211), .Z(n35203) );
  NOR U35150 ( .A(n35212), .B(n35213), .Z(n35211) );
  XNOR U35151 ( .A(n35210), .B(n35214), .Z(n35212) );
  XOR U35152 ( .A(n35215), .B(n35216), .Z(n35171) );
  NOR U35153 ( .A(n35217), .B(n35218), .Z(n35216) );
  XNOR U35154 ( .A(n35215), .B(n35219), .Z(n35217) );
  XNOR U35155 ( .A(n35116), .B(n35174), .Z(n35176) );
  XNOR U35156 ( .A(n35220), .B(n35221), .Z(n35116) );
  AND U35157 ( .A(n1282), .B(n35123), .Z(n35221) );
  XOR U35158 ( .A(n35220), .B(n35121), .Z(n35123) );
  AND U35159 ( .A(n35124), .B(n35127), .Z(n35174) );
  XOR U35160 ( .A(n35222), .B(n35202), .Z(n35127) );
  XNOR U35161 ( .A(p_input[1808]), .B(p_input[2048]), .Z(n35202) );
  XNOR U35162 ( .A(n35189), .B(n35188), .Z(n35222) );
  XNOR U35163 ( .A(n35223), .B(n35196), .Z(n35188) );
  XNOR U35164 ( .A(n35184), .B(n35183), .Z(n35196) );
  XNOR U35165 ( .A(n35224), .B(n35180), .Z(n35183) );
  XNOR U35166 ( .A(p_input[1818]), .B(p_input[2058]), .Z(n35180) );
  XOR U35167 ( .A(p_input[1819]), .B(n16732), .Z(n35224) );
  XOR U35168 ( .A(p_input[1820]), .B(p_input[2060]), .Z(n35184) );
  XOR U35169 ( .A(n35194), .B(n35225), .Z(n35223) );
  IV U35170 ( .A(n35185), .Z(n35225) );
  XOR U35171 ( .A(p_input[1809]), .B(p_input[2049]), .Z(n35185) );
  XNOR U35172 ( .A(n35226), .B(n35201), .Z(n35194) );
  XNOR U35173 ( .A(p_input[1823]), .B(n16735), .Z(n35201) );
  XOR U35174 ( .A(n35191), .B(n35200), .Z(n35226) );
  XOR U35175 ( .A(n35227), .B(n35197), .Z(n35200) );
  XOR U35176 ( .A(p_input[1821]), .B(p_input[2061]), .Z(n35197) );
  XOR U35177 ( .A(p_input[1822]), .B(n16737), .Z(n35227) );
  XOR U35178 ( .A(p_input[1817]), .B(p_input[2057]), .Z(n35191) );
  XOR U35179 ( .A(n35209), .B(n35207), .Z(n35189) );
  XNOR U35180 ( .A(n35228), .B(n35214), .Z(n35207) );
  XOR U35181 ( .A(p_input[1816]), .B(p_input[2056]), .Z(n35214) );
  XOR U35182 ( .A(n35204), .B(n35213), .Z(n35228) );
  XOR U35183 ( .A(n35229), .B(n35210), .Z(n35213) );
  XOR U35184 ( .A(p_input[1814]), .B(p_input[2054]), .Z(n35210) );
  XOR U35185 ( .A(p_input[1815]), .B(n17722), .Z(n35229) );
  XOR U35186 ( .A(p_input[1810]), .B(p_input[2050]), .Z(n35204) );
  XNOR U35187 ( .A(n35219), .B(n35218), .Z(n35209) );
  XOR U35188 ( .A(n35230), .B(n35215), .Z(n35218) );
  XOR U35189 ( .A(p_input[1811]), .B(p_input[2051]), .Z(n35215) );
  XOR U35190 ( .A(p_input[1812]), .B(n17724), .Z(n35230) );
  XOR U35191 ( .A(p_input[1813]), .B(p_input[2053]), .Z(n35219) );
  XNOR U35192 ( .A(n35231), .B(n35232), .Z(n35124) );
  AND U35193 ( .A(n1282), .B(n35233), .Z(n35232) );
  XNOR U35194 ( .A(n35234), .B(n35235), .Z(n1282) );
  AND U35195 ( .A(n35236), .B(n35237), .Z(n35235) );
  XOR U35196 ( .A(n35234), .B(n35134), .Z(n35237) );
  XNOR U35197 ( .A(n35234), .B(n35088), .Z(n35236) );
  XOR U35198 ( .A(n35238), .B(n35239), .Z(n35234) );
  AND U35199 ( .A(n35240), .B(n35241), .Z(n35239) );
  XOR U35200 ( .A(n35238), .B(n35098), .Z(n35240) );
  XOR U35201 ( .A(n35242), .B(n35243), .Z(n35077) );
  AND U35202 ( .A(n1286), .B(n35233), .Z(n35243) );
  XNOR U35203 ( .A(n35231), .B(n35242), .Z(n35233) );
  XNOR U35204 ( .A(n35244), .B(n35245), .Z(n1286) );
  AND U35205 ( .A(n35246), .B(n35247), .Z(n35245) );
  XNOR U35206 ( .A(n35248), .B(n35244), .Z(n35247) );
  IV U35207 ( .A(n35134), .Z(n35248) );
  XNOR U35208 ( .A(n35249), .B(n35250), .Z(n35134) );
  AND U35209 ( .A(n1289), .B(n35251), .Z(n35250) );
  XNOR U35210 ( .A(n35249), .B(n35252), .Z(n35251) );
  XNOR U35211 ( .A(n35088), .B(n35244), .Z(n35246) );
  XOR U35212 ( .A(n35253), .B(n35254), .Z(n35088) );
  AND U35213 ( .A(n1297), .B(n35255), .Z(n35254) );
  XOR U35214 ( .A(n35238), .B(n35256), .Z(n35244) );
  AND U35215 ( .A(n35257), .B(n35241), .Z(n35256) );
  XNOR U35216 ( .A(n35147), .B(n35238), .Z(n35241) );
  XNOR U35217 ( .A(n35258), .B(n35259), .Z(n35147) );
  AND U35218 ( .A(n1289), .B(n35260), .Z(n35259) );
  XOR U35219 ( .A(n35261), .B(n35258), .Z(n35260) );
  XNOR U35220 ( .A(n35262), .B(n35238), .Z(n35257) );
  IV U35221 ( .A(n35098), .Z(n35262) );
  XOR U35222 ( .A(n35263), .B(n35264), .Z(n35098) );
  AND U35223 ( .A(n1297), .B(n35265), .Z(n35264) );
  XOR U35224 ( .A(n35266), .B(n35267), .Z(n35238) );
  AND U35225 ( .A(n35268), .B(n35269), .Z(n35267) );
  XNOR U35226 ( .A(n35172), .B(n35266), .Z(n35269) );
  XNOR U35227 ( .A(n35270), .B(n35271), .Z(n35172) );
  AND U35228 ( .A(n1289), .B(n35272), .Z(n35271) );
  XNOR U35229 ( .A(n35273), .B(n35270), .Z(n35272) );
  XOR U35230 ( .A(n35266), .B(n35109), .Z(n35268) );
  XOR U35231 ( .A(n35274), .B(n35275), .Z(n35109) );
  AND U35232 ( .A(n1297), .B(n35276), .Z(n35275) );
  XOR U35233 ( .A(n35277), .B(n35278), .Z(n35266) );
  AND U35234 ( .A(n35279), .B(n35280), .Z(n35278) );
  XNOR U35235 ( .A(n35277), .B(n35220), .Z(n35280) );
  XNOR U35236 ( .A(n35281), .B(n35282), .Z(n35220) );
  AND U35237 ( .A(n1289), .B(n35283), .Z(n35282) );
  XOR U35238 ( .A(n35284), .B(n35281), .Z(n35283) );
  XNOR U35239 ( .A(n35285), .B(n35277), .Z(n35279) );
  IV U35240 ( .A(n35121), .Z(n35285) );
  XOR U35241 ( .A(n35286), .B(n35287), .Z(n35121) );
  AND U35242 ( .A(n1297), .B(n35288), .Z(n35287) );
  AND U35243 ( .A(n35242), .B(n35231), .Z(n35277) );
  XNOR U35244 ( .A(n35289), .B(n35290), .Z(n35231) );
  AND U35245 ( .A(n1289), .B(n35291), .Z(n35290) );
  XNOR U35246 ( .A(n35292), .B(n35289), .Z(n35291) );
  XNOR U35247 ( .A(n35293), .B(n35294), .Z(n1289) );
  AND U35248 ( .A(n35295), .B(n35296), .Z(n35294) );
  XOR U35249 ( .A(n35252), .B(n35293), .Z(n35296) );
  AND U35250 ( .A(n35297), .B(n35298), .Z(n35252) );
  XOR U35251 ( .A(n35293), .B(n35249), .Z(n35295) );
  XNOR U35252 ( .A(n35299), .B(n35300), .Z(n35249) );
  AND U35253 ( .A(n1293), .B(n35255), .Z(n35300) );
  XOR U35254 ( .A(n35253), .B(n35299), .Z(n35255) );
  XOR U35255 ( .A(n35301), .B(n35302), .Z(n35293) );
  AND U35256 ( .A(n35303), .B(n35304), .Z(n35302) );
  XNOR U35257 ( .A(n35301), .B(n35297), .Z(n35304) );
  IV U35258 ( .A(n35261), .Z(n35297) );
  XOR U35259 ( .A(n35305), .B(n35306), .Z(n35261) );
  XOR U35260 ( .A(n35307), .B(n35298), .Z(n35306) );
  AND U35261 ( .A(n35273), .B(n35308), .Z(n35298) );
  AND U35262 ( .A(n35309), .B(n35310), .Z(n35307) );
  XOR U35263 ( .A(n35311), .B(n35305), .Z(n35309) );
  XNOR U35264 ( .A(n35258), .B(n35301), .Z(n35303) );
  XNOR U35265 ( .A(n35312), .B(n35313), .Z(n35258) );
  AND U35266 ( .A(n1293), .B(n35265), .Z(n35313) );
  XOR U35267 ( .A(n35312), .B(n35263), .Z(n35265) );
  XOR U35268 ( .A(n35314), .B(n35315), .Z(n35301) );
  AND U35269 ( .A(n35316), .B(n35317), .Z(n35315) );
  XNOR U35270 ( .A(n35314), .B(n35273), .Z(n35317) );
  XOR U35271 ( .A(n35318), .B(n35310), .Z(n35273) );
  XNOR U35272 ( .A(n35319), .B(n35305), .Z(n35310) );
  XOR U35273 ( .A(n35320), .B(n35321), .Z(n35305) );
  AND U35274 ( .A(n35322), .B(n35323), .Z(n35321) );
  XOR U35275 ( .A(n35324), .B(n35320), .Z(n35322) );
  XNOR U35276 ( .A(n35325), .B(n35326), .Z(n35319) );
  AND U35277 ( .A(n35327), .B(n35328), .Z(n35326) );
  XOR U35278 ( .A(n35325), .B(n35329), .Z(n35327) );
  XNOR U35279 ( .A(n35311), .B(n35308), .Z(n35318) );
  AND U35280 ( .A(n35330), .B(n35331), .Z(n35308) );
  XOR U35281 ( .A(n35332), .B(n35333), .Z(n35311) );
  AND U35282 ( .A(n35334), .B(n35335), .Z(n35333) );
  XOR U35283 ( .A(n35332), .B(n35336), .Z(n35334) );
  XNOR U35284 ( .A(n35270), .B(n35314), .Z(n35316) );
  XNOR U35285 ( .A(n35337), .B(n35338), .Z(n35270) );
  AND U35286 ( .A(n1293), .B(n35276), .Z(n35338) );
  XOR U35287 ( .A(n35337), .B(n35274), .Z(n35276) );
  XOR U35288 ( .A(n35339), .B(n35340), .Z(n35314) );
  AND U35289 ( .A(n35341), .B(n35342), .Z(n35340) );
  XNOR U35290 ( .A(n35339), .B(n35330), .Z(n35342) );
  IV U35291 ( .A(n35284), .Z(n35330) );
  XNOR U35292 ( .A(n35343), .B(n35323), .Z(n35284) );
  XNOR U35293 ( .A(n35344), .B(n35329), .Z(n35323) );
  XNOR U35294 ( .A(n35345), .B(n35346), .Z(n35329) );
  NOR U35295 ( .A(n35347), .B(n35348), .Z(n35346) );
  XOR U35296 ( .A(n35345), .B(n35349), .Z(n35347) );
  XNOR U35297 ( .A(n35328), .B(n35320), .Z(n35344) );
  XOR U35298 ( .A(n35350), .B(n35351), .Z(n35320) );
  AND U35299 ( .A(n35352), .B(n35353), .Z(n35351) );
  XOR U35300 ( .A(n35350), .B(n35354), .Z(n35352) );
  XNOR U35301 ( .A(n35355), .B(n35325), .Z(n35328) );
  XOR U35302 ( .A(n35356), .B(n35357), .Z(n35325) );
  AND U35303 ( .A(n35358), .B(n35359), .Z(n35357) );
  XNOR U35304 ( .A(n35360), .B(n35361), .Z(n35358) );
  IV U35305 ( .A(n35356), .Z(n35360) );
  XNOR U35306 ( .A(n35362), .B(n35363), .Z(n35355) );
  NOR U35307 ( .A(n35364), .B(n35365), .Z(n35363) );
  XNOR U35308 ( .A(n35362), .B(n35366), .Z(n35364) );
  XNOR U35309 ( .A(n35324), .B(n35331), .Z(n35343) );
  NOR U35310 ( .A(n35292), .B(n35367), .Z(n35331) );
  XOR U35311 ( .A(n35336), .B(n35335), .Z(n35324) );
  XNOR U35312 ( .A(n35368), .B(n35332), .Z(n35335) );
  XOR U35313 ( .A(n35369), .B(n35370), .Z(n35332) );
  AND U35314 ( .A(n35371), .B(n35372), .Z(n35370) );
  XNOR U35315 ( .A(n35373), .B(n35374), .Z(n35371) );
  IV U35316 ( .A(n35369), .Z(n35373) );
  XNOR U35317 ( .A(n35375), .B(n35376), .Z(n35368) );
  NOR U35318 ( .A(n35377), .B(n35378), .Z(n35376) );
  XNOR U35319 ( .A(n35375), .B(n35379), .Z(n35377) );
  XOR U35320 ( .A(n35380), .B(n35381), .Z(n35336) );
  NOR U35321 ( .A(n35382), .B(n35383), .Z(n35381) );
  XNOR U35322 ( .A(n35380), .B(n35384), .Z(n35382) );
  XNOR U35323 ( .A(n35281), .B(n35339), .Z(n35341) );
  XNOR U35324 ( .A(n35385), .B(n35386), .Z(n35281) );
  AND U35325 ( .A(n1293), .B(n35288), .Z(n35386) );
  XOR U35326 ( .A(n35385), .B(n35286), .Z(n35288) );
  AND U35327 ( .A(n35289), .B(n35292), .Z(n35339) );
  XOR U35328 ( .A(n35387), .B(n35367), .Z(n35292) );
  XNOR U35329 ( .A(p_input[1824]), .B(p_input[2048]), .Z(n35367) );
  XNOR U35330 ( .A(n35354), .B(n35353), .Z(n35387) );
  XNOR U35331 ( .A(n35388), .B(n35361), .Z(n35353) );
  XNOR U35332 ( .A(n35349), .B(n35348), .Z(n35361) );
  XNOR U35333 ( .A(n35389), .B(n35345), .Z(n35348) );
  XNOR U35334 ( .A(p_input[1834]), .B(p_input[2058]), .Z(n35345) );
  XOR U35335 ( .A(p_input[1835]), .B(n16732), .Z(n35389) );
  XOR U35336 ( .A(p_input[1836]), .B(p_input[2060]), .Z(n35349) );
  XOR U35337 ( .A(n35359), .B(n35390), .Z(n35388) );
  IV U35338 ( .A(n35350), .Z(n35390) );
  XOR U35339 ( .A(p_input[1825]), .B(p_input[2049]), .Z(n35350) );
  XNOR U35340 ( .A(n35391), .B(n35366), .Z(n35359) );
  XNOR U35341 ( .A(p_input[1839]), .B(n16735), .Z(n35366) );
  XOR U35342 ( .A(n35356), .B(n35365), .Z(n35391) );
  XOR U35343 ( .A(n35392), .B(n35362), .Z(n35365) );
  XOR U35344 ( .A(p_input[1837]), .B(p_input[2061]), .Z(n35362) );
  XOR U35345 ( .A(p_input[1838]), .B(n16737), .Z(n35392) );
  XOR U35346 ( .A(p_input[1833]), .B(p_input[2057]), .Z(n35356) );
  XOR U35347 ( .A(n35374), .B(n35372), .Z(n35354) );
  XNOR U35348 ( .A(n35393), .B(n35379), .Z(n35372) );
  XOR U35349 ( .A(p_input[1832]), .B(p_input[2056]), .Z(n35379) );
  XOR U35350 ( .A(n35369), .B(n35378), .Z(n35393) );
  XOR U35351 ( .A(n35394), .B(n35375), .Z(n35378) );
  XOR U35352 ( .A(p_input[1830]), .B(p_input[2054]), .Z(n35375) );
  XOR U35353 ( .A(p_input[1831]), .B(n17722), .Z(n35394) );
  XOR U35354 ( .A(p_input[1826]), .B(p_input[2050]), .Z(n35369) );
  XNOR U35355 ( .A(n35384), .B(n35383), .Z(n35374) );
  XOR U35356 ( .A(n35395), .B(n35380), .Z(n35383) );
  XOR U35357 ( .A(p_input[1827]), .B(p_input[2051]), .Z(n35380) );
  XOR U35358 ( .A(p_input[1828]), .B(n17724), .Z(n35395) );
  XOR U35359 ( .A(p_input[1829]), .B(p_input[2053]), .Z(n35384) );
  XNOR U35360 ( .A(n35396), .B(n35397), .Z(n35289) );
  AND U35361 ( .A(n1293), .B(n35398), .Z(n35397) );
  XNOR U35362 ( .A(n35399), .B(n35400), .Z(n1293) );
  AND U35363 ( .A(n35401), .B(n35402), .Z(n35400) );
  XOR U35364 ( .A(n35399), .B(n35299), .Z(n35402) );
  XNOR U35365 ( .A(n35399), .B(n35253), .Z(n35401) );
  XOR U35366 ( .A(n35403), .B(n35404), .Z(n35399) );
  AND U35367 ( .A(n35405), .B(n35406), .Z(n35404) );
  XOR U35368 ( .A(n35403), .B(n35263), .Z(n35405) );
  XOR U35369 ( .A(n35407), .B(n35408), .Z(n35242) );
  AND U35370 ( .A(n1297), .B(n35398), .Z(n35408) );
  XNOR U35371 ( .A(n35396), .B(n35407), .Z(n35398) );
  XNOR U35372 ( .A(n35409), .B(n35410), .Z(n1297) );
  AND U35373 ( .A(n35411), .B(n35412), .Z(n35410) );
  XNOR U35374 ( .A(n35413), .B(n35409), .Z(n35412) );
  IV U35375 ( .A(n35299), .Z(n35413) );
  XNOR U35376 ( .A(n35414), .B(n35415), .Z(n35299) );
  AND U35377 ( .A(n1300), .B(n35416), .Z(n35415) );
  XNOR U35378 ( .A(n35414), .B(n35417), .Z(n35416) );
  XNOR U35379 ( .A(n35253), .B(n35409), .Z(n35411) );
  XOR U35380 ( .A(n35418), .B(n35419), .Z(n35253) );
  AND U35381 ( .A(n1308), .B(n35420), .Z(n35419) );
  XOR U35382 ( .A(n35403), .B(n35421), .Z(n35409) );
  AND U35383 ( .A(n35422), .B(n35406), .Z(n35421) );
  XNOR U35384 ( .A(n35312), .B(n35403), .Z(n35406) );
  XNOR U35385 ( .A(n35423), .B(n35424), .Z(n35312) );
  AND U35386 ( .A(n1300), .B(n35425), .Z(n35424) );
  XOR U35387 ( .A(n35426), .B(n35423), .Z(n35425) );
  XNOR U35388 ( .A(n35427), .B(n35403), .Z(n35422) );
  IV U35389 ( .A(n35263), .Z(n35427) );
  XOR U35390 ( .A(n35428), .B(n35429), .Z(n35263) );
  AND U35391 ( .A(n1308), .B(n35430), .Z(n35429) );
  XOR U35392 ( .A(n35431), .B(n35432), .Z(n35403) );
  AND U35393 ( .A(n35433), .B(n35434), .Z(n35432) );
  XNOR U35394 ( .A(n35337), .B(n35431), .Z(n35434) );
  XNOR U35395 ( .A(n35435), .B(n35436), .Z(n35337) );
  AND U35396 ( .A(n1300), .B(n35437), .Z(n35436) );
  XNOR U35397 ( .A(n35438), .B(n35435), .Z(n35437) );
  XOR U35398 ( .A(n35431), .B(n35274), .Z(n35433) );
  XOR U35399 ( .A(n35439), .B(n35440), .Z(n35274) );
  AND U35400 ( .A(n1308), .B(n35441), .Z(n35440) );
  XOR U35401 ( .A(n35442), .B(n35443), .Z(n35431) );
  AND U35402 ( .A(n35444), .B(n35445), .Z(n35443) );
  XNOR U35403 ( .A(n35442), .B(n35385), .Z(n35445) );
  XNOR U35404 ( .A(n35446), .B(n35447), .Z(n35385) );
  AND U35405 ( .A(n1300), .B(n35448), .Z(n35447) );
  XOR U35406 ( .A(n35449), .B(n35446), .Z(n35448) );
  XNOR U35407 ( .A(n35450), .B(n35442), .Z(n35444) );
  IV U35408 ( .A(n35286), .Z(n35450) );
  XOR U35409 ( .A(n35451), .B(n35452), .Z(n35286) );
  AND U35410 ( .A(n1308), .B(n35453), .Z(n35452) );
  AND U35411 ( .A(n35407), .B(n35396), .Z(n35442) );
  XNOR U35412 ( .A(n35454), .B(n35455), .Z(n35396) );
  AND U35413 ( .A(n1300), .B(n35456), .Z(n35455) );
  XNOR U35414 ( .A(n35457), .B(n35454), .Z(n35456) );
  XNOR U35415 ( .A(n35458), .B(n35459), .Z(n1300) );
  AND U35416 ( .A(n35460), .B(n35461), .Z(n35459) );
  XOR U35417 ( .A(n35417), .B(n35458), .Z(n35461) );
  AND U35418 ( .A(n35462), .B(n35463), .Z(n35417) );
  XOR U35419 ( .A(n35458), .B(n35414), .Z(n35460) );
  XNOR U35420 ( .A(n35464), .B(n35465), .Z(n35414) );
  AND U35421 ( .A(n1304), .B(n35420), .Z(n35465) );
  XOR U35422 ( .A(n35418), .B(n35464), .Z(n35420) );
  XOR U35423 ( .A(n35466), .B(n35467), .Z(n35458) );
  AND U35424 ( .A(n35468), .B(n35469), .Z(n35467) );
  XNOR U35425 ( .A(n35466), .B(n35462), .Z(n35469) );
  IV U35426 ( .A(n35426), .Z(n35462) );
  XOR U35427 ( .A(n35470), .B(n35471), .Z(n35426) );
  XOR U35428 ( .A(n35472), .B(n35463), .Z(n35471) );
  AND U35429 ( .A(n35438), .B(n35473), .Z(n35463) );
  AND U35430 ( .A(n35474), .B(n35475), .Z(n35472) );
  XOR U35431 ( .A(n35476), .B(n35470), .Z(n35474) );
  XNOR U35432 ( .A(n35423), .B(n35466), .Z(n35468) );
  XNOR U35433 ( .A(n35477), .B(n35478), .Z(n35423) );
  AND U35434 ( .A(n1304), .B(n35430), .Z(n35478) );
  XOR U35435 ( .A(n35477), .B(n35428), .Z(n35430) );
  XOR U35436 ( .A(n35479), .B(n35480), .Z(n35466) );
  AND U35437 ( .A(n35481), .B(n35482), .Z(n35480) );
  XNOR U35438 ( .A(n35479), .B(n35438), .Z(n35482) );
  XOR U35439 ( .A(n35483), .B(n35475), .Z(n35438) );
  XNOR U35440 ( .A(n35484), .B(n35470), .Z(n35475) );
  XOR U35441 ( .A(n35485), .B(n35486), .Z(n35470) );
  AND U35442 ( .A(n35487), .B(n35488), .Z(n35486) );
  XOR U35443 ( .A(n35489), .B(n35485), .Z(n35487) );
  XNOR U35444 ( .A(n35490), .B(n35491), .Z(n35484) );
  AND U35445 ( .A(n35492), .B(n35493), .Z(n35491) );
  XOR U35446 ( .A(n35490), .B(n35494), .Z(n35492) );
  XNOR U35447 ( .A(n35476), .B(n35473), .Z(n35483) );
  AND U35448 ( .A(n35495), .B(n35496), .Z(n35473) );
  XOR U35449 ( .A(n35497), .B(n35498), .Z(n35476) );
  AND U35450 ( .A(n35499), .B(n35500), .Z(n35498) );
  XOR U35451 ( .A(n35497), .B(n35501), .Z(n35499) );
  XNOR U35452 ( .A(n35435), .B(n35479), .Z(n35481) );
  XNOR U35453 ( .A(n35502), .B(n35503), .Z(n35435) );
  AND U35454 ( .A(n1304), .B(n35441), .Z(n35503) );
  XOR U35455 ( .A(n35502), .B(n35439), .Z(n35441) );
  XOR U35456 ( .A(n35504), .B(n35505), .Z(n35479) );
  AND U35457 ( .A(n35506), .B(n35507), .Z(n35505) );
  XNOR U35458 ( .A(n35504), .B(n35495), .Z(n35507) );
  IV U35459 ( .A(n35449), .Z(n35495) );
  XNOR U35460 ( .A(n35508), .B(n35488), .Z(n35449) );
  XNOR U35461 ( .A(n35509), .B(n35494), .Z(n35488) );
  XNOR U35462 ( .A(n35510), .B(n35511), .Z(n35494) );
  NOR U35463 ( .A(n35512), .B(n35513), .Z(n35511) );
  XOR U35464 ( .A(n35510), .B(n35514), .Z(n35512) );
  XNOR U35465 ( .A(n35493), .B(n35485), .Z(n35509) );
  XOR U35466 ( .A(n35515), .B(n35516), .Z(n35485) );
  AND U35467 ( .A(n35517), .B(n35518), .Z(n35516) );
  XOR U35468 ( .A(n35515), .B(n35519), .Z(n35517) );
  XNOR U35469 ( .A(n35520), .B(n35490), .Z(n35493) );
  XOR U35470 ( .A(n35521), .B(n35522), .Z(n35490) );
  AND U35471 ( .A(n35523), .B(n35524), .Z(n35522) );
  XNOR U35472 ( .A(n35525), .B(n35526), .Z(n35523) );
  IV U35473 ( .A(n35521), .Z(n35525) );
  XNOR U35474 ( .A(n35527), .B(n35528), .Z(n35520) );
  NOR U35475 ( .A(n35529), .B(n35530), .Z(n35528) );
  XNOR U35476 ( .A(n35527), .B(n35531), .Z(n35529) );
  XNOR U35477 ( .A(n35489), .B(n35496), .Z(n35508) );
  NOR U35478 ( .A(n35457), .B(n35532), .Z(n35496) );
  XOR U35479 ( .A(n35501), .B(n35500), .Z(n35489) );
  XNOR U35480 ( .A(n35533), .B(n35497), .Z(n35500) );
  XOR U35481 ( .A(n35534), .B(n35535), .Z(n35497) );
  AND U35482 ( .A(n35536), .B(n35537), .Z(n35535) );
  XNOR U35483 ( .A(n35538), .B(n35539), .Z(n35536) );
  IV U35484 ( .A(n35534), .Z(n35538) );
  XNOR U35485 ( .A(n35540), .B(n35541), .Z(n35533) );
  NOR U35486 ( .A(n35542), .B(n35543), .Z(n35541) );
  XNOR U35487 ( .A(n35540), .B(n35544), .Z(n35542) );
  XOR U35488 ( .A(n35545), .B(n35546), .Z(n35501) );
  NOR U35489 ( .A(n35547), .B(n35548), .Z(n35546) );
  XNOR U35490 ( .A(n35545), .B(n35549), .Z(n35547) );
  XNOR U35491 ( .A(n35446), .B(n35504), .Z(n35506) );
  XNOR U35492 ( .A(n35550), .B(n35551), .Z(n35446) );
  AND U35493 ( .A(n1304), .B(n35453), .Z(n35551) );
  XOR U35494 ( .A(n35550), .B(n35451), .Z(n35453) );
  AND U35495 ( .A(n35454), .B(n35457), .Z(n35504) );
  XOR U35496 ( .A(n35552), .B(n35532), .Z(n35457) );
  XNOR U35497 ( .A(p_input[1840]), .B(p_input[2048]), .Z(n35532) );
  XNOR U35498 ( .A(n35519), .B(n35518), .Z(n35552) );
  XNOR U35499 ( .A(n35553), .B(n35526), .Z(n35518) );
  XNOR U35500 ( .A(n35514), .B(n35513), .Z(n35526) );
  XNOR U35501 ( .A(n35554), .B(n35510), .Z(n35513) );
  XNOR U35502 ( .A(p_input[1850]), .B(p_input[2058]), .Z(n35510) );
  XOR U35503 ( .A(p_input[1851]), .B(n16732), .Z(n35554) );
  XOR U35504 ( .A(p_input[1852]), .B(p_input[2060]), .Z(n35514) );
  XOR U35505 ( .A(n35524), .B(n35555), .Z(n35553) );
  IV U35506 ( .A(n35515), .Z(n35555) );
  XOR U35507 ( .A(p_input[1841]), .B(p_input[2049]), .Z(n35515) );
  XNOR U35508 ( .A(n35556), .B(n35531), .Z(n35524) );
  XNOR U35509 ( .A(p_input[1855]), .B(n16735), .Z(n35531) );
  XOR U35510 ( .A(n35521), .B(n35530), .Z(n35556) );
  XOR U35511 ( .A(n35557), .B(n35527), .Z(n35530) );
  XOR U35512 ( .A(p_input[1853]), .B(p_input[2061]), .Z(n35527) );
  XOR U35513 ( .A(p_input[1854]), .B(n16737), .Z(n35557) );
  XOR U35514 ( .A(p_input[1849]), .B(p_input[2057]), .Z(n35521) );
  XOR U35515 ( .A(n35539), .B(n35537), .Z(n35519) );
  XNOR U35516 ( .A(n35558), .B(n35544), .Z(n35537) );
  XOR U35517 ( .A(p_input[1848]), .B(p_input[2056]), .Z(n35544) );
  XOR U35518 ( .A(n35534), .B(n35543), .Z(n35558) );
  XOR U35519 ( .A(n35559), .B(n35540), .Z(n35543) );
  XOR U35520 ( .A(p_input[1846]), .B(p_input[2054]), .Z(n35540) );
  XOR U35521 ( .A(p_input[1847]), .B(n17722), .Z(n35559) );
  XOR U35522 ( .A(p_input[1842]), .B(p_input[2050]), .Z(n35534) );
  XNOR U35523 ( .A(n35549), .B(n35548), .Z(n35539) );
  XOR U35524 ( .A(n35560), .B(n35545), .Z(n35548) );
  XOR U35525 ( .A(p_input[1843]), .B(p_input[2051]), .Z(n35545) );
  XOR U35526 ( .A(p_input[1844]), .B(n17724), .Z(n35560) );
  XOR U35527 ( .A(p_input[1845]), .B(p_input[2053]), .Z(n35549) );
  XNOR U35528 ( .A(n35561), .B(n35562), .Z(n35454) );
  AND U35529 ( .A(n1304), .B(n35563), .Z(n35562) );
  XNOR U35530 ( .A(n35564), .B(n35565), .Z(n1304) );
  AND U35531 ( .A(n35566), .B(n35567), .Z(n35565) );
  XOR U35532 ( .A(n35564), .B(n35464), .Z(n35567) );
  XNOR U35533 ( .A(n35564), .B(n35418), .Z(n35566) );
  XOR U35534 ( .A(n35568), .B(n35569), .Z(n35564) );
  AND U35535 ( .A(n35570), .B(n35571), .Z(n35569) );
  XOR U35536 ( .A(n35568), .B(n35428), .Z(n35570) );
  XOR U35537 ( .A(n35572), .B(n35573), .Z(n35407) );
  AND U35538 ( .A(n1308), .B(n35563), .Z(n35573) );
  XNOR U35539 ( .A(n35561), .B(n35572), .Z(n35563) );
  XNOR U35540 ( .A(n35574), .B(n35575), .Z(n1308) );
  AND U35541 ( .A(n35576), .B(n35577), .Z(n35575) );
  XNOR U35542 ( .A(n35578), .B(n35574), .Z(n35577) );
  IV U35543 ( .A(n35464), .Z(n35578) );
  XNOR U35544 ( .A(n35579), .B(n35580), .Z(n35464) );
  AND U35545 ( .A(n1311), .B(n35581), .Z(n35580) );
  XNOR U35546 ( .A(n35579), .B(n35582), .Z(n35581) );
  XNOR U35547 ( .A(n35418), .B(n35574), .Z(n35576) );
  XOR U35548 ( .A(n35583), .B(n35584), .Z(n35418) );
  AND U35549 ( .A(n1319), .B(n35585), .Z(n35584) );
  XOR U35550 ( .A(n35568), .B(n35586), .Z(n35574) );
  AND U35551 ( .A(n35587), .B(n35571), .Z(n35586) );
  XNOR U35552 ( .A(n35477), .B(n35568), .Z(n35571) );
  XNOR U35553 ( .A(n35588), .B(n35589), .Z(n35477) );
  AND U35554 ( .A(n1311), .B(n35590), .Z(n35589) );
  XOR U35555 ( .A(n35591), .B(n35588), .Z(n35590) );
  XNOR U35556 ( .A(n35592), .B(n35568), .Z(n35587) );
  IV U35557 ( .A(n35428), .Z(n35592) );
  XOR U35558 ( .A(n35593), .B(n35594), .Z(n35428) );
  AND U35559 ( .A(n1319), .B(n35595), .Z(n35594) );
  XOR U35560 ( .A(n35596), .B(n35597), .Z(n35568) );
  AND U35561 ( .A(n35598), .B(n35599), .Z(n35597) );
  XNOR U35562 ( .A(n35502), .B(n35596), .Z(n35599) );
  XNOR U35563 ( .A(n35600), .B(n35601), .Z(n35502) );
  AND U35564 ( .A(n1311), .B(n35602), .Z(n35601) );
  XNOR U35565 ( .A(n35603), .B(n35600), .Z(n35602) );
  XOR U35566 ( .A(n35596), .B(n35439), .Z(n35598) );
  XOR U35567 ( .A(n35604), .B(n35605), .Z(n35439) );
  AND U35568 ( .A(n1319), .B(n35606), .Z(n35605) );
  XOR U35569 ( .A(n35607), .B(n35608), .Z(n35596) );
  AND U35570 ( .A(n35609), .B(n35610), .Z(n35608) );
  XNOR U35571 ( .A(n35607), .B(n35550), .Z(n35610) );
  XNOR U35572 ( .A(n35611), .B(n35612), .Z(n35550) );
  AND U35573 ( .A(n1311), .B(n35613), .Z(n35612) );
  XOR U35574 ( .A(n35614), .B(n35611), .Z(n35613) );
  XNOR U35575 ( .A(n35615), .B(n35607), .Z(n35609) );
  IV U35576 ( .A(n35451), .Z(n35615) );
  XOR U35577 ( .A(n35616), .B(n35617), .Z(n35451) );
  AND U35578 ( .A(n1319), .B(n35618), .Z(n35617) );
  AND U35579 ( .A(n35572), .B(n35561), .Z(n35607) );
  XNOR U35580 ( .A(n35619), .B(n35620), .Z(n35561) );
  AND U35581 ( .A(n1311), .B(n35621), .Z(n35620) );
  XNOR U35582 ( .A(n35622), .B(n35619), .Z(n35621) );
  XNOR U35583 ( .A(n35623), .B(n35624), .Z(n1311) );
  AND U35584 ( .A(n35625), .B(n35626), .Z(n35624) );
  XOR U35585 ( .A(n35582), .B(n35623), .Z(n35626) );
  AND U35586 ( .A(n35627), .B(n35628), .Z(n35582) );
  XOR U35587 ( .A(n35623), .B(n35579), .Z(n35625) );
  XNOR U35588 ( .A(n35629), .B(n35630), .Z(n35579) );
  AND U35589 ( .A(n1315), .B(n35585), .Z(n35630) );
  XOR U35590 ( .A(n35583), .B(n35629), .Z(n35585) );
  XOR U35591 ( .A(n35631), .B(n35632), .Z(n35623) );
  AND U35592 ( .A(n35633), .B(n35634), .Z(n35632) );
  XNOR U35593 ( .A(n35631), .B(n35627), .Z(n35634) );
  IV U35594 ( .A(n35591), .Z(n35627) );
  XOR U35595 ( .A(n35635), .B(n35636), .Z(n35591) );
  XOR U35596 ( .A(n35637), .B(n35628), .Z(n35636) );
  AND U35597 ( .A(n35603), .B(n35638), .Z(n35628) );
  AND U35598 ( .A(n35639), .B(n35640), .Z(n35637) );
  XOR U35599 ( .A(n35641), .B(n35635), .Z(n35639) );
  XNOR U35600 ( .A(n35588), .B(n35631), .Z(n35633) );
  XNOR U35601 ( .A(n35642), .B(n35643), .Z(n35588) );
  AND U35602 ( .A(n1315), .B(n35595), .Z(n35643) );
  XOR U35603 ( .A(n35642), .B(n35593), .Z(n35595) );
  XOR U35604 ( .A(n35644), .B(n35645), .Z(n35631) );
  AND U35605 ( .A(n35646), .B(n35647), .Z(n35645) );
  XNOR U35606 ( .A(n35644), .B(n35603), .Z(n35647) );
  XOR U35607 ( .A(n35648), .B(n35640), .Z(n35603) );
  XNOR U35608 ( .A(n35649), .B(n35635), .Z(n35640) );
  XOR U35609 ( .A(n35650), .B(n35651), .Z(n35635) );
  AND U35610 ( .A(n35652), .B(n35653), .Z(n35651) );
  XOR U35611 ( .A(n35654), .B(n35650), .Z(n35652) );
  XNOR U35612 ( .A(n35655), .B(n35656), .Z(n35649) );
  AND U35613 ( .A(n35657), .B(n35658), .Z(n35656) );
  XOR U35614 ( .A(n35655), .B(n35659), .Z(n35657) );
  XNOR U35615 ( .A(n35641), .B(n35638), .Z(n35648) );
  AND U35616 ( .A(n35660), .B(n35661), .Z(n35638) );
  XOR U35617 ( .A(n35662), .B(n35663), .Z(n35641) );
  AND U35618 ( .A(n35664), .B(n35665), .Z(n35663) );
  XOR U35619 ( .A(n35662), .B(n35666), .Z(n35664) );
  XNOR U35620 ( .A(n35600), .B(n35644), .Z(n35646) );
  XNOR U35621 ( .A(n35667), .B(n35668), .Z(n35600) );
  AND U35622 ( .A(n1315), .B(n35606), .Z(n35668) );
  XOR U35623 ( .A(n35667), .B(n35604), .Z(n35606) );
  XOR U35624 ( .A(n35669), .B(n35670), .Z(n35644) );
  AND U35625 ( .A(n35671), .B(n35672), .Z(n35670) );
  XNOR U35626 ( .A(n35669), .B(n35660), .Z(n35672) );
  IV U35627 ( .A(n35614), .Z(n35660) );
  XNOR U35628 ( .A(n35673), .B(n35653), .Z(n35614) );
  XNOR U35629 ( .A(n35674), .B(n35659), .Z(n35653) );
  XNOR U35630 ( .A(n35675), .B(n35676), .Z(n35659) );
  NOR U35631 ( .A(n35677), .B(n35678), .Z(n35676) );
  XOR U35632 ( .A(n35675), .B(n35679), .Z(n35677) );
  XNOR U35633 ( .A(n35658), .B(n35650), .Z(n35674) );
  XOR U35634 ( .A(n35680), .B(n35681), .Z(n35650) );
  AND U35635 ( .A(n35682), .B(n35683), .Z(n35681) );
  XOR U35636 ( .A(n35680), .B(n35684), .Z(n35682) );
  XNOR U35637 ( .A(n35685), .B(n35655), .Z(n35658) );
  XOR U35638 ( .A(n35686), .B(n35687), .Z(n35655) );
  AND U35639 ( .A(n35688), .B(n35689), .Z(n35687) );
  XNOR U35640 ( .A(n35690), .B(n35691), .Z(n35688) );
  IV U35641 ( .A(n35686), .Z(n35690) );
  XNOR U35642 ( .A(n35692), .B(n35693), .Z(n35685) );
  NOR U35643 ( .A(n35694), .B(n35695), .Z(n35693) );
  XNOR U35644 ( .A(n35692), .B(n35696), .Z(n35694) );
  XNOR U35645 ( .A(n35654), .B(n35661), .Z(n35673) );
  NOR U35646 ( .A(n35622), .B(n35697), .Z(n35661) );
  XOR U35647 ( .A(n35666), .B(n35665), .Z(n35654) );
  XNOR U35648 ( .A(n35698), .B(n35662), .Z(n35665) );
  XOR U35649 ( .A(n35699), .B(n35700), .Z(n35662) );
  AND U35650 ( .A(n35701), .B(n35702), .Z(n35700) );
  XNOR U35651 ( .A(n35703), .B(n35704), .Z(n35701) );
  IV U35652 ( .A(n35699), .Z(n35703) );
  XNOR U35653 ( .A(n35705), .B(n35706), .Z(n35698) );
  NOR U35654 ( .A(n35707), .B(n35708), .Z(n35706) );
  XNOR U35655 ( .A(n35705), .B(n35709), .Z(n35707) );
  XOR U35656 ( .A(n35710), .B(n35711), .Z(n35666) );
  NOR U35657 ( .A(n35712), .B(n35713), .Z(n35711) );
  XNOR U35658 ( .A(n35710), .B(n35714), .Z(n35712) );
  XNOR U35659 ( .A(n35611), .B(n35669), .Z(n35671) );
  XNOR U35660 ( .A(n35715), .B(n35716), .Z(n35611) );
  AND U35661 ( .A(n1315), .B(n35618), .Z(n35716) );
  XOR U35662 ( .A(n35715), .B(n35616), .Z(n35618) );
  AND U35663 ( .A(n35619), .B(n35622), .Z(n35669) );
  XOR U35664 ( .A(n35717), .B(n35697), .Z(n35622) );
  XNOR U35665 ( .A(p_input[1856]), .B(p_input[2048]), .Z(n35697) );
  XNOR U35666 ( .A(n35684), .B(n35683), .Z(n35717) );
  XNOR U35667 ( .A(n35718), .B(n35691), .Z(n35683) );
  XNOR U35668 ( .A(n35679), .B(n35678), .Z(n35691) );
  XNOR U35669 ( .A(n35719), .B(n35675), .Z(n35678) );
  XNOR U35670 ( .A(p_input[1866]), .B(p_input[2058]), .Z(n35675) );
  XOR U35671 ( .A(p_input[1867]), .B(n16732), .Z(n35719) );
  XOR U35672 ( .A(p_input[1868]), .B(p_input[2060]), .Z(n35679) );
  XOR U35673 ( .A(n35689), .B(n35720), .Z(n35718) );
  IV U35674 ( .A(n35680), .Z(n35720) );
  XOR U35675 ( .A(p_input[1857]), .B(p_input[2049]), .Z(n35680) );
  XNOR U35676 ( .A(n35721), .B(n35696), .Z(n35689) );
  XNOR U35677 ( .A(p_input[1871]), .B(n16735), .Z(n35696) );
  XOR U35678 ( .A(n35686), .B(n35695), .Z(n35721) );
  XOR U35679 ( .A(n35722), .B(n35692), .Z(n35695) );
  XOR U35680 ( .A(p_input[1869]), .B(p_input[2061]), .Z(n35692) );
  XOR U35681 ( .A(p_input[1870]), .B(n16737), .Z(n35722) );
  XOR U35682 ( .A(p_input[1865]), .B(p_input[2057]), .Z(n35686) );
  XOR U35683 ( .A(n35704), .B(n35702), .Z(n35684) );
  XNOR U35684 ( .A(n35723), .B(n35709), .Z(n35702) );
  XOR U35685 ( .A(p_input[1864]), .B(p_input[2056]), .Z(n35709) );
  XOR U35686 ( .A(n35699), .B(n35708), .Z(n35723) );
  XOR U35687 ( .A(n35724), .B(n35705), .Z(n35708) );
  XOR U35688 ( .A(p_input[1862]), .B(p_input[2054]), .Z(n35705) );
  XOR U35689 ( .A(p_input[1863]), .B(n17722), .Z(n35724) );
  XOR U35690 ( .A(p_input[1858]), .B(p_input[2050]), .Z(n35699) );
  XNOR U35691 ( .A(n35714), .B(n35713), .Z(n35704) );
  XOR U35692 ( .A(n35725), .B(n35710), .Z(n35713) );
  XOR U35693 ( .A(p_input[1859]), .B(p_input[2051]), .Z(n35710) );
  XOR U35694 ( .A(p_input[1860]), .B(n17724), .Z(n35725) );
  XOR U35695 ( .A(p_input[1861]), .B(p_input[2053]), .Z(n35714) );
  XNOR U35696 ( .A(n35726), .B(n35727), .Z(n35619) );
  AND U35697 ( .A(n1315), .B(n35728), .Z(n35727) );
  XNOR U35698 ( .A(n35729), .B(n35730), .Z(n1315) );
  AND U35699 ( .A(n35731), .B(n35732), .Z(n35730) );
  XOR U35700 ( .A(n35729), .B(n35629), .Z(n35732) );
  XNOR U35701 ( .A(n35729), .B(n35583), .Z(n35731) );
  XOR U35702 ( .A(n35733), .B(n35734), .Z(n35729) );
  AND U35703 ( .A(n35735), .B(n35736), .Z(n35734) );
  XOR U35704 ( .A(n35733), .B(n35593), .Z(n35735) );
  XOR U35705 ( .A(n35737), .B(n35738), .Z(n35572) );
  AND U35706 ( .A(n1319), .B(n35728), .Z(n35738) );
  XNOR U35707 ( .A(n35726), .B(n35737), .Z(n35728) );
  XNOR U35708 ( .A(n35739), .B(n35740), .Z(n1319) );
  AND U35709 ( .A(n35741), .B(n35742), .Z(n35740) );
  XNOR U35710 ( .A(n35743), .B(n35739), .Z(n35742) );
  IV U35711 ( .A(n35629), .Z(n35743) );
  XNOR U35712 ( .A(n35744), .B(n35745), .Z(n35629) );
  AND U35713 ( .A(n1322), .B(n35746), .Z(n35745) );
  XNOR U35714 ( .A(n35744), .B(n35747), .Z(n35746) );
  XNOR U35715 ( .A(n35583), .B(n35739), .Z(n35741) );
  XOR U35716 ( .A(n35748), .B(n35749), .Z(n35583) );
  AND U35717 ( .A(n1330), .B(n35750), .Z(n35749) );
  XOR U35718 ( .A(n35733), .B(n35751), .Z(n35739) );
  AND U35719 ( .A(n35752), .B(n35736), .Z(n35751) );
  XNOR U35720 ( .A(n35642), .B(n35733), .Z(n35736) );
  XNOR U35721 ( .A(n35753), .B(n35754), .Z(n35642) );
  AND U35722 ( .A(n1322), .B(n35755), .Z(n35754) );
  XOR U35723 ( .A(n35756), .B(n35753), .Z(n35755) );
  XNOR U35724 ( .A(n35757), .B(n35733), .Z(n35752) );
  IV U35725 ( .A(n35593), .Z(n35757) );
  XOR U35726 ( .A(n35758), .B(n35759), .Z(n35593) );
  AND U35727 ( .A(n1330), .B(n35760), .Z(n35759) );
  XOR U35728 ( .A(n35761), .B(n35762), .Z(n35733) );
  AND U35729 ( .A(n35763), .B(n35764), .Z(n35762) );
  XNOR U35730 ( .A(n35667), .B(n35761), .Z(n35764) );
  XNOR U35731 ( .A(n35765), .B(n35766), .Z(n35667) );
  AND U35732 ( .A(n1322), .B(n35767), .Z(n35766) );
  XNOR U35733 ( .A(n35768), .B(n35765), .Z(n35767) );
  XOR U35734 ( .A(n35761), .B(n35604), .Z(n35763) );
  XOR U35735 ( .A(n35769), .B(n35770), .Z(n35604) );
  AND U35736 ( .A(n1330), .B(n35771), .Z(n35770) );
  XOR U35737 ( .A(n35772), .B(n35773), .Z(n35761) );
  AND U35738 ( .A(n35774), .B(n35775), .Z(n35773) );
  XNOR U35739 ( .A(n35772), .B(n35715), .Z(n35775) );
  XNOR U35740 ( .A(n35776), .B(n35777), .Z(n35715) );
  AND U35741 ( .A(n1322), .B(n35778), .Z(n35777) );
  XOR U35742 ( .A(n35779), .B(n35776), .Z(n35778) );
  XNOR U35743 ( .A(n35780), .B(n35772), .Z(n35774) );
  IV U35744 ( .A(n35616), .Z(n35780) );
  XOR U35745 ( .A(n35781), .B(n35782), .Z(n35616) );
  AND U35746 ( .A(n1330), .B(n35783), .Z(n35782) );
  AND U35747 ( .A(n35737), .B(n35726), .Z(n35772) );
  XNOR U35748 ( .A(n35784), .B(n35785), .Z(n35726) );
  AND U35749 ( .A(n1322), .B(n35786), .Z(n35785) );
  XNOR U35750 ( .A(n35787), .B(n35784), .Z(n35786) );
  XNOR U35751 ( .A(n35788), .B(n35789), .Z(n1322) );
  AND U35752 ( .A(n35790), .B(n35791), .Z(n35789) );
  XOR U35753 ( .A(n35747), .B(n35788), .Z(n35791) );
  AND U35754 ( .A(n35792), .B(n35793), .Z(n35747) );
  XOR U35755 ( .A(n35788), .B(n35744), .Z(n35790) );
  XNOR U35756 ( .A(n35794), .B(n35795), .Z(n35744) );
  AND U35757 ( .A(n1326), .B(n35750), .Z(n35795) );
  XOR U35758 ( .A(n35748), .B(n35794), .Z(n35750) );
  XOR U35759 ( .A(n35796), .B(n35797), .Z(n35788) );
  AND U35760 ( .A(n35798), .B(n35799), .Z(n35797) );
  XNOR U35761 ( .A(n35796), .B(n35792), .Z(n35799) );
  IV U35762 ( .A(n35756), .Z(n35792) );
  XOR U35763 ( .A(n35800), .B(n35801), .Z(n35756) );
  XOR U35764 ( .A(n35802), .B(n35793), .Z(n35801) );
  AND U35765 ( .A(n35768), .B(n35803), .Z(n35793) );
  AND U35766 ( .A(n35804), .B(n35805), .Z(n35802) );
  XOR U35767 ( .A(n35806), .B(n35800), .Z(n35804) );
  XNOR U35768 ( .A(n35753), .B(n35796), .Z(n35798) );
  XNOR U35769 ( .A(n35807), .B(n35808), .Z(n35753) );
  AND U35770 ( .A(n1326), .B(n35760), .Z(n35808) );
  XOR U35771 ( .A(n35807), .B(n35758), .Z(n35760) );
  XOR U35772 ( .A(n35809), .B(n35810), .Z(n35796) );
  AND U35773 ( .A(n35811), .B(n35812), .Z(n35810) );
  XNOR U35774 ( .A(n35809), .B(n35768), .Z(n35812) );
  XOR U35775 ( .A(n35813), .B(n35805), .Z(n35768) );
  XNOR U35776 ( .A(n35814), .B(n35800), .Z(n35805) );
  XOR U35777 ( .A(n35815), .B(n35816), .Z(n35800) );
  AND U35778 ( .A(n35817), .B(n35818), .Z(n35816) );
  XOR U35779 ( .A(n35819), .B(n35815), .Z(n35817) );
  XNOR U35780 ( .A(n35820), .B(n35821), .Z(n35814) );
  AND U35781 ( .A(n35822), .B(n35823), .Z(n35821) );
  XOR U35782 ( .A(n35820), .B(n35824), .Z(n35822) );
  XNOR U35783 ( .A(n35806), .B(n35803), .Z(n35813) );
  AND U35784 ( .A(n35825), .B(n35826), .Z(n35803) );
  XOR U35785 ( .A(n35827), .B(n35828), .Z(n35806) );
  AND U35786 ( .A(n35829), .B(n35830), .Z(n35828) );
  XOR U35787 ( .A(n35827), .B(n35831), .Z(n35829) );
  XNOR U35788 ( .A(n35765), .B(n35809), .Z(n35811) );
  XNOR U35789 ( .A(n35832), .B(n35833), .Z(n35765) );
  AND U35790 ( .A(n1326), .B(n35771), .Z(n35833) );
  XOR U35791 ( .A(n35832), .B(n35769), .Z(n35771) );
  XOR U35792 ( .A(n35834), .B(n35835), .Z(n35809) );
  AND U35793 ( .A(n35836), .B(n35837), .Z(n35835) );
  XNOR U35794 ( .A(n35834), .B(n35825), .Z(n35837) );
  IV U35795 ( .A(n35779), .Z(n35825) );
  XNOR U35796 ( .A(n35838), .B(n35818), .Z(n35779) );
  XNOR U35797 ( .A(n35839), .B(n35824), .Z(n35818) );
  XNOR U35798 ( .A(n35840), .B(n35841), .Z(n35824) );
  NOR U35799 ( .A(n35842), .B(n35843), .Z(n35841) );
  XOR U35800 ( .A(n35840), .B(n35844), .Z(n35842) );
  XNOR U35801 ( .A(n35823), .B(n35815), .Z(n35839) );
  XOR U35802 ( .A(n35845), .B(n35846), .Z(n35815) );
  AND U35803 ( .A(n35847), .B(n35848), .Z(n35846) );
  XOR U35804 ( .A(n35845), .B(n35849), .Z(n35847) );
  XNOR U35805 ( .A(n35850), .B(n35820), .Z(n35823) );
  XOR U35806 ( .A(n35851), .B(n35852), .Z(n35820) );
  AND U35807 ( .A(n35853), .B(n35854), .Z(n35852) );
  XNOR U35808 ( .A(n35855), .B(n35856), .Z(n35853) );
  IV U35809 ( .A(n35851), .Z(n35855) );
  XNOR U35810 ( .A(n35857), .B(n35858), .Z(n35850) );
  NOR U35811 ( .A(n35859), .B(n35860), .Z(n35858) );
  XNOR U35812 ( .A(n35857), .B(n35861), .Z(n35859) );
  XNOR U35813 ( .A(n35819), .B(n35826), .Z(n35838) );
  NOR U35814 ( .A(n35787), .B(n35862), .Z(n35826) );
  XOR U35815 ( .A(n35831), .B(n35830), .Z(n35819) );
  XNOR U35816 ( .A(n35863), .B(n35827), .Z(n35830) );
  XOR U35817 ( .A(n35864), .B(n35865), .Z(n35827) );
  AND U35818 ( .A(n35866), .B(n35867), .Z(n35865) );
  XNOR U35819 ( .A(n35868), .B(n35869), .Z(n35866) );
  IV U35820 ( .A(n35864), .Z(n35868) );
  XNOR U35821 ( .A(n35870), .B(n35871), .Z(n35863) );
  NOR U35822 ( .A(n35872), .B(n35873), .Z(n35871) );
  XNOR U35823 ( .A(n35870), .B(n35874), .Z(n35872) );
  XOR U35824 ( .A(n35875), .B(n35876), .Z(n35831) );
  NOR U35825 ( .A(n35877), .B(n35878), .Z(n35876) );
  XNOR U35826 ( .A(n35875), .B(n35879), .Z(n35877) );
  XNOR U35827 ( .A(n35776), .B(n35834), .Z(n35836) );
  XNOR U35828 ( .A(n35880), .B(n35881), .Z(n35776) );
  AND U35829 ( .A(n1326), .B(n35783), .Z(n35881) );
  XOR U35830 ( .A(n35880), .B(n35781), .Z(n35783) );
  AND U35831 ( .A(n35784), .B(n35787), .Z(n35834) );
  XOR U35832 ( .A(n35882), .B(n35862), .Z(n35787) );
  XNOR U35833 ( .A(p_input[1872]), .B(p_input[2048]), .Z(n35862) );
  XNOR U35834 ( .A(n35849), .B(n35848), .Z(n35882) );
  XNOR U35835 ( .A(n35883), .B(n35856), .Z(n35848) );
  XNOR U35836 ( .A(n35844), .B(n35843), .Z(n35856) );
  XNOR U35837 ( .A(n35884), .B(n35840), .Z(n35843) );
  XNOR U35838 ( .A(p_input[1882]), .B(p_input[2058]), .Z(n35840) );
  XOR U35839 ( .A(p_input[1883]), .B(n16732), .Z(n35884) );
  XOR U35840 ( .A(p_input[1884]), .B(p_input[2060]), .Z(n35844) );
  XOR U35841 ( .A(n35854), .B(n35885), .Z(n35883) );
  IV U35842 ( .A(n35845), .Z(n35885) );
  XOR U35843 ( .A(p_input[1873]), .B(p_input[2049]), .Z(n35845) );
  XNOR U35844 ( .A(n35886), .B(n35861), .Z(n35854) );
  XNOR U35845 ( .A(p_input[1887]), .B(n16735), .Z(n35861) );
  XOR U35846 ( .A(n35851), .B(n35860), .Z(n35886) );
  XOR U35847 ( .A(n35887), .B(n35857), .Z(n35860) );
  XOR U35848 ( .A(p_input[1885]), .B(p_input[2061]), .Z(n35857) );
  XOR U35849 ( .A(p_input[1886]), .B(n16737), .Z(n35887) );
  XOR U35850 ( .A(p_input[1881]), .B(p_input[2057]), .Z(n35851) );
  XOR U35851 ( .A(n35869), .B(n35867), .Z(n35849) );
  XNOR U35852 ( .A(n35888), .B(n35874), .Z(n35867) );
  XOR U35853 ( .A(p_input[1880]), .B(p_input[2056]), .Z(n35874) );
  XOR U35854 ( .A(n35864), .B(n35873), .Z(n35888) );
  XOR U35855 ( .A(n35889), .B(n35870), .Z(n35873) );
  XOR U35856 ( .A(p_input[1878]), .B(p_input[2054]), .Z(n35870) );
  XOR U35857 ( .A(p_input[1879]), .B(n17722), .Z(n35889) );
  XOR U35858 ( .A(p_input[1874]), .B(p_input[2050]), .Z(n35864) );
  XNOR U35859 ( .A(n35879), .B(n35878), .Z(n35869) );
  XOR U35860 ( .A(n35890), .B(n35875), .Z(n35878) );
  XOR U35861 ( .A(p_input[1875]), .B(p_input[2051]), .Z(n35875) );
  XOR U35862 ( .A(p_input[1876]), .B(n17724), .Z(n35890) );
  XOR U35863 ( .A(p_input[1877]), .B(p_input[2053]), .Z(n35879) );
  XNOR U35864 ( .A(n35891), .B(n35892), .Z(n35784) );
  AND U35865 ( .A(n1326), .B(n35893), .Z(n35892) );
  XNOR U35866 ( .A(n35894), .B(n35895), .Z(n1326) );
  AND U35867 ( .A(n35896), .B(n35897), .Z(n35895) );
  XOR U35868 ( .A(n35894), .B(n35794), .Z(n35897) );
  XNOR U35869 ( .A(n35894), .B(n35748), .Z(n35896) );
  XOR U35870 ( .A(n35898), .B(n35899), .Z(n35894) );
  AND U35871 ( .A(n35900), .B(n35901), .Z(n35899) );
  XOR U35872 ( .A(n35898), .B(n35758), .Z(n35900) );
  XOR U35873 ( .A(n35902), .B(n35903), .Z(n35737) );
  AND U35874 ( .A(n1330), .B(n35893), .Z(n35903) );
  XNOR U35875 ( .A(n35891), .B(n35902), .Z(n35893) );
  XNOR U35876 ( .A(n35904), .B(n35905), .Z(n1330) );
  AND U35877 ( .A(n35906), .B(n35907), .Z(n35905) );
  XNOR U35878 ( .A(n35908), .B(n35904), .Z(n35907) );
  IV U35879 ( .A(n35794), .Z(n35908) );
  XNOR U35880 ( .A(n35909), .B(n35910), .Z(n35794) );
  AND U35881 ( .A(n1333), .B(n35911), .Z(n35910) );
  XNOR U35882 ( .A(n35909), .B(n35912), .Z(n35911) );
  XNOR U35883 ( .A(n35748), .B(n35904), .Z(n35906) );
  XOR U35884 ( .A(n35913), .B(n35914), .Z(n35748) );
  AND U35885 ( .A(n1341), .B(n35915), .Z(n35914) );
  XOR U35886 ( .A(n35898), .B(n35916), .Z(n35904) );
  AND U35887 ( .A(n35917), .B(n35901), .Z(n35916) );
  XNOR U35888 ( .A(n35807), .B(n35898), .Z(n35901) );
  XNOR U35889 ( .A(n35918), .B(n35919), .Z(n35807) );
  AND U35890 ( .A(n1333), .B(n35920), .Z(n35919) );
  XOR U35891 ( .A(n35921), .B(n35918), .Z(n35920) );
  XNOR U35892 ( .A(n35922), .B(n35898), .Z(n35917) );
  IV U35893 ( .A(n35758), .Z(n35922) );
  XOR U35894 ( .A(n35923), .B(n35924), .Z(n35758) );
  AND U35895 ( .A(n1341), .B(n35925), .Z(n35924) );
  XOR U35896 ( .A(n35926), .B(n35927), .Z(n35898) );
  AND U35897 ( .A(n35928), .B(n35929), .Z(n35927) );
  XNOR U35898 ( .A(n35832), .B(n35926), .Z(n35929) );
  XNOR U35899 ( .A(n35930), .B(n35931), .Z(n35832) );
  AND U35900 ( .A(n1333), .B(n35932), .Z(n35931) );
  XNOR U35901 ( .A(n35933), .B(n35930), .Z(n35932) );
  XOR U35902 ( .A(n35926), .B(n35769), .Z(n35928) );
  XOR U35903 ( .A(n35934), .B(n35935), .Z(n35769) );
  AND U35904 ( .A(n1341), .B(n35936), .Z(n35935) );
  XOR U35905 ( .A(n35937), .B(n35938), .Z(n35926) );
  AND U35906 ( .A(n35939), .B(n35940), .Z(n35938) );
  XNOR U35907 ( .A(n35937), .B(n35880), .Z(n35940) );
  XNOR U35908 ( .A(n35941), .B(n35942), .Z(n35880) );
  AND U35909 ( .A(n1333), .B(n35943), .Z(n35942) );
  XOR U35910 ( .A(n35944), .B(n35941), .Z(n35943) );
  XNOR U35911 ( .A(n35945), .B(n35937), .Z(n35939) );
  IV U35912 ( .A(n35781), .Z(n35945) );
  XOR U35913 ( .A(n35946), .B(n35947), .Z(n35781) );
  AND U35914 ( .A(n1341), .B(n35948), .Z(n35947) );
  AND U35915 ( .A(n35902), .B(n35891), .Z(n35937) );
  XNOR U35916 ( .A(n35949), .B(n35950), .Z(n35891) );
  AND U35917 ( .A(n1333), .B(n35951), .Z(n35950) );
  XNOR U35918 ( .A(n35952), .B(n35949), .Z(n35951) );
  XNOR U35919 ( .A(n35953), .B(n35954), .Z(n1333) );
  AND U35920 ( .A(n35955), .B(n35956), .Z(n35954) );
  XOR U35921 ( .A(n35912), .B(n35953), .Z(n35956) );
  AND U35922 ( .A(n35957), .B(n35958), .Z(n35912) );
  XOR U35923 ( .A(n35953), .B(n35909), .Z(n35955) );
  XNOR U35924 ( .A(n35959), .B(n35960), .Z(n35909) );
  AND U35925 ( .A(n1337), .B(n35915), .Z(n35960) );
  XOR U35926 ( .A(n35913), .B(n35959), .Z(n35915) );
  XOR U35927 ( .A(n35961), .B(n35962), .Z(n35953) );
  AND U35928 ( .A(n35963), .B(n35964), .Z(n35962) );
  XNOR U35929 ( .A(n35961), .B(n35957), .Z(n35964) );
  IV U35930 ( .A(n35921), .Z(n35957) );
  XOR U35931 ( .A(n35965), .B(n35966), .Z(n35921) );
  XOR U35932 ( .A(n35967), .B(n35958), .Z(n35966) );
  AND U35933 ( .A(n35933), .B(n35968), .Z(n35958) );
  AND U35934 ( .A(n35969), .B(n35970), .Z(n35967) );
  XOR U35935 ( .A(n35971), .B(n35965), .Z(n35969) );
  XNOR U35936 ( .A(n35918), .B(n35961), .Z(n35963) );
  XNOR U35937 ( .A(n35972), .B(n35973), .Z(n35918) );
  AND U35938 ( .A(n1337), .B(n35925), .Z(n35973) );
  XOR U35939 ( .A(n35972), .B(n35923), .Z(n35925) );
  XOR U35940 ( .A(n35974), .B(n35975), .Z(n35961) );
  AND U35941 ( .A(n35976), .B(n35977), .Z(n35975) );
  XNOR U35942 ( .A(n35974), .B(n35933), .Z(n35977) );
  XOR U35943 ( .A(n35978), .B(n35970), .Z(n35933) );
  XNOR U35944 ( .A(n35979), .B(n35965), .Z(n35970) );
  XOR U35945 ( .A(n35980), .B(n35981), .Z(n35965) );
  AND U35946 ( .A(n35982), .B(n35983), .Z(n35981) );
  XOR U35947 ( .A(n35984), .B(n35980), .Z(n35982) );
  XNOR U35948 ( .A(n35985), .B(n35986), .Z(n35979) );
  AND U35949 ( .A(n35987), .B(n35988), .Z(n35986) );
  XOR U35950 ( .A(n35985), .B(n35989), .Z(n35987) );
  XNOR U35951 ( .A(n35971), .B(n35968), .Z(n35978) );
  AND U35952 ( .A(n35990), .B(n35991), .Z(n35968) );
  XOR U35953 ( .A(n35992), .B(n35993), .Z(n35971) );
  AND U35954 ( .A(n35994), .B(n35995), .Z(n35993) );
  XOR U35955 ( .A(n35992), .B(n35996), .Z(n35994) );
  XNOR U35956 ( .A(n35930), .B(n35974), .Z(n35976) );
  XNOR U35957 ( .A(n35997), .B(n35998), .Z(n35930) );
  AND U35958 ( .A(n1337), .B(n35936), .Z(n35998) );
  XOR U35959 ( .A(n35997), .B(n35934), .Z(n35936) );
  XOR U35960 ( .A(n35999), .B(n36000), .Z(n35974) );
  AND U35961 ( .A(n36001), .B(n36002), .Z(n36000) );
  XNOR U35962 ( .A(n35999), .B(n35990), .Z(n36002) );
  IV U35963 ( .A(n35944), .Z(n35990) );
  XNOR U35964 ( .A(n36003), .B(n35983), .Z(n35944) );
  XNOR U35965 ( .A(n36004), .B(n35989), .Z(n35983) );
  XNOR U35966 ( .A(n36005), .B(n36006), .Z(n35989) );
  NOR U35967 ( .A(n36007), .B(n36008), .Z(n36006) );
  XOR U35968 ( .A(n36005), .B(n36009), .Z(n36007) );
  XNOR U35969 ( .A(n35988), .B(n35980), .Z(n36004) );
  XOR U35970 ( .A(n36010), .B(n36011), .Z(n35980) );
  AND U35971 ( .A(n36012), .B(n36013), .Z(n36011) );
  XOR U35972 ( .A(n36010), .B(n36014), .Z(n36012) );
  XNOR U35973 ( .A(n36015), .B(n35985), .Z(n35988) );
  XOR U35974 ( .A(n36016), .B(n36017), .Z(n35985) );
  AND U35975 ( .A(n36018), .B(n36019), .Z(n36017) );
  XNOR U35976 ( .A(n36020), .B(n36021), .Z(n36018) );
  IV U35977 ( .A(n36016), .Z(n36020) );
  XNOR U35978 ( .A(n36022), .B(n36023), .Z(n36015) );
  NOR U35979 ( .A(n36024), .B(n36025), .Z(n36023) );
  XNOR U35980 ( .A(n36022), .B(n36026), .Z(n36024) );
  XNOR U35981 ( .A(n35984), .B(n35991), .Z(n36003) );
  NOR U35982 ( .A(n35952), .B(n36027), .Z(n35991) );
  XOR U35983 ( .A(n35996), .B(n35995), .Z(n35984) );
  XNOR U35984 ( .A(n36028), .B(n35992), .Z(n35995) );
  XOR U35985 ( .A(n36029), .B(n36030), .Z(n35992) );
  AND U35986 ( .A(n36031), .B(n36032), .Z(n36030) );
  XNOR U35987 ( .A(n36033), .B(n36034), .Z(n36031) );
  IV U35988 ( .A(n36029), .Z(n36033) );
  XNOR U35989 ( .A(n36035), .B(n36036), .Z(n36028) );
  NOR U35990 ( .A(n36037), .B(n36038), .Z(n36036) );
  XNOR U35991 ( .A(n36035), .B(n36039), .Z(n36037) );
  XOR U35992 ( .A(n36040), .B(n36041), .Z(n35996) );
  NOR U35993 ( .A(n36042), .B(n36043), .Z(n36041) );
  XNOR U35994 ( .A(n36040), .B(n36044), .Z(n36042) );
  XNOR U35995 ( .A(n35941), .B(n35999), .Z(n36001) );
  XNOR U35996 ( .A(n36045), .B(n36046), .Z(n35941) );
  AND U35997 ( .A(n1337), .B(n35948), .Z(n36046) );
  XOR U35998 ( .A(n36045), .B(n35946), .Z(n35948) );
  AND U35999 ( .A(n35949), .B(n35952), .Z(n35999) );
  XOR U36000 ( .A(n36047), .B(n36027), .Z(n35952) );
  XNOR U36001 ( .A(p_input[1888]), .B(p_input[2048]), .Z(n36027) );
  XNOR U36002 ( .A(n36014), .B(n36013), .Z(n36047) );
  XNOR U36003 ( .A(n36048), .B(n36021), .Z(n36013) );
  XNOR U36004 ( .A(n36009), .B(n36008), .Z(n36021) );
  XNOR U36005 ( .A(n36049), .B(n36005), .Z(n36008) );
  XNOR U36006 ( .A(p_input[1898]), .B(p_input[2058]), .Z(n36005) );
  XOR U36007 ( .A(p_input[1899]), .B(n16732), .Z(n36049) );
  XOR U36008 ( .A(p_input[1900]), .B(p_input[2060]), .Z(n36009) );
  XOR U36009 ( .A(n36019), .B(n36050), .Z(n36048) );
  IV U36010 ( .A(n36010), .Z(n36050) );
  XOR U36011 ( .A(p_input[1889]), .B(p_input[2049]), .Z(n36010) );
  XNOR U36012 ( .A(n36051), .B(n36026), .Z(n36019) );
  XNOR U36013 ( .A(p_input[1903]), .B(n16735), .Z(n36026) );
  XOR U36014 ( .A(n36016), .B(n36025), .Z(n36051) );
  XOR U36015 ( .A(n36052), .B(n36022), .Z(n36025) );
  XOR U36016 ( .A(p_input[1901]), .B(p_input[2061]), .Z(n36022) );
  XOR U36017 ( .A(p_input[1902]), .B(n16737), .Z(n36052) );
  XOR U36018 ( .A(p_input[1897]), .B(p_input[2057]), .Z(n36016) );
  XOR U36019 ( .A(n36034), .B(n36032), .Z(n36014) );
  XNOR U36020 ( .A(n36053), .B(n36039), .Z(n36032) );
  XOR U36021 ( .A(p_input[1896]), .B(p_input[2056]), .Z(n36039) );
  XOR U36022 ( .A(n36029), .B(n36038), .Z(n36053) );
  XOR U36023 ( .A(n36054), .B(n36035), .Z(n36038) );
  XOR U36024 ( .A(p_input[1894]), .B(p_input[2054]), .Z(n36035) );
  XOR U36025 ( .A(p_input[1895]), .B(n17722), .Z(n36054) );
  XOR U36026 ( .A(p_input[1890]), .B(p_input[2050]), .Z(n36029) );
  XNOR U36027 ( .A(n36044), .B(n36043), .Z(n36034) );
  XOR U36028 ( .A(n36055), .B(n36040), .Z(n36043) );
  XOR U36029 ( .A(p_input[1891]), .B(p_input[2051]), .Z(n36040) );
  XOR U36030 ( .A(p_input[1892]), .B(n17724), .Z(n36055) );
  XOR U36031 ( .A(p_input[1893]), .B(p_input[2053]), .Z(n36044) );
  XNOR U36032 ( .A(n36056), .B(n36057), .Z(n35949) );
  AND U36033 ( .A(n1337), .B(n36058), .Z(n36057) );
  XNOR U36034 ( .A(n36059), .B(n36060), .Z(n1337) );
  AND U36035 ( .A(n36061), .B(n36062), .Z(n36060) );
  XOR U36036 ( .A(n36059), .B(n35959), .Z(n36062) );
  XNOR U36037 ( .A(n36059), .B(n35913), .Z(n36061) );
  XOR U36038 ( .A(n36063), .B(n36064), .Z(n36059) );
  AND U36039 ( .A(n36065), .B(n36066), .Z(n36064) );
  XOR U36040 ( .A(n36063), .B(n35923), .Z(n36065) );
  XOR U36041 ( .A(n36067), .B(n36068), .Z(n35902) );
  AND U36042 ( .A(n1341), .B(n36058), .Z(n36068) );
  XNOR U36043 ( .A(n36056), .B(n36067), .Z(n36058) );
  XNOR U36044 ( .A(n36069), .B(n36070), .Z(n1341) );
  AND U36045 ( .A(n36071), .B(n36072), .Z(n36070) );
  XNOR U36046 ( .A(n36073), .B(n36069), .Z(n36072) );
  IV U36047 ( .A(n35959), .Z(n36073) );
  XNOR U36048 ( .A(n36074), .B(n36075), .Z(n35959) );
  AND U36049 ( .A(n1344), .B(n36076), .Z(n36075) );
  XNOR U36050 ( .A(n36074), .B(n36077), .Z(n36076) );
  XNOR U36051 ( .A(n35913), .B(n36069), .Z(n36071) );
  XOR U36052 ( .A(n36078), .B(n36079), .Z(n35913) );
  AND U36053 ( .A(n1352), .B(n36080), .Z(n36079) );
  XOR U36054 ( .A(n36063), .B(n36081), .Z(n36069) );
  AND U36055 ( .A(n36082), .B(n36066), .Z(n36081) );
  XNOR U36056 ( .A(n35972), .B(n36063), .Z(n36066) );
  XNOR U36057 ( .A(n36083), .B(n36084), .Z(n35972) );
  AND U36058 ( .A(n1344), .B(n36085), .Z(n36084) );
  XOR U36059 ( .A(n36086), .B(n36083), .Z(n36085) );
  XNOR U36060 ( .A(n36087), .B(n36063), .Z(n36082) );
  IV U36061 ( .A(n35923), .Z(n36087) );
  XOR U36062 ( .A(n36088), .B(n36089), .Z(n35923) );
  AND U36063 ( .A(n1352), .B(n36090), .Z(n36089) );
  XOR U36064 ( .A(n36091), .B(n36092), .Z(n36063) );
  AND U36065 ( .A(n36093), .B(n36094), .Z(n36092) );
  XNOR U36066 ( .A(n35997), .B(n36091), .Z(n36094) );
  XNOR U36067 ( .A(n36095), .B(n36096), .Z(n35997) );
  AND U36068 ( .A(n1344), .B(n36097), .Z(n36096) );
  XNOR U36069 ( .A(n36098), .B(n36095), .Z(n36097) );
  XOR U36070 ( .A(n36091), .B(n35934), .Z(n36093) );
  XOR U36071 ( .A(n36099), .B(n36100), .Z(n35934) );
  AND U36072 ( .A(n1352), .B(n36101), .Z(n36100) );
  XOR U36073 ( .A(n36102), .B(n36103), .Z(n36091) );
  AND U36074 ( .A(n36104), .B(n36105), .Z(n36103) );
  XNOR U36075 ( .A(n36102), .B(n36045), .Z(n36105) );
  XNOR U36076 ( .A(n36106), .B(n36107), .Z(n36045) );
  AND U36077 ( .A(n1344), .B(n36108), .Z(n36107) );
  XOR U36078 ( .A(n36109), .B(n36106), .Z(n36108) );
  XNOR U36079 ( .A(n36110), .B(n36102), .Z(n36104) );
  IV U36080 ( .A(n35946), .Z(n36110) );
  XOR U36081 ( .A(n36111), .B(n36112), .Z(n35946) );
  AND U36082 ( .A(n1352), .B(n36113), .Z(n36112) );
  AND U36083 ( .A(n36067), .B(n36056), .Z(n36102) );
  XNOR U36084 ( .A(n36114), .B(n36115), .Z(n36056) );
  AND U36085 ( .A(n1344), .B(n36116), .Z(n36115) );
  XNOR U36086 ( .A(n36117), .B(n36114), .Z(n36116) );
  XNOR U36087 ( .A(n36118), .B(n36119), .Z(n1344) );
  AND U36088 ( .A(n36120), .B(n36121), .Z(n36119) );
  XOR U36089 ( .A(n36077), .B(n36118), .Z(n36121) );
  AND U36090 ( .A(n36122), .B(n36123), .Z(n36077) );
  XOR U36091 ( .A(n36118), .B(n36074), .Z(n36120) );
  XNOR U36092 ( .A(n36124), .B(n36125), .Z(n36074) );
  AND U36093 ( .A(n1348), .B(n36080), .Z(n36125) );
  XOR U36094 ( .A(n36078), .B(n36124), .Z(n36080) );
  XOR U36095 ( .A(n36126), .B(n36127), .Z(n36118) );
  AND U36096 ( .A(n36128), .B(n36129), .Z(n36127) );
  XNOR U36097 ( .A(n36126), .B(n36122), .Z(n36129) );
  IV U36098 ( .A(n36086), .Z(n36122) );
  XOR U36099 ( .A(n36130), .B(n36131), .Z(n36086) );
  XOR U36100 ( .A(n36132), .B(n36123), .Z(n36131) );
  AND U36101 ( .A(n36098), .B(n36133), .Z(n36123) );
  AND U36102 ( .A(n36134), .B(n36135), .Z(n36132) );
  XOR U36103 ( .A(n36136), .B(n36130), .Z(n36134) );
  XNOR U36104 ( .A(n36083), .B(n36126), .Z(n36128) );
  XNOR U36105 ( .A(n36137), .B(n36138), .Z(n36083) );
  AND U36106 ( .A(n1348), .B(n36090), .Z(n36138) );
  XOR U36107 ( .A(n36137), .B(n36088), .Z(n36090) );
  XOR U36108 ( .A(n36139), .B(n36140), .Z(n36126) );
  AND U36109 ( .A(n36141), .B(n36142), .Z(n36140) );
  XNOR U36110 ( .A(n36139), .B(n36098), .Z(n36142) );
  XOR U36111 ( .A(n36143), .B(n36135), .Z(n36098) );
  XNOR U36112 ( .A(n36144), .B(n36130), .Z(n36135) );
  XOR U36113 ( .A(n36145), .B(n36146), .Z(n36130) );
  AND U36114 ( .A(n36147), .B(n36148), .Z(n36146) );
  XOR U36115 ( .A(n36149), .B(n36145), .Z(n36147) );
  XNOR U36116 ( .A(n36150), .B(n36151), .Z(n36144) );
  AND U36117 ( .A(n36152), .B(n36153), .Z(n36151) );
  XOR U36118 ( .A(n36150), .B(n36154), .Z(n36152) );
  XNOR U36119 ( .A(n36136), .B(n36133), .Z(n36143) );
  AND U36120 ( .A(n36155), .B(n36156), .Z(n36133) );
  XOR U36121 ( .A(n36157), .B(n36158), .Z(n36136) );
  AND U36122 ( .A(n36159), .B(n36160), .Z(n36158) );
  XOR U36123 ( .A(n36157), .B(n36161), .Z(n36159) );
  XNOR U36124 ( .A(n36095), .B(n36139), .Z(n36141) );
  XNOR U36125 ( .A(n36162), .B(n36163), .Z(n36095) );
  AND U36126 ( .A(n1348), .B(n36101), .Z(n36163) );
  XOR U36127 ( .A(n36162), .B(n36099), .Z(n36101) );
  XOR U36128 ( .A(n36164), .B(n36165), .Z(n36139) );
  AND U36129 ( .A(n36166), .B(n36167), .Z(n36165) );
  XNOR U36130 ( .A(n36164), .B(n36155), .Z(n36167) );
  IV U36131 ( .A(n36109), .Z(n36155) );
  XNOR U36132 ( .A(n36168), .B(n36148), .Z(n36109) );
  XNOR U36133 ( .A(n36169), .B(n36154), .Z(n36148) );
  XNOR U36134 ( .A(n36170), .B(n36171), .Z(n36154) );
  NOR U36135 ( .A(n36172), .B(n36173), .Z(n36171) );
  XOR U36136 ( .A(n36170), .B(n36174), .Z(n36172) );
  XNOR U36137 ( .A(n36153), .B(n36145), .Z(n36169) );
  XOR U36138 ( .A(n36175), .B(n36176), .Z(n36145) );
  AND U36139 ( .A(n36177), .B(n36178), .Z(n36176) );
  XOR U36140 ( .A(n36175), .B(n36179), .Z(n36177) );
  XNOR U36141 ( .A(n36180), .B(n36150), .Z(n36153) );
  XOR U36142 ( .A(n36181), .B(n36182), .Z(n36150) );
  AND U36143 ( .A(n36183), .B(n36184), .Z(n36182) );
  XNOR U36144 ( .A(n36185), .B(n36186), .Z(n36183) );
  IV U36145 ( .A(n36181), .Z(n36185) );
  XNOR U36146 ( .A(n36187), .B(n36188), .Z(n36180) );
  NOR U36147 ( .A(n36189), .B(n36190), .Z(n36188) );
  XNOR U36148 ( .A(n36187), .B(n36191), .Z(n36189) );
  XNOR U36149 ( .A(n36149), .B(n36156), .Z(n36168) );
  NOR U36150 ( .A(n36117), .B(n36192), .Z(n36156) );
  XOR U36151 ( .A(n36161), .B(n36160), .Z(n36149) );
  XNOR U36152 ( .A(n36193), .B(n36157), .Z(n36160) );
  XOR U36153 ( .A(n36194), .B(n36195), .Z(n36157) );
  AND U36154 ( .A(n36196), .B(n36197), .Z(n36195) );
  XNOR U36155 ( .A(n36198), .B(n36199), .Z(n36196) );
  IV U36156 ( .A(n36194), .Z(n36198) );
  XNOR U36157 ( .A(n36200), .B(n36201), .Z(n36193) );
  NOR U36158 ( .A(n36202), .B(n36203), .Z(n36201) );
  XNOR U36159 ( .A(n36200), .B(n36204), .Z(n36202) );
  XOR U36160 ( .A(n36205), .B(n36206), .Z(n36161) );
  NOR U36161 ( .A(n36207), .B(n36208), .Z(n36206) );
  XNOR U36162 ( .A(n36205), .B(n36209), .Z(n36207) );
  XNOR U36163 ( .A(n36106), .B(n36164), .Z(n36166) );
  XNOR U36164 ( .A(n36210), .B(n36211), .Z(n36106) );
  AND U36165 ( .A(n1348), .B(n36113), .Z(n36211) );
  XOR U36166 ( .A(n36210), .B(n36111), .Z(n36113) );
  AND U36167 ( .A(n36114), .B(n36117), .Z(n36164) );
  XOR U36168 ( .A(n36212), .B(n36192), .Z(n36117) );
  XNOR U36169 ( .A(p_input[1904]), .B(p_input[2048]), .Z(n36192) );
  XNOR U36170 ( .A(n36179), .B(n36178), .Z(n36212) );
  XNOR U36171 ( .A(n36213), .B(n36186), .Z(n36178) );
  XNOR U36172 ( .A(n36174), .B(n36173), .Z(n36186) );
  XNOR U36173 ( .A(n36214), .B(n36170), .Z(n36173) );
  XNOR U36174 ( .A(p_input[1914]), .B(p_input[2058]), .Z(n36170) );
  XOR U36175 ( .A(p_input[1915]), .B(n16732), .Z(n36214) );
  XOR U36176 ( .A(p_input[1916]), .B(p_input[2060]), .Z(n36174) );
  XOR U36177 ( .A(n36184), .B(n36215), .Z(n36213) );
  IV U36178 ( .A(n36175), .Z(n36215) );
  XOR U36179 ( .A(p_input[1905]), .B(p_input[2049]), .Z(n36175) );
  XNOR U36180 ( .A(n36216), .B(n36191), .Z(n36184) );
  XNOR U36181 ( .A(p_input[1919]), .B(n16735), .Z(n36191) );
  XOR U36182 ( .A(n36181), .B(n36190), .Z(n36216) );
  XOR U36183 ( .A(n36217), .B(n36187), .Z(n36190) );
  XOR U36184 ( .A(p_input[1917]), .B(p_input[2061]), .Z(n36187) );
  XOR U36185 ( .A(p_input[1918]), .B(n16737), .Z(n36217) );
  XOR U36186 ( .A(p_input[1913]), .B(p_input[2057]), .Z(n36181) );
  XOR U36187 ( .A(n36199), .B(n36197), .Z(n36179) );
  XNOR U36188 ( .A(n36218), .B(n36204), .Z(n36197) );
  XOR U36189 ( .A(p_input[1912]), .B(p_input[2056]), .Z(n36204) );
  XOR U36190 ( .A(n36194), .B(n36203), .Z(n36218) );
  XOR U36191 ( .A(n36219), .B(n36200), .Z(n36203) );
  XOR U36192 ( .A(p_input[1910]), .B(p_input[2054]), .Z(n36200) );
  XOR U36193 ( .A(p_input[1911]), .B(n17722), .Z(n36219) );
  XOR U36194 ( .A(p_input[1906]), .B(p_input[2050]), .Z(n36194) );
  XNOR U36195 ( .A(n36209), .B(n36208), .Z(n36199) );
  XOR U36196 ( .A(n36220), .B(n36205), .Z(n36208) );
  XOR U36197 ( .A(p_input[1907]), .B(p_input[2051]), .Z(n36205) );
  XOR U36198 ( .A(p_input[1908]), .B(n17724), .Z(n36220) );
  XOR U36199 ( .A(p_input[1909]), .B(p_input[2053]), .Z(n36209) );
  XNOR U36200 ( .A(n36221), .B(n36222), .Z(n36114) );
  AND U36201 ( .A(n1348), .B(n36223), .Z(n36222) );
  XNOR U36202 ( .A(n36224), .B(n36225), .Z(n1348) );
  AND U36203 ( .A(n36226), .B(n36227), .Z(n36225) );
  XOR U36204 ( .A(n36224), .B(n36124), .Z(n36227) );
  XNOR U36205 ( .A(n36224), .B(n36078), .Z(n36226) );
  XOR U36206 ( .A(n36228), .B(n36229), .Z(n36224) );
  AND U36207 ( .A(n36230), .B(n36231), .Z(n36229) );
  XOR U36208 ( .A(n36228), .B(n36088), .Z(n36230) );
  XOR U36209 ( .A(n36232), .B(n36233), .Z(n36067) );
  AND U36210 ( .A(n1352), .B(n36223), .Z(n36233) );
  XNOR U36211 ( .A(n36221), .B(n36232), .Z(n36223) );
  XNOR U36212 ( .A(n36234), .B(n36235), .Z(n1352) );
  AND U36213 ( .A(n36236), .B(n36237), .Z(n36235) );
  XNOR U36214 ( .A(n36238), .B(n36234), .Z(n36237) );
  IV U36215 ( .A(n36124), .Z(n36238) );
  XNOR U36216 ( .A(n36239), .B(n36240), .Z(n36124) );
  AND U36217 ( .A(n1355), .B(n36241), .Z(n36240) );
  XNOR U36218 ( .A(n36239), .B(n36242), .Z(n36241) );
  XNOR U36219 ( .A(n36078), .B(n36234), .Z(n36236) );
  XNOR U36220 ( .A(n36243), .B(n36244), .Z(n36078) );
  AND U36221 ( .A(n1363), .B(n36245), .Z(n36244) );
  XNOR U36222 ( .A(n36246), .B(n36247), .Z(n36245) );
  XOR U36223 ( .A(n36228), .B(n36248), .Z(n36234) );
  AND U36224 ( .A(n36249), .B(n36231), .Z(n36248) );
  XNOR U36225 ( .A(n36137), .B(n36228), .Z(n36231) );
  XNOR U36226 ( .A(n36250), .B(n36251), .Z(n36137) );
  AND U36227 ( .A(n1355), .B(n36252), .Z(n36251) );
  XOR U36228 ( .A(n36253), .B(n36250), .Z(n36252) );
  XNOR U36229 ( .A(n36254), .B(n36228), .Z(n36249) );
  IV U36230 ( .A(n36088), .Z(n36254) );
  XOR U36231 ( .A(n36255), .B(n36256), .Z(n36088) );
  AND U36232 ( .A(n1363), .B(n36257), .Z(n36256) );
  XOR U36233 ( .A(n36258), .B(n36259), .Z(n36228) );
  AND U36234 ( .A(n36260), .B(n36261), .Z(n36259) );
  XNOR U36235 ( .A(n36162), .B(n36258), .Z(n36261) );
  XNOR U36236 ( .A(n36262), .B(n36263), .Z(n36162) );
  AND U36237 ( .A(n1355), .B(n36264), .Z(n36263) );
  XNOR U36238 ( .A(n36265), .B(n36262), .Z(n36264) );
  XOR U36239 ( .A(n36258), .B(n36099), .Z(n36260) );
  XOR U36240 ( .A(n36266), .B(n36267), .Z(n36099) );
  AND U36241 ( .A(n1363), .B(n36268), .Z(n36267) );
  XOR U36242 ( .A(n36269), .B(n36270), .Z(n36258) );
  AND U36243 ( .A(n36271), .B(n36272), .Z(n36270) );
  XNOR U36244 ( .A(n36269), .B(n36210), .Z(n36272) );
  XNOR U36245 ( .A(n36273), .B(n36274), .Z(n36210) );
  AND U36246 ( .A(n1355), .B(n36275), .Z(n36274) );
  XOR U36247 ( .A(n36276), .B(n36273), .Z(n36275) );
  XNOR U36248 ( .A(n36277), .B(n36269), .Z(n36271) );
  IV U36249 ( .A(n36111), .Z(n36277) );
  XOR U36250 ( .A(n36278), .B(n36279), .Z(n36111) );
  AND U36251 ( .A(n1363), .B(n36280), .Z(n36279) );
  AND U36252 ( .A(n36232), .B(n36221), .Z(n36269) );
  XNOR U36253 ( .A(n36281), .B(n36282), .Z(n36221) );
  AND U36254 ( .A(n1355), .B(n36283), .Z(n36282) );
  XNOR U36255 ( .A(n36284), .B(n36281), .Z(n36283) );
  XNOR U36256 ( .A(n36285), .B(n36286), .Z(n1355) );
  AND U36257 ( .A(n36287), .B(n36288), .Z(n36286) );
  XOR U36258 ( .A(n36242), .B(n36285), .Z(n36288) );
  AND U36259 ( .A(n36289), .B(n36290), .Z(n36242) );
  XOR U36260 ( .A(n36285), .B(n36239), .Z(n36287) );
  XOR U36261 ( .A(n36246), .B(n36291), .Z(n36239) );
  AND U36262 ( .A(n1359), .B(n36292), .Z(n36291) );
  XOR U36263 ( .A(n36246), .B(n36243), .Z(n36292) );
  XOR U36264 ( .A(n36293), .B(n36294), .Z(n36285) );
  AND U36265 ( .A(n36295), .B(n36296), .Z(n36294) );
  XNOR U36266 ( .A(n36293), .B(n36289), .Z(n36296) );
  IV U36267 ( .A(n36253), .Z(n36289) );
  XOR U36268 ( .A(n36297), .B(n36298), .Z(n36253) );
  XOR U36269 ( .A(n36299), .B(n36290), .Z(n36298) );
  AND U36270 ( .A(n36265), .B(n36300), .Z(n36290) );
  AND U36271 ( .A(n36301), .B(n36302), .Z(n36299) );
  XOR U36272 ( .A(n36303), .B(n36297), .Z(n36301) );
  XNOR U36273 ( .A(n36250), .B(n36293), .Z(n36295) );
  XNOR U36274 ( .A(n36304), .B(n36305), .Z(n36250) );
  AND U36275 ( .A(n1359), .B(n36257), .Z(n36305) );
  XOR U36276 ( .A(n36304), .B(n36255), .Z(n36257) );
  XOR U36277 ( .A(n36306), .B(n36307), .Z(n36293) );
  AND U36278 ( .A(n36308), .B(n36309), .Z(n36307) );
  XNOR U36279 ( .A(n36306), .B(n36265), .Z(n36309) );
  XOR U36280 ( .A(n36310), .B(n36302), .Z(n36265) );
  XNOR U36281 ( .A(n36311), .B(n36297), .Z(n36302) );
  XOR U36282 ( .A(n36312), .B(n36313), .Z(n36297) );
  AND U36283 ( .A(n36314), .B(n36315), .Z(n36313) );
  XOR U36284 ( .A(n36316), .B(n36312), .Z(n36314) );
  XNOR U36285 ( .A(n36317), .B(n36318), .Z(n36311) );
  AND U36286 ( .A(n36319), .B(n36320), .Z(n36318) );
  XOR U36287 ( .A(n36317), .B(n36321), .Z(n36319) );
  XNOR U36288 ( .A(n36303), .B(n36300), .Z(n36310) );
  AND U36289 ( .A(n36322), .B(n36323), .Z(n36300) );
  XOR U36290 ( .A(n36324), .B(n36325), .Z(n36303) );
  AND U36291 ( .A(n36326), .B(n36327), .Z(n36325) );
  XOR U36292 ( .A(n36324), .B(n36328), .Z(n36326) );
  XNOR U36293 ( .A(n36262), .B(n36306), .Z(n36308) );
  XNOR U36294 ( .A(n36329), .B(n36330), .Z(n36262) );
  AND U36295 ( .A(n1359), .B(n36268), .Z(n36330) );
  XOR U36296 ( .A(n36329), .B(n36266), .Z(n36268) );
  XOR U36297 ( .A(n36331), .B(n36332), .Z(n36306) );
  AND U36298 ( .A(n36333), .B(n36334), .Z(n36332) );
  XNOR U36299 ( .A(n36331), .B(n36322), .Z(n36334) );
  IV U36300 ( .A(n36276), .Z(n36322) );
  XNOR U36301 ( .A(n36335), .B(n36315), .Z(n36276) );
  XNOR U36302 ( .A(n36336), .B(n36321), .Z(n36315) );
  XNOR U36303 ( .A(n36337), .B(n36338), .Z(n36321) );
  NOR U36304 ( .A(n36339), .B(n36340), .Z(n36338) );
  XOR U36305 ( .A(n36337), .B(n36341), .Z(n36339) );
  XNOR U36306 ( .A(n36320), .B(n36312), .Z(n36336) );
  XOR U36307 ( .A(n36342), .B(n36343), .Z(n36312) );
  AND U36308 ( .A(n36344), .B(n36345), .Z(n36343) );
  XOR U36309 ( .A(n36342), .B(n36346), .Z(n36344) );
  XNOR U36310 ( .A(n36347), .B(n36317), .Z(n36320) );
  XOR U36311 ( .A(n36348), .B(n36349), .Z(n36317) );
  AND U36312 ( .A(n36350), .B(n36351), .Z(n36349) );
  XNOR U36313 ( .A(n36352), .B(n36353), .Z(n36350) );
  IV U36314 ( .A(n36348), .Z(n36352) );
  XNOR U36315 ( .A(n36354), .B(n36355), .Z(n36347) );
  NOR U36316 ( .A(n36356), .B(n36357), .Z(n36355) );
  XNOR U36317 ( .A(n36354), .B(n36358), .Z(n36356) );
  XNOR U36318 ( .A(n36316), .B(n36323), .Z(n36335) );
  NOR U36319 ( .A(n36284), .B(n36359), .Z(n36323) );
  XOR U36320 ( .A(n36328), .B(n36327), .Z(n36316) );
  XNOR U36321 ( .A(n36360), .B(n36324), .Z(n36327) );
  XOR U36322 ( .A(n36361), .B(n36362), .Z(n36324) );
  AND U36323 ( .A(n36363), .B(n36364), .Z(n36362) );
  XNOR U36324 ( .A(n36365), .B(n36366), .Z(n36363) );
  IV U36325 ( .A(n36361), .Z(n36365) );
  XNOR U36326 ( .A(n36367), .B(n36368), .Z(n36360) );
  NOR U36327 ( .A(n36369), .B(n36370), .Z(n36368) );
  XNOR U36328 ( .A(n36367), .B(n36371), .Z(n36369) );
  XOR U36329 ( .A(n36372), .B(n36373), .Z(n36328) );
  NOR U36330 ( .A(n36374), .B(n36375), .Z(n36373) );
  XNOR U36331 ( .A(n36372), .B(n36376), .Z(n36374) );
  XNOR U36332 ( .A(n36273), .B(n36331), .Z(n36333) );
  XNOR U36333 ( .A(n36377), .B(n36378), .Z(n36273) );
  AND U36334 ( .A(n1359), .B(n36280), .Z(n36378) );
  XOR U36335 ( .A(n36377), .B(n36278), .Z(n36280) );
  AND U36336 ( .A(n36281), .B(n36284), .Z(n36331) );
  XOR U36337 ( .A(n36379), .B(n36359), .Z(n36284) );
  XNOR U36338 ( .A(p_input[1920]), .B(p_input[2048]), .Z(n36359) );
  XNOR U36339 ( .A(n36346), .B(n36345), .Z(n36379) );
  XNOR U36340 ( .A(n36380), .B(n36353), .Z(n36345) );
  XNOR U36341 ( .A(n36341), .B(n36340), .Z(n36353) );
  XNOR U36342 ( .A(n36381), .B(n36337), .Z(n36340) );
  XNOR U36343 ( .A(p_input[1930]), .B(p_input[2058]), .Z(n36337) );
  XOR U36344 ( .A(p_input[1931]), .B(n16732), .Z(n36381) );
  XOR U36345 ( .A(p_input[1932]), .B(p_input[2060]), .Z(n36341) );
  XOR U36346 ( .A(n36351), .B(n36382), .Z(n36380) );
  IV U36347 ( .A(n36342), .Z(n36382) );
  XOR U36348 ( .A(p_input[1921]), .B(p_input[2049]), .Z(n36342) );
  XNOR U36349 ( .A(n36383), .B(n36358), .Z(n36351) );
  XNOR U36350 ( .A(p_input[1935]), .B(n16735), .Z(n36358) );
  XOR U36351 ( .A(n36348), .B(n36357), .Z(n36383) );
  XOR U36352 ( .A(n36384), .B(n36354), .Z(n36357) );
  XOR U36353 ( .A(p_input[1933]), .B(p_input[2061]), .Z(n36354) );
  XOR U36354 ( .A(p_input[1934]), .B(n16737), .Z(n36384) );
  XOR U36355 ( .A(p_input[1929]), .B(p_input[2057]), .Z(n36348) );
  XOR U36356 ( .A(n36366), .B(n36364), .Z(n36346) );
  XNOR U36357 ( .A(n36385), .B(n36371), .Z(n36364) );
  XOR U36358 ( .A(p_input[1928]), .B(p_input[2056]), .Z(n36371) );
  XOR U36359 ( .A(n36361), .B(n36370), .Z(n36385) );
  XOR U36360 ( .A(n36386), .B(n36367), .Z(n36370) );
  XOR U36361 ( .A(p_input[1926]), .B(p_input[2054]), .Z(n36367) );
  XOR U36362 ( .A(p_input[1927]), .B(n17722), .Z(n36386) );
  XOR U36363 ( .A(p_input[1922]), .B(p_input[2050]), .Z(n36361) );
  XNOR U36364 ( .A(n36376), .B(n36375), .Z(n36366) );
  XOR U36365 ( .A(n36387), .B(n36372), .Z(n36375) );
  XOR U36366 ( .A(p_input[1923]), .B(p_input[2051]), .Z(n36372) );
  XOR U36367 ( .A(p_input[1924]), .B(n17724), .Z(n36387) );
  XOR U36368 ( .A(p_input[1925]), .B(p_input[2053]), .Z(n36376) );
  XNOR U36369 ( .A(n36388), .B(n36389), .Z(n36281) );
  AND U36370 ( .A(n1359), .B(n36390), .Z(n36389) );
  XNOR U36371 ( .A(n36391), .B(n36392), .Z(n1359) );
  AND U36372 ( .A(n36393), .B(n36394), .Z(n36392) );
  XNOR U36373 ( .A(n36391), .B(n36246), .Z(n36394) );
  XOR U36374 ( .A(n36391), .B(n36243), .Z(n36393) );
  XOR U36375 ( .A(n36395), .B(n36396), .Z(n36391) );
  AND U36376 ( .A(n36397), .B(n36398), .Z(n36396) );
  XOR U36377 ( .A(n36395), .B(n36255), .Z(n36397) );
  XOR U36378 ( .A(n36399), .B(n36400), .Z(n36232) );
  AND U36379 ( .A(n1363), .B(n36390), .Z(n36400) );
  XNOR U36380 ( .A(n36388), .B(n36399), .Z(n36390) );
  XNOR U36381 ( .A(n36401), .B(n36402), .Z(n1363) );
  AND U36382 ( .A(n36403), .B(n36404), .Z(n36402) );
  XNOR U36383 ( .A(n36246), .B(n36401), .Z(n36404) );
  XOR U36384 ( .A(n36405), .B(n36406), .Z(n36246) );
  AND U36385 ( .A(n36407), .B(n1366), .Z(n36406) );
  NOR U36386 ( .A(n36408), .B(n36405), .Z(n36407) );
  XOR U36387 ( .A(n36401), .B(n36243), .Z(n36403) );
  IV U36388 ( .A(n36247), .Z(n36243) );
  AND U36389 ( .A(n36409), .B(n36410), .Z(n36247) );
  XOR U36390 ( .A(n36395), .B(n36411), .Z(n36401) );
  AND U36391 ( .A(n36412), .B(n36398), .Z(n36411) );
  XNOR U36392 ( .A(n36304), .B(n36395), .Z(n36398) );
  XNOR U36393 ( .A(n36413), .B(n36414), .Z(n36304) );
  AND U36394 ( .A(n1366), .B(n36415), .Z(n36414) );
  XOR U36395 ( .A(n36416), .B(n36413), .Z(n36415) );
  XNOR U36396 ( .A(n36417), .B(n36395), .Z(n36412) );
  IV U36397 ( .A(n36255), .Z(n36417) );
  XOR U36398 ( .A(n36418), .B(n36419), .Z(n36255) );
  AND U36399 ( .A(n1374), .B(n36420), .Z(n36419) );
  XOR U36400 ( .A(n36421), .B(n36422), .Z(n36395) );
  AND U36401 ( .A(n36423), .B(n36424), .Z(n36422) );
  XNOR U36402 ( .A(n36329), .B(n36421), .Z(n36424) );
  XNOR U36403 ( .A(n36425), .B(n36426), .Z(n36329) );
  AND U36404 ( .A(n1366), .B(n36427), .Z(n36426) );
  XNOR U36405 ( .A(n36428), .B(n36425), .Z(n36427) );
  XOR U36406 ( .A(n36421), .B(n36266), .Z(n36423) );
  XOR U36407 ( .A(n36429), .B(n36430), .Z(n36266) );
  AND U36408 ( .A(n1374), .B(n36431), .Z(n36430) );
  XOR U36409 ( .A(n36432), .B(n36433), .Z(n36421) );
  AND U36410 ( .A(n36434), .B(n36435), .Z(n36433) );
  XNOR U36411 ( .A(n36432), .B(n36377), .Z(n36435) );
  XNOR U36412 ( .A(n36436), .B(n36437), .Z(n36377) );
  AND U36413 ( .A(n1366), .B(n36438), .Z(n36437) );
  XOR U36414 ( .A(n36439), .B(n36436), .Z(n36438) );
  XNOR U36415 ( .A(n36440), .B(n36432), .Z(n36434) );
  IV U36416 ( .A(n36278), .Z(n36440) );
  XOR U36417 ( .A(n36441), .B(n36442), .Z(n36278) );
  AND U36418 ( .A(n1374), .B(n36443), .Z(n36442) );
  AND U36419 ( .A(n36399), .B(n36388), .Z(n36432) );
  XNOR U36420 ( .A(n36444), .B(n36445), .Z(n36388) );
  AND U36421 ( .A(n1366), .B(n36446), .Z(n36445) );
  XNOR U36422 ( .A(n36447), .B(n36444), .Z(n36446) );
  XNOR U36423 ( .A(n36448), .B(n36449), .Z(n1366) );
  AND U36424 ( .A(n36450), .B(n36451), .Z(n36449) );
  XOR U36425 ( .A(n36408), .B(n36448), .Z(n36451) );
  AND U36426 ( .A(n36452), .B(n36453), .Z(n36408) );
  XOR U36427 ( .A(n36405), .B(n36448), .Z(n36450) );
  NOR U36428 ( .A(n36409), .B(n36410), .Z(n36405) );
  XOR U36429 ( .A(n36454), .B(n36455), .Z(n36448) );
  AND U36430 ( .A(n36456), .B(n36457), .Z(n36455) );
  XNOR U36431 ( .A(n36454), .B(n36452), .Z(n36457) );
  IV U36432 ( .A(n36416), .Z(n36452) );
  XOR U36433 ( .A(n36458), .B(n36459), .Z(n36416) );
  XOR U36434 ( .A(n36460), .B(n36453), .Z(n36459) );
  AND U36435 ( .A(n36428), .B(n36461), .Z(n36453) );
  AND U36436 ( .A(n36462), .B(n36463), .Z(n36460) );
  XOR U36437 ( .A(n36464), .B(n36458), .Z(n36462) );
  XNOR U36438 ( .A(n36413), .B(n36454), .Z(n36456) );
  XNOR U36439 ( .A(n36465), .B(n36466), .Z(n36413) );
  AND U36440 ( .A(n1370), .B(n36420), .Z(n36466) );
  XOR U36441 ( .A(n36465), .B(n36418), .Z(n36420) );
  XOR U36442 ( .A(n36467), .B(n36468), .Z(n36454) );
  AND U36443 ( .A(n36469), .B(n36470), .Z(n36468) );
  XNOR U36444 ( .A(n36467), .B(n36428), .Z(n36470) );
  XOR U36445 ( .A(n36471), .B(n36463), .Z(n36428) );
  XNOR U36446 ( .A(n36472), .B(n36458), .Z(n36463) );
  XOR U36447 ( .A(n36473), .B(n36474), .Z(n36458) );
  AND U36448 ( .A(n36475), .B(n36476), .Z(n36474) );
  XOR U36449 ( .A(n36477), .B(n36473), .Z(n36475) );
  XNOR U36450 ( .A(n36478), .B(n36479), .Z(n36472) );
  AND U36451 ( .A(n36480), .B(n36481), .Z(n36479) );
  XOR U36452 ( .A(n36478), .B(n36482), .Z(n36480) );
  XNOR U36453 ( .A(n36464), .B(n36461), .Z(n36471) );
  AND U36454 ( .A(n36483), .B(n36484), .Z(n36461) );
  XOR U36455 ( .A(n36485), .B(n36486), .Z(n36464) );
  AND U36456 ( .A(n36487), .B(n36488), .Z(n36486) );
  XOR U36457 ( .A(n36485), .B(n36489), .Z(n36487) );
  XNOR U36458 ( .A(n36425), .B(n36467), .Z(n36469) );
  XNOR U36459 ( .A(n36490), .B(n36491), .Z(n36425) );
  AND U36460 ( .A(n1370), .B(n36431), .Z(n36491) );
  XOR U36461 ( .A(n36490), .B(n36429), .Z(n36431) );
  XOR U36462 ( .A(n36492), .B(n36493), .Z(n36467) );
  AND U36463 ( .A(n36494), .B(n36495), .Z(n36493) );
  XNOR U36464 ( .A(n36492), .B(n36483), .Z(n36495) );
  IV U36465 ( .A(n36439), .Z(n36483) );
  XNOR U36466 ( .A(n36496), .B(n36476), .Z(n36439) );
  XNOR U36467 ( .A(n36497), .B(n36482), .Z(n36476) );
  XNOR U36468 ( .A(n36498), .B(n36499), .Z(n36482) );
  NOR U36469 ( .A(n36500), .B(n36501), .Z(n36499) );
  XOR U36470 ( .A(n36498), .B(n36502), .Z(n36500) );
  XNOR U36471 ( .A(n36481), .B(n36473), .Z(n36497) );
  XOR U36472 ( .A(n36503), .B(n36504), .Z(n36473) );
  AND U36473 ( .A(n36505), .B(n36506), .Z(n36504) );
  XOR U36474 ( .A(n36503), .B(n36507), .Z(n36505) );
  XNOR U36475 ( .A(n36508), .B(n36478), .Z(n36481) );
  XOR U36476 ( .A(n36509), .B(n36510), .Z(n36478) );
  AND U36477 ( .A(n36511), .B(n36512), .Z(n36510) );
  XNOR U36478 ( .A(n36513), .B(n36514), .Z(n36511) );
  IV U36479 ( .A(n36509), .Z(n36513) );
  XNOR U36480 ( .A(n36515), .B(n36516), .Z(n36508) );
  NOR U36481 ( .A(n36517), .B(n36518), .Z(n36516) );
  XNOR U36482 ( .A(n36515), .B(n36519), .Z(n36517) );
  XNOR U36483 ( .A(n36477), .B(n36484), .Z(n36496) );
  NOR U36484 ( .A(n36447), .B(n36520), .Z(n36484) );
  XOR U36485 ( .A(n36489), .B(n36488), .Z(n36477) );
  XNOR U36486 ( .A(n36521), .B(n36485), .Z(n36488) );
  XOR U36487 ( .A(n36522), .B(n36523), .Z(n36485) );
  AND U36488 ( .A(n36524), .B(n36525), .Z(n36523) );
  XNOR U36489 ( .A(n36526), .B(n36527), .Z(n36524) );
  IV U36490 ( .A(n36522), .Z(n36526) );
  XNOR U36491 ( .A(n36528), .B(n36529), .Z(n36521) );
  NOR U36492 ( .A(n36530), .B(n36531), .Z(n36529) );
  XNOR U36493 ( .A(n36528), .B(n36532), .Z(n36530) );
  XOR U36494 ( .A(n36533), .B(n36534), .Z(n36489) );
  NOR U36495 ( .A(n36535), .B(n36536), .Z(n36534) );
  XNOR U36496 ( .A(n36533), .B(n36537), .Z(n36535) );
  XNOR U36497 ( .A(n36436), .B(n36492), .Z(n36494) );
  XNOR U36498 ( .A(n36538), .B(n36539), .Z(n36436) );
  AND U36499 ( .A(n1370), .B(n36443), .Z(n36539) );
  XOR U36500 ( .A(n36538), .B(n36441), .Z(n36443) );
  AND U36501 ( .A(n36444), .B(n36447), .Z(n36492) );
  XOR U36502 ( .A(n36540), .B(n36520), .Z(n36447) );
  XNOR U36503 ( .A(p_input[1936]), .B(p_input[2048]), .Z(n36520) );
  XNOR U36504 ( .A(n36507), .B(n36506), .Z(n36540) );
  XNOR U36505 ( .A(n36541), .B(n36514), .Z(n36506) );
  XNOR U36506 ( .A(n36502), .B(n36501), .Z(n36514) );
  XNOR U36507 ( .A(n36542), .B(n36498), .Z(n36501) );
  XNOR U36508 ( .A(p_input[1946]), .B(p_input[2058]), .Z(n36498) );
  XOR U36509 ( .A(p_input[1947]), .B(n16732), .Z(n36542) );
  XOR U36510 ( .A(p_input[1948]), .B(p_input[2060]), .Z(n36502) );
  XOR U36511 ( .A(n36512), .B(n36543), .Z(n36541) );
  IV U36512 ( .A(n36503), .Z(n36543) );
  XOR U36513 ( .A(p_input[1937]), .B(p_input[2049]), .Z(n36503) );
  XNOR U36514 ( .A(n36544), .B(n36519), .Z(n36512) );
  XNOR U36515 ( .A(p_input[1951]), .B(n16735), .Z(n36519) );
  XOR U36516 ( .A(n36509), .B(n36518), .Z(n36544) );
  XOR U36517 ( .A(n36545), .B(n36515), .Z(n36518) );
  XOR U36518 ( .A(p_input[1949]), .B(p_input[2061]), .Z(n36515) );
  XOR U36519 ( .A(p_input[1950]), .B(n16737), .Z(n36545) );
  XOR U36520 ( .A(p_input[1945]), .B(p_input[2057]), .Z(n36509) );
  XOR U36521 ( .A(n36527), .B(n36525), .Z(n36507) );
  XNOR U36522 ( .A(n36546), .B(n36532), .Z(n36525) );
  XOR U36523 ( .A(p_input[1944]), .B(p_input[2056]), .Z(n36532) );
  XOR U36524 ( .A(n36522), .B(n36531), .Z(n36546) );
  XOR U36525 ( .A(n36547), .B(n36528), .Z(n36531) );
  XOR U36526 ( .A(p_input[1942]), .B(p_input[2054]), .Z(n36528) );
  XOR U36527 ( .A(p_input[1943]), .B(n17722), .Z(n36547) );
  XOR U36528 ( .A(p_input[1938]), .B(p_input[2050]), .Z(n36522) );
  XNOR U36529 ( .A(n36537), .B(n36536), .Z(n36527) );
  XOR U36530 ( .A(n36548), .B(n36533), .Z(n36536) );
  XOR U36531 ( .A(p_input[1939]), .B(p_input[2051]), .Z(n36533) );
  XOR U36532 ( .A(p_input[1940]), .B(n17724), .Z(n36548) );
  XOR U36533 ( .A(p_input[1941]), .B(p_input[2053]), .Z(n36537) );
  XNOR U36534 ( .A(n36549), .B(n36550), .Z(n36444) );
  AND U36535 ( .A(n1370), .B(n36551), .Z(n36550) );
  XNOR U36536 ( .A(n36552), .B(n36553), .Z(n1370) );
  NOR U36537 ( .A(n36554), .B(n36555), .Z(n36553) );
  XOR U36538 ( .A(n36410), .B(n36552), .Z(n36555) );
  NOR U36539 ( .A(n36552), .B(n36409), .Z(n36554) );
  XOR U36540 ( .A(n36556), .B(n36557), .Z(n36552) );
  AND U36541 ( .A(n36558), .B(n36559), .Z(n36557) );
  XOR U36542 ( .A(n36556), .B(n36418), .Z(n36558) );
  XOR U36543 ( .A(n36560), .B(n36561), .Z(n36399) );
  AND U36544 ( .A(n1374), .B(n36551), .Z(n36561) );
  XNOR U36545 ( .A(n36549), .B(n36560), .Z(n36551) );
  XNOR U36546 ( .A(n36562), .B(n36563), .Z(n1374) );
  NOR U36547 ( .A(n36564), .B(n36565), .Z(n36563) );
  XNOR U36548 ( .A(n36410), .B(n36566), .Z(n36565) );
  IV U36549 ( .A(n36562), .Z(n36566) );
  AND U36550 ( .A(n36567), .B(n36568), .Z(n36410) );
  NOR U36551 ( .A(n36562), .B(n36409), .Z(n36564) );
  AND U36552 ( .A(n36569), .B(n36570), .Z(n36409) );
  IV U36553 ( .A(n36571), .Z(n36569) );
  XOR U36554 ( .A(n36556), .B(n36572), .Z(n36562) );
  AND U36555 ( .A(n36573), .B(n36559), .Z(n36572) );
  XNOR U36556 ( .A(n36465), .B(n36556), .Z(n36559) );
  XNOR U36557 ( .A(n36574), .B(n36575), .Z(n36465) );
  AND U36558 ( .A(n1377), .B(n36576), .Z(n36575) );
  XOR U36559 ( .A(n36577), .B(n36574), .Z(n36576) );
  XNOR U36560 ( .A(n36578), .B(n36556), .Z(n36573) );
  IV U36561 ( .A(n36418), .Z(n36578) );
  XOR U36562 ( .A(n36579), .B(n36580), .Z(n36418) );
  AND U36563 ( .A(n1385), .B(n36581), .Z(n36580) );
  XOR U36564 ( .A(n36582), .B(n36583), .Z(n36556) );
  AND U36565 ( .A(n36584), .B(n36585), .Z(n36583) );
  XNOR U36566 ( .A(n36490), .B(n36582), .Z(n36585) );
  XNOR U36567 ( .A(n36586), .B(n36587), .Z(n36490) );
  AND U36568 ( .A(n1377), .B(n36588), .Z(n36587) );
  XNOR U36569 ( .A(n36589), .B(n36586), .Z(n36588) );
  XOR U36570 ( .A(n36582), .B(n36429), .Z(n36584) );
  XOR U36571 ( .A(n36590), .B(n36591), .Z(n36429) );
  AND U36572 ( .A(n1385), .B(n36592), .Z(n36591) );
  XOR U36573 ( .A(n36593), .B(n36594), .Z(n36582) );
  AND U36574 ( .A(n36595), .B(n36596), .Z(n36594) );
  XNOR U36575 ( .A(n36593), .B(n36538), .Z(n36596) );
  XNOR U36576 ( .A(n36597), .B(n36598), .Z(n36538) );
  AND U36577 ( .A(n1377), .B(n36599), .Z(n36598) );
  XOR U36578 ( .A(n36600), .B(n36597), .Z(n36599) );
  XNOR U36579 ( .A(n36601), .B(n36593), .Z(n36595) );
  IV U36580 ( .A(n36441), .Z(n36601) );
  XOR U36581 ( .A(n36602), .B(n36603), .Z(n36441) );
  AND U36582 ( .A(n1385), .B(n36604), .Z(n36603) );
  AND U36583 ( .A(n36560), .B(n36549), .Z(n36593) );
  XNOR U36584 ( .A(n36605), .B(n36606), .Z(n36549) );
  AND U36585 ( .A(n1377), .B(n36607), .Z(n36606) );
  XNOR U36586 ( .A(n36608), .B(n36605), .Z(n36607) );
  XNOR U36587 ( .A(n36609), .B(n36610), .Z(n1377) );
  NOR U36588 ( .A(n36611), .B(n36612), .Z(n36610) );
  XNOR U36589 ( .A(n36609), .B(n36571), .Z(n36612) );
  NOR U36590 ( .A(n36567), .B(n36568), .Z(n36571) );
  NOR U36591 ( .A(n36609), .B(n36570), .Z(n36611) );
  AND U36592 ( .A(n36613), .B(n36614), .Z(n36570) );
  XOR U36593 ( .A(n36615), .B(n36616), .Z(n36609) );
  AND U36594 ( .A(n36617), .B(n36618), .Z(n36616) );
  XNOR U36595 ( .A(n36615), .B(n36613), .Z(n36618) );
  IV U36596 ( .A(n36577), .Z(n36613) );
  XOR U36597 ( .A(n36619), .B(n36620), .Z(n36577) );
  XOR U36598 ( .A(n36621), .B(n36614), .Z(n36620) );
  AND U36599 ( .A(n36589), .B(n36622), .Z(n36614) );
  AND U36600 ( .A(n36623), .B(n36624), .Z(n36621) );
  XOR U36601 ( .A(n36625), .B(n36619), .Z(n36623) );
  XNOR U36602 ( .A(n36574), .B(n36615), .Z(n36617) );
  XNOR U36603 ( .A(n36626), .B(n36627), .Z(n36574) );
  AND U36604 ( .A(n1381), .B(n36581), .Z(n36627) );
  XOR U36605 ( .A(n36626), .B(n36579), .Z(n36581) );
  XOR U36606 ( .A(n36628), .B(n36629), .Z(n36615) );
  AND U36607 ( .A(n36630), .B(n36631), .Z(n36629) );
  XNOR U36608 ( .A(n36628), .B(n36589), .Z(n36631) );
  XOR U36609 ( .A(n36632), .B(n36624), .Z(n36589) );
  XNOR U36610 ( .A(n36633), .B(n36619), .Z(n36624) );
  XOR U36611 ( .A(n36634), .B(n36635), .Z(n36619) );
  AND U36612 ( .A(n36636), .B(n36637), .Z(n36635) );
  XOR U36613 ( .A(n36638), .B(n36634), .Z(n36636) );
  XNOR U36614 ( .A(n36639), .B(n36640), .Z(n36633) );
  AND U36615 ( .A(n36641), .B(n36642), .Z(n36640) );
  XOR U36616 ( .A(n36639), .B(n36643), .Z(n36641) );
  XNOR U36617 ( .A(n36625), .B(n36622), .Z(n36632) );
  AND U36618 ( .A(n36644), .B(n36645), .Z(n36622) );
  XOR U36619 ( .A(n36646), .B(n36647), .Z(n36625) );
  AND U36620 ( .A(n36648), .B(n36649), .Z(n36647) );
  XOR U36621 ( .A(n36646), .B(n36650), .Z(n36648) );
  XNOR U36622 ( .A(n36586), .B(n36628), .Z(n36630) );
  XNOR U36623 ( .A(n36651), .B(n36652), .Z(n36586) );
  AND U36624 ( .A(n1381), .B(n36592), .Z(n36652) );
  XOR U36625 ( .A(n36651), .B(n36590), .Z(n36592) );
  XOR U36626 ( .A(n36653), .B(n36654), .Z(n36628) );
  AND U36627 ( .A(n36655), .B(n36656), .Z(n36654) );
  XNOR U36628 ( .A(n36653), .B(n36644), .Z(n36656) );
  IV U36629 ( .A(n36600), .Z(n36644) );
  XNOR U36630 ( .A(n36657), .B(n36637), .Z(n36600) );
  XNOR U36631 ( .A(n36658), .B(n36643), .Z(n36637) );
  XNOR U36632 ( .A(n36659), .B(n36660), .Z(n36643) );
  NOR U36633 ( .A(n36661), .B(n36662), .Z(n36660) );
  XOR U36634 ( .A(n36659), .B(n36663), .Z(n36661) );
  XNOR U36635 ( .A(n36642), .B(n36634), .Z(n36658) );
  XOR U36636 ( .A(n36664), .B(n36665), .Z(n36634) );
  AND U36637 ( .A(n36666), .B(n36667), .Z(n36665) );
  XOR U36638 ( .A(n36664), .B(n36668), .Z(n36666) );
  XNOR U36639 ( .A(n36669), .B(n36639), .Z(n36642) );
  XOR U36640 ( .A(n36670), .B(n36671), .Z(n36639) );
  AND U36641 ( .A(n36672), .B(n36673), .Z(n36671) );
  XNOR U36642 ( .A(n36674), .B(n36675), .Z(n36672) );
  IV U36643 ( .A(n36670), .Z(n36674) );
  XNOR U36644 ( .A(n36676), .B(n36677), .Z(n36669) );
  NOR U36645 ( .A(n36678), .B(n36679), .Z(n36677) );
  XNOR U36646 ( .A(n36676), .B(n36680), .Z(n36678) );
  XNOR U36647 ( .A(n36638), .B(n36645), .Z(n36657) );
  NOR U36648 ( .A(n36608), .B(n36681), .Z(n36645) );
  XOR U36649 ( .A(n36650), .B(n36649), .Z(n36638) );
  XNOR U36650 ( .A(n36682), .B(n36646), .Z(n36649) );
  XOR U36651 ( .A(n36683), .B(n36684), .Z(n36646) );
  AND U36652 ( .A(n36685), .B(n36686), .Z(n36684) );
  XNOR U36653 ( .A(n36687), .B(n36688), .Z(n36685) );
  IV U36654 ( .A(n36683), .Z(n36687) );
  XNOR U36655 ( .A(n36689), .B(n36690), .Z(n36682) );
  NOR U36656 ( .A(n36691), .B(n36692), .Z(n36690) );
  XNOR U36657 ( .A(n36689), .B(n36693), .Z(n36691) );
  XOR U36658 ( .A(n36694), .B(n36695), .Z(n36650) );
  NOR U36659 ( .A(n36696), .B(n36697), .Z(n36695) );
  XNOR U36660 ( .A(n36694), .B(n36698), .Z(n36696) );
  XNOR U36661 ( .A(n36597), .B(n36653), .Z(n36655) );
  XNOR U36662 ( .A(n36699), .B(n36700), .Z(n36597) );
  AND U36663 ( .A(n1381), .B(n36604), .Z(n36700) );
  XOR U36664 ( .A(n36699), .B(n36602), .Z(n36604) );
  AND U36665 ( .A(n36605), .B(n36608), .Z(n36653) );
  XOR U36666 ( .A(n36701), .B(n36681), .Z(n36608) );
  XNOR U36667 ( .A(p_input[1952]), .B(p_input[2048]), .Z(n36681) );
  XNOR U36668 ( .A(n36668), .B(n36667), .Z(n36701) );
  XNOR U36669 ( .A(n36702), .B(n36675), .Z(n36667) );
  XNOR U36670 ( .A(n36663), .B(n36662), .Z(n36675) );
  XNOR U36671 ( .A(n36703), .B(n36659), .Z(n36662) );
  XNOR U36672 ( .A(p_input[1962]), .B(p_input[2058]), .Z(n36659) );
  XOR U36673 ( .A(p_input[1963]), .B(n16732), .Z(n36703) );
  XOR U36674 ( .A(p_input[1964]), .B(p_input[2060]), .Z(n36663) );
  XOR U36675 ( .A(n36673), .B(n36704), .Z(n36702) );
  IV U36676 ( .A(n36664), .Z(n36704) );
  XOR U36677 ( .A(p_input[1953]), .B(p_input[2049]), .Z(n36664) );
  XNOR U36678 ( .A(n36705), .B(n36680), .Z(n36673) );
  XNOR U36679 ( .A(p_input[1967]), .B(n16735), .Z(n36680) );
  XOR U36680 ( .A(n36670), .B(n36679), .Z(n36705) );
  XOR U36681 ( .A(n36706), .B(n36676), .Z(n36679) );
  XOR U36682 ( .A(p_input[1965]), .B(p_input[2061]), .Z(n36676) );
  XOR U36683 ( .A(p_input[1966]), .B(n16737), .Z(n36706) );
  XOR U36684 ( .A(p_input[1961]), .B(p_input[2057]), .Z(n36670) );
  XOR U36685 ( .A(n36688), .B(n36686), .Z(n36668) );
  XNOR U36686 ( .A(n36707), .B(n36693), .Z(n36686) );
  XOR U36687 ( .A(p_input[1960]), .B(p_input[2056]), .Z(n36693) );
  XOR U36688 ( .A(n36683), .B(n36692), .Z(n36707) );
  XOR U36689 ( .A(n36708), .B(n36689), .Z(n36692) );
  XOR U36690 ( .A(p_input[1958]), .B(p_input[2054]), .Z(n36689) );
  XOR U36691 ( .A(p_input[1959]), .B(n17722), .Z(n36708) );
  XOR U36692 ( .A(p_input[1954]), .B(p_input[2050]), .Z(n36683) );
  XNOR U36693 ( .A(n36698), .B(n36697), .Z(n36688) );
  XOR U36694 ( .A(n36709), .B(n36694), .Z(n36697) );
  XOR U36695 ( .A(p_input[1955]), .B(p_input[2051]), .Z(n36694) );
  XOR U36696 ( .A(p_input[1956]), .B(n17724), .Z(n36709) );
  XOR U36697 ( .A(p_input[1957]), .B(p_input[2053]), .Z(n36698) );
  XNOR U36698 ( .A(n36710), .B(n36711), .Z(n36605) );
  AND U36699 ( .A(n1381), .B(n36712), .Z(n36711) );
  XNOR U36700 ( .A(n36713), .B(n36714), .Z(n1381) );
  NOR U36701 ( .A(n36715), .B(n36716), .Z(n36714) );
  XOR U36702 ( .A(n36568), .B(n36713), .Z(n36716) );
  NOR U36703 ( .A(n36713), .B(n36567), .Z(n36715) );
  XOR U36704 ( .A(n36717), .B(n36718), .Z(n36713) );
  AND U36705 ( .A(n36719), .B(n36720), .Z(n36718) );
  XOR U36706 ( .A(n36717), .B(n36579), .Z(n36719) );
  XOR U36707 ( .A(n36721), .B(n36722), .Z(n36560) );
  AND U36708 ( .A(n1385), .B(n36712), .Z(n36722) );
  XNOR U36709 ( .A(n36710), .B(n36721), .Z(n36712) );
  XNOR U36710 ( .A(n36723), .B(n36724), .Z(n1385) );
  NOR U36711 ( .A(n36725), .B(n36726), .Z(n36724) );
  XNOR U36712 ( .A(n36568), .B(n36727), .Z(n36726) );
  IV U36713 ( .A(n36723), .Z(n36727) );
  AND U36714 ( .A(n36728), .B(n36729), .Z(n36568) );
  NOR U36715 ( .A(n36723), .B(n36567), .Z(n36725) );
  AND U36716 ( .A(n36730), .B(n36731), .Z(n36567) );
  IV U36717 ( .A(n36732), .Z(n36730) );
  XOR U36718 ( .A(n36717), .B(n36733), .Z(n36723) );
  AND U36719 ( .A(n36734), .B(n36720), .Z(n36733) );
  XNOR U36720 ( .A(n36626), .B(n36717), .Z(n36720) );
  XNOR U36721 ( .A(n36735), .B(n36736), .Z(n36626) );
  AND U36722 ( .A(n1388), .B(n36737), .Z(n36736) );
  XOR U36723 ( .A(n36738), .B(n36735), .Z(n36737) );
  XNOR U36724 ( .A(n36739), .B(n36717), .Z(n36734) );
  IV U36725 ( .A(n36579), .Z(n36739) );
  XOR U36726 ( .A(n36740), .B(n36741), .Z(n36579) );
  AND U36727 ( .A(n1396), .B(n36742), .Z(n36741) );
  XOR U36728 ( .A(n36743), .B(n36744), .Z(n36717) );
  AND U36729 ( .A(n36745), .B(n36746), .Z(n36744) );
  XNOR U36730 ( .A(n36651), .B(n36743), .Z(n36746) );
  XNOR U36731 ( .A(n36747), .B(n36748), .Z(n36651) );
  AND U36732 ( .A(n1388), .B(n36749), .Z(n36748) );
  XNOR U36733 ( .A(n36750), .B(n36747), .Z(n36749) );
  XOR U36734 ( .A(n36743), .B(n36590), .Z(n36745) );
  XOR U36735 ( .A(n36751), .B(n36752), .Z(n36590) );
  AND U36736 ( .A(n1396), .B(n36753), .Z(n36752) );
  XOR U36737 ( .A(n36754), .B(n36755), .Z(n36743) );
  AND U36738 ( .A(n36756), .B(n36757), .Z(n36755) );
  XNOR U36739 ( .A(n36754), .B(n36699), .Z(n36757) );
  XNOR U36740 ( .A(n36758), .B(n36759), .Z(n36699) );
  AND U36741 ( .A(n1388), .B(n36760), .Z(n36759) );
  XOR U36742 ( .A(n36761), .B(n36758), .Z(n36760) );
  XNOR U36743 ( .A(n36762), .B(n36754), .Z(n36756) );
  IV U36744 ( .A(n36602), .Z(n36762) );
  XOR U36745 ( .A(n36763), .B(n36764), .Z(n36602) );
  AND U36746 ( .A(n1396), .B(n36765), .Z(n36764) );
  AND U36747 ( .A(n36721), .B(n36710), .Z(n36754) );
  XNOR U36748 ( .A(n36766), .B(n36767), .Z(n36710) );
  AND U36749 ( .A(n1388), .B(n36768), .Z(n36767) );
  XNOR U36750 ( .A(n36769), .B(n36766), .Z(n36768) );
  XNOR U36751 ( .A(n36770), .B(n36771), .Z(n1388) );
  NOR U36752 ( .A(n36772), .B(n36773), .Z(n36771) );
  XNOR U36753 ( .A(n36770), .B(n36732), .Z(n36773) );
  NOR U36754 ( .A(n36728), .B(n36729), .Z(n36732) );
  NOR U36755 ( .A(n36770), .B(n36731), .Z(n36772) );
  AND U36756 ( .A(n36774), .B(n36775), .Z(n36731) );
  XOR U36757 ( .A(n36776), .B(n36777), .Z(n36770) );
  AND U36758 ( .A(n36778), .B(n36779), .Z(n36777) );
  XNOR U36759 ( .A(n36776), .B(n36774), .Z(n36779) );
  IV U36760 ( .A(n36738), .Z(n36774) );
  XOR U36761 ( .A(n36780), .B(n36781), .Z(n36738) );
  XOR U36762 ( .A(n36782), .B(n36775), .Z(n36781) );
  AND U36763 ( .A(n36750), .B(n36783), .Z(n36775) );
  AND U36764 ( .A(n36784), .B(n36785), .Z(n36782) );
  XOR U36765 ( .A(n36786), .B(n36780), .Z(n36784) );
  XNOR U36766 ( .A(n36735), .B(n36776), .Z(n36778) );
  XNOR U36767 ( .A(n36787), .B(n36788), .Z(n36735) );
  AND U36768 ( .A(n1392), .B(n36742), .Z(n36788) );
  XOR U36769 ( .A(n36787), .B(n36740), .Z(n36742) );
  XOR U36770 ( .A(n36789), .B(n36790), .Z(n36776) );
  AND U36771 ( .A(n36791), .B(n36792), .Z(n36790) );
  XNOR U36772 ( .A(n36789), .B(n36750), .Z(n36792) );
  XOR U36773 ( .A(n36793), .B(n36785), .Z(n36750) );
  XNOR U36774 ( .A(n36794), .B(n36780), .Z(n36785) );
  XOR U36775 ( .A(n36795), .B(n36796), .Z(n36780) );
  AND U36776 ( .A(n36797), .B(n36798), .Z(n36796) );
  XOR U36777 ( .A(n36799), .B(n36795), .Z(n36797) );
  XNOR U36778 ( .A(n36800), .B(n36801), .Z(n36794) );
  AND U36779 ( .A(n36802), .B(n36803), .Z(n36801) );
  XOR U36780 ( .A(n36800), .B(n36804), .Z(n36802) );
  XNOR U36781 ( .A(n36786), .B(n36783), .Z(n36793) );
  AND U36782 ( .A(n36805), .B(n36806), .Z(n36783) );
  XOR U36783 ( .A(n36807), .B(n36808), .Z(n36786) );
  AND U36784 ( .A(n36809), .B(n36810), .Z(n36808) );
  XOR U36785 ( .A(n36807), .B(n36811), .Z(n36809) );
  XNOR U36786 ( .A(n36747), .B(n36789), .Z(n36791) );
  XNOR U36787 ( .A(n36812), .B(n36813), .Z(n36747) );
  AND U36788 ( .A(n1392), .B(n36753), .Z(n36813) );
  XOR U36789 ( .A(n36812), .B(n36751), .Z(n36753) );
  XOR U36790 ( .A(n36814), .B(n36815), .Z(n36789) );
  AND U36791 ( .A(n36816), .B(n36817), .Z(n36815) );
  XNOR U36792 ( .A(n36814), .B(n36805), .Z(n36817) );
  IV U36793 ( .A(n36761), .Z(n36805) );
  XNOR U36794 ( .A(n36818), .B(n36798), .Z(n36761) );
  XNOR U36795 ( .A(n36819), .B(n36804), .Z(n36798) );
  XNOR U36796 ( .A(n36820), .B(n36821), .Z(n36804) );
  NOR U36797 ( .A(n36822), .B(n36823), .Z(n36821) );
  XOR U36798 ( .A(n36820), .B(n36824), .Z(n36822) );
  XNOR U36799 ( .A(n36803), .B(n36795), .Z(n36819) );
  XOR U36800 ( .A(n36825), .B(n36826), .Z(n36795) );
  AND U36801 ( .A(n36827), .B(n36828), .Z(n36826) );
  XOR U36802 ( .A(n36825), .B(n36829), .Z(n36827) );
  XNOR U36803 ( .A(n36830), .B(n36800), .Z(n36803) );
  XOR U36804 ( .A(n36831), .B(n36832), .Z(n36800) );
  AND U36805 ( .A(n36833), .B(n36834), .Z(n36832) );
  XNOR U36806 ( .A(n36835), .B(n36836), .Z(n36833) );
  IV U36807 ( .A(n36831), .Z(n36835) );
  XNOR U36808 ( .A(n36837), .B(n36838), .Z(n36830) );
  NOR U36809 ( .A(n36839), .B(n36840), .Z(n36838) );
  XNOR U36810 ( .A(n36837), .B(n36841), .Z(n36839) );
  XNOR U36811 ( .A(n36799), .B(n36806), .Z(n36818) );
  NOR U36812 ( .A(n36769), .B(n36842), .Z(n36806) );
  XOR U36813 ( .A(n36811), .B(n36810), .Z(n36799) );
  XNOR U36814 ( .A(n36843), .B(n36807), .Z(n36810) );
  XOR U36815 ( .A(n36844), .B(n36845), .Z(n36807) );
  AND U36816 ( .A(n36846), .B(n36847), .Z(n36845) );
  XNOR U36817 ( .A(n36848), .B(n36849), .Z(n36846) );
  IV U36818 ( .A(n36844), .Z(n36848) );
  XNOR U36819 ( .A(n36850), .B(n36851), .Z(n36843) );
  NOR U36820 ( .A(n36852), .B(n36853), .Z(n36851) );
  XNOR U36821 ( .A(n36850), .B(n36854), .Z(n36852) );
  XOR U36822 ( .A(n36855), .B(n36856), .Z(n36811) );
  NOR U36823 ( .A(n36857), .B(n36858), .Z(n36856) );
  XNOR U36824 ( .A(n36855), .B(n36859), .Z(n36857) );
  XNOR U36825 ( .A(n36758), .B(n36814), .Z(n36816) );
  XNOR U36826 ( .A(n36860), .B(n36861), .Z(n36758) );
  AND U36827 ( .A(n1392), .B(n36765), .Z(n36861) );
  XOR U36828 ( .A(n36860), .B(n36763), .Z(n36765) );
  AND U36829 ( .A(n36766), .B(n36769), .Z(n36814) );
  XOR U36830 ( .A(n36862), .B(n36842), .Z(n36769) );
  XNOR U36831 ( .A(p_input[1968]), .B(p_input[2048]), .Z(n36842) );
  XNOR U36832 ( .A(n36829), .B(n36828), .Z(n36862) );
  XNOR U36833 ( .A(n36863), .B(n36836), .Z(n36828) );
  XNOR U36834 ( .A(n36824), .B(n36823), .Z(n36836) );
  XNOR U36835 ( .A(n36864), .B(n36820), .Z(n36823) );
  XNOR U36836 ( .A(p_input[1978]), .B(p_input[2058]), .Z(n36820) );
  XOR U36837 ( .A(p_input[1979]), .B(n16732), .Z(n36864) );
  XOR U36838 ( .A(p_input[1980]), .B(p_input[2060]), .Z(n36824) );
  XOR U36839 ( .A(n36834), .B(n36865), .Z(n36863) );
  IV U36840 ( .A(n36825), .Z(n36865) );
  XOR U36841 ( .A(p_input[1969]), .B(p_input[2049]), .Z(n36825) );
  XNOR U36842 ( .A(n36866), .B(n36841), .Z(n36834) );
  XNOR U36843 ( .A(p_input[1983]), .B(n16735), .Z(n36841) );
  XOR U36844 ( .A(n36831), .B(n36840), .Z(n36866) );
  XOR U36845 ( .A(n36867), .B(n36837), .Z(n36840) );
  XOR U36846 ( .A(p_input[1981]), .B(p_input[2061]), .Z(n36837) );
  XOR U36847 ( .A(p_input[1982]), .B(n16737), .Z(n36867) );
  XOR U36848 ( .A(p_input[1977]), .B(p_input[2057]), .Z(n36831) );
  XOR U36849 ( .A(n36849), .B(n36847), .Z(n36829) );
  XNOR U36850 ( .A(n36868), .B(n36854), .Z(n36847) );
  XOR U36851 ( .A(p_input[1976]), .B(p_input[2056]), .Z(n36854) );
  XOR U36852 ( .A(n36844), .B(n36853), .Z(n36868) );
  XOR U36853 ( .A(n36869), .B(n36850), .Z(n36853) );
  XOR U36854 ( .A(p_input[1974]), .B(p_input[2054]), .Z(n36850) );
  XOR U36855 ( .A(p_input[1975]), .B(n17722), .Z(n36869) );
  XOR U36856 ( .A(p_input[1970]), .B(p_input[2050]), .Z(n36844) );
  XNOR U36857 ( .A(n36859), .B(n36858), .Z(n36849) );
  XOR U36858 ( .A(n36870), .B(n36855), .Z(n36858) );
  XOR U36859 ( .A(p_input[1971]), .B(p_input[2051]), .Z(n36855) );
  XOR U36860 ( .A(p_input[1972]), .B(n17724), .Z(n36870) );
  XOR U36861 ( .A(p_input[1973]), .B(p_input[2053]), .Z(n36859) );
  XNOR U36862 ( .A(n36871), .B(n36872), .Z(n36766) );
  AND U36863 ( .A(n1392), .B(n36873), .Z(n36872) );
  XNOR U36864 ( .A(n36874), .B(n36875), .Z(n1392) );
  NOR U36865 ( .A(n36876), .B(n36877), .Z(n36875) );
  XOR U36866 ( .A(n36729), .B(n36874), .Z(n36877) );
  NOR U36867 ( .A(n36874), .B(n36728), .Z(n36876) );
  XOR U36868 ( .A(n36878), .B(n36879), .Z(n36874) );
  AND U36869 ( .A(n36880), .B(n36881), .Z(n36879) );
  XOR U36870 ( .A(n36878), .B(n36740), .Z(n36880) );
  XOR U36871 ( .A(n36882), .B(n36883), .Z(n36721) );
  AND U36872 ( .A(n1396), .B(n36873), .Z(n36883) );
  XNOR U36873 ( .A(n36871), .B(n36882), .Z(n36873) );
  XNOR U36874 ( .A(n36884), .B(n36885), .Z(n1396) );
  NOR U36875 ( .A(n36886), .B(n36887), .Z(n36885) );
  XNOR U36876 ( .A(n36729), .B(n36888), .Z(n36887) );
  IV U36877 ( .A(n36884), .Z(n36888) );
  AND U36878 ( .A(n36889), .B(n36890), .Z(n36729) );
  NOR U36879 ( .A(n36884), .B(n36728), .Z(n36886) );
  AND U36880 ( .A(n36891), .B(n36892), .Z(n36728) );
  IV U36881 ( .A(n36893), .Z(n36891) );
  XOR U36882 ( .A(n36878), .B(n36894), .Z(n36884) );
  AND U36883 ( .A(n36895), .B(n36881), .Z(n36894) );
  XNOR U36884 ( .A(n36787), .B(n36878), .Z(n36881) );
  XNOR U36885 ( .A(n36896), .B(n36897), .Z(n36787) );
  AND U36886 ( .A(n1399), .B(n36898), .Z(n36897) );
  XOR U36887 ( .A(n36899), .B(n36896), .Z(n36898) );
  XNOR U36888 ( .A(n36900), .B(n36878), .Z(n36895) );
  IV U36889 ( .A(n36740), .Z(n36900) );
  XOR U36890 ( .A(n36901), .B(n36902), .Z(n36740) );
  AND U36891 ( .A(n1407), .B(n36903), .Z(n36902) );
  XOR U36892 ( .A(n36904), .B(n36905), .Z(n36878) );
  AND U36893 ( .A(n36906), .B(n36907), .Z(n36905) );
  XNOR U36894 ( .A(n36812), .B(n36904), .Z(n36907) );
  XNOR U36895 ( .A(n36908), .B(n36909), .Z(n36812) );
  AND U36896 ( .A(n1399), .B(n36910), .Z(n36909) );
  XNOR U36897 ( .A(n36911), .B(n36908), .Z(n36910) );
  XOR U36898 ( .A(n36904), .B(n36751), .Z(n36906) );
  XOR U36899 ( .A(n36912), .B(n36913), .Z(n36751) );
  AND U36900 ( .A(n1407), .B(n36914), .Z(n36913) );
  XOR U36901 ( .A(n36915), .B(n36916), .Z(n36904) );
  AND U36902 ( .A(n36917), .B(n36918), .Z(n36916) );
  XNOR U36903 ( .A(n36915), .B(n36860), .Z(n36918) );
  XNOR U36904 ( .A(n36919), .B(n36920), .Z(n36860) );
  AND U36905 ( .A(n1399), .B(n36921), .Z(n36920) );
  XOR U36906 ( .A(n36922), .B(n36919), .Z(n36921) );
  XNOR U36907 ( .A(n36923), .B(n36915), .Z(n36917) );
  IV U36908 ( .A(n36763), .Z(n36923) );
  XOR U36909 ( .A(n36924), .B(n36925), .Z(n36763) );
  AND U36910 ( .A(n1407), .B(n36926), .Z(n36925) );
  AND U36911 ( .A(n36882), .B(n36871), .Z(n36915) );
  XNOR U36912 ( .A(n36927), .B(n36928), .Z(n36871) );
  AND U36913 ( .A(n1399), .B(n36929), .Z(n36928) );
  XNOR U36914 ( .A(n36930), .B(n36927), .Z(n36929) );
  XNOR U36915 ( .A(n36931), .B(n36932), .Z(n1399) );
  NOR U36916 ( .A(n36933), .B(n36934), .Z(n36932) );
  XNOR U36917 ( .A(n36931), .B(n36893), .Z(n36934) );
  NOR U36918 ( .A(n36889), .B(n36890), .Z(n36893) );
  NOR U36919 ( .A(n36931), .B(n36892), .Z(n36933) );
  AND U36920 ( .A(n36935), .B(n36936), .Z(n36892) );
  XOR U36921 ( .A(n36937), .B(n36938), .Z(n36931) );
  AND U36922 ( .A(n36939), .B(n36940), .Z(n36938) );
  XNOR U36923 ( .A(n36937), .B(n36935), .Z(n36940) );
  IV U36924 ( .A(n36899), .Z(n36935) );
  XOR U36925 ( .A(n36941), .B(n36942), .Z(n36899) );
  XOR U36926 ( .A(n36943), .B(n36936), .Z(n36942) );
  AND U36927 ( .A(n36911), .B(n36944), .Z(n36936) );
  AND U36928 ( .A(n36945), .B(n36946), .Z(n36943) );
  XOR U36929 ( .A(n36947), .B(n36941), .Z(n36945) );
  XNOR U36930 ( .A(n36896), .B(n36937), .Z(n36939) );
  XNOR U36931 ( .A(n36948), .B(n36949), .Z(n36896) );
  AND U36932 ( .A(n1403), .B(n36903), .Z(n36949) );
  XOR U36933 ( .A(n36948), .B(n36901), .Z(n36903) );
  XOR U36934 ( .A(n36950), .B(n36951), .Z(n36937) );
  AND U36935 ( .A(n36952), .B(n36953), .Z(n36951) );
  XNOR U36936 ( .A(n36950), .B(n36911), .Z(n36953) );
  XOR U36937 ( .A(n36954), .B(n36946), .Z(n36911) );
  XNOR U36938 ( .A(n36955), .B(n36941), .Z(n36946) );
  XOR U36939 ( .A(n36956), .B(n36957), .Z(n36941) );
  AND U36940 ( .A(n36958), .B(n36959), .Z(n36957) );
  XOR U36941 ( .A(n36960), .B(n36956), .Z(n36958) );
  XNOR U36942 ( .A(n36961), .B(n36962), .Z(n36955) );
  AND U36943 ( .A(n36963), .B(n36964), .Z(n36962) );
  XOR U36944 ( .A(n36961), .B(n36965), .Z(n36963) );
  XNOR U36945 ( .A(n36947), .B(n36944), .Z(n36954) );
  AND U36946 ( .A(n36966), .B(n36967), .Z(n36944) );
  XOR U36947 ( .A(n36968), .B(n36969), .Z(n36947) );
  AND U36948 ( .A(n36970), .B(n36971), .Z(n36969) );
  XOR U36949 ( .A(n36968), .B(n36972), .Z(n36970) );
  XNOR U36950 ( .A(n36908), .B(n36950), .Z(n36952) );
  XNOR U36951 ( .A(n36973), .B(n36974), .Z(n36908) );
  AND U36952 ( .A(n1403), .B(n36914), .Z(n36974) );
  XOR U36953 ( .A(n36973), .B(n36912), .Z(n36914) );
  XOR U36954 ( .A(n36975), .B(n36976), .Z(n36950) );
  AND U36955 ( .A(n36977), .B(n36978), .Z(n36976) );
  XNOR U36956 ( .A(n36975), .B(n36966), .Z(n36978) );
  IV U36957 ( .A(n36922), .Z(n36966) );
  XNOR U36958 ( .A(n36979), .B(n36959), .Z(n36922) );
  XNOR U36959 ( .A(n36980), .B(n36965), .Z(n36959) );
  XNOR U36960 ( .A(n36981), .B(n36982), .Z(n36965) );
  NOR U36961 ( .A(n36983), .B(n36984), .Z(n36982) );
  XOR U36962 ( .A(n36981), .B(n36985), .Z(n36983) );
  XNOR U36963 ( .A(n36964), .B(n36956), .Z(n36980) );
  XOR U36964 ( .A(n36986), .B(n36987), .Z(n36956) );
  AND U36965 ( .A(n36988), .B(n36989), .Z(n36987) );
  XOR U36966 ( .A(n36986), .B(n36990), .Z(n36988) );
  XNOR U36967 ( .A(n36991), .B(n36961), .Z(n36964) );
  XOR U36968 ( .A(n36992), .B(n36993), .Z(n36961) );
  AND U36969 ( .A(n36994), .B(n36995), .Z(n36993) );
  XNOR U36970 ( .A(n36996), .B(n36997), .Z(n36994) );
  IV U36971 ( .A(n36992), .Z(n36996) );
  XNOR U36972 ( .A(n36998), .B(n36999), .Z(n36991) );
  NOR U36973 ( .A(n37000), .B(n37001), .Z(n36999) );
  XNOR U36974 ( .A(n36998), .B(n37002), .Z(n37000) );
  XNOR U36975 ( .A(n36960), .B(n36967), .Z(n36979) );
  NOR U36976 ( .A(n36930), .B(n37003), .Z(n36967) );
  XOR U36977 ( .A(n36972), .B(n36971), .Z(n36960) );
  XNOR U36978 ( .A(n37004), .B(n36968), .Z(n36971) );
  XOR U36979 ( .A(n37005), .B(n37006), .Z(n36968) );
  AND U36980 ( .A(n37007), .B(n37008), .Z(n37006) );
  XNOR U36981 ( .A(n37009), .B(n37010), .Z(n37007) );
  IV U36982 ( .A(n37005), .Z(n37009) );
  XNOR U36983 ( .A(n37011), .B(n37012), .Z(n37004) );
  NOR U36984 ( .A(n37013), .B(n37014), .Z(n37012) );
  XNOR U36985 ( .A(n37011), .B(n37015), .Z(n37013) );
  XOR U36986 ( .A(n37016), .B(n37017), .Z(n36972) );
  NOR U36987 ( .A(n37018), .B(n37019), .Z(n37017) );
  XNOR U36988 ( .A(n37016), .B(n37020), .Z(n37018) );
  XNOR U36989 ( .A(n36919), .B(n36975), .Z(n36977) );
  XNOR U36990 ( .A(n37021), .B(n37022), .Z(n36919) );
  AND U36991 ( .A(n1403), .B(n36926), .Z(n37022) );
  XOR U36992 ( .A(n37021), .B(n36924), .Z(n36926) );
  AND U36993 ( .A(n36927), .B(n36930), .Z(n36975) );
  XOR U36994 ( .A(n37023), .B(n37003), .Z(n36930) );
  XNOR U36995 ( .A(p_input[1984]), .B(p_input[2048]), .Z(n37003) );
  XNOR U36996 ( .A(n36990), .B(n36989), .Z(n37023) );
  XNOR U36997 ( .A(n37024), .B(n36997), .Z(n36989) );
  XNOR U36998 ( .A(n36985), .B(n36984), .Z(n36997) );
  XNOR U36999 ( .A(n37025), .B(n36981), .Z(n36984) );
  XNOR U37000 ( .A(p_input[1994]), .B(p_input[2058]), .Z(n36981) );
  XOR U37001 ( .A(p_input[1995]), .B(n16732), .Z(n37025) );
  XOR U37002 ( .A(p_input[1996]), .B(p_input[2060]), .Z(n36985) );
  XOR U37003 ( .A(n36995), .B(n37026), .Z(n37024) );
  IV U37004 ( .A(n36986), .Z(n37026) );
  XOR U37005 ( .A(p_input[1985]), .B(p_input[2049]), .Z(n36986) );
  XNOR U37006 ( .A(n37027), .B(n37002), .Z(n36995) );
  XNOR U37007 ( .A(p_input[1999]), .B(n16735), .Z(n37002) );
  XOR U37008 ( .A(n36992), .B(n37001), .Z(n37027) );
  XOR U37009 ( .A(n37028), .B(n36998), .Z(n37001) );
  XOR U37010 ( .A(p_input[1997]), .B(p_input[2061]), .Z(n36998) );
  XOR U37011 ( .A(p_input[1998]), .B(n16737), .Z(n37028) );
  XOR U37012 ( .A(p_input[1993]), .B(p_input[2057]), .Z(n36992) );
  XOR U37013 ( .A(n37010), .B(n37008), .Z(n36990) );
  XNOR U37014 ( .A(n37029), .B(n37015), .Z(n37008) );
  XOR U37015 ( .A(p_input[1992]), .B(p_input[2056]), .Z(n37015) );
  XOR U37016 ( .A(n37005), .B(n37014), .Z(n37029) );
  XOR U37017 ( .A(n37030), .B(n37011), .Z(n37014) );
  XOR U37018 ( .A(p_input[1990]), .B(p_input[2054]), .Z(n37011) );
  XOR U37019 ( .A(p_input[1991]), .B(n17722), .Z(n37030) );
  XOR U37020 ( .A(p_input[1986]), .B(p_input[2050]), .Z(n37005) );
  XNOR U37021 ( .A(n37020), .B(n37019), .Z(n37010) );
  XOR U37022 ( .A(n37031), .B(n37016), .Z(n37019) );
  XOR U37023 ( .A(p_input[1987]), .B(p_input[2051]), .Z(n37016) );
  XOR U37024 ( .A(p_input[1988]), .B(n17724), .Z(n37031) );
  XOR U37025 ( .A(p_input[1989]), .B(p_input[2053]), .Z(n37020) );
  XNOR U37026 ( .A(n37032), .B(n37033), .Z(n36927) );
  AND U37027 ( .A(n1403), .B(n37034), .Z(n37033) );
  XNOR U37028 ( .A(n37035), .B(n37036), .Z(n1403) );
  NOR U37029 ( .A(n37037), .B(n37038), .Z(n37036) );
  XOR U37030 ( .A(n36890), .B(n37035), .Z(n37038) );
  NOR U37031 ( .A(n37035), .B(n36889), .Z(n37037) );
  XOR U37032 ( .A(n37039), .B(n37040), .Z(n37035) );
  AND U37033 ( .A(n37041), .B(n37042), .Z(n37040) );
  XOR U37034 ( .A(n37039), .B(n36901), .Z(n37041) );
  XOR U37035 ( .A(n37043), .B(n37044), .Z(n36882) );
  AND U37036 ( .A(n1407), .B(n37034), .Z(n37044) );
  XNOR U37037 ( .A(n37032), .B(n37043), .Z(n37034) );
  XNOR U37038 ( .A(n37045), .B(n37046), .Z(n1407) );
  NOR U37039 ( .A(n37047), .B(n37048), .Z(n37046) );
  XNOR U37040 ( .A(n36890), .B(n37049), .Z(n37048) );
  IV U37041 ( .A(n37045), .Z(n37049) );
  AND U37042 ( .A(n37050), .B(n37051), .Z(n36890) );
  NOR U37043 ( .A(n37045), .B(n36889), .Z(n37047) );
  AND U37044 ( .A(n37052), .B(n37053), .Z(n36889) );
  IV U37045 ( .A(n37054), .Z(n37052) );
  XOR U37046 ( .A(n37039), .B(n37055), .Z(n37045) );
  AND U37047 ( .A(n37056), .B(n37042), .Z(n37055) );
  XNOR U37048 ( .A(n36948), .B(n37039), .Z(n37042) );
  XNOR U37049 ( .A(n37057), .B(n37058), .Z(n36948) );
  AND U37050 ( .A(n1410), .B(n37059), .Z(n37058) );
  XOR U37051 ( .A(n37060), .B(n37057), .Z(n37059) );
  XNOR U37052 ( .A(n37061), .B(n37039), .Z(n37056) );
  IV U37053 ( .A(n36901), .Z(n37061) );
  XOR U37054 ( .A(n37062), .B(n37063), .Z(n36901) );
  AND U37055 ( .A(n1417), .B(n37064), .Z(n37063) );
  XOR U37056 ( .A(n37065), .B(n37066), .Z(n37039) );
  AND U37057 ( .A(n37067), .B(n37068), .Z(n37066) );
  XNOR U37058 ( .A(n36973), .B(n37065), .Z(n37068) );
  XNOR U37059 ( .A(n37069), .B(n37070), .Z(n36973) );
  AND U37060 ( .A(n1410), .B(n37071), .Z(n37070) );
  XNOR U37061 ( .A(n37072), .B(n37069), .Z(n37071) );
  XOR U37062 ( .A(n37065), .B(n36912), .Z(n37067) );
  XOR U37063 ( .A(n37073), .B(n37074), .Z(n36912) );
  AND U37064 ( .A(n1417), .B(n37075), .Z(n37074) );
  XOR U37065 ( .A(n37076), .B(n37077), .Z(n37065) );
  AND U37066 ( .A(n37078), .B(n37079), .Z(n37077) );
  XNOR U37067 ( .A(n37076), .B(n37021), .Z(n37079) );
  XNOR U37068 ( .A(n37080), .B(n37081), .Z(n37021) );
  AND U37069 ( .A(n1410), .B(n37082), .Z(n37081) );
  XOR U37070 ( .A(n37083), .B(n37080), .Z(n37082) );
  XNOR U37071 ( .A(n37084), .B(n37076), .Z(n37078) );
  IV U37072 ( .A(n36924), .Z(n37084) );
  XOR U37073 ( .A(n37085), .B(n37086), .Z(n36924) );
  AND U37074 ( .A(n1417), .B(n37087), .Z(n37086) );
  AND U37075 ( .A(n37043), .B(n37032), .Z(n37076) );
  XNOR U37076 ( .A(n37088), .B(n37089), .Z(n37032) );
  AND U37077 ( .A(n1410), .B(n37090), .Z(n37089) );
  XNOR U37078 ( .A(n37091), .B(n37088), .Z(n37090) );
  XNOR U37079 ( .A(n37092), .B(n37093), .Z(n1410) );
  NOR U37080 ( .A(n37094), .B(n37095), .Z(n37093) );
  XNOR U37081 ( .A(n37092), .B(n37054), .Z(n37095) );
  NOR U37082 ( .A(n37050), .B(n37051), .Z(n37054) );
  NOR U37083 ( .A(n37092), .B(n37053), .Z(n37094) );
  AND U37084 ( .A(n37096), .B(n37097), .Z(n37053) );
  XOR U37085 ( .A(n37098), .B(n37099), .Z(n37092) );
  AND U37086 ( .A(n37100), .B(n37101), .Z(n37099) );
  XNOR U37087 ( .A(n37098), .B(n37096), .Z(n37101) );
  IV U37088 ( .A(n37060), .Z(n37096) );
  XOR U37089 ( .A(n37102), .B(n37103), .Z(n37060) );
  XOR U37090 ( .A(n37104), .B(n37097), .Z(n37103) );
  AND U37091 ( .A(n37072), .B(n37105), .Z(n37097) );
  AND U37092 ( .A(n37106), .B(n37107), .Z(n37104) );
  XOR U37093 ( .A(n37108), .B(n37102), .Z(n37106) );
  XNOR U37094 ( .A(n37057), .B(n37098), .Z(n37100) );
  XNOR U37095 ( .A(n37109), .B(n37110), .Z(n37057) );
  AND U37096 ( .A(n1414), .B(n37064), .Z(n37110) );
  XOR U37097 ( .A(n37109), .B(n37062), .Z(n37064) );
  XOR U37098 ( .A(n37111), .B(n37112), .Z(n37098) );
  AND U37099 ( .A(n37113), .B(n37114), .Z(n37112) );
  XNOR U37100 ( .A(n37111), .B(n37072), .Z(n37114) );
  XOR U37101 ( .A(n37115), .B(n37107), .Z(n37072) );
  XNOR U37102 ( .A(n37116), .B(n37102), .Z(n37107) );
  XOR U37103 ( .A(n37117), .B(n37118), .Z(n37102) );
  AND U37104 ( .A(n37119), .B(n37120), .Z(n37118) );
  XOR U37105 ( .A(n37121), .B(n37117), .Z(n37119) );
  XNOR U37106 ( .A(n37122), .B(n37123), .Z(n37116) );
  AND U37107 ( .A(n37124), .B(n37125), .Z(n37123) );
  XOR U37108 ( .A(n37122), .B(n37126), .Z(n37124) );
  XNOR U37109 ( .A(n37108), .B(n37105), .Z(n37115) );
  AND U37110 ( .A(n37127), .B(n37128), .Z(n37105) );
  XOR U37111 ( .A(n37129), .B(n37130), .Z(n37108) );
  AND U37112 ( .A(n37131), .B(n37132), .Z(n37130) );
  XOR U37113 ( .A(n37129), .B(n37133), .Z(n37131) );
  XNOR U37114 ( .A(n37069), .B(n37111), .Z(n37113) );
  XNOR U37115 ( .A(n37134), .B(n37135), .Z(n37069) );
  AND U37116 ( .A(n1414), .B(n37075), .Z(n37135) );
  XOR U37117 ( .A(n37134), .B(n37073), .Z(n37075) );
  XOR U37118 ( .A(n37136), .B(n37137), .Z(n37111) );
  AND U37119 ( .A(n37138), .B(n37139), .Z(n37137) );
  XNOR U37120 ( .A(n37136), .B(n37127), .Z(n37139) );
  IV U37121 ( .A(n37083), .Z(n37127) );
  XNOR U37122 ( .A(n37140), .B(n37120), .Z(n37083) );
  XNOR U37123 ( .A(n37141), .B(n37126), .Z(n37120) );
  XNOR U37124 ( .A(n37142), .B(n37143), .Z(n37126) );
  NOR U37125 ( .A(n37144), .B(n37145), .Z(n37143) );
  XOR U37126 ( .A(n37142), .B(n37146), .Z(n37144) );
  XNOR U37127 ( .A(n37125), .B(n37117), .Z(n37141) );
  XOR U37128 ( .A(n37147), .B(n37148), .Z(n37117) );
  AND U37129 ( .A(n37149), .B(n37150), .Z(n37148) );
  XOR U37130 ( .A(n37147), .B(n37151), .Z(n37149) );
  XNOR U37131 ( .A(n37152), .B(n37122), .Z(n37125) );
  XOR U37132 ( .A(n37153), .B(n37154), .Z(n37122) );
  AND U37133 ( .A(n37155), .B(n37156), .Z(n37154) );
  XNOR U37134 ( .A(n37157), .B(n37158), .Z(n37155) );
  IV U37135 ( .A(n37153), .Z(n37157) );
  XNOR U37136 ( .A(n37159), .B(n37160), .Z(n37152) );
  NOR U37137 ( .A(n37161), .B(n37162), .Z(n37160) );
  XNOR U37138 ( .A(n37159), .B(n37163), .Z(n37161) );
  XNOR U37139 ( .A(n37121), .B(n37128), .Z(n37140) );
  NOR U37140 ( .A(n37091), .B(n37164), .Z(n37128) );
  XOR U37141 ( .A(n37133), .B(n37132), .Z(n37121) );
  XNOR U37142 ( .A(n37165), .B(n37129), .Z(n37132) );
  XOR U37143 ( .A(n37166), .B(n37167), .Z(n37129) );
  AND U37144 ( .A(n37168), .B(n37169), .Z(n37167) );
  XNOR U37145 ( .A(n37170), .B(n37171), .Z(n37168) );
  IV U37146 ( .A(n37166), .Z(n37170) );
  XNOR U37147 ( .A(n37172), .B(n37173), .Z(n37165) );
  NOR U37148 ( .A(n37174), .B(n37175), .Z(n37173) );
  XNOR U37149 ( .A(n37172), .B(n37176), .Z(n37174) );
  XOR U37150 ( .A(n37177), .B(n37178), .Z(n37133) );
  NOR U37151 ( .A(n37179), .B(n37180), .Z(n37178) );
  XNOR U37152 ( .A(n37177), .B(n37181), .Z(n37179) );
  XNOR U37153 ( .A(n37080), .B(n37136), .Z(n37138) );
  XNOR U37154 ( .A(n37182), .B(n37183), .Z(n37080) );
  AND U37155 ( .A(n1414), .B(n37087), .Z(n37183) );
  XOR U37156 ( .A(n37182), .B(n37085), .Z(n37087) );
  AND U37157 ( .A(n37088), .B(n37091), .Z(n37136) );
  XOR U37158 ( .A(n37184), .B(n37164), .Z(n37091) );
  XNOR U37159 ( .A(p_input[2000]), .B(p_input[2048]), .Z(n37164) );
  XNOR U37160 ( .A(n37151), .B(n37150), .Z(n37184) );
  XNOR U37161 ( .A(n37185), .B(n37158), .Z(n37150) );
  XNOR U37162 ( .A(n37146), .B(n37145), .Z(n37158) );
  XNOR U37163 ( .A(n37186), .B(n37142), .Z(n37145) );
  XNOR U37164 ( .A(p_input[2010]), .B(p_input[2058]), .Z(n37142) );
  XOR U37165 ( .A(p_input[2011]), .B(n16732), .Z(n37186) );
  XOR U37166 ( .A(p_input[2012]), .B(p_input[2060]), .Z(n37146) );
  XOR U37167 ( .A(n37156), .B(n37187), .Z(n37185) );
  IV U37168 ( .A(n37147), .Z(n37187) );
  XOR U37169 ( .A(p_input[2001]), .B(p_input[2049]), .Z(n37147) );
  XNOR U37170 ( .A(n37188), .B(n37163), .Z(n37156) );
  XNOR U37171 ( .A(p_input[2015]), .B(n16735), .Z(n37163) );
  IV U37172 ( .A(p_input[2063]), .Z(n16735) );
  XOR U37173 ( .A(n37153), .B(n37162), .Z(n37188) );
  XOR U37174 ( .A(n37189), .B(n37159), .Z(n37162) );
  XOR U37175 ( .A(p_input[2013]), .B(p_input[2061]), .Z(n37159) );
  XOR U37176 ( .A(p_input[2014]), .B(n16737), .Z(n37189) );
  XOR U37177 ( .A(p_input[2009]), .B(p_input[2057]), .Z(n37153) );
  XOR U37178 ( .A(n37171), .B(n37169), .Z(n37151) );
  XNOR U37179 ( .A(n37190), .B(n37176), .Z(n37169) );
  XOR U37180 ( .A(p_input[2008]), .B(p_input[2056]), .Z(n37176) );
  XOR U37181 ( .A(n37166), .B(n37175), .Z(n37190) );
  XOR U37182 ( .A(n37191), .B(n37172), .Z(n37175) );
  XOR U37183 ( .A(p_input[2006]), .B(p_input[2054]), .Z(n37172) );
  XOR U37184 ( .A(p_input[2007]), .B(n17722), .Z(n37191) );
  XOR U37185 ( .A(p_input[2002]), .B(p_input[2050]), .Z(n37166) );
  XNOR U37186 ( .A(n37181), .B(n37180), .Z(n37171) );
  XOR U37187 ( .A(n37192), .B(n37177), .Z(n37180) );
  XOR U37188 ( .A(p_input[2003]), .B(p_input[2051]), .Z(n37177) );
  XOR U37189 ( .A(p_input[2004]), .B(n17724), .Z(n37192) );
  XOR U37190 ( .A(p_input[2005]), .B(p_input[2053]), .Z(n37181) );
  XNOR U37191 ( .A(n37193), .B(n37194), .Z(n37088) );
  AND U37192 ( .A(n1414), .B(n37195), .Z(n37194) );
  XNOR U37193 ( .A(n37196), .B(n37197), .Z(n1414) );
  NOR U37194 ( .A(n37198), .B(n37199), .Z(n37197) );
  XOR U37195 ( .A(n37051), .B(n37196), .Z(n37199) );
  NOR U37196 ( .A(n37196), .B(n37050), .Z(n37198) );
  XOR U37197 ( .A(n37200), .B(n37201), .Z(n37196) );
  AND U37198 ( .A(n37202), .B(n37203), .Z(n37201) );
  XOR U37199 ( .A(n37200), .B(n37062), .Z(n37202) );
  XOR U37200 ( .A(n37204), .B(n37205), .Z(n37043) );
  AND U37201 ( .A(n1417), .B(n37195), .Z(n37205) );
  XOR U37202 ( .A(n37206), .B(n37204), .Z(n37195) );
  XNOR U37203 ( .A(n37207), .B(n37208), .Z(n1417) );
  NOR U37204 ( .A(n37209), .B(n37210), .Z(n37208) );
  XNOR U37205 ( .A(n37051), .B(n37211), .Z(n37210) );
  IV U37206 ( .A(n37207), .Z(n37211) );
  AND U37207 ( .A(n37062), .B(n37212), .Z(n37051) );
  NOR U37208 ( .A(n37207), .B(n37050), .Z(n37209) );
  AND U37209 ( .A(n37109), .B(n37213), .Z(n37050) );
  XOR U37210 ( .A(n37200), .B(n37214), .Z(n37207) );
  AND U37211 ( .A(n37215), .B(n37203), .Z(n37214) );
  XNOR U37212 ( .A(n37109), .B(n37200), .Z(n37203) );
  XNOR U37213 ( .A(n37216), .B(n37217), .Z(n37109) );
  XOR U37214 ( .A(n37218), .B(n37213), .Z(n37217) );
  AND U37215 ( .A(n37134), .B(n37219), .Z(n37213) );
  AND U37216 ( .A(n37220), .B(n37221), .Z(n37218) );
  XOR U37217 ( .A(n37222), .B(n37216), .Z(n37220) );
  XNOR U37218 ( .A(n37223), .B(n37200), .Z(n37215) );
  IV U37219 ( .A(n37062), .Z(n37223) );
  XNOR U37220 ( .A(n37224), .B(n37225), .Z(n37062) );
  XOR U37221 ( .A(n37226), .B(n37212), .Z(n37225) );
  AND U37222 ( .A(n37073), .B(n37227), .Z(n37212) );
  AND U37223 ( .A(n37228), .B(n37229), .Z(n37226) );
  XNOR U37224 ( .A(n37224), .B(n37230), .Z(n37228) );
  XOR U37225 ( .A(n37231), .B(n37232), .Z(n37200) );
  AND U37226 ( .A(n37233), .B(n37234), .Z(n37232) );
  XNOR U37227 ( .A(n37134), .B(n37231), .Z(n37234) );
  XOR U37228 ( .A(n37235), .B(n37221), .Z(n37134) );
  XNOR U37229 ( .A(n37236), .B(n37216), .Z(n37221) );
  XOR U37230 ( .A(n37237), .B(n37238), .Z(n37216) );
  AND U37231 ( .A(n37239), .B(n37240), .Z(n37238) );
  XOR U37232 ( .A(n37241), .B(n37237), .Z(n37239) );
  XNOR U37233 ( .A(n37242), .B(n37243), .Z(n37236) );
  AND U37234 ( .A(n37244), .B(n37245), .Z(n37243) );
  XOR U37235 ( .A(n37242), .B(n37246), .Z(n37244) );
  XNOR U37236 ( .A(n37222), .B(n37219), .Z(n37235) );
  AND U37237 ( .A(n37182), .B(n37247), .Z(n37219) );
  XOR U37238 ( .A(n37248), .B(n37249), .Z(n37222) );
  AND U37239 ( .A(n37250), .B(n37251), .Z(n37249) );
  XOR U37240 ( .A(n37248), .B(n37252), .Z(n37250) );
  XOR U37241 ( .A(n37231), .B(n37073), .Z(n37233) );
  XNOR U37242 ( .A(n37253), .B(n37230), .Z(n37073) );
  XNOR U37243 ( .A(n37254), .B(n37255), .Z(n37230) );
  AND U37244 ( .A(n37256), .B(n37257), .Z(n37255) );
  XOR U37245 ( .A(n37254), .B(n37258), .Z(n37256) );
  XNOR U37246 ( .A(n37229), .B(n37227), .Z(n37253) );
  AND U37247 ( .A(n37085), .B(n37259), .Z(n37227) );
  XNOR U37248 ( .A(n37260), .B(n37224), .Z(n37229) );
  XOR U37249 ( .A(n37261), .B(n37262), .Z(n37224) );
  AND U37250 ( .A(n37263), .B(n37264), .Z(n37262) );
  XOR U37251 ( .A(n37261), .B(n37265), .Z(n37263) );
  XNOR U37252 ( .A(n37266), .B(n37267), .Z(n37260) );
  AND U37253 ( .A(n37268), .B(n37269), .Z(n37267) );
  XNOR U37254 ( .A(n37266), .B(n37270), .Z(n37268) );
  XOR U37255 ( .A(n37271), .B(n37272), .Z(n37231) );
  AND U37256 ( .A(n37273), .B(n37274), .Z(n37272) );
  XNOR U37257 ( .A(n37271), .B(n37182), .Z(n37274) );
  XOR U37258 ( .A(n37275), .B(n37240), .Z(n37182) );
  XNOR U37259 ( .A(n37276), .B(n37246), .Z(n37240) );
  XOR U37260 ( .A(n37277), .B(n37278), .Z(n37246) );
  NOR U37261 ( .A(n37279), .B(n37280), .Z(n37278) );
  XNOR U37262 ( .A(n37277), .B(n37281), .Z(n37279) );
  XNOR U37263 ( .A(n37245), .B(n37237), .Z(n37276) );
  XOR U37264 ( .A(n37282), .B(n37283), .Z(n37237) );
  AND U37265 ( .A(n37284), .B(n37285), .Z(n37283) );
  XNOR U37266 ( .A(n37282), .B(n37286), .Z(n37284) );
  XNOR U37267 ( .A(n37287), .B(n37242), .Z(n37245) );
  XOR U37268 ( .A(n37288), .B(n37289), .Z(n37242) );
  AND U37269 ( .A(n37290), .B(n37291), .Z(n37289) );
  XOR U37270 ( .A(n37288), .B(n37292), .Z(n37290) );
  XNOR U37271 ( .A(n37293), .B(n37294), .Z(n37287) );
  NOR U37272 ( .A(n37295), .B(n37296), .Z(n37294) );
  XOR U37273 ( .A(n37293), .B(n37297), .Z(n37295) );
  XNOR U37274 ( .A(n37241), .B(n37247), .Z(n37275) );
  AND U37275 ( .A(n37206), .B(n37298), .Z(n37247) );
  IV U37276 ( .A(n37193), .Z(n37206) );
  XOR U37277 ( .A(n37252), .B(n37251), .Z(n37241) );
  XNOR U37278 ( .A(n37299), .B(n37248), .Z(n37251) );
  XOR U37279 ( .A(n37300), .B(n37301), .Z(n37248) );
  AND U37280 ( .A(n37302), .B(n37303), .Z(n37301) );
  XOR U37281 ( .A(n37300), .B(n37304), .Z(n37302) );
  XNOR U37282 ( .A(n37305), .B(n37306), .Z(n37299) );
  NOR U37283 ( .A(n37307), .B(n37308), .Z(n37306) );
  XNOR U37284 ( .A(n37305), .B(n37309), .Z(n37307) );
  XOR U37285 ( .A(n37310), .B(n37311), .Z(n37252) );
  NOR U37286 ( .A(n37312), .B(n37313), .Z(n37311) );
  XNOR U37287 ( .A(n37310), .B(n37314), .Z(n37312) );
  XNOR U37288 ( .A(n37315), .B(n37271), .Z(n37273) );
  IV U37289 ( .A(n37085), .Z(n37315) );
  XOR U37290 ( .A(n37316), .B(n37265), .Z(n37085) );
  XOR U37291 ( .A(n37258), .B(n37257), .Z(n37265) );
  XNOR U37292 ( .A(n37317), .B(n37254), .Z(n37257) );
  XOR U37293 ( .A(n37318), .B(n37319), .Z(n37254) );
  AND U37294 ( .A(n37320), .B(n37321), .Z(n37319) );
  XOR U37295 ( .A(n37318), .B(n37322), .Z(n37320) );
  XNOR U37296 ( .A(n37323), .B(n37324), .Z(n37317) );
  NOR U37297 ( .A(n37325), .B(n37326), .Z(n37324) );
  XNOR U37298 ( .A(n37323), .B(n37327), .Z(n37325) );
  XOR U37299 ( .A(n37328), .B(n37329), .Z(n37258) );
  NOR U37300 ( .A(n37330), .B(n37331), .Z(n37329) );
  XNOR U37301 ( .A(n37328), .B(n37332), .Z(n37330) );
  XNOR U37302 ( .A(n37264), .B(n37259), .Z(n37316) );
  AND U37303 ( .A(n37204), .B(n37333), .Z(n37259) );
  XOR U37304 ( .A(n37334), .B(n37270), .Z(n37264) );
  XNOR U37305 ( .A(n37335), .B(n37336), .Z(n37270) );
  NOR U37306 ( .A(n37337), .B(n37338), .Z(n37336) );
  XNOR U37307 ( .A(n37335), .B(n37339), .Z(n37337) );
  XNOR U37308 ( .A(n37269), .B(n37261), .Z(n37334) );
  XOR U37309 ( .A(n37340), .B(n37341), .Z(n37261) );
  AND U37310 ( .A(n37342), .B(n37343), .Z(n37341) );
  XOR U37311 ( .A(n37340), .B(n37344), .Z(n37342) );
  XNOR U37312 ( .A(n37345), .B(n37266), .Z(n37269) );
  XOR U37313 ( .A(n37346), .B(n37347), .Z(n37266) );
  AND U37314 ( .A(n37348), .B(n37349), .Z(n37347) );
  XOR U37315 ( .A(n37346), .B(n37350), .Z(n37348) );
  XNOR U37316 ( .A(n37351), .B(n37352), .Z(n37345) );
  NOR U37317 ( .A(n37353), .B(n37354), .Z(n37352) );
  XOR U37318 ( .A(n37351), .B(n37355), .Z(n37353) );
  AND U37319 ( .A(n37204), .B(n37193), .Z(n37271) );
  XNOR U37320 ( .A(n37356), .B(n37298), .Z(n37193) );
  XOR U37321 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(
        p_input[2048]), .Z(n37298) );
  XOR U37322 ( .A(n37286), .B(n37285), .Z(n37356) );
  XNOR U37323 ( .A(n37357), .B(n37292), .Z(n37285) );
  XNOR U37324 ( .A(n37281), .B(n37280), .Z(n37292) );
  XOR U37325 ( .A(n37358), .B(n37277), .Z(n37280) );
  XNOR U37326 ( .A(n15566), .B(p_input[2058]), .Z(n37277) );
  IV U37327 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n15566)
         );
  XOR U37328 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n16732), 
        .Z(n37358) );
  XNOR U37329 ( .A(n13547), .B(p_input[2060]), .Z(n37281) );
  IV U37330 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n13547)
         );
  XNOR U37331 ( .A(n37291), .B(n37282), .Z(n37357) );
  XNOR U37332 ( .A(n9504), .B(p_input[2049]), .Z(n37282) );
  IV U37333 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n9504) );
  XOR U37334 ( .A(n37359), .B(n37297), .Z(n37291) );
  XNOR U37335 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(
        p_input[2063]), .Z(n37297) );
  XOR U37336 ( .A(n37288), .B(n37296), .Z(n37359) );
  XOR U37337 ( .A(n37360), .B(n37293), .Z(n37296) );
  XNOR U37338 ( .A(n12538), .B(p_input[2061]), .Z(n37293) );
  IV U37339 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n12538)
         );
  XOR U37340 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(n16737), 
        .Z(n37360) );
  XNOR U37341 ( .A(n1412), .B(p_input[2057]), .Z(n37288) );
  IV U37342 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .Z(n1412) );
  XNOR U37343 ( .A(n37304), .B(n37303), .Z(n37286) );
  XNOR U37344 ( .A(n37361), .B(n37309), .Z(n37303) );
  XNOR U37345 ( .A(n2425), .B(p_input[2056]), .Z(n37309) );
  IV U37346 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .Z(n2425) );
  XOR U37347 ( .A(n37300), .B(n37308), .Z(n37361) );
  XOR U37348 ( .A(n37362), .B(n37305), .Z(n37308) );
  XNOR U37349 ( .A(n4447), .B(p_input[2054]), .Z(n37305) );
  IV U37350 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .Z(n4447) );
  XOR U37351 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(n17722), 
        .Z(n37362) );
  XNOR U37352 ( .A(n8493), .B(p_input[2050]), .Z(n37300) );
  IV U37353 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n8493) );
  XNOR U37354 ( .A(n37314), .B(n37313), .Z(n37304) );
  XOR U37355 ( .A(n37363), .B(n37310), .Z(n37313) );
  XNOR U37356 ( .A(n7482), .B(p_input[2051]), .Z(n37310) );
  IV U37357 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .Z(n7482) );
  XOR U37358 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(n17724), 
        .Z(n37363) );
  XNOR U37359 ( .A(n5458), .B(p_input[2053]), .Z(n37314) );
  IV U37360 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .Z(n5458) );
  XOR U37361 ( .A(n37364), .B(n37344), .Z(n37204) );
  XOR U37362 ( .A(n37322), .B(n37321), .Z(n37344) );
  XNOR U37363 ( .A(n37365), .B(n37327), .Z(n37321) );
  XNOR U37364 ( .A(n2429), .B(p_input[2056]), .Z(n37327) );
  IV U37365 ( .A(\knn_comb_/min_val_out[0][8] ), .Z(n2429) );
  XOR U37366 ( .A(n37318), .B(n37326), .Z(n37365) );
  XOR U37367 ( .A(n37366), .B(n37323), .Z(n37326) );
  XNOR U37368 ( .A(n4451), .B(p_input[2054]), .Z(n37323) );
  IV U37369 ( .A(\knn_comb_/min_val_out[0][6] ), .Z(n4451) );
  XOR U37370 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n17722), .Z(n37366) );
  IV U37371 ( .A(p_input[2055]), .Z(n17722) );
  XNOR U37372 ( .A(n8497), .B(p_input[2050]), .Z(n37318) );
  IV U37373 ( .A(\knn_comb_/min_val_out[0][2] ), .Z(n8497) );
  XNOR U37374 ( .A(n37332), .B(n37331), .Z(n37322) );
  XOR U37375 ( .A(n37367), .B(n37328), .Z(n37331) );
  XNOR U37376 ( .A(n7486), .B(p_input[2051]), .Z(n37328) );
  IV U37377 ( .A(\knn_comb_/min_val_out[0][3] ), .Z(n7486) );
  XOR U37378 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n17724), .Z(n37367) );
  IV U37379 ( .A(p_input[2052]), .Z(n17724) );
  XNOR U37380 ( .A(n5462), .B(p_input[2053]), .Z(n37332) );
  IV U37381 ( .A(\knn_comb_/min_val_out[0][5] ), .Z(n5462) );
  XNOR U37382 ( .A(n37343), .B(n37333), .Z(n37364) );
  XOR U37383 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[2048]), .Z(n37333) );
  XNOR U37384 ( .A(n37368), .B(n37350), .Z(n37343) );
  XNOR U37385 ( .A(n37339), .B(n37338), .Z(n37350) );
  XOR U37386 ( .A(n37369), .B(n37335), .Z(n37338) );
  XNOR U37387 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n16904), .Z(n37335) );
  IV U37388 ( .A(p_input[2058]), .Z(n16904) );
  XOR U37389 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n16732), .Z(n37369) );
  IV U37390 ( .A(p_input[2059]), .Z(n16732) );
  XOR U37391 ( .A(\knn_comb_/min_val_out[0][12] ), .B(p_input[2060]), .Z(
        n37339) );
  XNOR U37392 ( .A(n37349), .B(n37340), .Z(n37368) );
  XNOR U37393 ( .A(n9508), .B(p_input[2049]), .Z(n37340) );
  IV U37394 ( .A(\knn_comb_/min_val_out[0][1] ), .Z(n9508) );
  XOR U37395 ( .A(n37370), .B(n37355), .Z(n37349) );
  XNOR U37396 ( .A(\knn_comb_/min_val_out[0][15] ), .B(p_input[2063]), .Z(
        n37355) );
  XOR U37397 ( .A(n37346), .B(n37354), .Z(n37370) );
  XOR U37398 ( .A(n37371), .B(n37351), .Z(n37354) );
  XOR U37399 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[2061]), .Z(
        n37351) );
  XOR U37400 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n16737), .Z(n37371) );
  IV U37401 ( .A(p_input[2062]), .Z(n16737) );
  XNOR U37402 ( .A(n1418), .B(p_input[2057]), .Z(n37346) );
  IV U37403 ( .A(\knn_comb_/min_val_out[0][9] ), .Z(n1418) );
endmodule

