
module knn_comb_BMR_W32_K1_N4 ( p_input, o );
  input [159:0] p_input;
  output [31:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/min_val_out[0][16] , \knn_comb_/min_val_out[0][17] ,
         \knn_comb_/min_val_out[0][18] , \knn_comb_/min_val_out[0][19] ,
         \knn_comb_/min_val_out[0][20] , \knn_comb_/min_val_out[0][21] ,
         \knn_comb_/min_val_out[0][22] , \knn_comb_/min_val_out[0][23] ,
         \knn_comb_/min_val_out[0][24] , \knn_comb_/min_val_out[0][25] ,
         \knn_comb_/min_val_out[0][26] , \knn_comb_/min_val_out[0][27] ,
         \knn_comb_/min_val_out[0][28] , \knn_comb_/min_val_out[0][29] ,
         \knn_comb_/min_val_out[0][30] , \knn_comb_/min_val_out[0][31] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064;
  assign \knn_comb_/min_val_out[0][0]  = p_input[96];
  assign \knn_comb_/min_val_out[0][1]  = p_input[97];
  assign \knn_comb_/min_val_out[0][2]  = p_input[98];
  assign \knn_comb_/min_val_out[0][3]  = p_input[99];
  assign \knn_comb_/min_val_out[0][4]  = p_input[100];
  assign \knn_comb_/min_val_out[0][5]  = p_input[101];
  assign \knn_comb_/min_val_out[0][6]  = p_input[102];
  assign \knn_comb_/min_val_out[0][7]  = p_input[103];
  assign \knn_comb_/min_val_out[0][8]  = p_input[104];
  assign \knn_comb_/min_val_out[0][9]  = p_input[105];
  assign \knn_comb_/min_val_out[0][10]  = p_input[106];
  assign \knn_comb_/min_val_out[0][11]  = p_input[107];
  assign \knn_comb_/min_val_out[0][12]  = p_input[108];
  assign \knn_comb_/min_val_out[0][13]  = p_input[109];
  assign \knn_comb_/min_val_out[0][14]  = p_input[110];
  assign \knn_comb_/min_val_out[0][15]  = p_input[111];
  assign \knn_comb_/min_val_out[0][16]  = p_input[112];
  assign \knn_comb_/min_val_out[0][17]  = p_input[113];
  assign \knn_comb_/min_val_out[0][18]  = p_input[114];
  assign \knn_comb_/min_val_out[0][19]  = p_input[115];
  assign \knn_comb_/min_val_out[0][20]  = p_input[116];
  assign \knn_comb_/min_val_out[0][21]  = p_input[117];
  assign \knn_comb_/min_val_out[0][22]  = p_input[118];
  assign \knn_comb_/min_val_out[0][23]  = p_input[119];
  assign \knn_comb_/min_val_out[0][24]  = p_input[120];
  assign \knn_comb_/min_val_out[0][25]  = p_input[121];
  assign \knn_comb_/min_val_out[0][26]  = p_input[122];
  assign \knn_comb_/min_val_out[0][27]  = p_input[123];
  assign \knn_comb_/min_val_out[0][28]  = p_input[124];
  assign \knn_comb_/min_val_out[0][29]  = p_input[125];
  assign \knn_comb_/min_val_out[0][30]  = p_input[126];
  assign \knn_comb_/min_val_out[0][31]  = p_input[127];

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(n3), .B(n4), .Z(n1) );
  XNOR U3 ( .A(p_input[9]), .B(n2), .Z(n4) );
  XNOR U4 ( .A(n5), .B(n6), .Z(n2) );
  AND U5 ( .A(n7), .B(n8), .Z(n6) );
  XOR U6 ( .A(p_input[41]), .B(n5), .Z(n8) );
  XOR U7 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n9), .Z(n5) );
  AND U8 ( .A(n10), .B(n11), .Z(n9) );
  XOR U9 ( .A(p_input[73]), .B(\knn_comb_/min_val_out[0][9] ), .Z(n11) );
  XNOR U10 ( .A(n12), .B(n13), .Z(o[8]) );
  AND U11 ( .A(n3), .B(n14), .Z(n12) );
  XNOR U12 ( .A(p_input[8]), .B(n13), .Z(n14) );
  XNOR U13 ( .A(n15), .B(n16), .Z(n13) );
  AND U14 ( .A(n7), .B(n17), .Z(n16) );
  XOR U15 ( .A(p_input[40]), .B(n15), .Z(n17) );
  XOR U16 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n18), .Z(n15) );
  AND U17 ( .A(n10), .B(n19), .Z(n18) );
  XOR U18 ( .A(p_input[72]), .B(\knn_comb_/min_val_out[0][8] ), .Z(n19) );
  XNOR U19 ( .A(n20), .B(n21), .Z(o[7]) );
  AND U20 ( .A(n3), .B(n22), .Z(n20) );
  XNOR U21 ( .A(p_input[7]), .B(n21), .Z(n22) );
  XNOR U22 ( .A(n23), .B(n24), .Z(n21) );
  AND U23 ( .A(n7), .B(n25), .Z(n24) );
  XOR U24 ( .A(p_input[39]), .B(n23), .Z(n25) );
  XOR U25 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n26), .Z(n23) );
  AND U26 ( .A(n10), .B(n27), .Z(n26) );
  XOR U27 ( .A(p_input[71]), .B(\knn_comb_/min_val_out[0][7] ), .Z(n27) );
  XNOR U28 ( .A(n28), .B(n29), .Z(o[6]) );
  AND U29 ( .A(n3), .B(n30), .Z(n28) );
  XNOR U30 ( .A(p_input[6]), .B(n29), .Z(n30) );
  XNOR U31 ( .A(n31), .B(n32), .Z(n29) );
  AND U32 ( .A(n7), .B(n33), .Z(n32) );
  XOR U33 ( .A(p_input[38]), .B(n31), .Z(n33) );
  XOR U34 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n34), .Z(n31) );
  AND U35 ( .A(n10), .B(n35), .Z(n34) );
  XOR U36 ( .A(p_input[70]), .B(\knn_comb_/min_val_out[0][6] ), .Z(n35) );
  XNOR U37 ( .A(n36), .B(n37), .Z(o[5]) );
  AND U38 ( .A(n3), .B(n38), .Z(n36) );
  XNOR U39 ( .A(p_input[5]), .B(n37), .Z(n38) );
  XNOR U40 ( .A(n39), .B(n40), .Z(n37) );
  AND U41 ( .A(n7), .B(n41), .Z(n40) );
  XOR U42 ( .A(p_input[37]), .B(n39), .Z(n41) );
  XOR U43 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n42), .Z(n39) );
  AND U44 ( .A(n10), .B(n43), .Z(n42) );
  XOR U45 ( .A(p_input[69]), .B(\knn_comb_/min_val_out[0][5] ), .Z(n43) );
  XNOR U46 ( .A(n44), .B(n45), .Z(o[4]) );
  AND U47 ( .A(n3), .B(n46), .Z(n44) );
  XNOR U48 ( .A(p_input[4]), .B(n45), .Z(n46) );
  XNOR U49 ( .A(n47), .B(n48), .Z(n45) );
  AND U50 ( .A(n7), .B(n49), .Z(n48) );
  XOR U51 ( .A(p_input[36]), .B(n47), .Z(n49) );
  XOR U52 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n50), .Z(n47) );
  AND U53 ( .A(n10), .B(n51), .Z(n50) );
  XOR U54 ( .A(p_input[68]), .B(\knn_comb_/min_val_out[0][4] ), .Z(n51) );
  XNOR U55 ( .A(n52), .B(n53), .Z(o[3]) );
  AND U56 ( .A(n3), .B(n54), .Z(n52) );
  XNOR U57 ( .A(p_input[3]), .B(n53), .Z(n54) );
  XNOR U58 ( .A(n55), .B(n56), .Z(n53) );
  AND U59 ( .A(n7), .B(n57), .Z(n56) );
  XOR U60 ( .A(p_input[35]), .B(n55), .Z(n57) );
  XOR U61 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n58), .Z(n55) );
  AND U62 ( .A(n10), .B(n59), .Z(n58) );
  XOR U63 ( .A(p_input[67]), .B(\knn_comb_/min_val_out[0][3] ), .Z(n59) );
  XNOR U64 ( .A(n60), .B(n61), .Z(o[31]) );
  AND U65 ( .A(n3), .B(n62), .Z(n60) );
  XNOR U66 ( .A(p_input[31]), .B(n61), .Z(n62) );
  XNOR U67 ( .A(n63), .B(n64), .Z(n61) );
  AND U68 ( .A(n7), .B(n65), .Z(n64) );
  XOR U69 ( .A(p_input[63]), .B(n63), .Z(n65) );
  XOR U70 ( .A(\knn_comb_/min_val_out[0][31] ), .B(n66), .Z(n63) );
  AND U71 ( .A(n10), .B(n67), .Z(n66) );
  XOR U72 ( .A(p_input[95]), .B(\knn_comb_/min_val_out[0][31] ), .Z(n67) );
  XNOR U73 ( .A(n68), .B(n69), .Z(o[30]) );
  AND U74 ( .A(n3), .B(n70), .Z(n68) );
  XNOR U75 ( .A(p_input[30]), .B(n69), .Z(n70) );
  XNOR U76 ( .A(n71), .B(n72), .Z(n69) );
  AND U77 ( .A(n7), .B(n73), .Z(n72) );
  XOR U78 ( .A(p_input[62]), .B(n71), .Z(n73) );
  XOR U79 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n74), .Z(n71) );
  AND U80 ( .A(n10), .B(n75), .Z(n74) );
  XOR U81 ( .A(p_input[94]), .B(\knn_comb_/min_val_out[0][30] ), .Z(n75) );
  XNOR U82 ( .A(n76), .B(n77), .Z(o[2]) );
  AND U83 ( .A(n3), .B(n78), .Z(n76) );
  XNOR U84 ( .A(p_input[2]), .B(n77), .Z(n78) );
  XNOR U85 ( .A(n79), .B(n80), .Z(n77) );
  AND U86 ( .A(n7), .B(n81), .Z(n80) );
  XOR U87 ( .A(p_input[34]), .B(n79), .Z(n81) );
  XOR U88 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n82), .Z(n79) );
  AND U89 ( .A(n10), .B(n83), .Z(n82) );
  XOR U90 ( .A(p_input[66]), .B(\knn_comb_/min_val_out[0][2] ), .Z(n83) );
  XNOR U91 ( .A(n84), .B(n85), .Z(o[29]) );
  AND U92 ( .A(n3), .B(n86), .Z(n84) );
  XNOR U93 ( .A(p_input[29]), .B(n85), .Z(n86) );
  XNOR U94 ( .A(n87), .B(n88), .Z(n85) );
  AND U95 ( .A(n7), .B(n89), .Z(n88) );
  XOR U96 ( .A(p_input[61]), .B(n87), .Z(n89) );
  XOR U97 ( .A(\knn_comb_/min_val_out[0][29] ), .B(n90), .Z(n87) );
  AND U98 ( .A(n10), .B(n91), .Z(n90) );
  XOR U99 ( .A(p_input[93]), .B(\knn_comb_/min_val_out[0][29] ), .Z(n91) );
  XNOR U100 ( .A(n92), .B(n93), .Z(o[28]) );
  AND U101 ( .A(n3), .B(n94), .Z(n92) );
  XNOR U102 ( .A(p_input[28]), .B(n93), .Z(n94) );
  XNOR U103 ( .A(n95), .B(n96), .Z(n93) );
  AND U104 ( .A(n7), .B(n97), .Z(n96) );
  XOR U105 ( .A(p_input[60]), .B(n95), .Z(n97) );
  XOR U106 ( .A(\knn_comb_/min_val_out[0][28] ), .B(n98), .Z(n95) );
  AND U107 ( .A(n10), .B(n99), .Z(n98) );
  XOR U108 ( .A(p_input[92]), .B(\knn_comb_/min_val_out[0][28] ), .Z(n99) );
  XNOR U109 ( .A(n100), .B(n101), .Z(o[27]) );
  AND U110 ( .A(n3), .B(n102), .Z(n100) );
  XNOR U111 ( .A(p_input[27]), .B(n101), .Z(n102) );
  XNOR U112 ( .A(n103), .B(n104), .Z(n101) );
  AND U113 ( .A(n7), .B(n105), .Z(n104) );
  XOR U114 ( .A(p_input[59]), .B(n103), .Z(n105) );
  XOR U115 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n106), .Z(n103) );
  AND U116 ( .A(n10), .B(n107), .Z(n106) );
  XOR U117 ( .A(p_input[91]), .B(\knn_comb_/min_val_out[0][27] ), .Z(n107) );
  XNOR U118 ( .A(n108), .B(n109), .Z(o[26]) );
  AND U119 ( .A(n3), .B(n110), .Z(n108) );
  XNOR U120 ( .A(p_input[26]), .B(n109), .Z(n110) );
  XNOR U121 ( .A(n111), .B(n112), .Z(n109) );
  AND U122 ( .A(n7), .B(n113), .Z(n112) );
  XOR U123 ( .A(p_input[58]), .B(n111), .Z(n113) );
  XOR U124 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n114), .Z(n111) );
  AND U125 ( .A(n10), .B(n115), .Z(n114) );
  XOR U126 ( .A(p_input[90]), .B(\knn_comb_/min_val_out[0][26] ), .Z(n115) );
  XNOR U127 ( .A(n116), .B(n117), .Z(o[25]) );
  AND U128 ( .A(n3), .B(n118), .Z(n116) );
  XNOR U129 ( .A(p_input[25]), .B(n117), .Z(n118) );
  XNOR U130 ( .A(n119), .B(n120), .Z(n117) );
  AND U131 ( .A(n7), .B(n121), .Z(n120) );
  XOR U132 ( .A(p_input[57]), .B(n119), .Z(n121) );
  XOR U133 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n122), .Z(n119) );
  AND U134 ( .A(n10), .B(n123), .Z(n122) );
  XOR U135 ( .A(p_input[89]), .B(\knn_comb_/min_val_out[0][25] ), .Z(n123) );
  XNOR U136 ( .A(n124), .B(n125), .Z(o[24]) );
  AND U137 ( .A(n3), .B(n126), .Z(n124) );
  XNOR U138 ( .A(p_input[24]), .B(n125), .Z(n126) );
  XNOR U139 ( .A(n127), .B(n128), .Z(n125) );
  AND U140 ( .A(n7), .B(n129), .Z(n128) );
  XOR U141 ( .A(p_input[56]), .B(n127), .Z(n129) );
  XOR U142 ( .A(\knn_comb_/min_val_out[0][24] ), .B(n130), .Z(n127) );
  AND U143 ( .A(n10), .B(n131), .Z(n130) );
  XOR U144 ( .A(p_input[88]), .B(\knn_comb_/min_val_out[0][24] ), .Z(n131) );
  XNOR U145 ( .A(n132), .B(n133), .Z(o[23]) );
  AND U146 ( .A(n3), .B(n134), .Z(n132) );
  XNOR U147 ( .A(p_input[23]), .B(n133), .Z(n134) );
  XNOR U148 ( .A(n135), .B(n136), .Z(n133) );
  AND U149 ( .A(n7), .B(n137), .Z(n136) );
  XOR U150 ( .A(p_input[55]), .B(n135), .Z(n137) );
  XOR U151 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n138), .Z(n135) );
  AND U152 ( .A(n10), .B(n139), .Z(n138) );
  XOR U153 ( .A(p_input[87]), .B(\knn_comb_/min_val_out[0][23] ), .Z(n139) );
  XNOR U154 ( .A(n140), .B(n141), .Z(o[22]) );
  AND U155 ( .A(n3), .B(n142), .Z(n140) );
  XNOR U156 ( .A(p_input[22]), .B(n141), .Z(n142) );
  XNOR U157 ( .A(n143), .B(n144), .Z(n141) );
  AND U158 ( .A(n7), .B(n145), .Z(n144) );
  XOR U159 ( .A(p_input[54]), .B(n143), .Z(n145) );
  XOR U160 ( .A(\knn_comb_/min_val_out[0][22] ), .B(n146), .Z(n143) );
  AND U161 ( .A(n10), .B(n147), .Z(n146) );
  XOR U162 ( .A(p_input[86]), .B(\knn_comb_/min_val_out[0][22] ), .Z(n147) );
  XNOR U163 ( .A(n148), .B(n149), .Z(o[21]) );
  AND U164 ( .A(n3), .B(n150), .Z(n148) );
  XNOR U165 ( .A(p_input[21]), .B(n149), .Z(n150) );
  XNOR U166 ( .A(n151), .B(n152), .Z(n149) );
  AND U167 ( .A(n7), .B(n153), .Z(n152) );
  XOR U168 ( .A(p_input[53]), .B(n151), .Z(n153) );
  XOR U169 ( .A(\knn_comb_/min_val_out[0][21] ), .B(n154), .Z(n151) );
  AND U170 ( .A(n10), .B(n155), .Z(n154) );
  XOR U171 ( .A(p_input[85]), .B(\knn_comb_/min_val_out[0][21] ), .Z(n155) );
  XNOR U172 ( .A(n156), .B(n157), .Z(o[20]) );
  AND U173 ( .A(n3), .B(n158), .Z(n156) );
  XNOR U174 ( .A(p_input[20]), .B(n157), .Z(n158) );
  XNOR U175 ( .A(n159), .B(n160), .Z(n157) );
  AND U176 ( .A(n7), .B(n161), .Z(n160) );
  XOR U177 ( .A(p_input[52]), .B(n159), .Z(n161) );
  XOR U178 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n162), .Z(n159) );
  AND U179 ( .A(n10), .B(n163), .Z(n162) );
  XOR U180 ( .A(p_input[84]), .B(\knn_comb_/min_val_out[0][20] ), .Z(n163) );
  XNOR U181 ( .A(n164), .B(n165), .Z(o[1]) );
  AND U182 ( .A(n3), .B(n166), .Z(n164) );
  XNOR U183 ( .A(p_input[1]), .B(n165), .Z(n166) );
  XNOR U184 ( .A(n167), .B(n168), .Z(n165) );
  AND U185 ( .A(n7), .B(n169), .Z(n168) );
  XOR U186 ( .A(p_input[33]), .B(n167), .Z(n169) );
  XOR U187 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n170), .Z(n167) );
  AND U188 ( .A(n10), .B(n171), .Z(n170) );
  XOR U189 ( .A(p_input[65]), .B(\knn_comb_/min_val_out[0][1] ), .Z(n171) );
  XNOR U190 ( .A(n172), .B(n173), .Z(o[19]) );
  AND U191 ( .A(n3), .B(n174), .Z(n172) );
  XNOR U192 ( .A(p_input[19]), .B(n173), .Z(n174) );
  XNOR U193 ( .A(n175), .B(n176), .Z(n173) );
  AND U194 ( .A(n7), .B(n177), .Z(n176) );
  XOR U195 ( .A(p_input[51]), .B(n175), .Z(n177) );
  XOR U196 ( .A(\knn_comb_/min_val_out[0][19] ), .B(n178), .Z(n175) );
  AND U197 ( .A(n10), .B(n179), .Z(n178) );
  XOR U198 ( .A(p_input[83]), .B(\knn_comb_/min_val_out[0][19] ), .Z(n179) );
  XNOR U199 ( .A(n180), .B(n181), .Z(o[18]) );
  AND U200 ( .A(n3), .B(n182), .Z(n180) );
  XNOR U201 ( .A(p_input[18]), .B(n181), .Z(n182) );
  XNOR U202 ( .A(n183), .B(n184), .Z(n181) );
  AND U203 ( .A(n7), .B(n185), .Z(n184) );
  XOR U204 ( .A(p_input[50]), .B(n183), .Z(n185) );
  XOR U205 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n186), .Z(n183) );
  AND U206 ( .A(n10), .B(n187), .Z(n186) );
  XOR U207 ( .A(p_input[82]), .B(\knn_comb_/min_val_out[0][18] ), .Z(n187) );
  XNOR U208 ( .A(n188), .B(n189), .Z(o[17]) );
  AND U209 ( .A(n3), .B(n190), .Z(n188) );
  XNOR U210 ( .A(p_input[17]), .B(n189), .Z(n190) );
  XNOR U211 ( .A(n191), .B(n192), .Z(n189) );
  AND U212 ( .A(n7), .B(n193), .Z(n192) );
  XOR U213 ( .A(p_input[49]), .B(n191), .Z(n193) );
  XOR U214 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n194), .Z(n191) );
  AND U215 ( .A(n10), .B(n195), .Z(n194) );
  XOR U216 ( .A(p_input[81]), .B(\knn_comb_/min_val_out[0][17] ), .Z(n195) );
  XNOR U217 ( .A(n196), .B(n197), .Z(o[16]) );
  AND U218 ( .A(n3), .B(n198), .Z(n196) );
  XNOR U219 ( .A(p_input[16]), .B(n197), .Z(n198) );
  XNOR U220 ( .A(n199), .B(n200), .Z(n197) );
  AND U221 ( .A(n7), .B(n201), .Z(n200) );
  XOR U222 ( .A(p_input[48]), .B(n199), .Z(n201) );
  XOR U223 ( .A(\knn_comb_/min_val_out[0][16] ), .B(n202), .Z(n199) );
  AND U224 ( .A(n10), .B(n203), .Z(n202) );
  XOR U225 ( .A(p_input[80]), .B(\knn_comb_/min_val_out[0][16] ), .Z(n203) );
  XNOR U226 ( .A(n204), .B(n205), .Z(o[15]) );
  AND U227 ( .A(n3), .B(n206), .Z(n204) );
  XNOR U228 ( .A(p_input[15]), .B(n205), .Z(n206) );
  XNOR U229 ( .A(n207), .B(n208), .Z(n205) );
  AND U230 ( .A(n7), .B(n209), .Z(n208) );
  XOR U231 ( .A(p_input[47]), .B(n207), .Z(n209) );
  XOR U232 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n210), .Z(n207) );
  AND U233 ( .A(n10), .B(n211), .Z(n210) );
  XOR U234 ( .A(p_input[79]), .B(\knn_comb_/min_val_out[0][15] ), .Z(n211) );
  XNOR U235 ( .A(n212), .B(n213), .Z(o[14]) );
  AND U236 ( .A(n3), .B(n214), .Z(n212) );
  XNOR U237 ( .A(p_input[14]), .B(n213), .Z(n214) );
  XNOR U238 ( .A(n215), .B(n216), .Z(n213) );
  AND U239 ( .A(n7), .B(n217), .Z(n216) );
  XOR U240 ( .A(p_input[46]), .B(n215), .Z(n217) );
  XOR U241 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n218), .Z(n215) );
  AND U242 ( .A(n10), .B(n219), .Z(n218) );
  XOR U243 ( .A(p_input[78]), .B(\knn_comb_/min_val_out[0][14] ), .Z(n219) );
  XNOR U244 ( .A(n220), .B(n221), .Z(o[13]) );
  AND U245 ( .A(n3), .B(n222), .Z(n220) );
  XNOR U246 ( .A(p_input[13]), .B(n221), .Z(n222) );
  XNOR U247 ( .A(n223), .B(n224), .Z(n221) );
  AND U248 ( .A(n7), .B(n225), .Z(n224) );
  XOR U249 ( .A(p_input[45]), .B(n223), .Z(n225) );
  XOR U250 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n226), .Z(n223) );
  AND U251 ( .A(n10), .B(n227), .Z(n226) );
  XOR U252 ( .A(p_input[77]), .B(\knn_comb_/min_val_out[0][13] ), .Z(n227) );
  XNOR U253 ( .A(n228), .B(n229), .Z(o[12]) );
  AND U254 ( .A(n3), .B(n230), .Z(n228) );
  XNOR U255 ( .A(p_input[12]), .B(n229), .Z(n230) );
  XNOR U256 ( .A(n231), .B(n232), .Z(n229) );
  AND U257 ( .A(n7), .B(n233), .Z(n232) );
  XOR U258 ( .A(p_input[44]), .B(n231), .Z(n233) );
  XOR U259 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n234), .Z(n231) );
  AND U260 ( .A(n10), .B(n235), .Z(n234) );
  XOR U261 ( .A(p_input[76]), .B(\knn_comb_/min_val_out[0][12] ), .Z(n235) );
  XNOR U262 ( .A(n236), .B(n237), .Z(o[11]) );
  AND U263 ( .A(n3), .B(n238), .Z(n236) );
  XNOR U264 ( .A(p_input[11]), .B(n237), .Z(n238) );
  XNOR U265 ( .A(n239), .B(n240), .Z(n237) );
  AND U266 ( .A(n7), .B(n241), .Z(n240) );
  XOR U267 ( .A(p_input[43]), .B(n239), .Z(n241) );
  XOR U268 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n242), .Z(n239) );
  AND U269 ( .A(n10), .B(n243), .Z(n242) );
  XOR U270 ( .A(p_input[75]), .B(\knn_comb_/min_val_out[0][11] ), .Z(n243) );
  XNOR U271 ( .A(n244), .B(n245), .Z(o[10]) );
  AND U272 ( .A(n3), .B(n246), .Z(n244) );
  XNOR U273 ( .A(p_input[10]), .B(n245), .Z(n246) );
  XNOR U274 ( .A(n247), .B(n248), .Z(n245) );
  AND U275 ( .A(n7), .B(n249), .Z(n248) );
  XOR U276 ( .A(p_input[42]), .B(n247), .Z(n249) );
  XOR U277 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n250), .Z(n247) );
  AND U278 ( .A(n10), .B(n251), .Z(n250) );
  XOR U279 ( .A(p_input[74]), .B(\knn_comb_/min_val_out[0][10] ), .Z(n251) );
  XNOR U280 ( .A(n252), .B(n253), .Z(o[0]) );
  AND U281 ( .A(n3), .B(n254), .Z(n252) );
  XNOR U282 ( .A(p_input[0]), .B(n253), .Z(n254) );
  XNOR U283 ( .A(n255), .B(n256), .Z(n253) );
  AND U284 ( .A(n7), .B(n257), .Z(n256) );
  XOR U285 ( .A(p_input[32]), .B(n255), .Z(n257) );
  XOR U286 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n258), .Z(n255) );
  AND U287 ( .A(n10), .B(n259), .Z(n258) );
  XOR U288 ( .A(p_input[64]), .B(\knn_comb_/min_val_out[0][0] ), .Z(n259) );
  XNOR U289 ( .A(n260), .B(n261), .Z(n3) );
  NOR U290 ( .A(n262), .B(n263), .Z(n261) );
  XOR U291 ( .A(n264), .B(n260), .Z(n263) );
  AND U292 ( .A(n265), .B(n266), .Z(n264) );
  NOR U293 ( .A(n267), .B(n260), .Z(n262) );
  AND U294 ( .A(n268), .B(n269), .Z(n267) );
  XOR U295 ( .A(n270), .B(n271), .Z(n260) );
  AND U296 ( .A(n272), .B(n273), .Z(n271) );
  XNOR U297 ( .A(n270), .B(n268), .Z(n273) );
  XNOR U298 ( .A(n274), .B(n275), .Z(n268) );
  XOR U299 ( .A(n276), .B(n269), .Z(n275) );
  AND U300 ( .A(n277), .B(n278), .Z(n269) );
  AND U301 ( .A(n279), .B(n280), .Z(n276) );
  XOR U302 ( .A(n281), .B(n274), .Z(n279) );
  XOR U303 ( .A(n282), .B(n270), .Z(n272) );
  XNOR U304 ( .A(n283), .B(n284), .Z(n282) );
  AND U305 ( .A(n7), .B(n285), .Z(n284) );
  XOR U306 ( .A(n286), .B(n283), .Z(n285) );
  XOR U307 ( .A(n287), .B(n288), .Z(n270) );
  AND U308 ( .A(n289), .B(n290), .Z(n288) );
  XNOR U309 ( .A(n287), .B(n277), .Z(n290) );
  XOR U310 ( .A(n291), .B(n280), .Z(n277) );
  XNOR U311 ( .A(n292), .B(n274), .Z(n280) );
  XOR U312 ( .A(n293), .B(n294), .Z(n274) );
  AND U313 ( .A(n295), .B(n296), .Z(n294) );
  XOR U314 ( .A(n297), .B(n293), .Z(n295) );
  XNOR U315 ( .A(n298), .B(n299), .Z(n292) );
  AND U316 ( .A(n300), .B(n301), .Z(n299) );
  XOR U317 ( .A(n298), .B(n302), .Z(n300) );
  XNOR U318 ( .A(n281), .B(n278), .Z(n291) );
  AND U319 ( .A(n303), .B(n304), .Z(n278) );
  XOR U320 ( .A(n305), .B(n306), .Z(n281) );
  AND U321 ( .A(n307), .B(n308), .Z(n306) );
  XOR U322 ( .A(n305), .B(n309), .Z(n307) );
  XOR U323 ( .A(n310), .B(n287), .Z(n289) );
  XNOR U324 ( .A(n311), .B(n312), .Z(n310) );
  AND U325 ( .A(n7), .B(n313), .Z(n312) );
  XNOR U326 ( .A(n314), .B(n311), .Z(n313) );
  XOR U327 ( .A(n315), .B(n316), .Z(n287) );
  AND U328 ( .A(n317), .B(n318), .Z(n316) );
  XNOR U329 ( .A(n315), .B(n303), .Z(n318) );
  XOR U330 ( .A(n319), .B(n296), .Z(n303) );
  XNOR U331 ( .A(n320), .B(n302), .Z(n296) );
  XOR U332 ( .A(n321), .B(n322), .Z(n302) );
  AND U333 ( .A(n323), .B(n324), .Z(n322) );
  XOR U334 ( .A(n321), .B(n325), .Z(n323) );
  XNOR U335 ( .A(n301), .B(n293), .Z(n320) );
  XOR U336 ( .A(n326), .B(n327), .Z(n293) );
  AND U337 ( .A(n328), .B(n329), .Z(n327) );
  XNOR U338 ( .A(n330), .B(n326), .Z(n328) );
  XNOR U339 ( .A(n331), .B(n298), .Z(n301) );
  XOR U340 ( .A(n332), .B(n333), .Z(n298) );
  AND U341 ( .A(n334), .B(n335), .Z(n333) );
  XOR U342 ( .A(n332), .B(n336), .Z(n334) );
  XNOR U343 ( .A(n337), .B(n338), .Z(n331) );
  AND U344 ( .A(n339), .B(n340), .Z(n338) );
  XNOR U345 ( .A(n337), .B(n341), .Z(n339) );
  XNOR U346 ( .A(n297), .B(n304), .Z(n319) );
  AND U347 ( .A(n342), .B(n343), .Z(n304) );
  XOR U348 ( .A(n309), .B(n308), .Z(n297) );
  XNOR U349 ( .A(n344), .B(n305), .Z(n308) );
  XOR U350 ( .A(n345), .B(n346), .Z(n305) );
  AND U351 ( .A(n347), .B(n348), .Z(n346) );
  XOR U352 ( .A(n345), .B(n349), .Z(n347) );
  XNOR U353 ( .A(n350), .B(n351), .Z(n344) );
  AND U354 ( .A(n352), .B(n353), .Z(n351) );
  XOR U355 ( .A(n350), .B(n354), .Z(n352) );
  XOR U356 ( .A(n355), .B(n356), .Z(n309) );
  AND U357 ( .A(n357), .B(n358), .Z(n356) );
  XOR U358 ( .A(n355), .B(n359), .Z(n357) );
  XOR U359 ( .A(n360), .B(n315), .Z(n317) );
  XNOR U360 ( .A(n361), .B(n362), .Z(n360) );
  AND U361 ( .A(n7), .B(n363), .Z(n362) );
  XOR U362 ( .A(n364), .B(n361), .Z(n363) );
  XOR U363 ( .A(n365), .B(n366), .Z(n315) );
  AND U364 ( .A(n367), .B(n368), .Z(n366) );
  XNOR U365 ( .A(n365), .B(n342), .Z(n368) );
  XOR U366 ( .A(n369), .B(n329), .Z(n342) );
  XNOR U367 ( .A(n370), .B(n336), .Z(n329) );
  XOR U368 ( .A(n325), .B(n324), .Z(n336) );
  XNOR U369 ( .A(n371), .B(n321), .Z(n324) );
  XOR U370 ( .A(n372), .B(n373), .Z(n321) );
  AND U371 ( .A(n374), .B(n375), .Z(n373) );
  XNOR U372 ( .A(n376), .B(n377), .Z(n374) );
  XNOR U373 ( .A(n378), .B(n379), .Z(n371) );
  NOR U374 ( .A(n380), .B(n381), .Z(n379) );
  XOR U375 ( .A(n378), .B(n382), .Z(n380) );
  XOR U376 ( .A(n383), .B(n384), .Z(n325) );
  NOR U377 ( .A(n385), .B(n386), .Z(n384) );
  XOR U378 ( .A(n383), .B(n387), .Z(n385) );
  XNOR U379 ( .A(n335), .B(n326), .Z(n370) );
  XOR U380 ( .A(n388), .B(n389), .Z(n326) );
  NOR U381 ( .A(n390), .B(n391), .Z(n389) );
  XOR U382 ( .A(n392), .B(n393), .Z(n390) );
  XOR U383 ( .A(n394), .B(n341), .Z(n335) );
  XOR U384 ( .A(n395), .B(n396), .Z(n341) );
  NOR U385 ( .A(n397), .B(n398), .Z(n396) );
  XNOR U386 ( .A(n395), .B(n399), .Z(n397) );
  XNOR U387 ( .A(n340), .B(n332), .Z(n394) );
  XOR U388 ( .A(n400), .B(n401), .Z(n332) );
  AND U389 ( .A(n402), .B(n403), .Z(n401) );
  XOR U390 ( .A(n400), .B(n404), .Z(n402) );
  XNOR U391 ( .A(n405), .B(n337), .Z(n340) );
  XOR U392 ( .A(n406), .B(n407), .Z(n337) );
  AND U393 ( .A(n408), .B(n409), .Z(n407) );
  XNOR U394 ( .A(n410), .B(n411), .Z(n408) );
  XNOR U395 ( .A(n412), .B(n413), .Z(n405) );
  NOR U396 ( .A(n414), .B(n415), .Z(n413) );
  XOR U397 ( .A(n412), .B(n416), .Z(n414) );
  XOR U398 ( .A(n330), .B(n343), .Z(n369) );
  NOR U399 ( .A(n417), .B(n418), .Z(n343) );
  XNOR U400 ( .A(n349), .B(n348), .Z(n330) );
  XNOR U401 ( .A(n419), .B(n354), .Z(n348) );
  XNOR U402 ( .A(n420), .B(n421), .Z(n354) );
  NOR U403 ( .A(n422), .B(n423), .Z(n421) );
  XOR U404 ( .A(n420), .B(n424), .Z(n422) );
  XNOR U405 ( .A(n353), .B(n345), .Z(n419) );
  XOR U406 ( .A(n425), .B(n426), .Z(n345) );
  AND U407 ( .A(n427), .B(n428), .Z(n426) );
  XNOR U408 ( .A(n425), .B(n429), .Z(n427) );
  XNOR U409 ( .A(n430), .B(n350), .Z(n353) );
  XOR U410 ( .A(n431), .B(n432), .Z(n350) );
  AND U411 ( .A(n433), .B(n434), .Z(n432) );
  XNOR U412 ( .A(n435), .B(n436), .Z(n433) );
  XNOR U413 ( .A(n437), .B(n438), .Z(n430) );
  NOR U414 ( .A(n439), .B(n440), .Z(n438) );
  XOR U415 ( .A(n437), .B(n441), .Z(n439) );
  XOR U416 ( .A(n359), .B(n358), .Z(n349) );
  XNOR U417 ( .A(n442), .B(n355), .Z(n358) );
  XOR U418 ( .A(n443), .B(n444), .Z(n355) );
  AND U419 ( .A(n445), .B(n446), .Z(n444) );
  XNOR U420 ( .A(n447), .B(n448), .Z(n445) );
  XNOR U421 ( .A(n449), .B(n450), .Z(n442) );
  NOR U422 ( .A(n451), .B(n452), .Z(n450) );
  XOR U423 ( .A(n449), .B(n453), .Z(n451) );
  XOR U424 ( .A(n454), .B(n455), .Z(n359) );
  NOR U425 ( .A(n456), .B(n457), .Z(n455) );
  XOR U426 ( .A(n454), .B(n458), .Z(n456) );
  XNOR U427 ( .A(n459), .B(n460), .Z(n367) );
  XOR U428 ( .A(n365), .B(n461), .Z(n460) );
  AND U429 ( .A(n7), .B(n462), .Z(n461) );
  XNOR U430 ( .A(n463), .B(n459), .Z(n462) );
  AND U431 ( .A(n464), .B(n417), .Z(n365) );
  XOR U432 ( .A(n465), .B(n418), .Z(n417) );
  XNOR U433 ( .A(p_input[0]), .B(p_input[128]), .Z(n418) );
  XOR U434 ( .A(n393), .B(n391), .Z(n465) );
  XOR U435 ( .A(n466), .B(n404), .Z(n391) );
  XOR U436 ( .A(n377), .B(n375), .Z(n404) );
  XOR U437 ( .A(n467), .B(n382), .Z(n375) );
  XNOR U438 ( .A(p_input[152]), .B(p_input[24]), .Z(n382) );
  XOR U439 ( .A(n372), .B(n381), .Z(n467) );
  XOR U440 ( .A(n468), .B(n378), .Z(n381) );
  XOR U441 ( .A(p_input[150]), .B(p_input[22]), .Z(n378) );
  XNOR U442 ( .A(p_input[151]), .B(p_input[23]), .Z(n468) );
  IV U443 ( .A(n376), .Z(n372) );
  XNOR U444 ( .A(p_input[146]), .B(p_input[18]), .Z(n376) );
  XOR U445 ( .A(n387), .B(n386), .Z(n377) );
  XOR U446 ( .A(n469), .B(n383), .Z(n386) );
  XOR U447 ( .A(p_input[147]), .B(p_input[19]), .Z(n383) );
  XNOR U448 ( .A(p_input[148]), .B(p_input[20]), .Z(n469) );
  XNOR U449 ( .A(p_input[149]), .B(p_input[21]), .Z(n387) );
  XOR U450 ( .A(n403), .B(n392), .Z(n466) );
  IV U451 ( .A(n388), .Z(n392) );
  XOR U452 ( .A(p_input[129]), .B(p_input[1]), .Z(n388) );
  XNOR U453 ( .A(n470), .B(n411), .Z(n403) );
  XOR U454 ( .A(n399), .B(n398), .Z(n411) );
  XNOR U455 ( .A(n471), .B(n395), .Z(n398) );
  XNOR U456 ( .A(p_input[154]), .B(p_input[26]), .Z(n395) );
  XNOR U457 ( .A(p_input[155]), .B(p_input[27]), .Z(n471) );
  XNOR U458 ( .A(p_input[156]), .B(p_input[28]), .Z(n399) );
  XOR U459 ( .A(n409), .B(n472), .Z(n470) );
  IV U460 ( .A(n400), .Z(n472) );
  XOR U461 ( .A(p_input[145]), .B(p_input[17]), .Z(n400) );
  XOR U462 ( .A(n473), .B(n416), .Z(n409) );
  XNOR U463 ( .A(p_input[159]), .B(p_input[31]), .Z(n416) );
  XOR U464 ( .A(n406), .B(n415), .Z(n473) );
  XOR U465 ( .A(n474), .B(n412), .Z(n415) );
  XOR U466 ( .A(p_input[157]), .B(p_input[29]), .Z(n412) );
  XNOR U467 ( .A(p_input[158]), .B(p_input[30]), .Z(n474) );
  IV U468 ( .A(n410), .Z(n406) );
  XNOR U469 ( .A(p_input[153]), .B(p_input[25]), .Z(n410) );
  XNOR U470 ( .A(n429), .B(n428), .Z(n393) );
  XNOR U471 ( .A(n475), .B(n436), .Z(n428) );
  XNOR U472 ( .A(n424), .B(n423), .Z(n436) );
  XOR U473 ( .A(n476), .B(n477), .Z(n423) );
  IV U474 ( .A(n420), .Z(n477) );
  XNOR U475 ( .A(p_input[11]), .B(p_input[139]), .Z(n420) );
  XOR U476 ( .A(p_input[12]), .B(n478), .Z(n476) );
  XOR U477 ( .A(p_input[13]), .B(p_input[141]), .Z(n424) );
  XOR U478 ( .A(n434), .B(n479), .Z(n475) );
  IV U479 ( .A(n425), .Z(n479) );
  XOR U480 ( .A(p_input[130]), .B(p_input[2]), .Z(n425) );
  XOR U481 ( .A(n480), .B(n441), .Z(n434) );
  XNOR U482 ( .A(p_input[144]), .B(p_input[16]), .Z(n441) );
  XOR U483 ( .A(n431), .B(n440), .Z(n480) );
  XOR U484 ( .A(n481), .B(n437), .Z(n440) );
  XOR U485 ( .A(p_input[142]), .B(p_input[14]), .Z(n437) );
  XNOR U486 ( .A(p_input[143]), .B(p_input[15]), .Z(n481) );
  IV U487 ( .A(n435), .Z(n431) );
  XNOR U488 ( .A(p_input[10]), .B(p_input[138]), .Z(n435) );
  XNOR U489 ( .A(n448), .B(n446), .Z(n429) );
  XOR U490 ( .A(n482), .B(n453), .Z(n446) );
  XNOR U491 ( .A(p_input[137]), .B(p_input[9]), .Z(n453) );
  XOR U492 ( .A(n443), .B(n452), .Z(n482) );
  XOR U493 ( .A(n483), .B(n449), .Z(n452) );
  XOR U494 ( .A(p_input[135]), .B(p_input[7]), .Z(n449) );
  XNOR U495 ( .A(p_input[136]), .B(p_input[8]), .Z(n483) );
  IV U496 ( .A(n447), .Z(n443) );
  XNOR U497 ( .A(p_input[131]), .B(p_input[3]), .Z(n447) );
  XOR U498 ( .A(n458), .B(n457), .Z(n448) );
  XOR U499 ( .A(n484), .B(n454), .Z(n457) );
  XOR U500 ( .A(p_input[132]), .B(p_input[4]), .Z(n454) );
  XNOR U501 ( .A(p_input[133]), .B(p_input[5]), .Z(n484) );
  XNOR U502 ( .A(p_input[134]), .B(p_input[6]), .Z(n458) );
  XNOR U503 ( .A(n485), .B(n486), .Z(n464) );
  AND U504 ( .A(n7), .B(n487), .Z(n486) );
  XNOR U505 ( .A(n488), .B(n489), .Z(n487) );
  XNOR U506 ( .A(n490), .B(n491), .Z(n7) );
  MUX U507 ( .IN0(n265), .IN1(n266), .SEL(n490), .F(n491) );
  AND U508 ( .A(n492), .B(n493), .Z(n266) );
  AND U509 ( .A(n494), .B(n495), .Z(n265) );
  XOR U510 ( .A(n496), .B(n497), .Z(n490) );
  AND U511 ( .A(n498), .B(n499), .Z(n497) );
  XNOR U512 ( .A(n496), .B(n494), .Z(n499) );
  IV U513 ( .A(n286), .Z(n494) );
  XOR U514 ( .A(n500), .B(n501), .Z(n286) );
  XOR U515 ( .A(n502), .B(n495), .Z(n501) );
  AND U516 ( .A(n314), .B(n503), .Z(n495) );
  AND U517 ( .A(n504), .B(n505), .Z(n502) );
  XOR U518 ( .A(n506), .B(n500), .Z(n504) );
  XNOR U519 ( .A(n283), .B(n496), .Z(n498) );
  XNOR U520 ( .A(n507), .B(n508), .Z(n283) );
  AND U521 ( .A(n10), .B(n509), .Z(n508) );
  XNOR U522 ( .A(n510), .B(n507), .Z(n509) );
  XOR U523 ( .A(n511), .B(n512), .Z(n496) );
  AND U524 ( .A(n513), .B(n514), .Z(n512) );
  XNOR U525 ( .A(n511), .B(n314), .Z(n514) );
  XOR U526 ( .A(n515), .B(n505), .Z(n314) );
  XNOR U527 ( .A(n516), .B(n500), .Z(n505) );
  XOR U528 ( .A(n517), .B(n518), .Z(n500) );
  AND U529 ( .A(n519), .B(n520), .Z(n518) );
  XOR U530 ( .A(n521), .B(n517), .Z(n519) );
  XNOR U531 ( .A(n522), .B(n523), .Z(n516) );
  AND U532 ( .A(n524), .B(n525), .Z(n523) );
  XOR U533 ( .A(n522), .B(n526), .Z(n524) );
  XNOR U534 ( .A(n506), .B(n503), .Z(n515) );
  AND U535 ( .A(n527), .B(n528), .Z(n503) );
  XOR U536 ( .A(n529), .B(n530), .Z(n506) );
  AND U537 ( .A(n531), .B(n532), .Z(n530) );
  XOR U538 ( .A(n529), .B(n533), .Z(n531) );
  XNOR U539 ( .A(n311), .B(n511), .Z(n513) );
  XNOR U540 ( .A(n534), .B(n535), .Z(n311) );
  AND U541 ( .A(n10), .B(n536), .Z(n535) );
  XOR U542 ( .A(n537), .B(n534), .Z(n536) );
  XOR U543 ( .A(n538), .B(n539), .Z(n511) );
  AND U544 ( .A(n540), .B(n541), .Z(n539) );
  XNOR U545 ( .A(n538), .B(n527), .Z(n541) );
  IV U546 ( .A(n364), .Z(n527) );
  XNOR U547 ( .A(n542), .B(n520), .Z(n364) );
  XNOR U548 ( .A(n543), .B(n526), .Z(n520) );
  XOR U549 ( .A(n544), .B(n545), .Z(n526) );
  AND U550 ( .A(n546), .B(n547), .Z(n545) );
  XOR U551 ( .A(n544), .B(n548), .Z(n546) );
  XNOR U552 ( .A(n525), .B(n517), .Z(n543) );
  XOR U553 ( .A(n549), .B(n550), .Z(n517) );
  AND U554 ( .A(n551), .B(n552), .Z(n550) );
  XNOR U555 ( .A(n553), .B(n549), .Z(n551) );
  XNOR U556 ( .A(n554), .B(n522), .Z(n525) );
  XOR U557 ( .A(n555), .B(n556), .Z(n522) );
  AND U558 ( .A(n557), .B(n558), .Z(n556) );
  XOR U559 ( .A(n555), .B(n559), .Z(n557) );
  XNOR U560 ( .A(n560), .B(n561), .Z(n554) );
  AND U561 ( .A(n562), .B(n563), .Z(n561) );
  XNOR U562 ( .A(n560), .B(n564), .Z(n562) );
  XNOR U563 ( .A(n521), .B(n528), .Z(n542) );
  AND U564 ( .A(n463), .B(n565), .Z(n528) );
  XOR U565 ( .A(n533), .B(n532), .Z(n521) );
  XNOR U566 ( .A(n566), .B(n529), .Z(n532) );
  XOR U567 ( .A(n567), .B(n568), .Z(n529) );
  AND U568 ( .A(n569), .B(n570), .Z(n568) );
  XOR U569 ( .A(n567), .B(n571), .Z(n569) );
  XNOR U570 ( .A(n572), .B(n573), .Z(n566) );
  AND U571 ( .A(n574), .B(n575), .Z(n573) );
  XOR U572 ( .A(n572), .B(n576), .Z(n574) );
  XOR U573 ( .A(n577), .B(n578), .Z(n533) );
  AND U574 ( .A(n579), .B(n580), .Z(n578) );
  XOR U575 ( .A(n577), .B(n581), .Z(n579) );
  XNOR U576 ( .A(n361), .B(n538), .Z(n540) );
  XNOR U577 ( .A(n582), .B(n583), .Z(n361) );
  AND U578 ( .A(n10), .B(n584), .Z(n583) );
  XNOR U579 ( .A(n585), .B(n582), .Z(n584) );
  XOR U580 ( .A(n586), .B(n587), .Z(n538) );
  AND U581 ( .A(n588), .B(n589), .Z(n587) );
  XNOR U582 ( .A(n586), .B(n463), .Z(n589) );
  XOR U583 ( .A(n590), .B(n552), .Z(n463) );
  XNOR U584 ( .A(n591), .B(n559), .Z(n552) );
  XOR U585 ( .A(n548), .B(n547), .Z(n559) );
  XNOR U586 ( .A(n592), .B(n544), .Z(n547) );
  XOR U587 ( .A(n593), .B(n594), .Z(n544) );
  AND U588 ( .A(n595), .B(n596), .Z(n594) );
  XOR U589 ( .A(n593), .B(n597), .Z(n595) );
  XNOR U590 ( .A(n598), .B(n599), .Z(n592) );
  NOR U591 ( .A(n600), .B(n601), .Z(n599) );
  XNOR U592 ( .A(n598), .B(n602), .Z(n600) );
  XOR U593 ( .A(n603), .B(n604), .Z(n548) );
  NOR U594 ( .A(n605), .B(n606), .Z(n604) );
  XNOR U595 ( .A(n603), .B(n607), .Z(n605) );
  XNOR U596 ( .A(n558), .B(n549), .Z(n591) );
  XOR U597 ( .A(n608), .B(n609), .Z(n549) );
  NOR U598 ( .A(n610), .B(n611), .Z(n609) );
  XNOR U599 ( .A(n608), .B(n612), .Z(n610) );
  XOR U600 ( .A(n613), .B(n564), .Z(n558) );
  XNOR U601 ( .A(n614), .B(n615), .Z(n564) );
  NOR U602 ( .A(n616), .B(n617), .Z(n615) );
  XNOR U603 ( .A(n614), .B(n618), .Z(n616) );
  XNOR U604 ( .A(n563), .B(n555), .Z(n613) );
  XOR U605 ( .A(n619), .B(n620), .Z(n555) );
  AND U606 ( .A(n621), .B(n622), .Z(n620) );
  XOR U607 ( .A(n619), .B(n623), .Z(n621) );
  XNOR U608 ( .A(n624), .B(n560), .Z(n563) );
  XOR U609 ( .A(n625), .B(n626), .Z(n560) );
  AND U610 ( .A(n627), .B(n628), .Z(n626) );
  XOR U611 ( .A(n625), .B(n629), .Z(n627) );
  XNOR U612 ( .A(n630), .B(n631), .Z(n624) );
  NOR U613 ( .A(n632), .B(n633), .Z(n631) );
  XOR U614 ( .A(n630), .B(n634), .Z(n632) );
  XOR U615 ( .A(n553), .B(n565), .Z(n590) );
  NOR U616 ( .A(n488), .B(n635), .Z(n565) );
  XNOR U617 ( .A(n571), .B(n570), .Z(n553) );
  XNOR U618 ( .A(n636), .B(n576), .Z(n570) );
  XOR U619 ( .A(n637), .B(n638), .Z(n576) );
  NOR U620 ( .A(n639), .B(n640), .Z(n638) );
  XNOR U621 ( .A(n637), .B(n641), .Z(n639) );
  XNOR U622 ( .A(n575), .B(n567), .Z(n636) );
  XOR U623 ( .A(n642), .B(n643), .Z(n567) );
  AND U624 ( .A(n644), .B(n645), .Z(n643) );
  XNOR U625 ( .A(n642), .B(n646), .Z(n644) );
  XNOR U626 ( .A(n647), .B(n572), .Z(n575) );
  XOR U627 ( .A(n648), .B(n649), .Z(n572) );
  AND U628 ( .A(n650), .B(n651), .Z(n649) );
  XOR U629 ( .A(n648), .B(n652), .Z(n650) );
  XNOR U630 ( .A(n653), .B(n654), .Z(n647) );
  NOR U631 ( .A(n655), .B(n656), .Z(n654) );
  XOR U632 ( .A(n653), .B(n657), .Z(n655) );
  XOR U633 ( .A(n581), .B(n580), .Z(n571) );
  XNOR U634 ( .A(n658), .B(n577), .Z(n580) );
  XOR U635 ( .A(n659), .B(n660), .Z(n577) );
  AND U636 ( .A(n661), .B(n662), .Z(n660) );
  XOR U637 ( .A(n659), .B(n663), .Z(n661) );
  XNOR U638 ( .A(n664), .B(n665), .Z(n658) );
  NOR U639 ( .A(n666), .B(n667), .Z(n665) );
  XNOR U640 ( .A(n664), .B(n668), .Z(n666) );
  XOR U641 ( .A(n669), .B(n670), .Z(n581) );
  NOR U642 ( .A(n671), .B(n672), .Z(n670) );
  XNOR U643 ( .A(n669), .B(n673), .Z(n671) );
  XNOR U644 ( .A(n459), .B(n586), .Z(n588) );
  XNOR U645 ( .A(n674), .B(n675), .Z(n459) );
  AND U646 ( .A(n10), .B(n676), .Z(n675) );
  XOR U647 ( .A(n677), .B(n674), .Z(n676) );
  AND U648 ( .A(n489), .B(n488), .Z(n586) );
  XOR U649 ( .A(n678), .B(n635), .Z(n488) );
  XNOR U650 ( .A(p_input[128]), .B(p_input[32]), .Z(n635) );
  XOR U651 ( .A(n612), .B(n611), .Z(n678) );
  XOR U652 ( .A(n679), .B(n623), .Z(n611) );
  XOR U653 ( .A(n597), .B(n596), .Z(n623) );
  XNOR U654 ( .A(n680), .B(n602), .Z(n596) );
  XNOR U655 ( .A(n681), .B(p_input[56]), .Z(n602) );
  XOR U656 ( .A(n593), .B(n601), .Z(n680) );
  XOR U657 ( .A(n682), .B(n598), .Z(n601) );
  XOR U658 ( .A(p_input[150]), .B(p_input[54]), .Z(n598) );
  XNOR U659 ( .A(p_input[151]), .B(p_input[55]), .Z(n682) );
  XOR U660 ( .A(p_input[146]), .B(p_input[50]), .Z(n593) );
  XNOR U661 ( .A(n607), .B(n606), .Z(n597) );
  XOR U662 ( .A(n683), .B(n603), .Z(n606) );
  XOR U663 ( .A(p_input[147]), .B(p_input[51]), .Z(n603) );
  XNOR U664 ( .A(p_input[148]), .B(p_input[52]), .Z(n683) );
  XNOR U665 ( .A(n684), .B(p_input[53]), .Z(n607) );
  XNOR U666 ( .A(n622), .B(n608), .Z(n679) );
  XNOR U667 ( .A(n685), .B(p_input[33]), .Z(n608) );
  XNOR U668 ( .A(n686), .B(n629), .Z(n622) );
  XNOR U669 ( .A(n618), .B(n617), .Z(n629) );
  XOR U670 ( .A(n687), .B(n614), .Z(n617) );
  XNOR U671 ( .A(n688), .B(p_input[58]), .Z(n614) );
  XNOR U672 ( .A(p_input[155]), .B(p_input[59]), .Z(n687) );
  XNOR U673 ( .A(n689), .B(p_input[60]), .Z(n618) );
  XNOR U674 ( .A(n628), .B(n619), .Z(n686) );
  XNOR U675 ( .A(n690), .B(p_input[49]), .Z(n619) );
  XOR U676 ( .A(n691), .B(n634), .Z(n628) );
  XNOR U677 ( .A(p_input[159]), .B(p_input[63]), .Z(n634) );
  XOR U678 ( .A(n625), .B(n633), .Z(n691) );
  XOR U679 ( .A(n692), .B(n630), .Z(n633) );
  XOR U680 ( .A(p_input[157]), .B(p_input[61]), .Z(n630) );
  XNOR U681 ( .A(p_input[158]), .B(p_input[62]), .Z(n692) );
  XOR U682 ( .A(p_input[153]), .B(p_input[57]), .Z(n625) );
  XNOR U683 ( .A(n646), .B(n645), .Z(n612) );
  XNOR U684 ( .A(n693), .B(n652), .Z(n645) );
  XNOR U685 ( .A(n641), .B(n640), .Z(n652) );
  XOR U686 ( .A(n694), .B(n637), .Z(n640) );
  XOR U687 ( .A(p_input[139]), .B(p_input[43]), .Z(n637) );
  XNOR U688 ( .A(p_input[140]), .B(p_input[44]), .Z(n694) );
  XOR U689 ( .A(p_input[141]), .B(p_input[45]), .Z(n641) );
  XNOR U690 ( .A(n651), .B(n642), .Z(n693) );
  XNOR U691 ( .A(n695), .B(p_input[34]), .Z(n642) );
  XOR U692 ( .A(n696), .B(n657), .Z(n651) );
  XNOR U693 ( .A(p_input[144]), .B(p_input[48]), .Z(n657) );
  XOR U694 ( .A(n648), .B(n656), .Z(n696) );
  XOR U695 ( .A(n697), .B(n653), .Z(n656) );
  XOR U696 ( .A(p_input[142]), .B(p_input[46]), .Z(n653) );
  XNOR U697 ( .A(p_input[143]), .B(p_input[47]), .Z(n697) );
  XOR U698 ( .A(p_input[138]), .B(p_input[42]), .Z(n648) );
  XNOR U699 ( .A(n663), .B(n662), .Z(n646) );
  XNOR U700 ( .A(n698), .B(n668), .Z(n662) );
  XNOR U701 ( .A(n699), .B(p_input[41]), .Z(n668) );
  XOR U702 ( .A(n659), .B(n667), .Z(n698) );
  XOR U703 ( .A(n700), .B(n664), .Z(n667) );
  XOR U704 ( .A(p_input[135]), .B(p_input[39]), .Z(n664) );
  XNOR U705 ( .A(p_input[136]), .B(p_input[40]), .Z(n700) );
  XOR U706 ( .A(p_input[131]), .B(p_input[35]), .Z(n659) );
  XNOR U707 ( .A(n673), .B(n672), .Z(n663) );
  XOR U708 ( .A(n701), .B(n669), .Z(n672) );
  XOR U709 ( .A(p_input[132]), .B(p_input[36]), .Z(n669) );
  XNOR U710 ( .A(p_input[133]), .B(p_input[37]), .Z(n701) );
  XNOR U711 ( .A(n702), .B(p_input[38]), .Z(n673) );
  IV U712 ( .A(n485), .Z(n489) );
  XNOR U713 ( .A(n703), .B(n704), .Z(n485) );
  AND U714 ( .A(n10), .B(n705), .Z(n704) );
  XNOR U715 ( .A(n706), .B(n703), .Z(n705) );
  XNOR U716 ( .A(n707), .B(n708), .Z(n10) );
  MUX U717 ( .IN0(n492), .IN1(n493), .SEL(n707), .F(n708) );
  AND U718 ( .A(n507), .B(n709), .Z(n493) );
  AND U719 ( .A(n710), .B(n711), .Z(n492) );
  XOR U720 ( .A(n712), .B(n713), .Z(n707) );
  AND U721 ( .A(n714), .B(n715), .Z(n713) );
  XNOR U722 ( .A(n712), .B(n710), .Z(n715) );
  IV U723 ( .A(n510), .Z(n710) );
  XOR U724 ( .A(n716), .B(n717), .Z(n510) );
  XOR U725 ( .A(n718), .B(n711), .Z(n717) );
  AND U726 ( .A(n537), .B(n719), .Z(n711) );
  AND U727 ( .A(n720), .B(n721), .Z(n718) );
  XOR U728 ( .A(n722), .B(n716), .Z(n720) );
  XNOR U729 ( .A(n723), .B(n712), .Z(n714) );
  IV U730 ( .A(n507), .Z(n723) );
  XNOR U731 ( .A(n724), .B(n725), .Z(n507) );
  XOR U732 ( .A(n726), .B(n709), .Z(n725) );
  AND U733 ( .A(n534), .B(n727), .Z(n709) );
  AND U734 ( .A(n728), .B(n729), .Z(n726) );
  XNOR U735 ( .A(n724), .B(n730), .Z(n728) );
  XOR U736 ( .A(n731), .B(n732), .Z(n712) );
  AND U737 ( .A(n733), .B(n734), .Z(n732) );
  XNOR U738 ( .A(n731), .B(n537), .Z(n734) );
  XOR U739 ( .A(n735), .B(n721), .Z(n537) );
  XNOR U740 ( .A(n736), .B(n716), .Z(n721) );
  XOR U741 ( .A(n737), .B(n738), .Z(n716) );
  AND U742 ( .A(n739), .B(n740), .Z(n738) );
  XOR U743 ( .A(n741), .B(n737), .Z(n739) );
  XNOR U744 ( .A(n742), .B(n743), .Z(n736) );
  AND U745 ( .A(n744), .B(n745), .Z(n743) );
  XOR U746 ( .A(n742), .B(n746), .Z(n744) );
  XNOR U747 ( .A(n722), .B(n719), .Z(n735) );
  AND U748 ( .A(n747), .B(n748), .Z(n719) );
  XOR U749 ( .A(n749), .B(n750), .Z(n722) );
  AND U750 ( .A(n751), .B(n752), .Z(n750) );
  XOR U751 ( .A(n749), .B(n753), .Z(n751) );
  XOR U752 ( .A(n534), .B(n731), .Z(n733) );
  XNOR U753 ( .A(n754), .B(n730), .Z(n534) );
  XNOR U754 ( .A(n755), .B(n756), .Z(n730) );
  AND U755 ( .A(n757), .B(n758), .Z(n756) );
  XOR U756 ( .A(n755), .B(n759), .Z(n757) );
  XNOR U757 ( .A(n729), .B(n727), .Z(n754) );
  AND U758 ( .A(n582), .B(n760), .Z(n727) );
  XNOR U759 ( .A(n761), .B(n724), .Z(n729) );
  XOR U760 ( .A(n762), .B(n763), .Z(n724) );
  AND U761 ( .A(n764), .B(n765), .Z(n763) );
  XOR U762 ( .A(n762), .B(n766), .Z(n764) );
  XNOR U763 ( .A(n767), .B(n768), .Z(n761) );
  AND U764 ( .A(n769), .B(n770), .Z(n768) );
  XNOR U765 ( .A(n767), .B(n771), .Z(n769) );
  XOR U766 ( .A(n772), .B(n773), .Z(n731) );
  AND U767 ( .A(n774), .B(n775), .Z(n773) );
  XNOR U768 ( .A(n772), .B(n747), .Z(n775) );
  IV U769 ( .A(n585), .Z(n747) );
  XNOR U770 ( .A(n776), .B(n740), .Z(n585) );
  XNOR U771 ( .A(n777), .B(n746), .Z(n740) );
  XOR U772 ( .A(n778), .B(n779), .Z(n746) );
  AND U773 ( .A(n780), .B(n781), .Z(n779) );
  XOR U774 ( .A(n778), .B(n782), .Z(n780) );
  XNOR U775 ( .A(n745), .B(n737), .Z(n777) );
  XOR U776 ( .A(n783), .B(n784), .Z(n737) );
  AND U777 ( .A(n785), .B(n786), .Z(n784) );
  XNOR U778 ( .A(n787), .B(n783), .Z(n785) );
  XNOR U779 ( .A(n788), .B(n742), .Z(n745) );
  XOR U780 ( .A(n789), .B(n790), .Z(n742) );
  AND U781 ( .A(n791), .B(n792), .Z(n790) );
  XOR U782 ( .A(n789), .B(n793), .Z(n791) );
  XNOR U783 ( .A(n794), .B(n795), .Z(n788) );
  AND U784 ( .A(n796), .B(n797), .Z(n795) );
  XNOR U785 ( .A(n794), .B(n798), .Z(n796) );
  XNOR U786 ( .A(n741), .B(n748), .Z(n776) );
  AND U787 ( .A(n677), .B(n799), .Z(n748) );
  XOR U788 ( .A(n753), .B(n752), .Z(n741) );
  XNOR U789 ( .A(n800), .B(n749), .Z(n752) );
  XOR U790 ( .A(n801), .B(n802), .Z(n749) );
  AND U791 ( .A(n803), .B(n804), .Z(n802) );
  XOR U792 ( .A(n801), .B(n805), .Z(n803) );
  XNOR U793 ( .A(n806), .B(n807), .Z(n800) );
  AND U794 ( .A(n808), .B(n809), .Z(n807) );
  XOR U795 ( .A(n806), .B(n810), .Z(n808) );
  XOR U796 ( .A(n811), .B(n812), .Z(n753) );
  AND U797 ( .A(n813), .B(n814), .Z(n812) );
  XOR U798 ( .A(n811), .B(n815), .Z(n813) );
  XNOR U799 ( .A(n816), .B(n772), .Z(n774) );
  IV U800 ( .A(n582), .Z(n816) );
  XOR U801 ( .A(n817), .B(n766), .Z(n582) );
  XOR U802 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U803 ( .A(n818), .B(n755), .Z(n758) );
  XOR U804 ( .A(n819), .B(n820), .Z(n755) );
  AND U805 ( .A(n821), .B(n822), .Z(n820) );
  XOR U806 ( .A(n819), .B(n823), .Z(n821) );
  XNOR U807 ( .A(n824), .B(n825), .Z(n818) );
  AND U808 ( .A(n826), .B(n827), .Z(n825) );
  XOR U809 ( .A(n824), .B(n828), .Z(n826) );
  XOR U810 ( .A(n829), .B(n830), .Z(n759) );
  AND U811 ( .A(n831), .B(n832), .Z(n830) );
  XOR U812 ( .A(n829), .B(n833), .Z(n831) );
  XNOR U813 ( .A(n765), .B(n760), .Z(n817) );
  AND U814 ( .A(n674), .B(n834), .Z(n760) );
  XOR U815 ( .A(n835), .B(n771), .Z(n765) );
  XNOR U816 ( .A(n836), .B(n837), .Z(n771) );
  AND U817 ( .A(n838), .B(n839), .Z(n837) );
  XOR U818 ( .A(n836), .B(n840), .Z(n838) );
  XNOR U819 ( .A(n770), .B(n762), .Z(n835) );
  XOR U820 ( .A(n841), .B(n842), .Z(n762) );
  AND U821 ( .A(n843), .B(n844), .Z(n842) );
  XOR U822 ( .A(n841), .B(n845), .Z(n843) );
  XNOR U823 ( .A(n846), .B(n767), .Z(n770) );
  XOR U824 ( .A(n847), .B(n848), .Z(n767) );
  AND U825 ( .A(n849), .B(n850), .Z(n848) );
  XOR U826 ( .A(n847), .B(n851), .Z(n849) );
  XNOR U827 ( .A(n852), .B(n853), .Z(n846) );
  AND U828 ( .A(n854), .B(n855), .Z(n853) );
  XNOR U829 ( .A(n852), .B(n856), .Z(n854) );
  XOR U830 ( .A(n857), .B(n858), .Z(n772) );
  AND U831 ( .A(n859), .B(n860), .Z(n858) );
  XNOR U832 ( .A(n857), .B(n677), .Z(n860) );
  XOR U833 ( .A(n861), .B(n786), .Z(n677) );
  XNOR U834 ( .A(n862), .B(n793), .Z(n786) );
  XOR U835 ( .A(n782), .B(n781), .Z(n793) );
  XNOR U836 ( .A(n863), .B(n778), .Z(n781) );
  XOR U837 ( .A(n864), .B(n865), .Z(n778) );
  AND U838 ( .A(n866), .B(n867), .Z(n865) );
  XOR U839 ( .A(n864), .B(n868), .Z(n866) );
  XNOR U840 ( .A(n869), .B(n870), .Z(n863) );
  NOR U841 ( .A(n871), .B(n872), .Z(n870) );
  XNOR U842 ( .A(n869), .B(n873), .Z(n871) );
  XOR U843 ( .A(n874), .B(n875), .Z(n782) );
  NOR U844 ( .A(n876), .B(n877), .Z(n875) );
  XNOR U845 ( .A(n874), .B(n878), .Z(n876) );
  XNOR U846 ( .A(n792), .B(n783), .Z(n862) );
  XOR U847 ( .A(n879), .B(n880), .Z(n783) );
  NOR U848 ( .A(n881), .B(n882), .Z(n880) );
  XNOR U849 ( .A(n879), .B(n883), .Z(n881) );
  XOR U850 ( .A(n884), .B(n798), .Z(n792) );
  XNOR U851 ( .A(n885), .B(n886), .Z(n798) );
  NOR U852 ( .A(n887), .B(n888), .Z(n886) );
  XNOR U853 ( .A(n885), .B(n889), .Z(n887) );
  XNOR U854 ( .A(n797), .B(n789), .Z(n884) );
  XOR U855 ( .A(n890), .B(n891), .Z(n789) );
  AND U856 ( .A(n892), .B(n893), .Z(n891) );
  XOR U857 ( .A(n890), .B(n894), .Z(n892) );
  XNOR U858 ( .A(n895), .B(n794), .Z(n797) );
  XOR U859 ( .A(n896), .B(n897), .Z(n794) );
  AND U860 ( .A(n898), .B(n899), .Z(n897) );
  XOR U861 ( .A(n896), .B(n900), .Z(n898) );
  XNOR U862 ( .A(n901), .B(n902), .Z(n895) );
  NOR U863 ( .A(n903), .B(n904), .Z(n902) );
  XOR U864 ( .A(n901), .B(n905), .Z(n903) );
  XOR U865 ( .A(n787), .B(n799), .Z(n861) );
  NOR U866 ( .A(n706), .B(n906), .Z(n799) );
  XNOR U867 ( .A(n805), .B(n804), .Z(n787) );
  XNOR U868 ( .A(n907), .B(n810), .Z(n804) );
  XOR U869 ( .A(n908), .B(n909), .Z(n810) );
  NOR U870 ( .A(n910), .B(n911), .Z(n909) );
  XNOR U871 ( .A(n908), .B(n912), .Z(n910) );
  XNOR U872 ( .A(n809), .B(n801), .Z(n907) );
  XOR U873 ( .A(n913), .B(n914), .Z(n801) );
  AND U874 ( .A(n915), .B(n916), .Z(n914) );
  XNOR U875 ( .A(n913), .B(n917), .Z(n915) );
  XNOR U876 ( .A(n918), .B(n806), .Z(n809) );
  XOR U877 ( .A(n919), .B(n920), .Z(n806) );
  AND U878 ( .A(n921), .B(n922), .Z(n920) );
  XOR U879 ( .A(n919), .B(n923), .Z(n921) );
  XNOR U880 ( .A(n924), .B(n925), .Z(n918) );
  NOR U881 ( .A(n926), .B(n927), .Z(n925) );
  XOR U882 ( .A(n924), .B(n928), .Z(n926) );
  XOR U883 ( .A(n815), .B(n814), .Z(n805) );
  XNOR U884 ( .A(n929), .B(n811), .Z(n814) );
  XOR U885 ( .A(n930), .B(n931), .Z(n811) );
  AND U886 ( .A(n932), .B(n933), .Z(n931) );
  XOR U887 ( .A(n930), .B(n934), .Z(n932) );
  XNOR U888 ( .A(n935), .B(n936), .Z(n929) );
  NOR U889 ( .A(n937), .B(n938), .Z(n936) );
  XNOR U890 ( .A(n935), .B(n939), .Z(n937) );
  XOR U891 ( .A(n940), .B(n941), .Z(n815) );
  NOR U892 ( .A(n942), .B(n943), .Z(n941) );
  XNOR U893 ( .A(n940), .B(n944), .Z(n942) );
  XNOR U894 ( .A(n945), .B(n857), .Z(n859) );
  IV U895 ( .A(n674), .Z(n945) );
  XOR U896 ( .A(n946), .B(n845), .Z(n674) );
  XOR U897 ( .A(n823), .B(n822), .Z(n845) );
  XNOR U898 ( .A(n947), .B(n828), .Z(n822) );
  XOR U899 ( .A(n948), .B(n949), .Z(n828) );
  NOR U900 ( .A(n950), .B(n951), .Z(n949) );
  XNOR U901 ( .A(n948), .B(n952), .Z(n950) );
  XNOR U902 ( .A(n827), .B(n819), .Z(n947) );
  XOR U903 ( .A(n953), .B(n954), .Z(n819) );
  AND U904 ( .A(n955), .B(n956), .Z(n954) );
  XNOR U905 ( .A(n953), .B(n957), .Z(n955) );
  XNOR U906 ( .A(n958), .B(n824), .Z(n827) );
  XOR U907 ( .A(n959), .B(n960), .Z(n824) );
  AND U908 ( .A(n961), .B(n962), .Z(n960) );
  XOR U909 ( .A(n959), .B(n963), .Z(n961) );
  XNOR U910 ( .A(n964), .B(n965), .Z(n958) );
  AND U911 ( .A(n966), .B(n967), .Z(n965) );
  XNOR U912 ( .A(n964), .B(n968), .Z(n966) );
  XOR U913 ( .A(n833), .B(n832), .Z(n823) );
  XNOR U914 ( .A(n969), .B(n829), .Z(n832) );
  XOR U915 ( .A(n970), .B(n971), .Z(n829) );
  AND U916 ( .A(n972), .B(n973), .Z(n971) );
  XNOR U917 ( .A(n974), .B(n975), .Z(n972) );
  IV U918 ( .A(n970), .Z(n974) );
  XNOR U919 ( .A(n976), .B(n977), .Z(n969) );
  AND U920 ( .A(n978), .B(n979), .Z(n977) );
  XNOR U921 ( .A(n976), .B(n980), .Z(n978) );
  XOR U922 ( .A(n981), .B(n982), .Z(n833) );
  AND U923 ( .A(n983), .B(n984), .Z(n982) );
  XOR U924 ( .A(n981), .B(n985), .Z(n983) );
  XNOR U925 ( .A(n844), .B(n834), .Z(n946) );
  AND U926 ( .A(n703), .B(n986), .Z(n834) );
  XNOR U927 ( .A(n987), .B(n851), .Z(n844) );
  XOR U928 ( .A(n840), .B(n839), .Z(n851) );
  XNOR U929 ( .A(n988), .B(n836), .Z(n839) );
  XOR U930 ( .A(n989), .B(n990), .Z(n836) );
  AND U931 ( .A(n991), .B(n992), .Z(n990) );
  XNOR U932 ( .A(n993), .B(n994), .Z(n991) );
  IV U933 ( .A(n989), .Z(n993) );
  XNOR U934 ( .A(n995), .B(n996), .Z(n988) );
  AND U935 ( .A(n997), .B(n998), .Z(n996) );
  XNOR U936 ( .A(n995), .B(n999), .Z(n997) );
  XOR U937 ( .A(n1000), .B(n1001), .Z(n840) );
  AND U938 ( .A(n1002), .B(n1003), .Z(n1001) );
  XOR U939 ( .A(n1000), .B(n1004), .Z(n1002) );
  XNOR U940 ( .A(n850), .B(n841), .Z(n987) );
  XOR U941 ( .A(n1005), .B(n1006), .Z(n841) );
  NOR U942 ( .A(n1007), .B(n1008), .Z(n1006) );
  XNOR U943 ( .A(n1005), .B(n1009), .Z(n1007) );
  XOR U944 ( .A(n1010), .B(n856), .Z(n850) );
  XNOR U945 ( .A(n1011), .B(n1012), .Z(n856) );
  AND U946 ( .A(n1013), .B(n1014), .Z(n1012) );
  XOR U947 ( .A(n1011), .B(n1015), .Z(n1013) );
  XNOR U948 ( .A(n855), .B(n847), .Z(n1010) );
  XOR U949 ( .A(n1016), .B(n1017), .Z(n847) );
  AND U950 ( .A(n1018), .B(n1019), .Z(n1017) );
  XOR U951 ( .A(n1016), .B(n1020), .Z(n1018) );
  XNOR U952 ( .A(n1021), .B(n852), .Z(n855) );
  XOR U953 ( .A(n1022), .B(n1023), .Z(n852) );
  AND U954 ( .A(n1024), .B(n1025), .Z(n1023) );
  XNOR U955 ( .A(n1026), .B(n1027), .Z(n1024) );
  IV U956 ( .A(n1022), .Z(n1026) );
  XNOR U957 ( .A(n1028), .B(n1029), .Z(n1021) );
  AND U958 ( .A(n1030), .B(n1031), .Z(n1029) );
  XNOR U959 ( .A(n1028), .B(n1032), .Z(n1030) );
  AND U960 ( .A(n703), .B(n706), .Z(n857) );
  XOR U961 ( .A(n1033), .B(n906), .Z(n706) );
  XNOR U962 ( .A(p_input[128]), .B(p_input[64]), .Z(n906) );
  XOR U963 ( .A(n883), .B(n882), .Z(n1033) );
  XOR U964 ( .A(n1034), .B(n894), .Z(n882) );
  XOR U965 ( .A(n868), .B(n867), .Z(n894) );
  XNOR U966 ( .A(n1035), .B(n873), .Z(n867) );
  XNOR U967 ( .A(n681), .B(p_input[88]), .Z(n873) );
  IV U968 ( .A(p_input[152]), .Z(n681) );
  XOR U969 ( .A(n864), .B(n872), .Z(n1035) );
  XOR U970 ( .A(n1036), .B(n869), .Z(n872) );
  XOR U971 ( .A(p_input[150]), .B(p_input[86]), .Z(n869) );
  XNOR U972 ( .A(p_input[151]), .B(p_input[87]), .Z(n1036) );
  XOR U973 ( .A(p_input[146]), .B(p_input[82]), .Z(n864) );
  XNOR U974 ( .A(n878), .B(n877), .Z(n868) );
  XOR U975 ( .A(n1037), .B(n874), .Z(n877) );
  XOR U976 ( .A(p_input[147]), .B(p_input[83]), .Z(n874) );
  XNOR U977 ( .A(p_input[148]), .B(p_input[84]), .Z(n1037) );
  XNOR U978 ( .A(n684), .B(p_input[85]), .Z(n878) );
  IV U979 ( .A(p_input[149]), .Z(n684) );
  XNOR U980 ( .A(n893), .B(n879), .Z(n1034) );
  XNOR U981 ( .A(n685), .B(p_input[65]), .Z(n879) );
  IV U982 ( .A(p_input[129]), .Z(n685) );
  XNOR U983 ( .A(n1038), .B(n900), .Z(n893) );
  XNOR U984 ( .A(n889), .B(n888), .Z(n900) );
  XOR U985 ( .A(n1039), .B(n885), .Z(n888) );
  XNOR U986 ( .A(n688), .B(p_input[90]), .Z(n885) );
  IV U987 ( .A(p_input[154]), .Z(n688) );
  XNOR U988 ( .A(p_input[155]), .B(p_input[91]), .Z(n1039) );
  XNOR U989 ( .A(n689), .B(p_input[92]), .Z(n889) );
  IV U990 ( .A(p_input[156]), .Z(n689) );
  XNOR U991 ( .A(n899), .B(n890), .Z(n1038) );
  XNOR U992 ( .A(n690), .B(p_input[81]), .Z(n890) );
  IV U993 ( .A(p_input[145]), .Z(n690) );
  XOR U994 ( .A(n1040), .B(n905), .Z(n899) );
  XNOR U995 ( .A(p_input[159]), .B(p_input[95]), .Z(n905) );
  XOR U996 ( .A(n896), .B(n904), .Z(n1040) );
  XOR U997 ( .A(n1041), .B(n901), .Z(n904) );
  XOR U998 ( .A(p_input[157]), .B(p_input[93]), .Z(n901) );
  XNOR U999 ( .A(p_input[158]), .B(p_input[94]), .Z(n1041) );
  XOR U1000 ( .A(p_input[153]), .B(p_input[89]), .Z(n896) );
  XNOR U1001 ( .A(n917), .B(n916), .Z(n883) );
  XNOR U1002 ( .A(n1042), .B(n923), .Z(n916) );
  XNOR U1003 ( .A(n912), .B(n911), .Z(n923) );
  XOR U1004 ( .A(n1043), .B(n908), .Z(n911) );
  XOR U1005 ( .A(p_input[139]), .B(p_input[75]), .Z(n908) );
  XNOR U1006 ( .A(p_input[140]), .B(p_input[76]), .Z(n1043) );
  XOR U1007 ( .A(p_input[141]), .B(p_input[77]), .Z(n912) );
  XNOR U1008 ( .A(n922), .B(n913), .Z(n1042) );
  XNOR U1009 ( .A(n695), .B(p_input[66]), .Z(n913) );
  IV U1010 ( .A(p_input[130]), .Z(n695) );
  XOR U1011 ( .A(n1044), .B(n928), .Z(n922) );
  XNOR U1012 ( .A(p_input[144]), .B(p_input[80]), .Z(n928) );
  XOR U1013 ( .A(n919), .B(n927), .Z(n1044) );
  XOR U1014 ( .A(n1045), .B(n924), .Z(n927) );
  XOR U1015 ( .A(p_input[142]), .B(p_input[78]), .Z(n924) );
  XNOR U1016 ( .A(p_input[143]), .B(p_input[79]), .Z(n1045) );
  XOR U1017 ( .A(p_input[138]), .B(p_input[74]), .Z(n919) );
  XNOR U1018 ( .A(n934), .B(n933), .Z(n917) );
  XNOR U1019 ( .A(n1046), .B(n939), .Z(n933) );
  XNOR U1020 ( .A(n699), .B(p_input[73]), .Z(n939) );
  IV U1021 ( .A(p_input[137]), .Z(n699) );
  XOR U1022 ( .A(n930), .B(n938), .Z(n1046) );
  XOR U1023 ( .A(n1047), .B(n935), .Z(n938) );
  XOR U1024 ( .A(p_input[135]), .B(p_input[71]), .Z(n935) );
  XNOR U1025 ( .A(p_input[136]), .B(p_input[72]), .Z(n1047) );
  XOR U1026 ( .A(p_input[131]), .B(p_input[67]), .Z(n930) );
  XNOR U1027 ( .A(n944), .B(n943), .Z(n934) );
  XOR U1028 ( .A(n1048), .B(n940), .Z(n943) );
  XOR U1029 ( .A(p_input[132]), .B(p_input[68]), .Z(n940) );
  XNOR U1030 ( .A(p_input[133]), .B(p_input[69]), .Z(n1048) );
  XNOR U1031 ( .A(n702), .B(p_input[70]), .Z(n944) );
  IV U1032 ( .A(p_input[134]), .Z(n702) );
  XOR U1033 ( .A(n1049), .B(n1009), .Z(n703) );
  XNOR U1034 ( .A(n957), .B(n956), .Z(n1009) );
  XNOR U1035 ( .A(n1050), .B(n963), .Z(n956) );
  XNOR U1036 ( .A(n952), .B(n951), .Z(n963) );
  XOR U1037 ( .A(n1051), .B(n948), .Z(n951) );
  XOR U1038 ( .A(\knn_comb_/min_val_out[0][11] ), .B(p_input[139]), .Z(n948)
         );
  XOR U1039 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n478), .Z(n1051) );
  IV U1040 ( .A(p_input[140]), .Z(n478) );
  XOR U1041 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[141]), .Z(n952)
         );
  XNOR U1042 ( .A(n962), .B(n953), .Z(n1050) );
  XOR U1043 ( .A(\knn_comb_/min_val_out[0][2] ), .B(p_input[130]), .Z(n953) );
  XOR U1044 ( .A(n1052), .B(n968), .Z(n962) );
  XNOR U1045 ( .A(\knn_comb_/min_val_out[0][16] ), .B(p_input[144]), .Z(n968)
         );
  XNOR U1046 ( .A(n959), .B(n967), .Z(n1052) );
  XNOR U1047 ( .A(n1053), .B(n964), .Z(n967) );
  XOR U1048 ( .A(\knn_comb_/min_val_out[0][14] ), .B(p_input[142]), .Z(n964)
         );
  XNOR U1049 ( .A(\knn_comb_/min_val_out[0][15] ), .B(p_input[143]), .Z(n1053)
         );
  XOR U1050 ( .A(\knn_comb_/min_val_out[0][10] ), .B(p_input[138]), .Z(n959)
         );
  XNOR U1051 ( .A(n975), .B(n973), .Z(n957) );
  XOR U1052 ( .A(n1054), .B(n980), .Z(n973) );
  XNOR U1053 ( .A(\knn_comb_/min_val_out[0][9] ), .B(p_input[137]), .Z(n980)
         );
  XNOR U1054 ( .A(n970), .B(n979), .Z(n1054) );
  XNOR U1055 ( .A(n1055), .B(n976), .Z(n979) );
  XOR U1056 ( .A(\knn_comb_/min_val_out[0][7] ), .B(p_input[135]), .Z(n976) );
  XNOR U1057 ( .A(\knn_comb_/min_val_out[0][8] ), .B(p_input[136]), .Z(n1055)
         );
  XOR U1058 ( .A(\knn_comb_/min_val_out[0][3] ), .B(p_input[131]), .Z(n970) );
  XOR U1059 ( .A(n985), .B(n984), .Z(n975) );
  XNOR U1060 ( .A(n1056), .B(n981), .Z(n984) );
  XOR U1061 ( .A(\knn_comb_/min_val_out[0][4] ), .B(p_input[132]), .Z(n981) );
  XNOR U1062 ( .A(\knn_comb_/min_val_out[0][5] ), .B(p_input[133]), .Z(n1056)
         );
  XOR U1063 ( .A(\knn_comb_/min_val_out[0][6] ), .B(p_input[134]), .Z(n985) );
  XOR U1064 ( .A(n1008), .B(n986), .Z(n1049) );
  XOR U1065 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[128]), .Z(n986) );
  XOR U1066 ( .A(n1057), .B(n1020), .Z(n1008) );
  XOR U1067 ( .A(n994), .B(n992), .Z(n1020) );
  XOR U1068 ( .A(n1058), .B(n999), .Z(n992) );
  XNOR U1069 ( .A(\knn_comb_/min_val_out[0][24] ), .B(p_input[152]), .Z(n999)
         );
  XNOR U1070 ( .A(n989), .B(n998), .Z(n1058) );
  XNOR U1071 ( .A(n1059), .B(n995), .Z(n998) );
  XOR U1072 ( .A(\knn_comb_/min_val_out[0][22] ), .B(p_input[150]), .Z(n995)
         );
  XNOR U1073 ( .A(\knn_comb_/min_val_out[0][23] ), .B(p_input[151]), .Z(n1059)
         );
  XOR U1074 ( .A(\knn_comb_/min_val_out[0][18] ), .B(p_input[146]), .Z(n989)
         );
  XOR U1075 ( .A(n1004), .B(n1003), .Z(n994) );
  XNOR U1076 ( .A(n1060), .B(n1000), .Z(n1003) );
  XOR U1077 ( .A(\knn_comb_/min_val_out[0][19] ), .B(p_input[147]), .Z(n1000)
         );
  XNOR U1078 ( .A(\knn_comb_/min_val_out[0][20] ), .B(p_input[148]), .Z(n1060)
         );
  XOR U1079 ( .A(\knn_comb_/min_val_out[0][21] ), .B(p_input[149]), .Z(n1004)
         );
  XNOR U1080 ( .A(n1019), .B(n1005), .Z(n1057) );
  XOR U1081 ( .A(\knn_comb_/min_val_out[0][1] ), .B(p_input[129]), .Z(n1005)
         );
  XNOR U1082 ( .A(n1061), .B(n1027), .Z(n1019) );
  XOR U1083 ( .A(n1015), .B(n1014), .Z(n1027) );
  XNOR U1084 ( .A(n1062), .B(n1011), .Z(n1014) );
  XOR U1085 ( .A(\knn_comb_/min_val_out[0][26] ), .B(p_input[154]), .Z(n1011)
         );
  XNOR U1086 ( .A(\knn_comb_/min_val_out[0][27] ), .B(p_input[155]), .Z(n1062)
         );
  XOR U1087 ( .A(\knn_comb_/min_val_out[0][28] ), .B(p_input[156]), .Z(n1015)
         );
  XNOR U1088 ( .A(n1025), .B(n1016), .Z(n1061) );
  XOR U1089 ( .A(\knn_comb_/min_val_out[0][17] ), .B(p_input[145]), .Z(n1016)
         );
  XOR U1090 ( .A(n1063), .B(n1032), .Z(n1025) );
  XNOR U1091 ( .A(\knn_comb_/min_val_out[0][31] ), .B(p_input[159]), .Z(n1032)
         );
  XNOR U1092 ( .A(n1022), .B(n1031), .Z(n1063) );
  XNOR U1093 ( .A(n1064), .B(n1028), .Z(n1031) );
  XOR U1094 ( .A(\knn_comb_/min_val_out[0][29] ), .B(p_input[157]), .Z(n1028)
         );
  XNOR U1095 ( .A(\knn_comb_/min_val_out[0][30] ), .B(p_input[158]), .Z(n1064)
         );
  XOR U1096 ( .A(\knn_comb_/min_val_out[0][25] ), .B(p_input[153]), .Z(n1022)
         );
endmodule

