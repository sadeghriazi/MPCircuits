
module voting_N1_M4 ( p_input, o );
  input [15:0] p_input;
  output [0:0] o;
  wire   \dV[15][1] , \dV[14][1] , \dV[13][1] , \dV[12][1] , \dV[11][1] ,
         \dV[10][1] , \dV[9][1] , \dV[8][1] , \dV[7][1] , \dV[6][1] ,
         \dV[5][1] , \dV[4][1] , \dV[3][1] , \dV[2][1] , \dV[1][1] ,
         \dV[0][1] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204;
  assign \dV[15][1]  = p_input[15];
  assign \dV[14][1]  = p_input[14];
  assign \dV[13][1]  = p_input[13];
  assign \dV[12][1]  = p_input[12];
  assign \dV[11][1]  = p_input[11];
  assign \dV[10][1]  = p_input[10];
  assign \dV[9][1]  = p_input[9];
  assign \dV[8][1]  = p_input[8];
  assign \dV[7][1]  = p_input[7];
  assign \dV[6][1]  = p_input[6];
  assign \dV[5][1]  = p_input[5];
  assign \dV[4][1]  = p_input[4];
  assign \dV[3][1]  = p_input[3];
  assign \dV[2][1]  = p_input[2];
  assign \dV[1][1]  = p_input[1];
  assign \dV[0][1]  = p_input[0];

  XOR U2 ( .A(n1), .B(n2), .Z(o[0]) );
  AND U3 ( .A(n3), .B(n4), .Z(n2) );
  XOR U4 ( .A(n5), .B(n6), .Z(n4) );
  XNOR U5 ( .A(n7), .B(n1), .Z(n6) );
  AND U6 ( .A(n8), .B(n9), .Z(n7) );
  XOR U7 ( .A(n10), .B(n11), .Z(n5) );
  AND U8 ( .A(n12), .B(n13), .Z(n11) );
  NOR U9 ( .A(n14), .B(n15), .Z(n13) );
  NOR U10 ( .A(n16), .B(n17), .Z(n12) );
  AND U11 ( .A(n18), .B(n19), .Z(n17) );
  AND U12 ( .A(n20), .B(n21), .Z(n10) );
  NOR U13 ( .A(n22), .B(n23), .Z(n21) );
  AND U14 ( .A(n16), .B(n24), .Z(n23) );
  AND U15 ( .A(n14), .B(n25), .Z(n22) );
  NOR U16 ( .A(n26), .B(n27), .Z(n20) );
  AND U17 ( .A(n28), .B(n29), .Z(n27) );
  AND U18 ( .A(n30), .B(n31), .Z(n29) );
  NOR U19 ( .A(n32), .B(n33), .Z(n30) );
  NOR U20 ( .A(n34), .B(n35), .Z(n28) );
  AND U21 ( .A(n15), .B(n36), .Z(n26) );
  XOR U22 ( .A(n37), .B(n38), .Z(n3) );
  XOR U23 ( .A(n39), .B(n40), .Z(n38) );
  XOR U24 ( .A(n41), .B(n42), .Z(n40) );
  NOR U25 ( .A(n43), .B(n44), .Z(n42) );
  NOR U26 ( .A(n45), .B(n46), .Z(n41) );
  AND U27 ( .A(n47), .B(n48), .Z(n46) );
  IV U28 ( .A(n49), .Z(n45) );
  NOR U29 ( .A(n50), .B(n51), .Z(n49) );
  AND U30 ( .A(n43), .B(n52), .Z(n51) );
  AND U31 ( .A(n44), .B(n53), .Z(n50) );
  IV U32 ( .A(n54), .Z(n53) );
  AND U33 ( .A(n55), .B(n56), .Z(n39) );
  AND U34 ( .A(n57), .B(n58), .Z(n56) );
  NOR U35 ( .A(n59), .B(n60), .Z(n57) );
  NOR U36 ( .A(n61), .B(n62), .Z(n55) );
  XNOR U37 ( .A(n63), .B(n1), .Z(n37) );
  XNOR U38 ( .A(n64), .B(n65), .Z(n63) );
  AND U39 ( .A(n66), .B(n67), .Z(n65) );
  AND U40 ( .A(n68), .B(n69), .Z(n64) );
  XOR U41 ( .A(n70), .B(n71), .Z(n1) );
  AND U42 ( .A(n72), .B(n73), .Z(n71) );
  XOR U43 ( .A(n70), .B(n8), .Z(n73) );
  XOR U44 ( .A(n18), .B(n9), .Z(n8) );
  AND U45 ( .A(n74), .B(n75), .Z(n9) );
  XNOR U46 ( .A(n25), .B(n19), .Z(n18) );
  AND U47 ( .A(n76), .B(n77), .Z(n19) );
  XOR U48 ( .A(n24), .B(n14), .Z(n25) );
  AND U49 ( .A(n78), .B(n79), .Z(n14) );
  XOR U50 ( .A(n36), .B(n16), .Z(n24) );
  AND U51 ( .A(n80), .B(n81), .Z(n16) );
  XNOR U52 ( .A(n82), .B(n83), .Z(n36) );
  XOR U53 ( .A(n34), .B(n84), .Z(n83) );
  XNOR U54 ( .A(n32), .B(n31), .Z(n84) );
  IV U55 ( .A(n85), .Z(n31) );
  AND U56 ( .A(n86), .B(n87), .Z(n85) );
  AND U57 ( .A(n88), .B(n89), .Z(n32) );
  AND U58 ( .A(n90), .B(n91), .Z(n34) );
  XNOR U59 ( .A(n92), .B(n33), .Z(n82) );
  XOR U60 ( .A(n93), .B(n94), .Z(n33) );
  XOR U61 ( .A(n95), .B(n96), .Z(n94) );
  AND U62 ( .A(n97), .B(n98), .Z(n96) );
  XNOR U63 ( .A(n99), .B(n100), .Z(n93) );
  NOR U64 ( .A(n101), .B(n102), .Z(n100) );
  NOR U65 ( .A(n103), .B(n104), .Z(n102) );
  IV U66 ( .A(n105), .Z(n101) );
  NOR U67 ( .A(n95), .B(n106), .Z(n105) );
  AND U68 ( .A(n107), .B(n108), .Z(n106) );
  NOR U69 ( .A(n97), .B(n107), .Z(n99) );
  XNOR U70 ( .A(n35), .B(n15), .Z(n92) );
  AND U71 ( .A(n109), .B(n110), .Z(n15) );
  AND U72 ( .A(n111), .B(n112), .Z(n35) );
  XNOR U73 ( .A(n66), .B(n70), .Z(n72) );
  XOR U74 ( .A(n68), .B(n67), .Z(n66) );
  AND U75 ( .A(n113), .B(n114), .Z(n67) );
  XOR U76 ( .A(n54), .B(n69), .Z(n68) );
  AND U77 ( .A(n115), .B(n116), .Z(n69) );
  XNOR U78 ( .A(n52), .B(n44), .Z(n54) );
  AND U79 ( .A(n117), .B(n118), .Z(n44) );
  XNOR U80 ( .A(n47), .B(n43), .Z(n52) );
  AND U81 ( .A(n119), .B(n120), .Z(n43) );
  XOR U82 ( .A(n121), .B(n122), .Z(n47) );
  XOR U83 ( .A(n61), .B(n123), .Z(n122) );
  XNOR U84 ( .A(n59), .B(n58), .Z(n123) );
  IV U85 ( .A(n124), .Z(n58) );
  AND U86 ( .A(n125), .B(n126), .Z(n124) );
  AND U87 ( .A(n127), .B(n128), .Z(n59) );
  AND U88 ( .A(n129), .B(n130), .Z(n61) );
  XNOR U89 ( .A(n131), .B(n60), .Z(n121) );
  XOR U90 ( .A(n132), .B(n133), .Z(n60) );
  XOR U91 ( .A(n134), .B(n135), .Z(n133) );
  AND U92 ( .A(n136), .B(n137), .Z(n135) );
  XNOR U93 ( .A(n138), .B(n139), .Z(n132) );
  NOR U94 ( .A(n140), .B(n141), .Z(n139) );
  NOR U95 ( .A(n142), .B(n143), .Z(n141) );
  IV U96 ( .A(n144), .Z(n140) );
  NOR U97 ( .A(n134), .B(n145), .Z(n144) );
  AND U98 ( .A(n146), .B(n147), .Z(n145) );
  NOR U99 ( .A(n136), .B(n146), .Z(n138) );
  XNOR U100 ( .A(n62), .B(n48), .Z(n131) );
  AND U101 ( .A(n148), .B(n149), .Z(n48) );
  AND U102 ( .A(n150), .B(n151), .Z(n62) );
  XNOR U103 ( .A(n152), .B(n153), .Z(n70) );
  AND U104 ( .A(n154), .B(n155), .Z(n153) );
  XNOR U105 ( .A(n74), .B(n152), .Z(n155) );
  XOR U106 ( .A(n76), .B(n75), .Z(n74) );
  NOR U107 ( .A(n156), .B(n157), .Z(n75) );
  XOR U108 ( .A(n78), .B(n77), .Z(n76) );
  AND U109 ( .A(\dV[14][1] ), .B(n158), .Z(n77) );
  XOR U110 ( .A(n80), .B(n79), .Z(n78) );
  AND U111 ( .A(\dV[13][1] ), .B(n159), .Z(n79) );
  XOR U112 ( .A(n109), .B(n81), .Z(n80) );
  NOR U113 ( .A(n160), .B(n161), .Z(n81) );
  XOR U114 ( .A(n111), .B(n110), .Z(n109) );
  AND U115 ( .A(\dV[11][1] ), .B(n162), .Z(n110) );
  XOR U116 ( .A(n90), .B(n112), .Z(n111) );
  NOR U117 ( .A(n163), .B(n164), .Z(n112) );
  XOR U118 ( .A(n86), .B(n91), .Z(n90) );
  AND U119 ( .A(\dV[9][1] ), .B(n165), .Z(n91) );
  XOR U120 ( .A(n88), .B(n87), .Z(n86) );
  NOR U121 ( .A(n166), .B(n167), .Z(n87) );
  XNOR U122 ( .A(n98), .B(n89), .Z(n88) );
  AND U123 ( .A(\dV[7][1] ), .B(n168), .Z(n89) );
  XOR U124 ( .A(n108), .B(n97), .Z(n98) );
  NOR U125 ( .A(n169), .B(n170), .Z(n97) );
  XOR U126 ( .A(n171), .B(n103), .Z(n108) );
  XOR U127 ( .A(n104), .B(n172), .Z(n103) );
  NOR U128 ( .A(n173), .B(n174), .Z(n172) );
  XNOR U129 ( .A(n175), .B(n176), .Z(n104) );
  NOR U130 ( .A(n177), .B(n178), .Z(n176) );
  AND U131 ( .A(\dV[0][1] ), .B(\dV[1][1] ), .Z(n178) );
  AND U132 ( .A(\dV[2][1] ), .B(n179), .Z(n177) );
  XNOR U133 ( .A(n95), .B(n107), .Z(n171) );
  AND U134 ( .A(\dV[5][1] ), .B(n180), .Z(n107) );
  NOR U135 ( .A(n181), .B(n182), .Z(n95) );
  XOR U136 ( .A(n152), .B(n113), .Z(n154) );
  XOR U137 ( .A(n115), .B(n114), .Z(n113) );
  AND U138 ( .A(n183), .B(n156), .Z(n114) );
  IV U139 ( .A(\dV[15][1] ), .Z(n156) );
  XOR U140 ( .A(n117), .B(n116), .Z(n115) );
  NOR U141 ( .A(n184), .B(\dV[14][1] ), .Z(n116) );
  XOR U142 ( .A(n119), .B(n118), .Z(n117) );
  NOR U143 ( .A(n185), .B(\dV[13][1] ), .Z(n118) );
  XOR U144 ( .A(n148), .B(n120), .Z(n119) );
  NOR U145 ( .A(n186), .B(\dV[12][1] ), .Z(n120) );
  XOR U146 ( .A(n150), .B(n149), .Z(n148) );
  NOR U147 ( .A(n187), .B(\dV[11][1] ), .Z(n149) );
  XOR U148 ( .A(n129), .B(n151), .Z(n150) );
  NOR U149 ( .A(n188), .B(\dV[10][1] ), .Z(n151) );
  XOR U150 ( .A(n125), .B(n130), .Z(n129) );
  NOR U151 ( .A(n189), .B(\dV[9][1] ), .Z(n130) );
  XOR U152 ( .A(n127), .B(n126), .Z(n125) );
  NOR U153 ( .A(n190), .B(\dV[8][1] ), .Z(n126) );
  XNOR U154 ( .A(n137), .B(n128), .Z(n127) );
  NOR U155 ( .A(n191), .B(\dV[7][1] ), .Z(n128) );
  XOR U156 ( .A(n147), .B(n136), .Z(n137) );
  NOR U157 ( .A(n192), .B(\dV[6][1] ), .Z(n136) );
  XOR U158 ( .A(n193), .B(n142), .Z(n147) );
  XOR U159 ( .A(n143), .B(n194), .Z(n142) );
  AND U160 ( .A(n195), .B(n173), .Z(n194) );
  XNOR U161 ( .A(n175), .B(n196), .Z(n143) );
  NOR U162 ( .A(n197), .B(n198), .Z(n196) );
  NOR U163 ( .A(\dV[1][1] ), .B(\dV[0][1] ), .Z(n198) );
  NOR U164 ( .A(n175), .B(\dV[2][1] ), .Z(n197) );
  XNOR U165 ( .A(n134), .B(n146), .Z(n193) );
  NOR U166 ( .A(n199), .B(\dV[5][1] ), .Z(n146) );
  AND U167 ( .A(n200), .B(n181), .Z(n134) );
  AND U168 ( .A(n201), .B(n202), .Z(n152) );
  XNOR U169 ( .A(\dV[15][1] ), .B(n157), .Z(n202) );
  XNOR U170 ( .A(n158), .B(\dV[14][1] ), .Z(n157) );
  XOR U171 ( .A(n159), .B(\dV[13][1] ), .Z(n158) );
  XOR U172 ( .A(n161), .B(n160), .Z(n159) );
  IV U173 ( .A(\dV[12][1] ), .Z(n160) );
  XNOR U174 ( .A(n162), .B(\dV[11][1] ), .Z(n161) );
  XOR U175 ( .A(n164), .B(n163), .Z(n162) );
  IV U176 ( .A(\dV[10][1] ), .Z(n163) );
  XNOR U177 ( .A(n165), .B(\dV[9][1] ), .Z(n164) );
  XOR U178 ( .A(n167), .B(n166), .Z(n165) );
  IV U179 ( .A(\dV[8][1] ), .Z(n166) );
  XNOR U180 ( .A(n168), .B(\dV[7][1] ), .Z(n167) );
  XOR U181 ( .A(n170), .B(n169), .Z(n168) );
  IV U182 ( .A(\dV[6][1] ), .Z(n169) );
  XNOR U183 ( .A(n180), .B(\dV[5][1] ), .Z(n170) );
  XOR U184 ( .A(n182), .B(n181), .Z(n180) );
  IV U185 ( .A(\dV[4][1] ), .Z(n181) );
  XNOR U186 ( .A(n174), .B(n173), .Z(n182) );
  XNOR U187 ( .A(\dV[2][1] ), .B(n179), .Z(n174) );
  XOR U188 ( .A(\dV[0][1] ), .B(\dV[1][1] ), .Z(n179) );
  XOR U189 ( .A(n183), .B(\dV[15][1] ), .Z(n201) );
  XOR U190 ( .A(n184), .B(\dV[14][1] ), .Z(n183) );
  XNOR U191 ( .A(n185), .B(\dV[13][1] ), .Z(n184) );
  XNOR U192 ( .A(n186), .B(\dV[12][1] ), .Z(n185) );
  XNOR U193 ( .A(n187), .B(\dV[11][1] ), .Z(n186) );
  XNOR U194 ( .A(n188), .B(\dV[10][1] ), .Z(n187) );
  XNOR U195 ( .A(n189), .B(\dV[9][1] ), .Z(n188) );
  XNOR U196 ( .A(n190), .B(\dV[8][1] ), .Z(n189) );
  XNOR U197 ( .A(n191), .B(\dV[7][1] ), .Z(n190) );
  XNOR U198 ( .A(n192), .B(\dV[6][1] ), .Z(n191) );
  XNOR U199 ( .A(n199), .B(\dV[5][1] ), .Z(n192) );
  XOR U200 ( .A(n200), .B(\dV[4][1] ), .Z(n199) );
  XNOR U201 ( .A(n203), .B(n173), .Z(n200) );
  IV U202 ( .A(\dV[3][1] ), .Z(n173) );
  IV U203 ( .A(n195), .Z(n203) );
  XOR U204 ( .A(\dV[2][1] ), .B(n175), .Z(n195) );
  XOR U205 ( .A(\dV[0][1] ), .B(n204), .Z(n175) );
  IV U206 ( .A(\dV[1][1] ), .Z(n204) );
endmodule

