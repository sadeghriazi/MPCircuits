
module knn_comb_BMR_W16_K3_N16 ( p_input, o );
  input [271:0] p_input;
  output [47:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][15] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427;
  assign \knn_comb_/min_val_out[0][0]  = p_input[240];
  assign \knn_comb_/min_val_out[0][1]  = p_input[241];
  assign \knn_comb_/min_val_out[0][2]  = p_input[242];
  assign \knn_comb_/min_val_out[0][3]  = p_input[243];
  assign \knn_comb_/min_val_out[0][4]  = p_input[244];
  assign \knn_comb_/min_val_out[0][5]  = p_input[245];
  assign \knn_comb_/min_val_out[0][6]  = p_input[246];
  assign \knn_comb_/min_val_out[0][7]  = p_input[247];
  assign \knn_comb_/min_val_out[0][8]  = p_input[248];
  assign \knn_comb_/min_val_out[0][9]  = p_input[249];
  assign \knn_comb_/min_val_out[0][10]  = p_input[250];
  assign \knn_comb_/min_val_out[0][11]  = p_input[251];
  assign \knn_comb_/min_val_out[0][12]  = p_input[252];
  assign \knn_comb_/min_val_out[0][13]  = p_input[253];
  assign \knn_comb_/min_val_out[0][14]  = p_input[254];
  assign \knn_comb_/min_val_out[0][15]  = p_input[255];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][0]  = p_input[208];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][1]  = p_input[209];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][2]  = p_input[210];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][3]  = p_input[211];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][4]  = p_input[212];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][5]  = p_input[213];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][6]  = p_input[214];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][7]  = p_input[215];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][8]  = p_input[216];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][9]  = p_input[217];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][10]  = p_input[218];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][11]  = p_input[219];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][12]  = p_input[220];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][13]  = p_input[221];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][14]  = p_input[222];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][15]  = p_input[223];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][0]  = p_input[224];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][1]  = p_input[225];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][2]  = p_input[226];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][3]  = p_input[227];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][4]  = p_input[228];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][5]  = p_input[229];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][6]  = p_input[230];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][7]  = p_input[231];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][8]  = p_input[232];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][9]  = p_input[233];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][10]  = p_input[234];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][11]  = p_input[235];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][12]  = p_input[236];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][13]  = p_input[237];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][14]  = p_input[238];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][15]  = p_input[239];

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  XOR U2 ( .A(n3), .B(n4), .Z(o[8]) );
  XOR U3 ( .A(n5), .B(n6), .Z(o[7]) );
  XOR U4 ( .A(n7), .B(n8), .Z(o[6]) );
  XOR U5 ( .A(n9), .B(n10), .Z(o[5]) );
  XOR U6 ( .A(n11), .B(n12), .Z(o[4]) );
  XOR U7 ( .A(n13), .B(n14), .Z(o[47]) );
  XOR U8 ( .A(n15), .B(n16), .Z(o[46]) );
  XOR U9 ( .A(n17), .B(n18), .Z(o[45]) );
  XOR U10 ( .A(n19), .B(n20), .Z(o[44]) );
  XOR U11 ( .A(n21), .B(n22), .Z(o[43]) );
  XOR U12 ( .A(n23), .B(n24), .Z(o[42]) );
  XOR U13 ( .A(n25), .B(n26), .Z(o[41]) );
  XOR U14 ( .A(n27), .B(n28), .Z(o[40]) );
  XOR U15 ( .A(n29), .B(n30), .Z(o[3]) );
  XOR U16 ( .A(n31), .B(n32), .Z(o[39]) );
  XOR U17 ( .A(n33), .B(n34), .Z(o[38]) );
  XOR U18 ( .A(n35), .B(n36), .Z(o[37]) );
  XOR U19 ( .A(n37), .B(n38), .Z(o[36]) );
  XOR U20 ( .A(n39), .B(n40), .Z(o[35]) );
  XOR U21 ( .A(n41), .B(n42), .Z(o[34]) );
  XOR U22 ( .A(n43), .B(n44), .Z(o[33]) );
  XOR U23 ( .A(n45), .B(n46), .Z(o[32]) );
  XOR U24 ( .A(n47), .B(n48), .Z(o[31]) );
  XOR U25 ( .A(n49), .B(n50), .Z(o[30]) );
  XOR U26 ( .A(n51), .B(n52), .Z(o[2]) );
  XOR U27 ( .A(n53), .B(n54), .Z(o[29]) );
  XOR U28 ( .A(n55), .B(n56), .Z(o[28]) );
  XOR U29 ( .A(n57), .B(n58), .Z(o[27]) );
  XOR U30 ( .A(n59), .B(n60), .Z(o[26]) );
  XOR U31 ( .A(n1), .B(n61), .Z(o[25]) );
  AND U32 ( .A(n62), .B(n63), .Z(n1) );
  XOR U33 ( .A(n2), .B(n61), .Z(n63) );
  XOR U34 ( .A(n64), .B(n25), .Z(n61) );
  AND U35 ( .A(n65), .B(n66), .Z(n25) );
  XNOR U36 ( .A(n67), .B(n26), .Z(n66) );
  XOR U37 ( .A(n68), .B(n69), .Z(n26) );
  AND U38 ( .A(n70), .B(n71), .Z(n69) );
  XOR U39 ( .A(p_input[9]), .B(n68), .Z(n71) );
  XOR U40 ( .A(n72), .B(n73), .Z(n68) );
  AND U41 ( .A(n74), .B(n75), .Z(n73) );
  IV U42 ( .A(n64), .Z(n67) );
  XOR U43 ( .A(n76), .B(n77), .Z(n64) );
  AND U44 ( .A(n78), .B(n79), .Z(n77) );
  XOR U45 ( .A(n80), .B(n81), .Z(n2) );
  AND U46 ( .A(n82), .B(n79), .Z(n81) );
  XNOR U47 ( .A(n83), .B(n76), .Z(n79) );
  XOR U48 ( .A(n84), .B(n85), .Z(n76) );
  AND U49 ( .A(n86), .B(n75), .Z(n85) );
  XNOR U50 ( .A(n87), .B(n72), .Z(n75) );
  XOR U51 ( .A(n88), .B(n89), .Z(n72) );
  AND U52 ( .A(n90), .B(n91), .Z(n89) );
  XOR U53 ( .A(p_input[25]), .B(n88), .Z(n91) );
  XOR U54 ( .A(n92), .B(n93), .Z(n88) );
  AND U55 ( .A(n94), .B(n95), .Z(n93) );
  IV U56 ( .A(n84), .Z(n87) );
  XOR U57 ( .A(n96), .B(n97), .Z(n84) );
  AND U58 ( .A(n98), .B(n99), .Z(n97) );
  IV U59 ( .A(n80), .Z(n83) );
  XNOR U60 ( .A(n100), .B(n101), .Z(n80) );
  AND U61 ( .A(n102), .B(n99), .Z(n101) );
  XNOR U62 ( .A(n100), .B(n96), .Z(n99) );
  XOR U63 ( .A(n103), .B(n104), .Z(n96) );
  AND U64 ( .A(n105), .B(n95), .Z(n104) );
  XNOR U65 ( .A(n106), .B(n92), .Z(n95) );
  XOR U66 ( .A(n107), .B(n108), .Z(n92) );
  AND U67 ( .A(n109), .B(n110), .Z(n108) );
  XOR U68 ( .A(p_input[41]), .B(n107), .Z(n110) );
  XOR U69 ( .A(n111), .B(n112), .Z(n107) );
  AND U70 ( .A(n113), .B(n114), .Z(n112) );
  IV U71 ( .A(n103), .Z(n106) );
  XOR U72 ( .A(n115), .B(n116), .Z(n103) );
  AND U73 ( .A(n117), .B(n118), .Z(n116) );
  XOR U74 ( .A(n119), .B(n120), .Z(n100) );
  AND U75 ( .A(n121), .B(n118), .Z(n120) );
  XNOR U76 ( .A(n119), .B(n115), .Z(n118) );
  XOR U77 ( .A(n122), .B(n123), .Z(n115) );
  AND U78 ( .A(n124), .B(n114), .Z(n123) );
  XNOR U79 ( .A(n125), .B(n111), .Z(n114) );
  XOR U80 ( .A(n126), .B(n127), .Z(n111) );
  AND U81 ( .A(n128), .B(n129), .Z(n127) );
  XOR U82 ( .A(p_input[57]), .B(n126), .Z(n129) );
  XOR U83 ( .A(n130), .B(n131), .Z(n126) );
  AND U84 ( .A(n132), .B(n133), .Z(n131) );
  IV U85 ( .A(n122), .Z(n125) );
  XOR U86 ( .A(n134), .B(n135), .Z(n122) );
  AND U87 ( .A(n136), .B(n137), .Z(n135) );
  XOR U88 ( .A(n138), .B(n139), .Z(n119) );
  AND U89 ( .A(n140), .B(n137), .Z(n139) );
  XNOR U90 ( .A(n138), .B(n134), .Z(n137) );
  XOR U91 ( .A(n141), .B(n142), .Z(n134) );
  AND U92 ( .A(n143), .B(n133), .Z(n142) );
  XNOR U93 ( .A(n144), .B(n130), .Z(n133) );
  XOR U94 ( .A(n145), .B(n146), .Z(n130) );
  AND U95 ( .A(n147), .B(n148), .Z(n146) );
  XOR U96 ( .A(p_input[73]), .B(n145), .Z(n148) );
  XOR U97 ( .A(n149), .B(n150), .Z(n145) );
  AND U98 ( .A(n151), .B(n152), .Z(n150) );
  IV U99 ( .A(n141), .Z(n144) );
  XOR U100 ( .A(n153), .B(n154), .Z(n141) );
  AND U101 ( .A(n155), .B(n156), .Z(n154) );
  XOR U102 ( .A(n157), .B(n158), .Z(n138) );
  AND U103 ( .A(n159), .B(n156), .Z(n158) );
  XNOR U104 ( .A(n157), .B(n153), .Z(n156) );
  XOR U105 ( .A(n160), .B(n161), .Z(n153) );
  AND U106 ( .A(n162), .B(n152), .Z(n161) );
  XNOR U107 ( .A(n163), .B(n149), .Z(n152) );
  XOR U108 ( .A(n164), .B(n165), .Z(n149) );
  AND U109 ( .A(n166), .B(n167), .Z(n165) );
  XOR U110 ( .A(p_input[89]), .B(n164), .Z(n167) );
  XOR U111 ( .A(n168), .B(n169), .Z(n164) );
  AND U112 ( .A(n170), .B(n171), .Z(n169) );
  IV U113 ( .A(n160), .Z(n163) );
  XOR U114 ( .A(n172), .B(n173), .Z(n160) );
  AND U115 ( .A(n174), .B(n175), .Z(n173) );
  XOR U116 ( .A(n176), .B(n177), .Z(n157) );
  AND U117 ( .A(n178), .B(n175), .Z(n177) );
  XNOR U118 ( .A(n176), .B(n172), .Z(n175) );
  XOR U119 ( .A(n179), .B(n180), .Z(n172) );
  AND U120 ( .A(n181), .B(n171), .Z(n180) );
  XNOR U121 ( .A(n182), .B(n168), .Z(n171) );
  XOR U122 ( .A(n183), .B(n184), .Z(n168) );
  AND U123 ( .A(n185), .B(n186), .Z(n184) );
  XOR U124 ( .A(p_input[105]), .B(n183), .Z(n186) );
  XOR U125 ( .A(n187), .B(n188), .Z(n183) );
  AND U126 ( .A(n189), .B(n190), .Z(n188) );
  IV U127 ( .A(n179), .Z(n182) );
  XOR U128 ( .A(n191), .B(n192), .Z(n179) );
  AND U129 ( .A(n193), .B(n194), .Z(n192) );
  XOR U130 ( .A(n195), .B(n196), .Z(n176) );
  AND U131 ( .A(n197), .B(n194), .Z(n196) );
  XNOR U132 ( .A(n195), .B(n191), .Z(n194) );
  XOR U133 ( .A(n198), .B(n199), .Z(n191) );
  AND U134 ( .A(n200), .B(n190), .Z(n199) );
  XNOR U135 ( .A(n201), .B(n187), .Z(n190) );
  XOR U136 ( .A(n202), .B(n203), .Z(n187) );
  AND U137 ( .A(n204), .B(n205), .Z(n203) );
  XOR U138 ( .A(p_input[121]), .B(n202), .Z(n205) );
  XOR U139 ( .A(n206), .B(n207), .Z(n202) );
  AND U140 ( .A(n208), .B(n209), .Z(n207) );
  IV U141 ( .A(n198), .Z(n201) );
  XOR U142 ( .A(n210), .B(n211), .Z(n198) );
  AND U143 ( .A(n212), .B(n213), .Z(n211) );
  XOR U144 ( .A(n214), .B(n215), .Z(n195) );
  AND U145 ( .A(n216), .B(n213), .Z(n215) );
  XNOR U146 ( .A(n214), .B(n210), .Z(n213) );
  XOR U147 ( .A(n217), .B(n218), .Z(n210) );
  AND U148 ( .A(n219), .B(n209), .Z(n218) );
  XNOR U149 ( .A(n220), .B(n206), .Z(n209) );
  XOR U150 ( .A(n221), .B(n222), .Z(n206) );
  AND U151 ( .A(n223), .B(n224), .Z(n222) );
  XOR U152 ( .A(p_input[137]), .B(n221), .Z(n224) );
  XOR U153 ( .A(n225), .B(n226), .Z(n221) );
  AND U154 ( .A(n227), .B(n228), .Z(n226) );
  IV U155 ( .A(n217), .Z(n220) );
  XOR U156 ( .A(n229), .B(n230), .Z(n217) );
  AND U157 ( .A(n231), .B(n232), .Z(n230) );
  XOR U158 ( .A(n233), .B(n234), .Z(n214) );
  AND U159 ( .A(n235), .B(n232), .Z(n234) );
  XNOR U160 ( .A(n233), .B(n229), .Z(n232) );
  XOR U161 ( .A(n236), .B(n237), .Z(n229) );
  AND U162 ( .A(n238), .B(n228), .Z(n237) );
  XNOR U163 ( .A(n239), .B(n225), .Z(n228) );
  XOR U164 ( .A(n240), .B(n241), .Z(n225) );
  AND U165 ( .A(n242), .B(n243), .Z(n241) );
  XOR U166 ( .A(p_input[153]), .B(n240), .Z(n243) );
  XOR U167 ( .A(n244), .B(n245), .Z(n240) );
  AND U168 ( .A(n246), .B(n247), .Z(n245) );
  IV U169 ( .A(n236), .Z(n239) );
  XOR U170 ( .A(n248), .B(n249), .Z(n236) );
  AND U171 ( .A(n250), .B(n251), .Z(n249) );
  XOR U172 ( .A(n252), .B(n253), .Z(n233) );
  AND U173 ( .A(n254), .B(n251), .Z(n253) );
  XNOR U174 ( .A(n252), .B(n248), .Z(n251) );
  XOR U175 ( .A(n255), .B(n256), .Z(n248) );
  AND U176 ( .A(n257), .B(n247), .Z(n256) );
  XNOR U177 ( .A(n258), .B(n244), .Z(n247) );
  XOR U178 ( .A(n259), .B(n260), .Z(n244) );
  AND U179 ( .A(n261), .B(n262), .Z(n260) );
  XOR U180 ( .A(p_input[169]), .B(n259), .Z(n262) );
  XOR U181 ( .A(n263), .B(n264), .Z(n259) );
  AND U182 ( .A(n265), .B(n266), .Z(n264) );
  IV U183 ( .A(n255), .Z(n258) );
  XOR U184 ( .A(n267), .B(n268), .Z(n255) );
  AND U185 ( .A(n269), .B(n270), .Z(n268) );
  XOR U186 ( .A(n271), .B(n272), .Z(n252) );
  AND U187 ( .A(n273), .B(n270), .Z(n272) );
  XNOR U188 ( .A(n271), .B(n267), .Z(n270) );
  XOR U189 ( .A(n274), .B(n275), .Z(n267) );
  AND U190 ( .A(n276), .B(n266), .Z(n275) );
  XNOR U191 ( .A(n277), .B(n263), .Z(n266) );
  XOR U192 ( .A(n278), .B(n279), .Z(n263) );
  AND U193 ( .A(n280), .B(n281), .Z(n279) );
  XOR U194 ( .A(p_input[185]), .B(n278), .Z(n281) );
  XOR U195 ( .A(n282), .B(n283), .Z(n278) );
  AND U196 ( .A(n284), .B(n285), .Z(n283) );
  IV U197 ( .A(n274), .Z(n277) );
  XOR U198 ( .A(n286), .B(n287), .Z(n274) );
  AND U199 ( .A(n288), .B(n289), .Z(n287) );
  XOR U200 ( .A(n290), .B(n291), .Z(n271) );
  AND U201 ( .A(n292), .B(n289), .Z(n291) );
  XNOR U202 ( .A(n290), .B(n286), .Z(n289) );
  XOR U203 ( .A(n293), .B(n294), .Z(n286) );
  AND U204 ( .A(n295), .B(n285), .Z(n294) );
  XNOR U205 ( .A(n296), .B(n282), .Z(n285) );
  XOR U206 ( .A(n297), .B(n298), .Z(n282) );
  AND U207 ( .A(n299), .B(n300), .Z(n298) );
  XOR U208 ( .A(p_input[201]), .B(n297), .Z(n300) );
  XOR U209 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n301), .Z(
        n297) );
  AND U210 ( .A(n302), .B(n303), .Z(n301) );
  IV U211 ( .A(n293), .Z(n296) );
  XOR U212 ( .A(n304), .B(n305), .Z(n293) );
  AND U213 ( .A(n306), .B(n307), .Z(n305) );
  XOR U214 ( .A(n308), .B(n309), .Z(n290) );
  AND U215 ( .A(n310), .B(n307), .Z(n309) );
  XNOR U216 ( .A(n308), .B(n304), .Z(n307) );
  XNOR U217 ( .A(n311), .B(n312), .Z(n304) );
  AND U218 ( .A(n313), .B(n303), .Z(n312) );
  XNOR U219 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n311), .Z(
        n303) );
  XNOR U220 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .B(n314), .Z(
        n311) );
  AND U221 ( .A(n315), .B(n316), .Z(n314) );
  XNOR U222 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n317), .Z(n308) );
  AND U223 ( .A(n318), .B(n316), .Z(n317) );
  XOR U224 ( .A(n319), .B(n320), .Z(n316) );
  XOR U225 ( .A(n3), .B(n321), .Z(o[24]) );
  AND U226 ( .A(n62), .B(n322), .Z(n3) );
  XOR U227 ( .A(n4), .B(n321), .Z(n322) );
  XOR U228 ( .A(n323), .B(n27), .Z(n321) );
  AND U229 ( .A(n65), .B(n324), .Z(n27) );
  XNOR U230 ( .A(n325), .B(n28), .Z(n324) );
  XOR U231 ( .A(n326), .B(n327), .Z(n28) );
  AND U232 ( .A(n70), .B(n328), .Z(n327) );
  XOR U233 ( .A(p_input[8]), .B(n326), .Z(n328) );
  XOR U234 ( .A(n329), .B(n330), .Z(n326) );
  AND U235 ( .A(n74), .B(n331), .Z(n330) );
  IV U236 ( .A(n323), .Z(n325) );
  XOR U237 ( .A(n332), .B(n333), .Z(n323) );
  AND U238 ( .A(n78), .B(n334), .Z(n333) );
  XOR U239 ( .A(n335), .B(n336), .Z(n4) );
  AND U240 ( .A(n82), .B(n334), .Z(n336) );
  XNOR U241 ( .A(n337), .B(n332), .Z(n334) );
  XOR U242 ( .A(n338), .B(n339), .Z(n332) );
  AND U243 ( .A(n86), .B(n331), .Z(n339) );
  XNOR U244 ( .A(n340), .B(n329), .Z(n331) );
  XOR U245 ( .A(n341), .B(n342), .Z(n329) );
  AND U246 ( .A(n90), .B(n343), .Z(n342) );
  XOR U247 ( .A(p_input[24]), .B(n341), .Z(n343) );
  XOR U248 ( .A(n344), .B(n345), .Z(n341) );
  AND U249 ( .A(n94), .B(n346), .Z(n345) );
  IV U250 ( .A(n338), .Z(n340) );
  XOR U251 ( .A(n347), .B(n348), .Z(n338) );
  AND U252 ( .A(n98), .B(n349), .Z(n348) );
  IV U253 ( .A(n335), .Z(n337) );
  XNOR U254 ( .A(n350), .B(n351), .Z(n335) );
  AND U255 ( .A(n102), .B(n349), .Z(n351) );
  XNOR U256 ( .A(n350), .B(n347), .Z(n349) );
  XOR U257 ( .A(n352), .B(n353), .Z(n347) );
  AND U258 ( .A(n105), .B(n346), .Z(n353) );
  XNOR U259 ( .A(n354), .B(n344), .Z(n346) );
  XOR U260 ( .A(n355), .B(n356), .Z(n344) );
  AND U261 ( .A(n109), .B(n357), .Z(n356) );
  XOR U262 ( .A(p_input[40]), .B(n355), .Z(n357) );
  XOR U263 ( .A(n358), .B(n359), .Z(n355) );
  AND U264 ( .A(n113), .B(n360), .Z(n359) );
  IV U265 ( .A(n352), .Z(n354) );
  XOR U266 ( .A(n361), .B(n362), .Z(n352) );
  AND U267 ( .A(n117), .B(n363), .Z(n362) );
  XOR U268 ( .A(n364), .B(n365), .Z(n350) );
  AND U269 ( .A(n121), .B(n363), .Z(n365) );
  XNOR U270 ( .A(n364), .B(n361), .Z(n363) );
  XOR U271 ( .A(n366), .B(n367), .Z(n361) );
  AND U272 ( .A(n124), .B(n360), .Z(n367) );
  XNOR U273 ( .A(n368), .B(n358), .Z(n360) );
  XOR U274 ( .A(n369), .B(n370), .Z(n358) );
  AND U275 ( .A(n128), .B(n371), .Z(n370) );
  XOR U276 ( .A(p_input[56]), .B(n369), .Z(n371) );
  XOR U277 ( .A(n372), .B(n373), .Z(n369) );
  AND U278 ( .A(n132), .B(n374), .Z(n373) );
  IV U279 ( .A(n366), .Z(n368) );
  XOR U280 ( .A(n375), .B(n376), .Z(n366) );
  AND U281 ( .A(n136), .B(n377), .Z(n376) );
  XOR U282 ( .A(n378), .B(n379), .Z(n364) );
  AND U283 ( .A(n140), .B(n377), .Z(n379) );
  XNOR U284 ( .A(n378), .B(n375), .Z(n377) );
  XOR U285 ( .A(n380), .B(n381), .Z(n375) );
  AND U286 ( .A(n143), .B(n374), .Z(n381) );
  XNOR U287 ( .A(n382), .B(n372), .Z(n374) );
  XOR U288 ( .A(n383), .B(n384), .Z(n372) );
  AND U289 ( .A(n147), .B(n385), .Z(n384) );
  XOR U290 ( .A(p_input[72]), .B(n383), .Z(n385) );
  XOR U291 ( .A(n386), .B(n387), .Z(n383) );
  AND U292 ( .A(n151), .B(n388), .Z(n387) );
  IV U293 ( .A(n380), .Z(n382) );
  XOR U294 ( .A(n389), .B(n390), .Z(n380) );
  AND U295 ( .A(n155), .B(n391), .Z(n390) );
  XOR U296 ( .A(n392), .B(n393), .Z(n378) );
  AND U297 ( .A(n159), .B(n391), .Z(n393) );
  XNOR U298 ( .A(n392), .B(n389), .Z(n391) );
  XOR U299 ( .A(n394), .B(n395), .Z(n389) );
  AND U300 ( .A(n162), .B(n388), .Z(n395) );
  XNOR U301 ( .A(n396), .B(n386), .Z(n388) );
  XOR U302 ( .A(n397), .B(n398), .Z(n386) );
  AND U303 ( .A(n166), .B(n399), .Z(n398) );
  XOR U304 ( .A(p_input[88]), .B(n397), .Z(n399) );
  XOR U305 ( .A(n400), .B(n401), .Z(n397) );
  AND U306 ( .A(n170), .B(n402), .Z(n401) );
  IV U307 ( .A(n394), .Z(n396) );
  XOR U308 ( .A(n403), .B(n404), .Z(n394) );
  AND U309 ( .A(n174), .B(n405), .Z(n404) );
  XOR U310 ( .A(n406), .B(n407), .Z(n392) );
  AND U311 ( .A(n178), .B(n405), .Z(n407) );
  XNOR U312 ( .A(n406), .B(n403), .Z(n405) );
  XOR U313 ( .A(n408), .B(n409), .Z(n403) );
  AND U314 ( .A(n181), .B(n402), .Z(n409) );
  XNOR U315 ( .A(n410), .B(n400), .Z(n402) );
  XOR U316 ( .A(n411), .B(n412), .Z(n400) );
  AND U317 ( .A(n185), .B(n413), .Z(n412) );
  XOR U318 ( .A(p_input[104]), .B(n411), .Z(n413) );
  XOR U319 ( .A(n414), .B(n415), .Z(n411) );
  AND U320 ( .A(n189), .B(n416), .Z(n415) );
  IV U321 ( .A(n408), .Z(n410) );
  XOR U322 ( .A(n417), .B(n418), .Z(n408) );
  AND U323 ( .A(n193), .B(n419), .Z(n418) );
  XOR U324 ( .A(n420), .B(n421), .Z(n406) );
  AND U325 ( .A(n197), .B(n419), .Z(n421) );
  XNOR U326 ( .A(n420), .B(n417), .Z(n419) );
  XOR U327 ( .A(n422), .B(n423), .Z(n417) );
  AND U328 ( .A(n200), .B(n416), .Z(n423) );
  XNOR U329 ( .A(n424), .B(n414), .Z(n416) );
  XOR U330 ( .A(n425), .B(n426), .Z(n414) );
  AND U331 ( .A(n204), .B(n427), .Z(n426) );
  XOR U332 ( .A(p_input[120]), .B(n425), .Z(n427) );
  XOR U333 ( .A(n428), .B(n429), .Z(n425) );
  AND U334 ( .A(n208), .B(n430), .Z(n429) );
  IV U335 ( .A(n422), .Z(n424) );
  XOR U336 ( .A(n431), .B(n432), .Z(n422) );
  AND U337 ( .A(n212), .B(n433), .Z(n432) );
  XOR U338 ( .A(n434), .B(n435), .Z(n420) );
  AND U339 ( .A(n216), .B(n433), .Z(n435) );
  XNOR U340 ( .A(n434), .B(n431), .Z(n433) );
  XOR U341 ( .A(n436), .B(n437), .Z(n431) );
  AND U342 ( .A(n219), .B(n430), .Z(n437) );
  XNOR U343 ( .A(n438), .B(n428), .Z(n430) );
  XOR U344 ( .A(n439), .B(n440), .Z(n428) );
  AND U345 ( .A(n223), .B(n441), .Z(n440) );
  XOR U346 ( .A(p_input[136]), .B(n439), .Z(n441) );
  XOR U347 ( .A(n442), .B(n443), .Z(n439) );
  AND U348 ( .A(n227), .B(n444), .Z(n443) );
  IV U349 ( .A(n436), .Z(n438) );
  XOR U350 ( .A(n445), .B(n446), .Z(n436) );
  AND U351 ( .A(n231), .B(n447), .Z(n446) );
  XOR U352 ( .A(n448), .B(n449), .Z(n434) );
  AND U353 ( .A(n235), .B(n447), .Z(n449) );
  XNOR U354 ( .A(n448), .B(n445), .Z(n447) );
  XOR U355 ( .A(n450), .B(n451), .Z(n445) );
  AND U356 ( .A(n238), .B(n444), .Z(n451) );
  XNOR U357 ( .A(n452), .B(n442), .Z(n444) );
  XOR U358 ( .A(n453), .B(n454), .Z(n442) );
  AND U359 ( .A(n242), .B(n455), .Z(n454) );
  XOR U360 ( .A(p_input[152]), .B(n453), .Z(n455) );
  XOR U361 ( .A(n456), .B(n457), .Z(n453) );
  AND U362 ( .A(n246), .B(n458), .Z(n457) );
  IV U363 ( .A(n450), .Z(n452) );
  XOR U364 ( .A(n459), .B(n460), .Z(n450) );
  AND U365 ( .A(n250), .B(n461), .Z(n460) );
  XOR U366 ( .A(n462), .B(n463), .Z(n448) );
  AND U367 ( .A(n254), .B(n461), .Z(n463) );
  XNOR U368 ( .A(n462), .B(n459), .Z(n461) );
  XOR U369 ( .A(n464), .B(n465), .Z(n459) );
  AND U370 ( .A(n257), .B(n458), .Z(n465) );
  XNOR U371 ( .A(n466), .B(n456), .Z(n458) );
  XOR U372 ( .A(n467), .B(n468), .Z(n456) );
  AND U373 ( .A(n261), .B(n469), .Z(n468) );
  XOR U374 ( .A(p_input[168]), .B(n467), .Z(n469) );
  XOR U375 ( .A(n470), .B(n471), .Z(n467) );
  AND U376 ( .A(n265), .B(n472), .Z(n471) );
  IV U377 ( .A(n464), .Z(n466) );
  XOR U378 ( .A(n473), .B(n474), .Z(n464) );
  AND U379 ( .A(n269), .B(n475), .Z(n474) );
  XOR U380 ( .A(n476), .B(n477), .Z(n462) );
  AND U381 ( .A(n273), .B(n475), .Z(n477) );
  XNOR U382 ( .A(n476), .B(n473), .Z(n475) );
  XOR U383 ( .A(n478), .B(n479), .Z(n473) );
  AND U384 ( .A(n276), .B(n472), .Z(n479) );
  XNOR U385 ( .A(n480), .B(n470), .Z(n472) );
  XOR U386 ( .A(n481), .B(n482), .Z(n470) );
  AND U387 ( .A(n280), .B(n483), .Z(n482) );
  XOR U388 ( .A(p_input[184]), .B(n481), .Z(n483) );
  XOR U389 ( .A(n484), .B(n485), .Z(n481) );
  AND U390 ( .A(n284), .B(n486), .Z(n485) );
  IV U391 ( .A(n478), .Z(n480) );
  XOR U392 ( .A(n487), .B(n488), .Z(n478) );
  AND U393 ( .A(n288), .B(n489), .Z(n488) );
  XOR U394 ( .A(n490), .B(n491), .Z(n476) );
  AND U395 ( .A(n292), .B(n489), .Z(n491) );
  XNOR U396 ( .A(n490), .B(n487), .Z(n489) );
  XOR U397 ( .A(n492), .B(n493), .Z(n487) );
  AND U398 ( .A(n295), .B(n486), .Z(n493) );
  XNOR U399 ( .A(n494), .B(n484), .Z(n486) );
  XOR U400 ( .A(n495), .B(n496), .Z(n484) );
  AND U401 ( .A(n299), .B(n497), .Z(n496) );
  XOR U402 ( .A(p_input[200]), .B(n495), .Z(n497) );
  XOR U403 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n498), .Z(
        n495) );
  AND U404 ( .A(n302), .B(n499), .Z(n498) );
  IV U405 ( .A(n492), .Z(n494) );
  XOR U406 ( .A(n500), .B(n501), .Z(n492) );
  AND U407 ( .A(n306), .B(n502), .Z(n501) );
  XOR U408 ( .A(n503), .B(n504), .Z(n490) );
  AND U409 ( .A(n310), .B(n502), .Z(n504) );
  XNOR U410 ( .A(n503), .B(n500), .Z(n502) );
  XNOR U411 ( .A(n505), .B(n506), .Z(n500) );
  AND U412 ( .A(n313), .B(n499), .Z(n506) );
  XNOR U413 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n505), .Z(
        n499) );
  XNOR U414 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(n507), .Z(
        n505) );
  AND U415 ( .A(n315), .B(n508), .Z(n507) );
  XNOR U416 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n509), .Z(n503) );
  AND U417 ( .A(n318), .B(n508), .Z(n509) );
  XOR U418 ( .A(n510), .B(n511), .Z(n508) );
  XOR U419 ( .A(n5), .B(n512), .Z(o[23]) );
  AND U420 ( .A(n62), .B(n513), .Z(n5) );
  XOR U421 ( .A(n6), .B(n512), .Z(n513) );
  XOR U422 ( .A(n514), .B(n31), .Z(n512) );
  AND U423 ( .A(n65), .B(n515), .Z(n31) );
  XNOR U424 ( .A(n516), .B(n32), .Z(n515) );
  XOR U425 ( .A(n517), .B(n518), .Z(n32) );
  AND U426 ( .A(n70), .B(n519), .Z(n518) );
  XOR U427 ( .A(p_input[7]), .B(n517), .Z(n519) );
  XOR U428 ( .A(n520), .B(n521), .Z(n517) );
  AND U429 ( .A(n74), .B(n522), .Z(n521) );
  IV U430 ( .A(n514), .Z(n516) );
  XOR U431 ( .A(n523), .B(n524), .Z(n514) );
  AND U432 ( .A(n78), .B(n525), .Z(n524) );
  XOR U433 ( .A(n526), .B(n527), .Z(n6) );
  AND U434 ( .A(n82), .B(n525), .Z(n527) );
  XNOR U435 ( .A(n528), .B(n523), .Z(n525) );
  XOR U436 ( .A(n529), .B(n530), .Z(n523) );
  AND U437 ( .A(n86), .B(n522), .Z(n530) );
  XNOR U438 ( .A(n531), .B(n520), .Z(n522) );
  XOR U439 ( .A(n532), .B(n533), .Z(n520) );
  AND U440 ( .A(n90), .B(n534), .Z(n533) );
  XOR U441 ( .A(p_input[23]), .B(n532), .Z(n534) );
  XOR U442 ( .A(n535), .B(n536), .Z(n532) );
  AND U443 ( .A(n94), .B(n537), .Z(n536) );
  IV U444 ( .A(n529), .Z(n531) );
  XOR U445 ( .A(n538), .B(n539), .Z(n529) );
  AND U446 ( .A(n98), .B(n540), .Z(n539) );
  IV U447 ( .A(n526), .Z(n528) );
  XNOR U448 ( .A(n541), .B(n542), .Z(n526) );
  AND U449 ( .A(n102), .B(n540), .Z(n542) );
  XNOR U450 ( .A(n541), .B(n538), .Z(n540) );
  XOR U451 ( .A(n543), .B(n544), .Z(n538) );
  AND U452 ( .A(n105), .B(n537), .Z(n544) );
  XNOR U453 ( .A(n545), .B(n535), .Z(n537) );
  XOR U454 ( .A(n546), .B(n547), .Z(n535) );
  AND U455 ( .A(n109), .B(n548), .Z(n547) );
  XOR U456 ( .A(p_input[39]), .B(n546), .Z(n548) );
  XOR U457 ( .A(n549), .B(n550), .Z(n546) );
  AND U458 ( .A(n113), .B(n551), .Z(n550) );
  IV U459 ( .A(n543), .Z(n545) );
  XOR U460 ( .A(n552), .B(n553), .Z(n543) );
  AND U461 ( .A(n117), .B(n554), .Z(n553) );
  XOR U462 ( .A(n555), .B(n556), .Z(n541) );
  AND U463 ( .A(n121), .B(n554), .Z(n556) );
  XNOR U464 ( .A(n555), .B(n552), .Z(n554) );
  XOR U465 ( .A(n557), .B(n558), .Z(n552) );
  AND U466 ( .A(n124), .B(n551), .Z(n558) );
  XNOR U467 ( .A(n559), .B(n549), .Z(n551) );
  XOR U468 ( .A(n560), .B(n561), .Z(n549) );
  AND U469 ( .A(n128), .B(n562), .Z(n561) );
  XOR U470 ( .A(p_input[55]), .B(n560), .Z(n562) );
  XOR U471 ( .A(n563), .B(n564), .Z(n560) );
  AND U472 ( .A(n132), .B(n565), .Z(n564) );
  IV U473 ( .A(n557), .Z(n559) );
  XOR U474 ( .A(n566), .B(n567), .Z(n557) );
  AND U475 ( .A(n136), .B(n568), .Z(n567) );
  XOR U476 ( .A(n569), .B(n570), .Z(n555) );
  AND U477 ( .A(n140), .B(n568), .Z(n570) );
  XNOR U478 ( .A(n569), .B(n566), .Z(n568) );
  XOR U479 ( .A(n571), .B(n572), .Z(n566) );
  AND U480 ( .A(n143), .B(n565), .Z(n572) );
  XNOR U481 ( .A(n573), .B(n563), .Z(n565) );
  XOR U482 ( .A(n574), .B(n575), .Z(n563) );
  AND U483 ( .A(n147), .B(n576), .Z(n575) );
  XOR U484 ( .A(p_input[71]), .B(n574), .Z(n576) );
  XOR U485 ( .A(n577), .B(n578), .Z(n574) );
  AND U486 ( .A(n151), .B(n579), .Z(n578) );
  IV U487 ( .A(n571), .Z(n573) );
  XOR U488 ( .A(n580), .B(n581), .Z(n571) );
  AND U489 ( .A(n155), .B(n582), .Z(n581) );
  XOR U490 ( .A(n583), .B(n584), .Z(n569) );
  AND U491 ( .A(n159), .B(n582), .Z(n584) );
  XNOR U492 ( .A(n583), .B(n580), .Z(n582) );
  XOR U493 ( .A(n585), .B(n586), .Z(n580) );
  AND U494 ( .A(n162), .B(n579), .Z(n586) );
  XNOR U495 ( .A(n587), .B(n577), .Z(n579) );
  XOR U496 ( .A(n588), .B(n589), .Z(n577) );
  AND U497 ( .A(n166), .B(n590), .Z(n589) );
  XOR U498 ( .A(p_input[87]), .B(n588), .Z(n590) );
  XOR U499 ( .A(n591), .B(n592), .Z(n588) );
  AND U500 ( .A(n170), .B(n593), .Z(n592) );
  IV U501 ( .A(n585), .Z(n587) );
  XOR U502 ( .A(n594), .B(n595), .Z(n585) );
  AND U503 ( .A(n174), .B(n596), .Z(n595) );
  XOR U504 ( .A(n597), .B(n598), .Z(n583) );
  AND U505 ( .A(n178), .B(n596), .Z(n598) );
  XNOR U506 ( .A(n597), .B(n594), .Z(n596) );
  XOR U507 ( .A(n599), .B(n600), .Z(n594) );
  AND U508 ( .A(n181), .B(n593), .Z(n600) );
  XNOR U509 ( .A(n601), .B(n591), .Z(n593) );
  XOR U510 ( .A(n602), .B(n603), .Z(n591) );
  AND U511 ( .A(n185), .B(n604), .Z(n603) );
  XOR U512 ( .A(p_input[103]), .B(n602), .Z(n604) );
  XOR U513 ( .A(n605), .B(n606), .Z(n602) );
  AND U514 ( .A(n189), .B(n607), .Z(n606) );
  IV U515 ( .A(n599), .Z(n601) );
  XOR U516 ( .A(n608), .B(n609), .Z(n599) );
  AND U517 ( .A(n193), .B(n610), .Z(n609) );
  XOR U518 ( .A(n611), .B(n612), .Z(n597) );
  AND U519 ( .A(n197), .B(n610), .Z(n612) );
  XNOR U520 ( .A(n611), .B(n608), .Z(n610) );
  XOR U521 ( .A(n613), .B(n614), .Z(n608) );
  AND U522 ( .A(n200), .B(n607), .Z(n614) );
  XNOR U523 ( .A(n615), .B(n605), .Z(n607) );
  XOR U524 ( .A(n616), .B(n617), .Z(n605) );
  AND U525 ( .A(n204), .B(n618), .Z(n617) );
  XOR U526 ( .A(p_input[119]), .B(n616), .Z(n618) );
  XOR U527 ( .A(n619), .B(n620), .Z(n616) );
  AND U528 ( .A(n208), .B(n621), .Z(n620) );
  IV U529 ( .A(n613), .Z(n615) );
  XOR U530 ( .A(n622), .B(n623), .Z(n613) );
  AND U531 ( .A(n212), .B(n624), .Z(n623) );
  XOR U532 ( .A(n625), .B(n626), .Z(n611) );
  AND U533 ( .A(n216), .B(n624), .Z(n626) );
  XNOR U534 ( .A(n625), .B(n622), .Z(n624) );
  XOR U535 ( .A(n627), .B(n628), .Z(n622) );
  AND U536 ( .A(n219), .B(n621), .Z(n628) );
  XNOR U537 ( .A(n629), .B(n619), .Z(n621) );
  XOR U538 ( .A(n630), .B(n631), .Z(n619) );
  AND U539 ( .A(n223), .B(n632), .Z(n631) );
  XOR U540 ( .A(p_input[135]), .B(n630), .Z(n632) );
  XOR U541 ( .A(n633), .B(n634), .Z(n630) );
  AND U542 ( .A(n227), .B(n635), .Z(n634) );
  IV U543 ( .A(n627), .Z(n629) );
  XOR U544 ( .A(n636), .B(n637), .Z(n627) );
  AND U545 ( .A(n231), .B(n638), .Z(n637) );
  XOR U546 ( .A(n639), .B(n640), .Z(n625) );
  AND U547 ( .A(n235), .B(n638), .Z(n640) );
  XNOR U548 ( .A(n639), .B(n636), .Z(n638) );
  XOR U549 ( .A(n641), .B(n642), .Z(n636) );
  AND U550 ( .A(n238), .B(n635), .Z(n642) );
  XNOR U551 ( .A(n643), .B(n633), .Z(n635) );
  XOR U552 ( .A(n644), .B(n645), .Z(n633) );
  AND U553 ( .A(n242), .B(n646), .Z(n645) );
  XOR U554 ( .A(p_input[151]), .B(n644), .Z(n646) );
  XOR U555 ( .A(n647), .B(n648), .Z(n644) );
  AND U556 ( .A(n246), .B(n649), .Z(n648) );
  IV U557 ( .A(n641), .Z(n643) );
  XOR U558 ( .A(n650), .B(n651), .Z(n641) );
  AND U559 ( .A(n250), .B(n652), .Z(n651) );
  XOR U560 ( .A(n653), .B(n654), .Z(n639) );
  AND U561 ( .A(n254), .B(n652), .Z(n654) );
  XNOR U562 ( .A(n653), .B(n650), .Z(n652) );
  XOR U563 ( .A(n655), .B(n656), .Z(n650) );
  AND U564 ( .A(n257), .B(n649), .Z(n656) );
  XNOR U565 ( .A(n657), .B(n647), .Z(n649) );
  XOR U566 ( .A(n658), .B(n659), .Z(n647) );
  AND U567 ( .A(n261), .B(n660), .Z(n659) );
  XOR U568 ( .A(p_input[167]), .B(n658), .Z(n660) );
  XOR U569 ( .A(n661), .B(n662), .Z(n658) );
  AND U570 ( .A(n265), .B(n663), .Z(n662) );
  IV U571 ( .A(n655), .Z(n657) );
  XOR U572 ( .A(n664), .B(n665), .Z(n655) );
  AND U573 ( .A(n269), .B(n666), .Z(n665) );
  XOR U574 ( .A(n667), .B(n668), .Z(n653) );
  AND U575 ( .A(n273), .B(n666), .Z(n668) );
  XNOR U576 ( .A(n667), .B(n664), .Z(n666) );
  XOR U577 ( .A(n669), .B(n670), .Z(n664) );
  AND U578 ( .A(n276), .B(n663), .Z(n670) );
  XNOR U579 ( .A(n671), .B(n661), .Z(n663) );
  XOR U580 ( .A(n672), .B(n673), .Z(n661) );
  AND U581 ( .A(n280), .B(n674), .Z(n673) );
  XOR U582 ( .A(p_input[183]), .B(n672), .Z(n674) );
  XOR U583 ( .A(n675), .B(n676), .Z(n672) );
  AND U584 ( .A(n284), .B(n677), .Z(n676) );
  IV U585 ( .A(n669), .Z(n671) );
  XOR U586 ( .A(n678), .B(n679), .Z(n669) );
  AND U587 ( .A(n288), .B(n680), .Z(n679) );
  XOR U588 ( .A(n681), .B(n682), .Z(n667) );
  AND U589 ( .A(n292), .B(n680), .Z(n682) );
  XNOR U590 ( .A(n681), .B(n678), .Z(n680) );
  XOR U591 ( .A(n683), .B(n684), .Z(n678) );
  AND U592 ( .A(n295), .B(n677), .Z(n684) );
  XNOR U593 ( .A(n685), .B(n675), .Z(n677) );
  XOR U594 ( .A(n686), .B(n687), .Z(n675) );
  AND U595 ( .A(n299), .B(n688), .Z(n687) );
  XOR U596 ( .A(p_input[199]), .B(n686), .Z(n688) );
  XOR U597 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n689), .Z(
        n686) );
  AND U598 ( .A(n302), .B(n690), .Z(n689) );
  IV U599 ( .A(n683), .Z(n685) );
  XOR U600 ( .A(n691), .B(n692), .Z(n683) );
  AND U601 ( .A(n306), .B(n693), .Z(n692) );
  XOR U602 ( .A(n694), .B(n695), .Z(n681) );
  AND U603 ( .A(n310), .B(n693), .Z(n695) );
  XNOR U604 ( .A(n694), .B(n691), .Z(n693) );
  XNOR U605 ( .A(n696), .B(n697), .Z(n691) );
  AND U606 ( .A(n313), .B(n690), .Z(n697) );
  XNOR U607 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n696), .Z(
        n690) );
  XNOR U608 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(n698), .Z(
        n696) );
  AND U609 ( .A(n315), .B(n699), .Z(n698) );
  XNOR U610 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n700), .Z(n694) );
  AND U611 ( .A(n318), .B(n699), .Z(n700) );
  XOR U612 ( .A(n701), .B(n702), .Z(n699) );
  IV U613 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .Z(n702) );
  IV U614 ( .A(\knn_comb_/min_val_out[0][7] ), .Z(n701) );
  XOR U615 ( .A(n7), .B(n703), .Z(o[22]) );
  AND U616 ( .A(n62), .B(n704), .Z(n7) );
  XOR U617 ( .A(n8), .B(n703), .Z(n704) );
  XOR U618 ( .A(n705), .B(n33), .Z(n703) );
  AND U619 ( .A(n65), .B(n706), .Z(n33) );
  XNOR U620 ( .A(n707), .B(n34), .Z(n706) );
  XOR U621 ( .A(n708), .B(n709), .Z(n34) );
  AND U622 ( .A(n70), .B(n710), .Z(n709) );
  XOR U623 ( .A(p_input[6]), .B(n708), .Z(n710) );
  XOR U624 ( .A(n711), .B(n712), .Z(n708) );
  AND U625 ( .A(n74), .B(n713), .Z(n712) );
  IV U626 ( .A(n705), .Z(n707) );
  XOR U627 ( .A(n714), .B(n715), .Z(n705) );
  AND U628 ( .A(n78), .B(n716), .Z(n715) );
  XOR U629 ( .A(n717), .B(n718), .Z(n8) );
  AND U630 ( .A(n82), .B(n716), .Z(n718) );
  XNOR U631 ( .A(n719), .B(n714), .Z(n716) );
  XOR U632 ( .A(n720), .B(n721), .Z(n714) );
  AND U633 ( .A(n86), .B(n713), .Z(n721) );
  XNOR U634 ( .A(n722), .B(n711), .Z(n713) );
  XOR U635 ( .A(n723), .B(n724), .Z(n711) );
  AND U636 ( .A(n90), .B(n725), .Z(n724) );
  XOR U637 ( .A(p_input[22]), .B(n723), .Z(n725) );
  XOR U638 ( .A(n726), .B(n727), .Z(n723) );
  AND U639 ( .A(n94), .B(n728), .Z(n727) );
  IV U640 ( .A(n720), .Z(n722) );
  XOR U641 ( .A(n729), .B(n730), .Z(n720) );
  AND U642 ( .A(n98), .B(n731), .Z(n730) );
  IV U643 ( .A(n717), .Z(n719) );
  XNOR U644 ( .A(n732), .B(n733), .Z(n717) );
  AND U645 ( .A(n102), .B(n731), .Z(n733) );
  XNOR U646 ( .A(n732), .B(n729), .Z(n731) );
  XOR U647 ( .A(n734), .B(n735), .Z(n729) );
  AND U648 ( .A(n105), .B(n728), .Z(n735) );
  XNOR U649 ( .A(n736), .B(n726), .Z(n728) );
  XOR U650 ( .A(n737), .B(n738), .Z(n726) );
  AND U651 ( .A(n109), .B(n739), .Z(n738) );
  XOR U652 ( .A(p_input[38]), .B(n737), .Z(n739) );
  XOR U653 ( .A(n740), .B(n741), .Z(n737) );
  AND U654 ( .A(n113), .B(n742), .Z(n741) );
  IV U655 ( .A(n734), .Z(n736) );
  XOR U656 ( .A(n743), .B(n744), .Z(n734) );
  AND U657 ( .A(n117), .B(n745), .Z(n744) );
  XOR U658 ( .A(n746), .B(n747), .Z(n732) );
  AND U659 ( .A(n121), .B(n745), .Z(n747) );
  XNOR U660 ( .A(n746), .B(n743), .Z(n745) );
  XOR U661 ( .A(n748), .B(n749), .Z(n743) );
  AND U662 ( .A(n124), .B(n742), .Z(n749) );
  XNOR U663 ( .A(n750), .B(n740), .Z(n742) );
  XOR U664 ( .A(n751), .B(n752), .Z(n740) );
  AND U665 ( .A(n128), .B(n753), .Z(n752) );
  XOR U666 ( .A(p_input[54]), .B(n751), .Z(n753) );
  XOR U667 ( .A(n754), .B(n755), .Z(n751) );
  AND U668 ( .A(n132), .B(n756), .Z(n755) );
  IV U669 ( .A(n748), .Z(n750) );
  XOR U670 ( .A(n757), .B(n758), .Z(n748) );
  AND U671 ( .A(n136), .B(n759), .Z(n758) );
  XOR U672 ( .A(n760), .B(n761), .Z(n746) );
  AND U673 ( .A(n140), .B(n759), .Z(n761) );
  XNOR U674 ( .A(n760), .B(n757), .Z(n759) );
  XOR U675 ( .A(n762), .B(n763), .Z(n757) );
  AND U676 ( .A(n143), .B(n756), .Z(n763) );
  XNOR U677 ( .A(n764), .B(n754), .Z(n756) );
  XOR U678 ( .A(n765), .B(n766), .Z(n754) );
  AND U679 ( .A(n147), .B(n767), .Z(n766) );
  XOR U680 ( .A(p_input[70]), .B(n765), .Z(n767) );
  XOR U681 ( .A(n768), .B(n769), .Z(n765) );
  AND U682 ( .A(n151), .B(n770), .Z(n769) );
  IV U683 ( .A(n762), .Z(n764) );
  XOR U684 ( .A(n771), .B(n772), .Z(n762) );
  AND U685 ( .A(n155), .B(n773), .Z(n772) );
  XOR U686 ( .A(n774), .B(n775), .Z(n760) );
  AND U687 ( .A(n159), .B(n773), .Z(n775) );
  XNOR U688 ( .A(n774), .B(n771), .Z(n773) );
  XOR U689 ( .A(n776), .B(n777), .Z(n771) );
  AND U690 ( .A(n162), .B(n770), .Z(n777) );
  XNOR U691 ( .A(n778), .B(n768), .Z(n770) );
  XOR U692 ( .A(n779), .B(n780), .Z(n768) );
  AND U693 ( .A(n166), .B(n781), .Z(n780) );
  XOR U694 ( .A(p_input[86]), .B(n779), .Z(n781) );
  XOR U695 ( .A(n782), .B(n783), .Z(n779) );
  AND U696 ( .A(n170), .B(n784), .Z(n783) );
  IV U697 ( .A(n776), .Z(n778) );
  XOR U698 ( .A(n785), .B(n786), .Z(n776) );
  AND U699 ( .A(n174), .B(n787), .Z(n786) );
  XOR U700 ( .A(n788), .B(n789), .Z(n774) );
  AND U701 ( .A(n178), .B(n787), .Z(n789) );
  XNOR U702 ( .A(n788), .B(n785), .Z(n787) );
  XOR U703 ( .A(n790), .B(n791), .Z(n785) );
  AND U704 ( .A(n181), .B(n784), .Z(n791) );
  XNOR U705 ( .A(n792), .B(n782), .Z(n784) );
  XOR U706 ( .A(n793), .B(n794), .Z(n782) );
  AND U707 ( .A(n185), .B(n795), .Z(n794) );
  XOR U708 ( .A(p_input[102]), .B(n793), .Z(n795) );
  XOR U709 ( .A(n796), .B(n797), .Z(n793) );
  AND U710 ( .A(n189), .B(n798), .Z(n797) );
  IV U711 ( .A(n790), .Z(n792) );
  XOR U712 ( .A(n799), .B(n800), .Z(n790) );
  AND U713 ( .A(n193), .B(n801), .Z(n800) );
  XOR U714 ( .A(n802), .B(n803), .Z(n788) );
  AND U715 ( .A(n197), .B(n801), .Z(n803) );
  XNOR U716 ( .A(n802), .B(n799), .Z(n801) );
  XOR U717 ( .A(n804), .B(n805), .Z(n799) );
  AND U718 ( .A(n200), .B(n798), .Z(n805) );
  XNOR U719 ( .A(n806), .B(n796), .Z(n798) );
  XOR U720 ( .A(n807), .B(n808), .Z(n796) );
  AND U721 ( .A(n204), .B(n809), .Z(n808) );
  XOR U722 ( .A(p_input[118]), .B(n807), .Z(n809) );
  XOR U723 ( .A(n810), .B(n811), .Z(n807) );
  AND U724 ( .A(n208), .B(n812), .Z(n811) );
  IV U725 ( .A(n804), .Z(n806) );
  XOR U726 ( .A(n813), .B(n814), .Z(n804) );
  AND U727 ( .A(n212), .B(n815), .Z(n814) );
  XOR U728 ( .A(n816), .B(n817), .Z(n802) );
  AND U729 ( .A(n216), .B(n815), .Z(n817) );
  XNOR U730 ( .A(n816), .B(n813), .Z(n815) );
  XOR U731 ( .A(n818), .B(n819), .Z(n813) );
  AND U732 ( .A(n219), .B(n812), .Z(n819) );
  XNOR U733 ( .A(n820), .B(n810), .Z(n812) );
  XOR U734 ( .A(n821), .B(n822), .Z(n810) );
  AND U735 ( .A(n223), .B(n823), .Z(n822) );
  XOR U736 ( .A(p_input[134]), .B(n821), .Z(n823) );
  XOR U737 ( .A(n824), .B(n825), .Z(n821) );
  AND U738 ( .A(n227), .B(n826), .Z(n825) );
  IV U739 ( .A(n818), .Z(n820) );
  XOR U740 ( .A(n827), .B(n828), .Z(n818) );
  AND U741 ( .A(n231), .B(n829), .Z(n828) );
  XOR U742 ( .A(n830), .B(n831), .Z(n816) );
  AND U743 ( .A(n235), .B(n829), .Z(n831) );
  XNOR U744 ( .A(n830), .B(n827), .Z(n829) );
  XOR U745 ( .A(n832), .B(n833), .Z(n827) );
  AND U746 ( .A(n238), .B(n826), .Z(n833) );
  XNOR U747 ( .A(n834), .B(n824), .Z(n826) );
  XOR U748 ( .A(n835), .B(n836), .Z(n824) );
  AND U749 ( .A(n242), .B(n837), .Z(n836) );
  XOR U750 ( .A(p_input[150]), .B(n835), .Z(n837) );
  XOR U751 ( .A(n838), .B(n839), .Z(n835) );
  AND U752 ( .A(n246), .B(n840), .Z(n839) );
  IV U753 ( .A(n832), .Z(n834) );
  XOR U754 ( .A(n841), .B(n842), .Z(n832) );
  AND U755 ( .A(n250), .B(n843), .Z(n842) );
  XOR U756 ( .A(n844), .B(n845), .Z(n830) );
  AND U757 ( .A(n254), .B(n843), .Z(n845) );
  XNOR U758 ( .A(n844), .B(n841), .Z(n843) );
  XOR U759 ( .A(n846), .B(n847), .Z(n841) );
  AND U760 ( .A(n257), .B(n840), .Z(n847) );
  XNOR U761 ( .A(n848), .B(n838), .Z(n840) );
  XOR U762 ( .A(n849), .B(n850), .Z(n838) );
  AND U763 ( .A(n261), .B(n851), .Z(n850) );
  XOR U764 ( .A(p_input[166]), .B(n849), .Z(n851) );
  XOR U765 ( .A(n852), .B(n853), .Z(n849) );
  AND U766 ( .A(n265), .B(n854), .Z(n853) );
  IV U767 ( .A(n846), .Z(n848) );
  XOR U768 ( .A(n855), .B(n856), .Z(n846) );
  AND U769 ( .A(n269), .B(n857), .Z(n856) );
  XOR U770 ( .A(n858), .B(n859), .Z(n844) );
  AND U771 ( .A(n273), .B(n857), .Z(n859) );
  XNOR U772 ( .A(n858), .B(n855), .Z(n857) );
  XOR U773 ( .A(n860), .B(n861), .Z(n855) );
  AND U774 ( .A(n276), .B(n854), .Z(n861) );
  XNOR U775 ( .A(n862), .B(n852), .Z(n854) );
  XOR U776 ( .A(n863), .B(n864), .Z(n852) );
  AND U777 ( .A(n280), .B(n865), .Z(n864) );
  XOR U778 ( .A(p_input[182]), .B(n863), .Z(n865) );
  XOR U779 ( .A(n866), .B(n867), .Z(n863) );
  AND U780 ( .A(n284), .B(n868), .Z(n867) );
  IV U781 ( .A(n860), .Z(n862) );
  XOR U782 ( .A(n869), .B(n870), .Z(n860) );
  AND U783 ( .A(n288), .B(n871), .Z(n870) );
  XOR U784 ( .A(n872), .B(n873), .Z(n858) );
  AND U785 ( .A(n292), .B(n871), .Z(n873) );
  XNOR U786 ( .A(n872), .B(n869), .Z(n871) );
  XOR U787 ( .A(n874), .B(n875), .Z(n869) );
  AND U788 ( .A(n295), .B(n868), .Z(n875) );
  XNOR U789 ( .A(n876), .B(n866), .Z(n868) );
  XOR U790 ( .A(n877), .B(n878), .Z(n866) );
  AND U791 ( .A(n299), .B(n879), .Z(n878) );
  XOR U792 ( .A(p_input[198]), .B(n877), .Z(n879) );
  XOR U793 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(n880), .Z(
        n877) );
  AND U794 ( .A(n302), .B(n881), .Z(n880) );
  IV U795 ( .A(n874), .Z(n876) );
  XOR U796 ( .A(n882), .B(n883), .Z(n874) );
  AND U797 ( .A(n306), .B(n884), .Z(n883) );
  XOR U798 ( .A(n885), .B(n886), .Z(n872) );
  AND U799 ( .A(n310), .B(n884), .Z(n886) );
  XNOR U800 ( .A(n885), .B(n882), .Z(n884) );
  XNOR U801 ( .A(n887), .B(n888), .Z(n882) );
  AND U802 ( .A(n313), .B(n881), .Z(n888) );
  XNOR U803 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(n887), .Z(
        n881) );
  XNOR U804 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .B(n889), .Z(
        n887) );
  AND U805 ( .A(n315), .B(n890), .Z(n889) );
  XNOR U806 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n891), .Z(n885) );
  AND U807 ( .A(n318), .B(n890), .Z(n891) );
  XOR U808 ( .A(n892), .B(n893), .Z(n890) );
  XOR U809 ( .A(n9), .B(n894), .Z(o[21]) );
  AND U810 ( .A(n62), .B(n895), .Z(n9) );
  XOR U811 ( .A(n10), .B(n894), .Z(n895) );
  XOR U812 ( .A(n896), .B(n35), .Z(n894) );
  AND U813 ( .A(n65), .B(n897), .Z(n35) );
  XNOR U814 ( .A(n898), .B(n36), .Z(n897) );
  XOR U815 ( .A(n899), .B(n900), .Z(n36) );
  AND U816 ( .A(n70), .B(n901), .Z(n900) );
  XOR U817 ( .A(p_input[5]), .B(n899), .Z(n901) );
  XOR U818 ( .A(n902), .B(n903), .Z(n899) );
  AND U819 ( .A(n74), .B(n904), .Z(n903) );
  IV U820 ( .A(n896), .Z(n898) );
  XOR U821 ( .A(n905), .B(n906), .Z(n896) );
  AND U822 ( .A(n78), .B(n907), .Z(n906) );
  XOR U823 ( .A(n908), .B(n909), .Z(n10) );
  AND U824 ( .A(n82), .B(n907), .Z(n909) );
  XNOR U825 ( .A(n910), .B(n905), .Z(n907) );
  XOR U826 ( .A(n911), .B(n912), .Z(n905) );
  AND U827 ( .A(n86), .B(n904), .Z(n912) );
  XNOR U828 ( .A(n913), .B(n902), .Z(n904) );
  XOR U829 ( .A(n914), .B(n915), .Z(n902) );
  AND U830 ( .A(n90), .B(n916), .Z(n915) );
  XOR U831 ( .A(p_input[21]), .B(n914), .Z(n916) );
  XOR U832 ( .A(n917), .B(n918), .Z(n914) );
  AND U833 ( .A(n94), .B(n919), .Z(n918) );
  IV U834 ( .A(n911), .Z(n913) );
  XOR U835 ( .A(n920), .B(n921), .Z(n911) );
  AND U836 ( .A(n98), .B(n922), .Z(n921) );
  IV U837 ( .A(n908), .Z(n910) );
  XNOR U838 ( .A(n923), .B(n924), .Z(n908) );
  AND U839 ( .A(n102), .B(n922), .Z(n924) );
  XNOR U840 ( .A(n923), .B(n920), .Z(n922) );
  XOR U841 ( .A(n925), .B(n926), .Z(n920) );
  AND U842 ( .A(n105), .B(n919), .Z(n926) );
  XNOR U843 ( .A(n927), .B(n917), .Z(n919) );
  XOR U844 ( .A(n928), .B(n929), .Z(n917) );
  AND U845 ( .A(n109), .B(n930), .Z(n929) );
  XOR U846 ( .A(p_input[37]), .B(n928), .Z(n930) );
  XOR U847 ( .A(n931), .B(n932), .Z(n928) );
  AND U848 ( .A(n113), .B(n933), .Z(n932) );
  IV U849 ( .A(n925), .Z(n927) );
  XOR U850 ( .A(n934), .B(n935), .Z(n925) );
  AND U851 ( .A(n117), .B(n936), .Z(n935) );
  XOR U852 ( .A(n937), .B(n938), .Z(n923) );
  AND U853 ( .A(n121), .B(n936), .Z(n938) );
  XNOR U854 ( .A(n937), .B(n934), .Z(n936) );
  XOR U855 ( .A(n939), .B(n940), .Z(n934) );
  AND U856 ( .A(n124), .B(n933), .Z(n940) );
  XNOR U857 ( .A(n941), .B(n931), .Z(n933) );
  XOR U858 ( .A(n942), .B(n943), .Z(n931) );
  AND U859 ( .A(n128), .B(n944), .Z(n943) );
  XOR U860 ( .A(p_input[53]), .B(n942), .Z(n944) );
  XOR U861 ( .A(n945), .B(n946), .Z(n942) );
  AND U862 ( .A(n132), .B(n947), .Z(n946) );
  IV U863 ( .A(n939), .Z(n941) );
  XOR U864 ( .A(n948), .B(n949), .Z(n939) );
  AND U865 ( .A(n136), .B(n950), .Z(n949) );
  XOR U866 ( .A(n951), .B(n952), .Z(n937) );
  AND U867 ( .A(n140), .B(n950), .Z(n952) );
  XNOR U868 ( .A(n951), .B(n948), .Z(n950) );
  XOR U869 ( .A(n953), .B(n954), .Z(n948) );
  AND U870 ( .A(n143), .B(n947), .Z(n954) );
  XNOR U871 ( .A(n955), .B(n945), .Z(n947) );
  XOR U872 ( .A(n956), .B(n957), .Z(n945) );
  AND U873 ( .A(n147), .B(n958), .Z(n957) );
  XOR U874 ( .A(p_input[69]), .B(n956), .Z(n958) );
  XOR U875 ( .A(n959), .B(n960), .Z(n956) );
  AND U876 ( .A(n151), .B(n961), .Z(n960) );
  IV U877 ( .A(n953), .Z(n955) );
  XOR U878 ( .A(n962), .B(n963), .Z(n953) );
  AND U879 ( .A(n155), .B(n964), .Z(n963) );
  XOR U880 ( .A(n965), .B(n966), .Z(n951) );
  AND U881 ( .A(n159), .B(n964), .Z(n966) );
  XNOR U882 ( .A(n965), .B(n962), .Z(n964) );
  XOR U883 ( .A(n967), .B(n968), .Z(n962) );
  AND U884 ( .A(n162), .B(n961), .Z(n968) );
  XNOR U885 ( .A(n969), .B(n959), .Z(n961) );
  XOR U886 ( .A(n970), .B(n971), .Z(n959) );
  AND U887 ( .A(n166), .B(n972), .Z(n971) );
  XOR U888 ( .A(p_input[85]), .B(n970), .Z(n972) );
  XOR U889 ( .A(n973), .B(n974), .Z(n970) );
  AND U890 ( .A(n170), .B(n975), .Z(n974) );
  IV U891 ( .A(n967), .Z(n969) );
  XOR U892 ( .A(n976), .B(n977), .Z(n967) );
  AND U893 ( .A(n174), .B(n978), .Z(n977) );
  XOR U894 ( .A(n979), .B(n980), .Z(n965) );
  AND U895 ( .A(n178), .B(n978), .Z(n980) );
  XNOR U896 ( .A(n979), .B(n976), .Z(n978) );
  XOR U897 ( .A(n981), .B(n982), .Z(n976) );
  AND U898 ( .A(n181), .B(n975), .Z(n982) );
  XNOR U899 ( .A(n983), .B(n973), .Z(n975) );
  XOR U900 ( .A(n984), .B(n985), .Z(n973) );
  AND U901 ( .A(n185), .B(n986), .Z(n985) );
  XOR U902 ( .A(p_input[101]), .B(n984), .Z(n986) );
  XOR U903 ( .A(n987), .B(n988), .Z(n984) );
  AND U904 ( .A(n189), .B(n989), .Z(n988) );
  IV U905 ( .A(n981), .Z(n983) );
  XOR U906 ( .A(n990), .B(n991), .Z(n981) );
  AND U907 ( .A(n193), .B(n992), .Z(n991) );
  XOR U908 ( .A(n993), .B(n994), .Z(n979) );
  AND U909 ( .A(n197), .B(n992), .Z(n994) );
  XNOR U910 ( .A(n993), .B(n990), .Z(n992) );
  XOR U911 ( .A(n995), .B(n996), .Z(n990) );
  AND U912 ( .A(n200), .B(n989), .Z(n996) );
  XNOR U913 ( .A(n997), .B(n987), .Z(n989) );
  XOR U914 ( .A(n998), .B(n999), .Z(n987) );
  AND U915 ( .A(n204), .B(n1000), .Z(n999) );
  XOR U916 ( .A(p_input[117]), .B(n998), .Z(n1000) );
  XOR U917 ( .A(n1001), .B(n1002), .Z(n998) );
  AND U918 ( .A(n208), .B(n1003), .Z(n1002) );
  IV U919 ( .A(n995), .Z(n997) );
  XOR U920 ( .A(n1004), .B(n1005), .Z(n995) );
  AND U921 ( .A(n212), .B(n1006), .Z(n1005) );
  XOR U922 ( .A(n1007), .B(n1008), .Z(n993) );
  AND U923 ( .A(n216), .B(n1006), .Z(n1008) );
  XNOR U924 ( .A(n1007), .B(n1004), .Z(n1006) );
  XOR U925 ( .A(n1009), .B(n1010), .Z(n1004) );
  AND U926 ( .A(n219), .B(n1003), .Z(n1010) );
  XNOR U927 ( .A(n1011), .B(n1001), .Z(n1003) );
  XOR U928 ( .A(n1012), .B(n1013), .Z(n1001) );
  AND U929 ( .A(n223), .B(n1014), .Z(n1013) );
  XOR U930 ( .A(p_input[133]), .B(n1012), .Z(n1014) );
  XOR U931 ( .A(n1015), .B(n1016), .Z(n1012) );
  AND U932 ( .A(n227), .B(n1017), .Z(n1016) );
  IV U933 ( .A(n1009), .Z(n1011) );
  XOR U934 ( .A(n1018), .B(n1019), .Z(n1009) );
  AND U935 ( .A(n231), .B(n1020), .Z(n1019) );
  XOR U936 ( .A(n1021), .B(n1022), .Z(n1007) );
  AND U937 ( .A(n235), .B(n1020), .Z(n1022) );
  XNOR U938 ( .A(n1021), .B(n1018), .Z(n1020) );
  XOR U939 ( .A(n1023), .B(n1024), .Z(n1018) );
  AND U940 ( .A(n238), .B(n1017), .Z(n1024) );
  XNOR U941 ( .A(n1025), .B(n1015), .Z(n1017) );
  XOR U942 ( .A(n1026), .B(n1027), .Z(n1015) );
  AND U943 ( .A(n242), .B(n1028), .Z(n1027) );
  XOR U944 ( .A(p_input[149]), .B(n1026), .Z(n1028) );
  XOR U945 ( .A(n1029), .B(n1030), .Z(n1026) );
  AND U946 ( .A(n246), .B(n1031), .Z(n1030) );
  IV U947 ( .A(n1023), .Z(n1025) );
  XOR U948 ( .A(n1032), .B(n1033), .Z(n1023) );
  AND U949 ( .A(n250), .B(n1034), .Z(n1033) );
  XOR U950 ( .A(n1035), .B(n1036), .Z(n1021) );
  AND U951 ( .A(n254), .B(n1034), .Z(n1036) );
  XNOR U952 ( .A(n1035), .B(n1032), .Z(n1034) );
  XOR U953 ( .A(n1037), .B(n1038), .Z(n1032) );
  AND U954 ( .A(n257), .B(n1031), .Z(n1038) );
  XNOR U955 ( .A(n1039), .B(n1029), .Z(n1031) );
  XOR U956 ( .A(n1040), .B(n1041), .Z(n1029) );
  AND U957 ( .A(n261), .B(n1042), .Z(n1041) );
  XOR U958 ( .A(p_input[165]), .B(n1040), .Z(n1042) );
  XOR U959 ( .A(n1043), .B(n1044), .Z(n1040) );
  AND U960 ( .A(n265), .B(n1045), .Z(n1044) );
  IV U961 ( .A(n1037), .Z(n1039) );
  XOR U962 ( .A(n1046), .B(n1047), .Z(n1037) );
  AND U963 ( .A(n269), .B(n1048), .Z(n1047) );
  XOR U964 ( .A(n1049), .B(n1050), .Z(n1035) );
  AND U965 ( .A(n273), .B(n1048), .Z(n1050) );
  XNOR U966 ( .A(n1049), .B(n1046), .Z(n1048) );
  XOR U967 ( .A(n1051), .B(n1052), .Z(n1046) );
  AND U968 ( .A(n276), .B(n1045), .Z(n1052) );
  XNOR U969 ( .A(n1053), .B(n1043), .Z(n1045) );
  XOR U970 ( .A(n1054), .B(n1055), .Z(n1043) );
  AND U971 ( .A(n280), .B(n1056), .Z(n1055) );
  XOR U972 ( .A(p_input[181]), .B(n1054), .Z(n1056) );
  XOR U973 ( .A(n1057), .B(n1058), .Z(n1054) );
  AND U974 ( .A(n284), .B(n1059), .Z(n1058) );
  IV U975 ( .A(n1051), .Z(n1053) );
  XOR U976 ( .A(n1060), .B(n1061), .Z(n1051) );
  AND U977 ( .A(n288), .B(n1062), .Z(n1061) );
  XOR U978 ( .A(n1063), .B(n1064), .Z(n1049) );
  AND U979 ( .A(n292), .B(n1062), .Z(n1064) );
  XNOR U980 ( .A(n1063), .B(n1060), .Z(n1062) );
  XOR U981 ( .A(n1065), .B(n1066), .Z(n1060) );
  AND U982 ( .A(n295), .B(n1059), .Z(n1066) );
  XNOR U983 ( .A(n1067), .B(n1057), .Z(n1059) );
  XOR U984 ( .A(n1068), .B(n1069), .Z(n1057) );
  AND U985 ( .A(n299), .B(n1070), .Z(n1069) );
  XOR U986 ( .A(p_input[197]), .B(n1068), .Z(n1070) );
  XOR U987 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n1071), .Z(
        n1068) );
  AND U988 ( .A(n302), .B(n1072), .Z(n1071) );
  IV U989 ( .A(n1065), .Z(n1067) );
  XOR U990 ( .A(n1073), .B(n1074), .Z(n1065) );
  AND U991 ( .A(n306), .B(n1075), .Z(n1074) );
  XOR U992 ( .A(n1076), .B(n1077), .Z(n1063) );
  AND U993 ( .A(n310), .B(n1075), .Z(n1077) );
  XNOR U994 ( .A(n1076), .B(n1073), .Z(n1075) );
  XNOR U995 ( .A(n1078), .B(n1079), .Z(n1073) );
  AND U996 ( .A(n313), .B(n1072), .Z(n1079) );
  XNOR U997 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n1078), 
        .Z(n1072) );
  XNOR U998 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(n1080), 
        .Z(n1078) );
  AND U999 ( .A(n315), .B(n1081), .Z(n1080) );
  XNOR U1000 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n1082), .Z(n1076) );
  AND U1001 ( .A(n318), .B(n1081), .Z(n1082) );
  XOR U1002 ( .A(n1083), .B(n1084), .Z(n1081) );
  XOR U1003 ( .A(n11), .B(n1085), .Z(o[20]) );
  AND U1004 ( .A(n62), .B(n1086), .Z(n11) );
  XOR U1005 ( .A(n12), .B(n1085), .Z(n1086) );
  XOR U1006 ( .A(n1087), .B(n37), .Z(n1085) );
  AND U1007 ( .A(n65), .B(n1088), .Z(n37) );
  XNOR U1008 ( .A(n1089), .B(n38), .Z(n1088) );
  XOR U1009 ( .A(n1090), .B(n1091), .Z(n38) );
  AND U1010 ( .A(n70), .B(n1092), .Z(n1091) );
  XOR U1011 ( .A(p_input[4]), .B(n1090), .Z(n1092) );
  XOR U1012 ( .A(n1093), .B(n1094), .Z(n1090) );
  AND U1013 ( .A(n74), .B(n1095), .Z(n1094) );
  IV U1014 ( .A(n1087), .Z(n1089) );
  XOR U1015 ( .A(n1096), .B(n1097), .Z(n1087) );
  AND U1016 ( .A(n78), .B(n1098), .Z(n1097) );
  XOR U1017 ( .A(n1099), .B(n1100), .Z(n12) );
  AND U1018 ( .A(n82), .B(n1098), .Z(n1100) );
  XNOR U1019 ( .A(n1101), .B(n1096), .Z(n1098) );
  XOR U1020 ( .A(n1102), .B(n1103), .Z(n1096) );
  AND U1021 ( .A(n86), .B(n1095), .Z(n1103) );
  XNOR U1022 ( .A(n1104), .B(n1093), .Z(n1095) );
  XOR U1023 ( .A(n1105), .B(n1106), .Z(n1093) );
  AND U1024 ( .A(n90), .B(n1107), .Z(n1106) );
  XOR U1025 ( .A(p_input[20]), .B(n1105), .Z(n1107) );
  XOR U1026 ( .A(n1108), .B(n1109), .Z(n1105) );
  AND U1027 ( .A(n94), .B(n1110), .Z(n1109) );
  IV U1028 ( .A(n1102), .Z(n1104) );
  XOR U1029 ( .A(n1111), .B(n1112), .Z(n1102) );
  AND U1030 ( .A(n98), .B(n1113), .Z(n1112) );
  IV U1031 ( .A(n1099), .Z(n1101) );
  XNOR U1032 ( .A(n1114), .B(n1115), .Z(n1099) );
  AND U1033 ( .A(n102), .B(n1113), .Z(n1115) );
  XNOR U1034 ( .A(n1114), .B(n1111), .Z(n1113) );
  XOR U1035 ( .A(n1116), .B(n1117), .Z(n1111) );
  AND U1036 ( .A(n105), .B(n1110), .Z(n1117) );
  XNOR U1037 ( .A(n1118), .B(n1108), .Z(n1110) );
  XOR U1038 ( .A(n1119), .B(n1120), .Z(n1108) );
  AND U1039 ( .A(n109), .B(n1121), .Z(n1120) );
  XOR U1040 ( .A(p_input[36]), .B(n1119), .Z(n1121) );
  XOR U1041 ( .A(n1122), .B(n1123), .Z(n1119) );
  AND U1042 ( .A(n113), .B(n1124), .Z(n1123) );
  IV U1043 ( .A(n1116), .Z(n1118) );
  XOR U1044 ( .A(n1125), .B(n1126), .Z(n1116) );
  AND U1045 ( .A(n117), .B(n1127), .Z(n1126) );
  XOR U1046 ( .A(n1128), .B(n1129), .Z(n1114) );
  AND U1047 ( .A(n121), .B(n1127), .Z(n1129) );
  XNOR U1048 ( .A(n1128), .B(n1125), .Z(n1127) );
  XOR U1049 ( .A(n1130), .B(n1131), .Z(n1125) );
  AND U1050 ( .A(n124), .B(n1124), .Z(n1131) );
  XNOR U1051 ( .A(n1132), .B(n1122), .Z(n1124) );
  XOR U1052 ( .A(n1133), .B(n1134), .Z(n1122) );
  AND U1053 ( .A(n128), .B(n1135), .Z(n1134) );
  XOR U1054 ( .A(p_input[52]), .B(n1133), .Z(n1135) );
  XOR U1055 ( .A(n1136), .B(n1137), .Z(n1133) );
  AND U1056 ( .A(n132), .B(n1138), .Z(n1137) );
  IV U1057 ( .A(n1130), .Z(n1132) );
  XOR U1058 ( .A(n1139), .B(n1140), .Z(n1130) );
  AND U1059 ( .A(n136), .B(n1141), .Z(n1140) );
  XOR U1060 ( .A(n1142), .B(n1143), .Z(n1128) );
  AND U1061 ( .A(n140), .B(n1141), .Z(n1143) );
  XNOR U1062 ( .A(n1142), .B(n1139), .Z(n1141) );
  XOR U1063 ( .A(n1144), .B(n1145), .Z(n1139) );
  AND U1064 ( .A(n143), .B(n1138), .Z(n1145) );
  XNOR U1065 ( .A(n1146), .B(n1136), .Z(n1138) );
  XOR U1066 ( .A(n1147), .B(n1148), .Z(n1136) );
  AND U1067 ( .A(n147), .B(n1149), .Z(n1148) );
  XOR U1068 ( .A(p_input[68]), .B(n1147), .Z(n1149) );
  XOR U1069 ( .A(n1150), .B(n1151), .Z(n1147) );
  AND U1070 ( .A(n151), .B(n1152), .Z(n1151) );
  IV U1071 ( .A(n1144), .Z(n1146) );
  XOR U1072 ( .A(n1153), .B(n1154), .Z(n1144) );
  AND U1073 ( .A(n155), .B(n1155), .Z(n1154) );
  XOR U1074 ( .A(n1156), .B(n1157), .Z(n1142) );
  AND U1075 ( .A(n159), .B(n1155), .Z(n1157) );
  XNOR U1076 ( .A(n1156), .B(n1153), .Z(n1155) );
  XOR U1077 ( .A(n1158), .B(n1159), .Z(n1153) );
  AND U1078 ( .A(n162), .B(n1152), .Z(n1159) );
  XNOR U1079 ( .A(n1160), .B(n1150), .Z(n1152) );
  XOR U1080 ( .A(n1161), .B(n1162), .Z(n1150) );
  AND U1081 ( .A(n166), .B(n1163), .Z(n1162) );
  XOR U1082 ( .A(p_input[84]), .B(n1161), .Z(n1163) );
  XOR U1083 ( .A(n1164), .B(n1165), .Z(n1161) );
  AND U1084 ( .A(n170), .B(n1166), .Z(n1165) );
  IV U1085 ( .A(n1158), .Z(n1160) );
  XOR U1086 ( .A(n1167), .B(n1168), .Z(n1158) );
  AND U1087 ( .A(n174), .B(n1169), .Z(n1168) );
  XOR U1088 ( .A(n1170), .B(n1171), .Z(n1156) );
  AND U1089 ( .A(n178), .B(n1169), .Z(n1171) );
  XNOR U1090 ( .A(n1170), .B(n1167), .Z(n1169) );
  XOR U1091 ( .A(n1172), .B(n1173), .Z(n1167) );
  AND U1092 ( .A(n181), .B(n1166), .Z(n1173) );
  XNOR U1093 ( .A(n1174), .B(n1164), .Z(n1166) );
  XOR U1094 ( .A(n1175), .B(n1176), .Z(n1164) );
  AND U1095 ( .A(n185), .B(n1177), .Z(n1176) );
  XOR U1096 ( .A(p_input[100]), .B(n1175), .Z(n1177) );
  XOR U1097 ( .A(n1178), .B(n1179), .Z(n1175) );
  AND U1098 ( .A(n189), .B(n1180), .Z(n1179) );
  IV U1099 ( .A(n1172), .Z(n1174) );
  XOR U1100 ( .A(n1181), .B(n1182), .Z(n1172) );
  AND U1101 ( .A(n193), .B(n1183), .Z(n1182) );
  XOR U1102 ( .A(n1184), .B(n1185), .Z(n1170) );
  AND U1103 ( .A(n197), .B(n1183), .Z(n1185) );
  XNOR U1104 ( .A(n1184), .B(n1181), .Z(n1183) );
  XOR U1105 ( .A(n1186), .B(n1187), .Z(n1181) );
  AND U1106 ( .A(n200), .B(n1180), .Z(n1187) );
  XNOR U1107 ( .A(n1188), .B(n1178), .Z(n1180) );
  XOR U1108 ( .A(n1189), .B(n1190), .Z(n1178) );
  AND U1109 ( .A(n204), .B(n1191), .Z(n1190) );
  XOR U1110 ( .A(p_input[116]), .B(n1189), .Z(n1191) );
  XOR U1111 ( .A(n1192), .B(n1193), .Z(n1189) );
  AND U1112 ( .A(n208), .B(n1194), .Z(n1193) );
  IV U1113 ( .A(n1186), .Z(n1188) );
  XOR U1114 ( .A(n1195), .B(n1196), .Z(n1186) );
  AND U1115 ( .A(n212), .B(n1197), .Z(n1196) );
  XOR U1116 ( .A(n1198), .B(n1199), .Z(n1184) );
  AND U1117 ( .A(n216), .B(n1197), .Z(n1199) );
  XNOR U1118 ( .A(n1198), .B(n1195), .Z(n1197) );
  XOR U1119 ( .A(n1200), .B(n1201), .Z(n1195) );
  AND U1120 ( .A(n219), .B(n1194), .Z(n1201) );
  XNOR U1121 ( .A(n1202), .B(n1192), .Z(n1194) );
  XOR U1122 ( .A(n1203), .B(n1204), .Z(n1192) );
  AND U1123 ( .A(n223), .B(n1205), .Z(n1204) );
  XOR U1124 ( .A(p_input[132]), .B(n1203), .Z(n1205) );
  XOR U1125 ( .A(n1206), .B(n1207), .Z(n1203) );
  AND U1126 ( .A(n227), .B(n1208), .Z(n1207) );
  IV U1127 ( .A(n1200), .Z(n1202) );
  XOR U1128 ( .A(n1209), .B(n1210), .Z(n1200) );
  AND U1129 ( .A(n231), .B(n1211), .Z(n1210) );
  XOR U1130 ( .A(n1212), .B(n1213), .Z(n1198) );
  AND U1131 ( .A(n235), .B(n1211), .Z(n1213) );
  XNOR U1132 ( .A(n1212), .B(n1209), .Z(n1211) );
  XOR U1133 ( .A(n1214), .B(n1215), .Z(n1209) );
  AND U1134 ( .A(n238), .B(n1208), .Z(n1215) );
  XNOR U1135 ( .A(n1216), .B(n1206), .Z(n1208) );
  XOR U1136 ( .A(n1217), .B(n1218), .Z(n1206) );
  AND U1137 ( .A(n242), .B(n1219), .Z(n1218) );
  XOR U1138 ( .A(p_input[148]), .B(n1217), .Z(n1219) );
  XOR U1139 ( .A(n1220), .B(n1221), .Z(n1217) );
  AND U1140 ( .A(n246), .B(n1222), .Z(n1221) );
  IV U1141 ( .A(n1214), .Z(n1216) );
  XOR U1142 ( .A(n1223), .B(n1224), .Z(n1214) );
  AND U1143 ( .A(n250), .B(n1225), .Z(n1224) );
  XOR U1144 ( .A(n1226), .B(n1227), .Z(n1212) );
  AND U1145 ( .A(n254), .B(n1225), .Z(n1227) );
  XNOR U1146 ( .A(n1226), .B(n1223), .Z(n1225) );
  XOR U1147 ( .A(n1228), .B(n1229), .Z(n1223) );
  AND U1148 ( .A(n257), .B(n1222), .Z(n1229) );
  XNOR U1149 ( .A(n1230), .B(n1220), .Z(n1222) );
  XOR U1150 ( .A(n1231), .B(n1232), .Z(n1220) );
  AND U1151 ( .A(n261), .B(n1233), .Z(n1232) );
  XOR U1152 ( .A(p_input[164]), .B(n1231), .Z(n1233) );
  XOR U1153 ( .A(n1234), .B(n1235), .Z(n1231) );
  AND U1154 ( .A(n265), .B(n1236), .Z(n1235) );
  IV U1155 ( .A(n1228), .Z(n1230) );
  XOR U1156 ( .A(n1237), .B(n1238), .Z(n1228) );
  AND U1157 ( .A(n269), .B(n1239), .Z(n1238) );
  XOR U1158 ( .A(n1240), .B(n1241), .Z(n1226) );
  AND U1159 ( .A(n273), .B(n1239), .Z(n1241) );
  XNOR U1160 ( .A(n1240), .B(n1237), .Z(n1239) );
  XOR U1161 ( .A(n1242), .B(n1243), .Z(n1237) );
  AND U1162 ( .A(n276), .B(n1236), .Z(n1243) );
  XNOR U1163 ( .A(n1244), .B(n1234), .Z(n1236) );
  XOR U1164 ( .A(n1245), .B(n1246), .Z(n1234) );
  AND U1165 ( .A(n280), .B(n1247), .Z(n1246) );
  XOR U1166 ( .A(p_input[180]), .B(n1245), .Z(n1247) );
  XOR U1167 ( .A(n1248), .B(n1249), .Z(n1245) );
  AND U1168 ( .A(n284), .B(n1250), .Z(n1249) );
  IV U1169 ( .A(n1242), .Z(n1244) );
  XOR U1170 ( .A(n1251), .B(n1252), .Z(n1242) );
  AND U1171 ( .A(n288), .B(n1253), .Z(n1252) );
  XOR U1172 ( .A(n1254), .B(n1255), .Z(n1240) );
  AND U1173 ( .A(n292), .B(n1253), .Z(n1255) );
  XNOR U1174 ( .A(n1254), .B(n1251), .Z(n1253) );
  XOR U1175 ( .A(n1256), .B(n1257), .Z(n1251) );
  AND U1176 ( .A(n295), .B(n1250), .Z(n1257) );
  XNOR U1177 ( .A(n1258), .B(n1248), .Z(n1250) );
  XOR U1178 ( .A(n1259), .B(n1260), .Z(n1248) );
  AND U1179 ( .A(n299), .B(n1261), .Z(n1260) );
  XOR U1180 ( .A(p_input[196]), .B(n1259), .Z(n1261) );
  XOR U1181 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n1262), 
        .Z(n1259) );
  AND U1182 ( .A(n302), .B(n1263), .Z(n1262) );
  IV U1183 ( .A(n1256), .Z(n1258) );
  XOR U1184 ( .A(n1264), .B(n1265), .Z(n1256) );
  AND U1185 ( .A(n306), .B(n1266), .Z(n1265) );
  XOR U1186 ( .A(n1267), .B(n1268), .Z(n1254) );
  AND U1187 ( .A(n310), .B(n1266), .Z(n1268) );
  XNOR U1188 ( .A(n1267), .B(n1264), .Z(n1266) );
  XNOR U1189 ( .A(n1269), .B(n1270), .Z(n1264) );
  AND U1190 ( .A(n313), .B(n1263), .Z(n1270) );
  XNOR U1191 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n1269), 
        .Z(n1263) );
  XNOR U1192 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(n1271), 
        .Z(n1269) );
  AND U1193 ( .A(n315), .B(n1272), .Z(n1271) );
  XNOR U1194 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n1273), .Z(n1267) );
  AND U1195 ( .A(n318), .B(n1272), .Z(n1273) );
  XOR U1196 ( .A(n1274), .B(n1275), .Z(n1272) );
  IV U1197 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .Z(n1275) );
  IV U1198 ( .A(\knn_comb_/min_val_out[0][4] ), .Z(n1274) );
  XOR U1199 ( .A(n1276), .B(n1277), .Z(o[1]) );
  XOR U1200 ( .A(n29), .B(n1278), .Z(o[19]) );
  AND U1201 ( .A(n62), .B(n1279), .Z(n29) );
  XOR U1202 ( .A(n30), .B(n1278), .Z(n1279) );
  XOR U1203 ( .A(n1280), .B(n39), .Z(n1278) );
  AND U1204 ( .A(n65), .B(n1281), .Z(n39) );
  XNOR U1205 ( .A(n1282), .B(n40), .Z(n1281) );
  XOR U1206 ( .A(n1283), .B(n1284), .Z(n40) );
  AND U1207 ( .A(n70), .B(n1285), .Z(n1284) );
  XOR U1208 ( .A(p_input[3]), .B(n1283), .Z(n1285) );
  XOR U1209 ( .A(n1286), .B(n1287), .Z(n1283) );
  AND U1210 ( .A(n74), .B(n1288), .Z(n1287) );
  IV U1211 ( .A(n1280), .Z(n1282) );
  XOR U1212 ( .A(n1289), .B(n1290), .Z(n1280) );
  AND U1213 ( .A(n78), .B(n1291), .Z(n1290) );
  XOR U1214 ( .A(n1292), .B(n1293), .Z(n30) );
  AND U1215 ( .A(n82), .B(n1291), .Z(n1293) );
  XNOR U1216 ( .A(n1294), .B(n1289), .Z(n1291) );
  XOR U1217 ( .A(n1295), .B(n1296), .Z(n1289) );
  AND U1218 ( .A(n86), .B(n1288), .Z(n1296) );
  XNOR U1219 ( .A(n1297), .B(n1286), .Z(n1288) );
  XOR U1220 ( .A(n1298), .B(n1299), .Z(n1286) );
  AND U1221 ( .A(n90), .B(n1300), .Z(n1299) );
  XOR U1222 ( .A(p_input[19]), .B(n1298), .Z(n1300) );
  XOR U1223 ( .A(n1301), .B(n1302), .Z(n1298) );
  AND U1224 ( .A(n94), .B(n1303), .Z(n1302) );
  IV U1225 ( .A(n1295), .Z(n1297) );
  XOR U1226 ( .A(n1304), .B(n1305), .Z(n1295) );
  AND U1227 ( .A(n98), .B(n1306), .Z(n1305) );
  IV U1228 ( .A(n1292), .Z(n1294) );
  XNOR U1229 ( .A(n1307), .B(n1308), .Z(n1292) );
  AND U1230 ( .A(n102), .B(n1306), .Z(n1308) );
  XNOR U1231 ( .A(n1307), .B(n1304), .Z(n1306) );
  XOR U1232 ( .A(n1309), .B(n1310), .Z(n1304) );
  AND U1233 ( .A(n105), .B(n1303), .Z(n1310) );
  XNOR U1234 ( .A(n1311), .B(n1301), .Z(n1303) );
  XOR U1235 ( .A(n1312), .B(n1313), .Z(n1301) );
  AND U1236 ( .A(n109), .B(n1314), .Z(n1313) );
  XOR U1237 ( .A(p_input[35]), .B(n1312), .Z(n1314) );
  XOR U1238 ( .A(n1315), .B(n1316), .Z(n1312) );
  AND U1239 ( .A(n113), .B(n1317), .Z(n1316) );
  IV U1240 ( .A(n1309), .Z(n1311) );
  XOR U1241 ( .A(n1318), .B(n1319), .Z(n1309) );
  AND U1242 ( .A(n117), .B(n1320), .Z(n1319) );
  XOR U1243 ( .A(n1321), .B(n1322), .Z(n1307) );
  AND U1244 ( .A(n121), .B(n1320), .Z(n1322) );
  XNOR U1245 ( .A(n1321), .B(n1318), .Z(n1320) );
  XOR U1246 ( .A(n1323), .B(n1324), .Z(n1318) );
  AND U1247 ( .A(n124), .B(n1317), .Z(n1324) );
  XNOR U1248 ( .A(n1325), .B(n1315), .Z(n1317) );
  XOR U1249 ( .A(n1326), .B(n1327), .Z(n1315) );
  AND U1250 ( .A(n128), .B(n1328), .Z(n1327) );
  XOR U1251 ( .A(p_input[51]), .B(n1326), .Z(n1328) );
  XOR U1252 ( .A(n1329), .B(n1330), .Z(n1326) );
  AND U1253 ( .A(n132), .B(n1331), .Z(n1330) );
  IV U1254 ( .A(n1323), .Z(n1325) );
  XOR U1255 ( .A(n1332), .B(n1333), .Z(n1323) );
  AND U1256 ( .A(n136), .B(n1334), .Z(n1333) );
  XOR U1257 ( .A(n1335), .B(n1336), .Z(n1321) );
  AND U1258 ( .A(n140), .B(n1334), .Z(n1336) );
  XNOR U1259 ( .A(n1335), .B(n1332), .Z(n1334) );
  XOR U1260 ( .A(n1337), .B(n1338), .Z(n1332) );
  AND U1261 ( .A(n143), .B(n1331), .Z(n1338) );
  XNOR U1262 ( .A(n1339), .B(n1329), .Z(n1331) );
  XOR U1263 ( .A(n1340), .B(n1341), .Z(n1329) );
  AND U1264 ( .A(n147), .B(n1342), .Z(n1341) );
  XOR U1265 ( .A(p_input[67]), .B(n1340), .Z(n1342) );
  XOR U1266 ( .A(n1343), .B(n1344), .Z(n1340) );
  AND U1267 ( .A(n151), .B(n1345), .Z(n1344) );
  IV U1268 ( .A(n1337), .Z(n1339) );
  XOR U1269 ( .A(n1346), .B(n1347), .Z(n1337) );
  AND U1270 ( .A(n155), .B(n1348), .Z(n1347) );
  XOR U1271 ( .A(n1349), .B(n1350), .Z(n1335) );
  AND U1272 ( .A(n159), .B(n1348), .Z(n1350) );
  XNOR U1273 ( .A(n1349), .B(n1346), .Z(n1348) );
  XOR U1274 ( .A(n1351), .B(n1352), .Z(n1346) );
  AND U1275 ( .A(n162), .B(n1345), .Z(n1352) );
  XNOR U1276 ( .A(n1353), .B(n1343), .Z(n1345) );
  XOR U1277 ( .A(n1354), .B(n1355), .Z(n1343) );
  AND U1278 ( .A(n166), .B(n1356), .Z(n1355) );
  XOR U1279 ( .A(p_input[83]), .B(n1354), .Z(n1356) );
  XOR U1280 ( .A(n1357), .B(n1358), .Z(n1354) );
  AND U1281 ( .A(n170), .B(n1359), .Z(n1358) );
  IV U1282 ( .A(n1351), .Z(n1353) );
  XOR U1283 ( .A(n1360), .B(n1361), .Z(n1351) );
  AND U1284 ( .A(n174), .B(n1362), .Z(n1361) );
  XOR U1285 ( .A(n1363), .B(n1364), .Z(n1349) );
  AND U1286 ( .A(n178), .B(n1362), .Z(n1364) );
  XNOR U1287 ( .A(n1363), .B(n1360), .Z(n1362) );
  XOR U1288 ( .A(n1365), .B(n1366), .Z(n1360) );
  AND U1289 ( .A(n181), .B(n1359), .Z(n1366) );
  XNOR U1290 ( .A(n1367), .B(n1357), .Z(n1359) );
  XOR U1291 ( .A(n1368), .B(n1369), .Z(n1357) );
  AND U1292 ( .A(n185), .B(n1370), .Z(n1369) );
  XOR U1293 ( .A(p_input[99]), .B(n1368), .Z(n1370) );
  XOR U1294 ( .A(n1371), .B(n1372), .Z(n1368) );
  AND U1295 ( .A(n189), .B(n1373), .Z(n1372) );
  IV U1296 ( .A(n1365), .Z(n1367) );
  XOR U1297 ( .A(n1374), .B(n1375), .Z(n1365) );
  AND U1298 ( .A(n193), .B(n1376), .Z(n1375) );
  XOR U1299 ( .A(n1377), .B(n1378), .Z(n1363) );
  AND U1300 ( .A(n197), .B(n1376), .Z(n1378) );
  XNOR U1301 ( .A(n1377), .B(n1374), .Z(n1376) );
  XOR U1302 ( .A(n1379), .B(n1380), .Z(n1374) );
  AND U1303 ( .A(n200), .B(n1373), .Z(n1380) );
  XNOR U1304 ( .A(n1381), .B(n1371), .Z(n1373) );
  XOR U1305 ( .A(n1382), .B(n1383), .Z(n1371) );
  AND U1306 ( .A(n204), .B(n1384), .Z(n1383) );
  XOR U1307 ( .A(p_input[115]), .B(n1382), .Z(n1384) );
  XOR U1308 ( .A(n1385), .B(n1386), .Z(n1382) );
  AND U1309 ( .A(n208), .B(n1387), .Z(n1386) );
  IV U1310 ( .A(n1379), .Z(n1381) );
  XOR U1311 ( .A(n1388), .B(n1389), .Z(n1379) );
  AND U1312 ( .A(n212), .B(n1390), .Z(n1389) );
  XOR U1313 ( .A(n1391), .B(n1392), .Z(n1377) );
  AND U1314 ( .A(n216), .B(n1390), .Z(n1392) );
  XNOR U1315 ( .A(n1391), .B(n1388), .Z(n1390) );
  XOR U1316 ( .A(n1393), .B(n1394), .Z(n1388) );
  AND U1317 ( .A(n219), .B(n1387), .Z(n1394) );
  XNOR U1318 ( .A(n1395), .B(n1385), .Z(n1387) );
  XOR U1319 ( .A(n1396), .B(n1397), .Z(n1385) );
  AND U1320 ( .A(n223), .B(n1398), .Z(n1397) );
  XOR U1321 ( .A(p_input[131]), .B(n1396), .Z(n1398) );
  XOR U1322 ( .A(n1399), .B(n1400), .Z(n1396) );
  AND U1323 ( .A(n227), .B(n1401), .Z(n1400) );
  IV U1324 ( .A(n1393), .Z(n1395) );
  XOR U1325 ( .A(n1402), .B(n1403), .Z(n1393) );
  AND U1326 ( .A(n231), .B(n1404), .Z(n1403) );
  XOR U1327 ( .A(n1405), .B(n1406), .Z(n1391) );
  AND U1328 ( .A(n235), .B(n1404), .Z(n1406) );
  XNOR U1329 ( .A(n1405), .B(n1402), .Z(n1404) );
  XOR U1330 ( .A(n1407), .B(n1408), .Z(n1402) );
  AND U1331 ( .A(n238), .B(n1401), .Z(n1408) );
  XNOR U1332 ( .A(n1409), .B(n1399), .Z(n1401) );
  XOR U1333 ( .A(n1410), .B(n1411), .Z(n1399) );
  AND U1334 ( .A(n242), .B(n1412), .Z(n1411) );
  XOR U1335 ( .A(p_input[147]), .B(n1410), .Z(n1412) );
  XOR U1336 ( .A(n1413), .B(n1414), .Z(n1410) );
  AND U1337 ( .A(n246), .B(n1415), .Z(n1414) );
  IV U1338 ( .A(n1407), .Z(n1409) );
  XOR U1339 ( .A(n1416), .B(n1417), .Z(n1407) );
  AND U1340 ( .A(n250), .B(n1418), .Z(n1417) );
  XOR U1341 ( .A(n1419), .B(n1420), .Z(n1405) );
  AND U1342 ( .A(n254), .B(n1418), .Z(n1420) );
  XNOR U1343 ( .A(n1419), .B(n1416), .Z(n1418) );
  XOR U1344 ( .A(n1421), .B(n1422), .Z(n1416) );
  AND U1345 ( .A(n257), .B(n1415), .Z(n1422) );
  XNOR U1346 ( .A(n1423), .B(n1413), .Z(n1415) );
  XOR U1347 ( .A(n1424), .B(n1425), .Z(n1413) );
  AND U1348 ( .A(n261), .B(n1426), .Z(n1425) );
  XOR U1349 ( .A(p_input[163]), .B(n1424), .Z(n1426) );
  XOR U1350 ( .A(n1427), .B(n1428), .Z(n1424) );
  AND U1351 ( .A(n265), .B(n1429), .Z(n1428) );
  IV U1352 ( .A(n1421), .Z(n1423) );
  XOR U1353 ( .A(n1430), .B(n1431), .Z(n1421) );
  AND U1354 ( .A(n269), .B(n1432), .Z(n1431) );
  XOR U1355 ( .A(n1433), .B(n1434), .Z(n1419) );
  AND U1356 ( .A(n273), .B(n1432), .Z(n1434) );
  XNOR U1357 ( .A(n1433), .B(n1430), .Z(n1432) );
  XOR U1358 ( .A(n1435), .B(n1436), .Z(n1430) );
  AND U1359 ( .A(n276), .B(n1429), .Z(n1436) );
  XNOR U1360 ( .A(n1437), .B(n1427), .Z(n1429) );
  XOR U1361 ( .A(n1438), .B(n1439), .Z(n1427) );
  AND U1362 ( .A(n280), .B(n1440), .Z(n1439) );
  XOR U1363 ( .A(p_input[179]), .B(n1438), .Z(n1440) );
  XOR U1364 ( .A(n1441), .B(n1442), .Z(n1438) );
  AND U1365 ( .A(n284), .B(n1443), .Z(n1442) );
  IV U1366 ( .A(n1435), .Z(n1437) );
  XOR U1367 ( .A(n1444), .B(n1445), .Z(n1435) );
  AND U1368 ( .A(n288), .B(n1446), .Z(n1445) );
  XOR U1369 ( .A(n1447), .B(n1448), .Z(n1433) );
  AND U1370 ( .A(n292), .B(n1446), .Z(n1448) );
  XNOR U1371 ( .A(n1447), .B(n1444), .Z(n1446) );
  XOR U1372 ( .A(n1449), .B(n1450), .Z(n1444) );
  AND U1373 ( .A(n295), .B(n1443), .Z(n1450) );
  XNOR U1374 ( .A(n1451), .B(n1441), .Z(n1443) );
  XOR U1375 ( .A(n1452), .B(n1453), .Z(n1441) );
  AND U1376 ( .A(n299), .B(n1454), .Z(n1453) );
  XOR U1377 ( .A(p_input[195]), .B(n1452), .Z(n1454) );
  XOR U1378 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n1455), 
        .Z(n1452) );
  AND U1379 ( .A(n302), .B(n1456), .Z(n1455) );
  IV U1380 ( .A(n1449), .Z(n1451) );
  XOR U1381 ( .A(n1457), .B(n1458), .Z(n1449) );
  AND U1382 ( .A(n306), .B(n1459), .Z(n1458) );
  XOR U1383 ( .A(n1460), .B(n1461), .Z(n1447) );
  AND U1384 ( .A(n310), .B(n1459), .Z(n1461) );
  XNOR U1385 ( .A(n1460), .B(n1457), .Z(n1459) );
  XNOR U1386 ( .A(n1462), .B(n1463), .Z(n1457) );
  AND U1387 ( .A(n313), .B(n1456), .Z(n1463) );
  XNOR U1388 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n1462), 
        .Z(n1456) );
  XNOR U1389 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .B(n1464), 
        .Z(n1462) );
  AND U1390 ( .A(n315), .B(n1465), .Z(n1464) );
  XNOR U1391 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n1466), .Z(n1460) );
  AND U1392 ( .A(n318), .B(n1465), .Z(n1466) );
  XOR U1393 ( .A(n1467), .B(n1468), .Z(n1465) );
  XOR U1394 ( .A(n51), .B(n1469), .Z(o[18]) );
  AND U1395 ( .A(n62), .B(n1470), .Z(n51) );
  XOR U1396 ( .A(n52), .B(n1469), .Z(n1470) );
  XOR U1397 ( .A(n1471), .B(n41), .Z(n1469) );
  AND U1398 ( .A(n65), .B(n1472), .Z(n41) );
  XOR U1399 ( .A(n42), .B(n1471), .Z(n1472) );
  XOR U1400 ( .A(n1473), .B(n1474), .Z(n42) );
  AND U1401 ( .A(n70), .B(n1475), .Z(n1474) );
  XOR U1402 ( .A(p_input[2]), .B(n1473), .Z(n1475) );
  XNOR U1403 ( .A(n1476), .B(n1477), .Z(n1473) );
  AND U1404 ( .A(n74), .B(n1478), .Z(n1477) );
  XOR U1405 ( .A(n1479), .B(n1480), .Z(n1471) );
  AND U1406 ( .A(n78), .B(n1481), .Z(n1480) );
  XOR U1407 ( .A(n1482), .B(n1483), .Z(n52) );
  AND U1408 ( .A(n82), .B(n1481), .Z(n1483) );
  XNOR U1409 ( .A(n1484), .B(n1482), .Z(n1481) );
  IV U1410 ( .A(n1479), .Z(n1484) );
  XOR U1411 ( .A(n1485), .B(n1486), .Z(n1479) );
  AND U1412 ( .A(n86), .B(n1478), .Z(n1486) );
  XNOR U1413 ( .A(n1476), .B(n1485), .Z(n1478) );
  XNOR U1414 ( .A(n1487), .B(n1488), .Z(n1476) );
  AND U1415 ( .A(n90), .B(n1489), .Z(n1488) );
  XOR U1416 ( .A(p_input[18]), .B(n1487), .Z(n1489) );
  XNOR U1417 ( .A(n1490), .B(n1491), .Z(n1487) );
  AND U1418 ( .A(n94), .B(n1492), .Z(n1491) );
  XOR U1419 ( .A(n1493), .B(n1494), .Z(n1485) );
  AND U1420 ( .A(n98), .B(n1495), .Z(n1494) );
  XOR U1421 ( .A(n1496), .B(n1497), .Z(n1482) );
  AND U1422 ( .A(n102), .B(n1495), .Z(n1497) );
  XNOR U1423 ( .A(n1498), .B(n1496), .Z(n1495) );
  IV U1424 ( .A(n1493), .Z(n1498) );
  XOR U1425 ( .A(n1499), .B(n1500), .Z(n1493) );
  AND U1426 ( .A(n105), .B(n1492), .Z(n1500) );
  XNOR U1427 ( .A(n1490), .B(n1499), .Z(n1492) );
  XNOR U1428 ( .A(n1501), .B(n1502), .Z(n1490) );
  AND U1429 ( .A(n109), .B(n1503), .Z(n1502) );
  XOR U1430 ( .A(p_input[34]), .B(n1501), .Z(n1503) );
  XNOR U1431 ( .A(n1504), .B(n1505), .Z(n1501) );
  AND U1432 ( .A(n113), .B(n1506), .Z(n1505) );
  XOR U1433 ( .A(n1507), .B(n1508), .Z(n1499) );
  AND U1434 ( .A(n117), .B(n1509), .Z(n1508) );
  XOR U1435 ( .A(n1510), .B(n1511), .Z(n1496) );
  AND U1436 ( .A(n121), .B(n1509), .Z(n1511) );
  XNOR U1437 ( .A(n1512), .B(n1510), .Z(n1509) );
  IV U1438 ( .A(n1507), .Z(n1512) );
  XOR U1439 ( .A(n1513), .B(n1514), .Z(n1507) );
  AND U1440 ( .A(n124), .B(n1506), .Z(n1514) );
  XNOR U1441 ( .A(n1504), .B(n1513), .Z(n1506) );
  XNOR U1442 ( .A(n1515), .B(n1516), .Z(n1504) );
  AND U1443 ( .A(n128), .B(n1517), .Z(n1516) );
  XOR U1444 ( .A(p_input[50]), .B(n1515), .Z(n1517) );
  XNOR U1445 ( .A(n1518), .B(n1519), .Z(n1515) );
  AND U1446 ( .A(n132), .B(n1520), .Z(n1519) );
  XOR U1447 ( .A(n1521), .B(n1522), .Z(n1513) );
  AND U1448 ( .A(n136), .B(n1523), .Z(n1522) );
  XOR U1449 ( .A(n1524), .B(n1525), .Z(n1510) );
  AND U1450 ( .A(n140), .B(n1523), .Z(n1525) );
  XNOR U1451 ( .A(n1526), .B(n1524), .Z(n1523) );
  IV U1452 ( .A(n1521), .Z(n1526) );
  XOR U1453 ( .A(n1527), .B(n1528), .Z(n1521) );
  AND U1454 ( .A(n143), .B(n1520), .Z(n1528) );
  XNOR U1455 ( .A(n1518), .B(n1527), .Z(n1520) );
  XNOR U1456 ( .A(n1529), .B(n1530), .Z(n1518) );
  AND U1457 ( .A(n147), .B(n1531), .Z(n1530) );
  XOR U1458 ( .A(p_input[66]), .B(n1529), .Z(n1531) );
  XNOR U1459 ( .A(n1532), .B(n1533), .Z(n1529) );
  AND U1460 ( .A(n151), .B(n1534), .Z(n1533) );
  XOR U1461 ( .A(n1535), .B(n1536), .Z(n1527) );
  AND U1462 ( .A(n155), .B(n1537), .Z(n1536) );
  XOR U1463 ( .A(n1538), .B(n1539), .Z(n1524) );
  AND U1464 ( .A(n159), .B(n1537), .Z(n1539) );
  XNOR U1465 ( .A(n1540), .B(n1538), .Z(n1537) );
  IV U1466 ( .A(n1535), .Z(n1540) );
  XOR U1467 ( .A(n1541), .B(n1542), .Z(n1535) );
  AND U1468 ( .A(n162), .B(n1534), .Z(n1542) );
  XNOR U1469 ( .A(n1532), .B(n1541), .Z(n1534) );
  XNOR U1470 ( .A(n1543), .B(n1544), .Z(n1532) );
  AND U1471 ( .A(n166), .B(n1545), .Z(n1544) );
  XOR U1472 ( .A(p_input[82]), .B(n1543), .Z(n1545) );
  XNOR U1473 ( .A(n1546), .B(n1547), .Z(n1543) );
  AND U1474 ( .A(n170), .B(n1548), .Z(n1547) );
  XOR U1475 ( .A(n1549), .B(n1550), .Z(n1541) );
  AND U1476 ( .A(n174), .B(n1551), .Z(n1550) );
  XOR U1477 ( .A(n1552), .B(n1553), .Z(n1538) );
  AND U1478 ( .A(n178), .B(n1551), .Z(n1553) );
  XNOR U1479 ( .A(n1554), .B(n1552), .Z(n1551) );
  IV U1480 ( .A(n1549), .Z(n1554) );
  XOR U1481 ( .A(n1555), .B(n1556), .Z(n1549) );
  AND U1482 ( .A(n181), .B(n1548), .Z(n1556) );
  XNOR U1483 ( .A(n1546), .B(n1555), .Z(n1548) );
  XNOR U1484 ( .A(n1557), .B(n1558), .Z(n1546) );
  AND U1485 ( .A(n185), .B(n1559), .Z(n1558) );
  XOR U1486 ( .A(p_input[98]), .B(n1557), .Z(n1559) );
  XNOR U1487 ( .A(n1560), .B(n1561), .Z(n1557) );
  AND U1488 ( .A(n189), .B(n1562), .Z(n1561) );
  XOR U1489 ( .A(n1563), .B(n1564), .Z(n1555) );
  AND U1490 ( .A(n193), .B(n1565), .Z(n1564) );
  XOR U1491 ( .A(n1566), .B(n1567), .Z(n1552) );
  AND U1492 ( .A(n197), .B(n1565), .Z(n1567) );
  XNOR U1493 ( .A(n1568), .B(n1566), .Z(n1565) );
  IV U1494 ( .A(n1563), .Z(n1568) );
  XOR U1495 ( .A(n1569), .B(n1570), .Z(n1563) );
  AND U1496 ( .A(n200), .B(n1562), .Z(n1570) );
  XNOR U1497 ( .A(n1560), .B(n1569), .Z(n1562) );
  XNOR U1498 ( .A(n1571), .B(n1572), .Z(n1560) );
  AND U1499 ( .A(n204), .B(n1573), .Z(n1572) );
  XOR U1500 ( .A(p_input[114]), .B(n1571), .Z(n1573) );
  XNOR U1501 ( .A(n1574), .B(n1575), .Z(n1571) );
  AND U1502 ( .A(n208), .B(n1576), .Z(n1575) );
  XOR U1503 ( .A(n1577), .B(n1578), .Z(n1569) );
  AND U1504 ( .A(n212), .B(n1579), .Z(n1578) );
  XOR U1505 ( .A(n1580), .B(n1581), .Z(n1566) );
  AND U1506 ( .A(n216), .B(n1579), .Z(n1581) );
  XNOR U1507 ( .A(n1582), .B(n1580), .Z(n1579) );
  IV U1508 ( .A(n1577), .Z(n1582) );
  XOR U1509 ( .A(n1583), .B(n1584), .Z(n1577) );
  AND U1510 ( .A(n219), .B(n1576), .Z(n1584) );
  XNOR U1511 ( .A(n1574), .B(n1583), .Z(n1576) );
  XNOR U1512 ( .A(n1585), .B(n1586), .Z(n1574) );
  AND U1513 ( .A(n223), .B(n1587), .Z(n1586) );
  XOR U1514 ( .A(p_input[130]), .B(n1585), .Z(n1587) );
  XNOR U1515 ( .A(n1588), .B(n1589), .Z(n1585) );
  AND U1516 ( .A(n227), .B(n1590), .Z(n1589) );
  XOR U1517 ( .A(n1591), .B(n1592), .Z(n1583) );
  AND U1518 ( .A(n231), .B(n1593), .Z(n1592) );
  XOR U1519 ( .A(n1594), .B(n1595), .Z(n1580) );
  AND U1520 ( .A(n235), .B(n1593), .Z(n1595) );
  XNOR U1521 ( .A(n1596), .B(n1594), .Z(n1593) );
  IV U1522 ( .A(n1591), .Z(n1596) );
  XOR U1523 ( .A(n1597), .B(n1598), .Z(n1591) );
  AND U1524 ( .A(n238), .B(n1590), .Z(n1598) );
  XNOR U1525 ( .A(n1588), .B(n1597), .Z(n1590) );
  XNOR U1526 ( .A(n1599), .B(n1600), .Z(n1588) );
  AND U1527 ( .A(n242), .B(n1601), .Z(n1600) );
  XOR U1528 ( .A(p_input[146]), .B(n1599), .Z(n1601) );
  XNOR U1529 ( .A(n1602), .B(n1603), .Z(n1599) );
  AND U1530 ( .A(n246), .B(n1604), .Z(n1603) );
  XOR U1531 ( .A(n1605), .B(n1606), .Z(n1597) );
  AND U1532 ( .A(n250), .B(n1607), .Z(n1606) );
  XOR U1533 ( .A(n1608), .B(n1609), .Z(n1594) );
  AND U1534 ( .A(n254), .B(n1607), .Z(n1609) );
  XNOR U1535 ( .A(n1610), .B(n1608), .Z(n1607) );
  IV U1536 ( .A(n1605), .Z(n1610) );
  XOR U1537 ( .A(n1611), .B(n1612), .Z(n1605) );
  AND U1538 ( .A(n257), .B(n1604), .Z(n1612) );
  XNOR U1539 ( .A(n1602), .B(n1611), .Z(n1604) );
  XNOR U1540 ( .A(n1613), .B(n1614), .Z(n1602) );
  AND U1541 ( .A(n261), .B(n1615), .Z(n1614) );
  XOR U1542 ( .A(p_input[162]), .B(n1613), .Z(n1615) );
  XNOR U1543 ( .A(n1616), .B(n1617), .Z(n1613) );
  AND U1544 ( .A(n265), .B(n1618), .Z(n1617) );
  XOR U1545 ( .A(n1619), .B(n1620), .Z(n1611) );
  AND U1546 ( .A(n269), .B(n1621), .Z(n1620) );
  XOR U1547 ( .A(n1622), .B(n1623), .Z(n1608) );
  AND U1548 ( .A(n273), .B(n1621), .Z(n1623) );
  XNOR U1549 ( .A(n1624), .B(n1622), .Z(n1621) );
  IV U1550 ( .A(n1619), .Z(n1624) );
  XOR U1551 ( .A(n1625), .B(n1626), .Z(n1619) );
  AND U1552 ( .A(n276), .B(n1618), .Z(n1626) );
  XNOR U1553 ( .A(n1616), .B(n1625), .Z(n1618) );
  XNOR U1554 ( .A(n1627), .B(n1628), .Z(n1616) );
  AND U1555 ( .A(n280), .B(n1629), .Z(n1628) );
  XOR U1556 ( .A(p_input[178]), .B(n1627), .Z(n1629) );
  XNOR U1557 ( .A(n1630), .B(n1631), .Z(n1627) );
  AND U1558 ( .A(n284), .B(n1632), .Z(n1631) );
  XOR U1559 ( .A(n1633), .B(n1634), .Z(n1625) );
  AND U1560 ( .A(n288), .B(n1635), .Z(n1634) );
  XOR U1561 ( .A(n1636), .B(n1637), .Z(n1622) );
  AND U1562 ( .A(n292), .B(n1635), .Z(n1637) );
  XNOR U1563 ( .A(n1638), .B(n1636), .Z(n1635) );
  IV U1564 ( .A(n1633), .Z(n1638) );
  XOR U1565 ( .A(n1639), .B(n1640), .Z(n1633) );
  AND U1566 ( .A(n295), .B(n1632), .Z(n1640) );
  XNOR U1567 ( .A(n1630), .B(n1639), .Z(n1632) );
  XNOR U1568 ( .A(n1641), .B(n1642), .Z(n1630) );
  AND U1569 ( .A(n299), .B(n1643), .Z(n1642) );
  XOR U1570 ( .A(p_input[194]), .B(n1641), .Z(n1643) );
  XOR U1571 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n1644), 
        .Z(n1641) );
  AND U1572 ( .A(n302), .B(n1645), .Z(n1644) );
  XOR U1573 ( .A(n1646), .B(n1647), .Z(n1639) );
  AND U1574 ( .A(n306), .B(n1648), .Z(n1647) );
  XOR U1575 ( .A(n1649), .B(n1650), .Z(n1636) );
  AND U1576 ( .A(n310), .B(n1648), .Z(n1650) );
  XNOR U1577 ( .A(n1651), .B(n1649), .Z(n1648) );
  IV U1578 ( .A(n1646), .Z(n1651) );
  XOR U1579 ( .A(n1652), .B(n1653), .Z(n1646) );
  AND U1580 ( .A(n313), .B(n1645), .Z(n1653) );
  XOR U1581 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n1652), 
        .Z(n1645) );
  XOR U1582 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .B(n1654), 
        .Z(n1652) );
  AND U1583 ( .A(n315), .B(n1655), .Z(n1654) );
  XOR U1584 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n1656), .Z(n1649) );
  AND U1585 ( .A(n318), .B(n1655), .Z(n1656) );
  XOR U1586 ( .A(\knn_comb_/min_val_out[0][2] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n1655) );
  XOR U1587 ( .A(n1276), .B(n1657), .Z(o[17]) );
  AND U1588 ( .A(n62), .B(n1658), .Z(n1276) );
  XOR U1589 ( .A(n1277), .B(n1657), .Z(n1658) );
  XOR U1590 ( .A(n1659), .B(n43), .Z(n1657) );
  AND U1591 ( .A(n65), .B(n1660), .Z(n43) );
  XOR U1592 ( .A(n44), .B(n1659), .Z(n1660) );
  XOR U1593 ( .A(n1661), .B(n1662), .Z(n44) );
  AND U1594 ( .A(n70), .B(n1663), .Z(n1662) );
  XOR U1595 ( .A(p_input[1]), .B(n1661), .Z(n1663) );
  XNOR U1596 ( .A(n1664), .B(n1665), .Z(n1661) );
  AND U1597 ( .A(n74), .B(n1666), .Z(n1665) );
  XOR U1598 ( .A(n1667), .B(n1668), .Z(n1659) );
  AND U1599 ( .A(n78), .B(n1669), .Z(n1668) );
  XOR U1600 ( .A(n1670), .B(n1671), .Z(n1277) );
  AND U1601 ( .A(n82), .B(n1669), .Z(n1671) );
  XNOR U1602 ( .A(n1672), .B(n1670), .Z(n1669) );
  IV U1603 ( .A(n1667), .Z(n1672) );
  XOR U1604 ( .A(n1673), .B(n1674), .Z(n1667) );
  AND U1605 ( .A(n86), .B(n1666), .Z(n1674) );
  XNOR U1606 ( .A(n1664), .B(n1673), .Z(n1666) );
  XNOR U1607 ( .A(n1675), .B(n1676), .Z(n1664) );
  AND U1608 ( .A(n90), .B(n1677), .Z(n1676) );
  XOR U1609 ( .A(p_input[17]), .B(n1675), .Z(n1677) );
  XNOR U1610 ( .A(n1678), .B(n1679), .Z(n1675) );
  AND U1611 ( .A(n94), .B(n1680), .Z(n1679) );
  XOR U1612 ( .A(n1681), .B(n1682), .Z(n1673) );
  AND U1613 ( .A(n98), .B(n1683), .Z(n1682) );
  XOR U1614 ( .A(n1684), .B(n1685), .Z(n1670) );
  AND U1615 ( .A(n102), .B(n1683), .Z(n1685) );
  XNOR U1616 ( .A(n1686), .B(n1684), .Z(n1683) );
  IV U1617 ( .A(n1681), .Z(n1686) );
  XOR U1618 ( .A(n1687), .B(n1688), .Z(n1681) );
  AND U1619 ( .A(n105), .B(n1680), .Z(n1688) );
  XNOR U1620 ( .A(n1678), .B(n1687), .Z(n1680) );
  XNOR U1621 ( .A(n1689), .B(n1690), .Z(n1678) );
  AND U1622 ( .A(n109), .B(n1691), .Z(n1690) );
  XOR U1623 ( .A(p_input[33]), .B(n1689), .Z(n1691) );
  XNOR U1624 ( .A(n1692), .B(n1693), .Z(n1689) );
  AND U1625 ( .A(n113), .B(n1694), .Z(n1693) );
  XOR U1626 ( .A(n1695), .B(n1696), .Z(n1687) );
  AND U1627 ( .A(n117), .B(n1697), .Z(n1696) );
  XOR U1628 ( .A(n1698), .B(n1699), .Z(n1684) );
  AND U1629 ( .A(n121), .B(n1697), .Z(n1699) );
  XNOR U1630 ( .A(n1700), .B(n1698), .Z(n1697) );
  IV U1631 ( .A(n1695), .Z(n1700) );
  XOR U1632 ( .A(n1701), .B(n1702), .Z(n1695) );
  AND U1633 ( .A(n124), .B(n1694), .Z(n1702) );
  XNOR U1634 ( .A(n1692), .B(n1701), .Z(n1694) );
  XNOR U1635 ( .A(n1703), .B(n1704), .Z(n1692) );
  AND U1636 ( .A(n128), .B(n1705), .Z(n1704) );
  XOR U1637 ( .A(p_input[49]), .B(n1703), .Z(n1705) );
  XNOR U1638 ( .A(n1706), .B(n1707), .Z(n1703) );
  AND U1639 ( .A(n132), .B(n1708), .Z(n1707) );
  XOR U1640 ( .A(n1709), .B(n1710), .Z(n1701) );
  AND U1641 ( .A(n136), .B(n1711), .Z(n1710) );
  XOR U1642 ( .A(n1712), .B(n1713), .Z(n1698) );
  AND U1643 ( .A(n140), .B(n1711), .Z(n1713) );
  XNOR U1644 ( .A(n1714), .B(n1712), .Z(n1711) );
  IV U1645 ( .A(n1709), .Z(n1714) );
  XOR U1646 ( .A(n1715), .B(n1716), .Z(n1709) );
  AND U1647 ( .A(n143), .B(n1708), .Z(n1716) );
  XNOR U1648 ( .A(n1706), .B(n1715), .Z(n1708) );
  XNOR U1649 ( .A(n1717), .B(n1718), .Z(n1706) );
  AND U1650 ( .A(n147), .B(n1719), .Z(n1718) );
  XOR U1651 ( .A(p_input[65]), .B(n1717), .Z(n1719) );
  XNOR U1652 ( .A(n1720), .B(n1721), .Z(n1717) );
  AND U1653 ( .A(n151), .B(n1722), .Z(n1721) );
  XOR U1654 ( .A(n1723), .B(n1724), .Z(n1715) );
  AND U1655 ( .A(n155), .B(n1725), .Z(n1724) );
  XOR U1656 ( .A(n1726), .B(n1727), .Z(n1712) );
  AND U1657 ( .A(n159), .B(n1725), .Z(n1727) );
  XNOR U1658 ( .A(n1728), .B(n1726), .Z(n1725) );
  IV U1659 ( .A(n1723), .Z(n1728) );
  XOR U1660 ( .A(n1729), .B(n1730), .Z(n1723) );
  AND U1661 ( .A(n162), .B(n1722), .Z(n1730) );
  XNOR U1662 ( .A(n1720), .B(n1729), .Z(n1722) );
  XNOR U1663 ( .A(n1731), .B(n1732), .Z(n1720) );
  AND U1664 ( .A(n166), .B(n1733), .Z(n1732) );
  XOR U1665 ( .A(p_input[81]), .B(n1731), .Z(n1733) );
  XNOR U1666 ( .A(n1734), .B(n1735), .Z(n1731) );
  AND U1667 ( .A(n170), .B(n1736), .Z(n1735) );
  XOR U1668 ( .A(n1737), .B(n1738), .Z(n1729) );
  AND U1669 ( .A(n174), .B(n1739), .Z(n1738) );
  XOR U1670 ( .A(n1740), .B(n1741), .Z(n1726) );
  AND U1671 ( .A(n178), .B(n1739), .Z(n1741) );
  XNOR U1672 ( .A(n1742), .B(n1740), .Z(n1739) );
  IV U1673 ( .A(n1737), .Z(n1742) );
  XOR U1674 ( .A(n1743), .B(n1744), .Z(n1737) );
  AND U1675 ( .A(n181), .B(n1736), .Z(n1744) );
  XNOR U1676 ( .A(n1734), .B(n1743), .Z(n1736) );
  XNOR U1677 ( .A(n1745), .B(n1746), .Z(n1734) );
  AND U1678 ( .A(n185), .B(n1747), .Z(n1746) );
  XOR U1679 ( .A(p_input[97]), .B(n1745), .Z(n1747) );
  XNOR U1680 ( .A(n1748), .B(n1749), .Z(n1745) );
  AND U1681 ( .A(n189), .B(n1750), .Z(n1749) );
  XOR U1682 ( .A(n1751), .B(n1752), .Z(n1743) );
  AND U1683 ( .A(n193), .B(n1753), .Z(n1752) );
  XOR U1684 ( .A(n1754), .B(n1755), .Z(n1740) );
  AND U1685 ( .A(n197), .B(n1753), .Z(n1755) );
  XNOR U1686 ( .A(n1756), .B(n1754), .Z(n1753) );
  IV U1687 ( .A(n1751), .Z(n1756) );
  XOR U1688 ( .A(n1757), .B(n1758), .Z(n1751) );
  AND U1689 ( .A(n200), .B(n1750), .Z(n1758) );
  XNOR U1690 ( .A(n1748), .B(n1757), .Z(n1750) );
  XNOR U1691 ( .A(n1759), .B(n1760), .Z(n1748) );
  AND U1692 ( .A(n204), .B(n1761), .Z(n1760) );
  XOR U1693 ( .A(p_input[113]), .B(n1759), .Z(n1761) );
  XNOR U1694 ( .A(n1762), .B(n1763), .Z(n1759) );
  AND U1695 ( .A(n208), .B(n1764), .Z(n1763) );
  XOR U1696 ( .A(n1765), .B(n1766), .Z(n1757) );
  AND U1697 ( .A(n212), .B(n1767), .Z(n1766) );
  XOR U1698 ( .A(n1768), .B(n1769), .Z(n1754) );
  AND U1699 ( .A(n216), .B(n1767), .Z(n1769) );
  XNOR U1700 ( .A(n1770), .B(n1768), .Z(n1767) );
  IV U1701 ( .A(n1765), .Z(n1770) );
  XOR U1702 ( .A(n1771), .B(n1772), .Z(n1765) );
  AND U1703 ( .A(n219), .B(n1764), .Z(n1772) );
  XNOR U1704 ( .A(n1762), .B(n1771), .Z(n1764) );
  XNOR U1705 ( .A(n1773), .B(n1774), .Z(n1762) );
  AND U1706 ( .A(n223), .B(n1775), .Z(n1774) );
  XOR U1707 ( .A(p_input[129]), .B(n1773), .Z(n1775) );
  XNOR U1708 ( .A(n1776), .B(n1777), .Z(n1773) );
  AND U1709 ( .A(n227), .B(n1778), .Z(n1777) );
  XOR U1710 ( .A(n1779), .B(n1780), .Z(n1771) );
  AND U1711 ( .A(n231), .B(n1781), .Z(n1780) );
  XOR U1712 ( .A(n1782), .B(n1783), .Z(n1768) );
  AND U1713 ( .A(n235), .B(n1781), .Z(n1783) );
  XNOR U1714 ( .A(n1784), .B(n1782), .Z(n1781) );
  IV U1715 ( .A(n1779), .Z(n1784) );
  XOR U1716 ( .A(n1785), .B(n1786), .Z(n1779) );
  AND U1717 ( .A(n238), .B(n1778), .Z(n1786) );
  XNOR U1718 ( .A(n1776), .B(n1785), .Z(n1778) );
  XNOR U1719 ( .A(n1787), .B(n1788), .Z(n1776) );
  AND U1720 ( .A(n242), .B(n1789), .Z(n1788) );
  XOR U1721 ( .A(p_input[145]), .B(n1787), .Z(n1789) );
  XNOR U1722 ( .A(n1790), .B(n1791), .Z(n1787) );
  AND U1723 ( .A(n246), .B(n1792), .Z(n1791) );
  XOR U1724 ( .A(n1793), .B(n1794), .Z(n1785) );
  AND U1725 ( .A(n250), .B(n1795), .Z(n1794) );
  XOR U1726 ( .A(n1796), .B(n1797), .Z(n1782) );
  AND U1727 ( .A(n254), .B(n1795), .Z(n1797) );
  XNOR U1728 ( .A(n1798), .B(n1796), .Z(n1795) );
  IV U1729 ( .A(n1793), .Z(n1798) );
  XOR U1730 ( .A(n1799), .B(n1800), .Z(n1793) );
  AND U1731 ( .A(n257), .B(n1792), .Z(n1800) );
  XNOR U1732 ( .A(n1790), .B(n1799), .Z(n1792) );
  XNOR U1733 ( .A(n1801), .B(n1802), .Z(n1790) );
  AND U1734 ( .A(n261), .B(n1803), .Z(n1802) );
  XOR U1735 ( .A(p_input[161]), .B(n1801), .Z(n1803) );
  XNOR U1736 ( .A(n1804), .B(n1805), .Z(n1801) );
  AND U1737 ( .A(n265), .B(n1806), .Z(n1805) );
  XOR U1738 ( .A(n1807), .B(n1808), .Z(n1799) );
  AND U1739 ( .A(n269), .B(n1809), .Z(n1808) );
  XOR U1740 ( .A(n1810), .B(n1811), .Z(n1796) );
  AND U1741 ( .A(n273), .B(n1809), .Z(n1811) );
  XNOR U1742 ( .A(n1812), .B(n1810), .Z(n1809) );
  IV U1743 ( .A(n1807), .Z(n1812) );
  XOR U1744 ( .A(n1813), .B(n1814), .Z(n1807) );
  AND U1745 ( .A(n276), .B(n1806), .Z(n1814) );
  XNOR U1746 ( .A(n1804), .B(n1813), .Z(n1806) );
  XNOR U1747 ( .A(n1815), .B(n1816), .Z(n1804) );
  AND U1748 ( .A(n280), .B(n1817), .Z(n1816) );
  XOR U1749 ( .A(p_input[177]), .B(n1815), .Z(n1817) );
  XNOR U1750 ( .A(n1818), .B(n1819), .Z(n1815) );
  AND U1751 ( .A(n284), .B(n1820), .Z(n1819) );
  XOR U1752 ( .A(n1821), .B(n1822), .Z(n1813) );
  AND U1753 ( .A(n288), .B(n1823), .Z(n1822) );
  XOR U1754 ( .A(n1824), .B(n1825), .Z(n1810) );
  AND U1755 ( .A(n292), .B(n1823), .Z(n1825) );
  XNOR U1756 ( .A(n1826), .B(n1824), .Z(n1823) );
  IV U1757 ( .A(n1821), .Z(n1826) );
  XOR U1758 ( .A(n1827), .B(n1828), .Z(n1821) );
  AND U1759 ( .A(n295), .B(n1820), .Z(n1828) );
  XNOR U1760 ( .A(n1818), .B(n1827), .Z(n1820) );
  XNOR U1761 ( .A(n1829), .B(n1830), .Z(n1818) );
  AND U1762 ( .A(n299), .B(n1831), .Z(n1830) );
  XOR U1763 ( .A(p_input[193]), .B(n1829), .Z(n1831) );
  XOR U1764 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n1832), 
        .Z(n1829) );
  AND U1765 ( .A(n302), .B(n1833), .Z(n1832) );
  XOR U1766 ( .A(n1834), .B(n1835), .Z(n1827) );
  AND U1767 ( .A(n306), .B(n1836), .Z(n1835) );
  XOR U1768 ( .A(n1837), .B(n1838), .Z(n1824) );
  AND U1769 ( .A(n310), .B(n1836), .Z(n1838) );
  XNOR U1770 ( .A(n1839), .B(n1837), .Z(n1836) );
  IV U1771 ( .A(n1834), .Z(n1839) );
  XOR U1772 ( .A(n1840), .B(n1841), .Z(n1834) );
  AND U1773 ( .A(n313), .B(n1833), .Z(n1841) );
  XOR U1774 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n1840), 
        .Z(n1833) );
  XOR U1775 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(n1842), 
        .Z(n1840) );
  AND U1776 ( .A(n315), .B(n1843), .Z(n1842) );
  XOR U1777 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n1844), .Z(n1837) );
  AND U1778 ( .A(n318), .B(n1843), .Z(n1844) );
  XOR U1779 ( .A(\knn_comb_/min_val_out[0][1] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n1843) );
  XOR U1780 ( .A(n1845), .B(n1846), .Z(o[16]) );
  XOR U1781 ( .A(n47), .B(n1847), .Z(o[15]) );
  AND U1782 ( .A(n62), .B(n1848), .Z(n47) );
  XOR U1783 ( .A(n48), .B(n1847), .Z(n1848) );
  XOR U1784 ( .A(n1849), .B(n1850), .Z(n1847) );
  AND U1785 ( .A(n82), .B(n1851), .Z(n1850) );
  XOR U1786 ( .A(n1852), .B(n13), .Z(n48) );
  AND U1787 ( .A(n65), .B(n1853), .Z(n13) );
  XOR U1788 ( .A(n14), .B(n1852), .Z(n1853) );
  XOR U1789 ( .A(n1854), .B(n1855), .Z(n14) );
  AND U1790 ( .A(n70), .B(n1856), .Z(n1855) );
  XOR U1791 ( .A(p_input[15]), .B(n1854), .Z(n1856) );
  XNOR U1792 ( .A(n1857), .B(n1858), .Z(n1854) );
  AND U1793 ( .A(n74), .B(n1859), .Z(n1858) );
  XOR U1794 ( .A(n1860), .B(n1861), .Z(n1852) );
  AND U1795 ( .A(n78), .B(n1851), .Z(n1861) );
  XNOR U1796 ( .A(n1862), .B(n1849), .Z(n1851) );
  XOR U1797 ( .A(n1863), .B(n1864), .Z(n1849) );
  AND U1798 ( .A(n102), .B(n1865), .Z(n1864) );
  IV U1799 ( .A(n1860), .Z(n1862) );
  XOR U1800 ( .A(n1866), .B(n1867), .Z(n1860) );
  AND U1801 ( .A(n86), .B(n1859), .Z(n1867) );
  XNOR U1802 ( .A(n1857), .B(n1866), .Z(n1859) );
  XNOR U1803 ( .A(n1868), .B(n1869), .Z(n1857) );
  AND U1804 ( .A(n90), .B(n1870), .Z(n1869) );
  XOR U1805 ( .A(p_input[31]), .B(n1868), .Z(n1870) );
  XNOR U1806 ( .A(n1871), .B(n1872), .Z(n1868) );
  AND U1807 ( .A(n94), .B(n1873), .Z(n1872) );
  XOR U1808 ( .A(n1874), .B(n1875), .Z(n1866) );
  AND U1809 ( .A(n98), .B(n1865), .Z(n1875) );
  XNOR U1810 ( .A(n1876), .B(n1863), .Z(n1865) );
  XOR U1811 ( .A(n1877), .B(n1878), .Z(n1863) );
  AND U1812 ( .A(n121), .B(n1879), .Z(n1878) );
  IV U1813 ( .A(n1874), .Z(n1876) );
  XOR U1814 ( .A(n1880), .B(n1881), .Z(n1874) );
  AND U1815 ( .A(n105), .B(n1873), .Z(n1881) );
  XNOR U1816 ( .A(n1871), .B(n1880), .Z(n1873) );
  XNOR U1817 ( .A(n1882), .B(n1883), .Z(n1871) );
  AND U1818 ( .A(n109), .B(n1884), .Z(n1883) );
  XOR U1819 ( .A(p_input[47]), .B(n1882), .Z(n1884) );
  XNOR U1820 ( .A(n1885), .B(n1886), .Z(n1882) );
  AND U1821 ( .A(n113), .B(n1887), .Z(n1886) );
  XOR U1822 ( .A(n1888), .B(n1889), .Z(n1880) );
  AND U1823 ( .A(n117), .B(n1879), .Z(n1889) );
  XNOR U1824 ( .A(n1890), .B(n1877), .Z(n1879) );
  XOR U1825 ( .A(n1891), .B(n1892), .Z(n1877) );
  AND U1826 ( .A(n140), .B(n1893), .Z(n1892) );
  IV U1827 ( .A(n1888), .Z(n1890) );
  XOR U1828 ( .A(n1894), .B(n1895), .Z(n1888) );
  AND U1829 ( .A(n124), .B(n1887), .Z(n1895) );
  XNOR U1830 ( .A(n1885), .B(n1894), .Z(n1887) );
  XNOR U1831 ( .A(n1896), .B(n1897), .Z(n1885) );
  AND U1832 ( .A(n128), .B(n1898), .Z(n1897) );
  XOR U1833 ( .A(p_input[63]), .B(n1896), .Z(n1898) );
  XNOR U1834 ( .A(n1899), .B(n1900), .Z(n1896) );
  AND U1835 ( .A(n132), .B(n1901), .Z(n1900) );
  XOR U1836 ( .A(n1902), .B(n1903), .Z(n1894) );
  AND U1837 ( .A(n136), .B(n1893), .Z(n1903) );
  XNOR U1838 ( .A(n1904), .B(n1891), .Z(n1893) );
  XOR U1839 ( .A(n1905), .B(n1906), .Z(n1891) );
  AND U1840 ( .A(n159), .B(n1907), .Z(n1906) );
  IV U1841 ( .A(n1902), .Z(n1904) );
  XOR U1842 ( .A(n1908), .B(n1909), .Z(n1902) );
  AND U1843 ( .A(n143), .B(n1901), .Z(n1909) );
  XNOR U1844 ( .A(n1899), .B(n1908), .Z(n1901) );
  XNOR U1845 ( .A(n1910), .B(n1911), .Z(n1899) );
  AND U1846 ( .A(n147), .B(n1912), .Z(n1911) );
  XOR U1847 ( .A(p_input[79]), .B(n1910), .Z(n1912) );
  XNOR U1848 ( .A(n1913), .B(n1914), .Z(n1910) );
  AND U1849 ( .A(n151), .B(n1915), .Z(n1914) );
  XOR U1850 ( .A(n1916), .B(n1917), .Z(n1908) );
  AND U1851 ( .A(n155), .B(n1907), .Z(n1917) );
  XNOR U1852 ( .A(n1918), .B(n1905), .Z(n1907) );
  XOR U1853 ( .A(n1919), .B(n1920), .Z(n1905) );
  AND U1854 ( .A(n178), .B(n1921), .Z(n1920) );
  IV U1855 ( .A(n1916), .Z(n1918) );
  XOR U1856 ( .A(n1922), .B(n1923), .Z(n1916) );
  AND U1857 ( .A(n162), .B(n1915), .Z(n1923) );
  XNOR U1858 ( .A(n1913), .B(n1922), .Z(n1915) );
  XNOR U1859 ( .A(n1924), .B(n1925), .Z(n1913) );
  AND U1860 ( .A(n166), .B(n1926), .Z(n1925) );
  XOR U1861 ( .A(p_input[95]), .B(n1924), .Z(n1926) );
  XNOR U1862 ( .A(n1927), .B(n1928), .Z(n1924) );
  AND U1863 ( .A(n170), .B(n1929), .Z(n1928) );
  XOR U1864 ( .A(n1930), .B(n1931), .Z(n1922) );
  AND U1865 ( .A(n174), .B(n1921), .Z(n1931) );
  XNOR U1866 ( .A(n1932), .B(n1919), .Z(n1921) );
  XOR U1867 ( .A(n1933), .B(n1934), .Z(n1919) );
  AND U1868 ( .A(n197), .B(n1935), .Z(n1934) );
  IV U1869 ( .A(n1930), .Z(n1932) );
  XOR U1870 ( .A(n1936), .B(n1937), .Z(n1930) );
  AND U1871 ( .A(n181), .B(n1929), .Z(n1937) );
  XNOR U1872 ( .A(n1927), .B(n1936), .Z(n1929) );
  XNOR U1873 ( .A(n1938), .B(n1939), .Z(n1927) );
  AND U1874 ( .A(n185), .B(n1940), .Z(n1939) );
  XOR U1875 ( .A(p_input[111]), .B(n1938), .Z(n1940) );
  XNOR U1876 ( .A(n1941), .B(n1942), .Z(n1938) );
  AND U1877 ( .A(n189), .B(n1943), .Z(n1942) );
  XOR U1878 ( .A(n1944), .B(n1945), .Z(n1936) );
  AND U1879 ( .A(n193), .B(n1935), .Z(n1945) );
  XNOR U1880 ( .A(n1946), .B(n1933), .Z(n1935) );
  XOR U1881 ( .A(n1947), .B(n1948), .Z(n1933) );
  AND U1882 ( .A(n216), .B(n1949), .Z(n1948) );
  IV U1883 ( .A(n1944), .Z(n1946) );
  XOR U1884 ( .A(n1950), .B(n1951), .Z(n1944) );
  AND U1885 ( .A(n200), .B(n1943), .Z(n1951) );
  XNOR U1886 ( .A(n1941), .B(n1950), .Z(n1943) );
  XNOR U1887 ( .A(n1952), .B(n1953), .Z(n1941) );
  AND U1888 ( .A(n204), .B(n1954), .Z(n1953) );
  XOR U1889 ( .A(p_input[127]), .B(n1952), .Z(n1954) );
  XNOR U1890 ( .A(n1955), .B(n1956), .Z(n1952) );
  AND U1891 ( .A(n208), .B(n1957), .Z(n1956) );
  XOR U1892 ( .A(n1958), .B(n1959), .Z(n1950) );
  AND U1893 ( .A(n212), .B(n1949), .Z(n1959) );
  XNOR U1894 ( .A(n1960), .B(n1947), .Z(n1949) );
  XOR U1895 ( .A(n1961), .B(n1962), .Z(n1947) );
  AND U1896 ( .A(n235), .B(n1963), .Z(n1962) );
  IV U1897 ( .A(n1958), .Z(n1960) );
  XOR U1898 ( .A(n1964), .B(n1965), .Z(n1958) );
  AND U1899 ( .A(n219), .B(n1957), .Z(n1965) );
  XNOR U1900 ( .A(n1955), .B(n1964), .Z(n1957) );
  XNOR U1901 ( .A(n1966), .B(n1967), .Z(n1955) );
  AND U1902 ( .A(n223), .B(n1968), .Z(n1967) );
  XOR U1903 ( .A(p_input[143]), .B(n1966), .Z(n1968) );
  XNOR U1904 ( .A(n1969), .B(n1970), .Z(n1966) );
  AND U1905 ( .A(n227), .B(n1971), .Z(n1970) );
  XOR U1906 ( .A(n1972), .B(n1973), .Z(n1964) );
  AND U1907 ( .A(n231), .B(n1963), .Z(n1973) );
  XNOR U1908 ( .A(n1974), .B(n1961), .Z(n1963) );
  XOR U1909 ( .A(n1975), .B(n1976), .Z(n1961) );
  AND U1910 ( .A(n254), .B(n1977), .Z(n1976) );
  IV U1911 ( .A(n1972), .Z(n1974) );
  XOR U1912 ( .A(n1978), .B(n1979), .Z(n1972) );
  AND U1913 ( .A(n238), .B(n1971), .Z(n1979) );
  XNOR U1914 ( .A(n1969), .B(n1978), .Z(n1971) );
  XNOR U1915 ( .A(n1980), .B(n1981), .Z(n1969) );
  AND U1916 ( .A(n242), .B(n1982), .Z(n1981) );
  XOR U1917 ( .A(p_input[159]), .B(n1980), .Z(n1982) );
  XNOR U1918 ( .A(n1983), .B(n1984), .Z(n1980) );
  AND U1919 ( .A(n246), .B(n1985), .Z(n1984) );
  XOR U1920 ( .A(n1986), .B(n1987), .Z(n1978) );
  AND U1921 ( .A(n250), .B(n1977), .Z(n1987) );
  XNOR U1922 ( .A(n1988), .B(n1975), .Z(n1977) );
  XOR U1923 ( .A(n1989), .B(n1990), .Z(n1975) );
  AND U1924 ( .A(n273), .B(n1991), .Z(n1990) );
  IV U1925 ( .A(n1986), .Z(n1988) );
  XOR U1926 ( .A(n1992), .B(n1993), .Z(n1986) );
  AND U1927 ( .A(n257), .B(n1985), .Z(n1993) );
  XNOR U1928 ( .A(n1983), .B(n1992), .Z(n1985) );
  XNOR U1929 ( .A(n1994), .B(n1995), .Z(n1983) );
  AND U1930 ( .A(n261), .B(n1996), .Z(n1995) );
  XOR U1931 ( .A(p_input[175]), .B(n1994), .Z(n1996) );
  XNOR U1932 ( .A(n1997), .B(n1998), .Z(n1994) );
  AND U1933 ( .A(n265), .B(n1999), .Z(n1998) );
  XOR U1934 ( .A(n2000), .B(n2001), .Z(n1992) );
  AND U1935 ( .A(n269), .B(n1991), .Z(n2001) );
  XNOR U1936 ( .A(n2002), .B(n1989), .Z(n1991) );
  XOR U1937 ( .A(n2003), .B(n2004), .Z(n1989) );
  AND U1938 ( .A(n292), .B(n2005), .Z(n2004) );
  IV U1939 ( .A(n2000), .Z(n2002) );
  XOR U1940 ( .A(n2006), .B(n2007), .Z(n2000) );
  AND U1941 ( .A(n276), .B(n1999), .Z(n2007) );
  XNOR U1942 ( .A(n1997), .B(n2006), .Z(n1999) );
  XNOR U1943 ( .A(n2008), .B(n2009), .Z(n1997) );
  AND U1944 ( .A(n280), .B(n2010), .Z(n2009) );
  XOR U1945 ( .A(p_input[191]), .B(n2008), .Z(n2010) );
  XNOR U1946 ( .A(n2011), .B(n2012), .Z(n2008) );
  AND U1947 ( .A(n284), .B(n2013), .Z(n2012) );
  XOR U1948 ( .A(n2014), .B(n2015), .Z(n2006) );
  AND U1949 ( .A(n288), .B(n2005), .Z(n2015) );
  XNOR U1950 ( .A(n2016), .B(n2003), .Z(n2005) );
  XOR U1951 ( .A(n2017), .B(n2018), .Z(n2003) );
  AND U1952 ( .A(n310), .B(n2019), .Z(n2018) );
  IV U1953 ( .A(n2014), .Z(n2016) );
  XOR U1954 ( .A(n2020), .B(n2021), .Z(n2014) );
  AND U1955 ( .A(n295), .B(n2013), .Z(n2021) );
  XNOR U1956 ( .A(n2011), .B(n2020), .Z(n2013) );
  XNOR U1957 ( .A(n2022), .B(n2023), .Z(n2011) );
  AND U1958 ( .A(n299), .B(n2024), .Z(n2023) );
  XOR U1959 ( .A(p_input[207]), .B(n2022), .Z(n2024) );
  XOR U1960 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n2025), 
        .Z(n2022) );
  AND U1961 ( .A(n302), .B(n2026), .Z(n2025) );
  XOR U1962 ( .A(n2027), .B(n2028), .Z(n2020) );
  AND U1963 ( .A(n306), .B(n2019), .Z(n2028) );
  XNOR U1964 ( .A(n2029), .B(n2017), .Z(n2019) );
  XOR U1965 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n2030), .Z(n2017) );
  AND U1966 ( .A(n318), .B(n2031), .Z(n2030) );
  IV U1967 ( .A(n2027), .Z(n2029) );
  XOR U1968 ( .A(n2032), .B(n2033), .Z(n2027) );
  AND U1969 ( .A(n313), .B(n2026), .Z(n2033) );
  XOR U1970 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n2032), 
        .Z(n2026) );
  XOR U1971 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(n2034), 
        .Z(n2032) );
  AND U1972 ( .A(n315), .B(n2031), .Z(n2034) );
  XOR U1973 ( .A(n2035), .B(n2036), .Z(n2031) );
  IV U1974 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .Z(n2036) );
  IV U1975 ( .A(\knn_comb_/min_val_out[0][15] ), .Z(n2035) );
  XOR U1976 ( .A(n49), .B(n2037), .Z(o[14]) );
  AND U1977 ( .A(n62), .B(n2038), .Z(n49) );
  XOR U1978 ( .A(n50), .B(n2037), .Z(n2038) );
  XOR U1979 ( .A(n2039), .B(n2040), .Z(n2037) );
  AND U1980 ( .A(n82), .B(n2041), .Z(n2040) );
  XOR U1981 ( .A(n2042), .B(n15), .Z(n50) );
  AND U1982 ( .A(n65), .B(n2043), .Z(n15) );
  XOR U1983 ( .A(n16), .B(n2042), .Z(n2043) );
  XOR U1984 ( .A(n2044), .B(n2045), .Z(n16) );
  AND U1985 ( .A(n70), .B(n2046), .Z(n2045) );
  XOR U1986 ( .A(p_input[14]), .B(n2044), .Z(n2046) );
  XNOR U1987 ( .A(n2047), .B(n2048), .Z(n2044) );
  AND U1988 ( .A(n74), .B(n2049), .Z(n2048) );
  XOR U1989 ( .A(n2050), .B(n2051), .Z(n2042) );
  AND U1990 ( .A(n78), .B(n2041), .Z(n2051) );
  XNOR U1991 ( .A(n2052), .B(n2039), .Z(n2041) );
  XOR U1992 ( .A(n2053), .B(n2054), .Z(n2039) );
  AND U1993 ( .A(n102), .B(n2055), .Z(n2054) );
  IV U1994 ( .A(n2050), .Z(n2052) );
  XOR U1995 ( .A(n2056), .B(n2057), .Z(n2050) );
  AND U1996 ( .A(n86), .B(n2049), .Z(n2057) );
  XNOR U1997 ( .A(n2047), .B(n2056), .Z(n2049) );
  XNOR U1998 ( .A(n2058), .B(n2059), .Z(n2047) );
  AND U1999 ( .A(n90), .B(n2060), .Z(n2059) );
  XOR U2000 ( .A(p_input[30]), .B(n2058), .Z(n2060) );
  XNOR U2001 ( .A(n2061), .B(n2062), .Z(n2058) );
  AND U2002 ( .A(n94), .B(n2063), .Z(n2062) );
  XOR U2003 ( .A(n2064), .B(n2065), .Z(n2056) );
  AND U2004 ( .A(n98), .B(n2055), .Z(n2065) );
  XNOR U2005 ( .A(n2066), .B(n2053), .Z(n2055) );
  XOR U2006 ( .A(n2067), .B(n2068), .Z(n2053) );
  AND U2007 ( .A(n121), .B(n2069), .Z(n2068) );
  IV U2008 ( .A(n2064), .Z(n2066) );
  XOR U2009 ( .A(n2070), .B(n2071), .Z(n2064) );
  AND U2010 ( .A(n105), .B(n2063), .Z(n2071) );
  XNOR U2011 ( .A(n2061), .B(n2070), .Z(n2063) );
  XNOR U2012 ( .A(n2072), .B(n2073), .Z(n2061) );
  AND U2013 ( .A(n109), .B(n2074), .Z(n2073) );
  XOR U2014 ( .A(p_input[46]), .B(n2072), .Z(n2074) );
  XNOR U2015 ( .A(n2075), .B(n2076), .Z(n2072) );
  AND U2016 ( .A(n113), .B(n2077), .Z(n2076) );
  XOR U2017 ( .A(n2078), .B(n2079), .Z(n2070) );
  AND U2018 ( .A(n117), .B(n2069), .Z(n2079) );
  XNOR U2019 ( .A(n2080), .B(n2067), .Z(n2069) );
  XOR U2020 ( .A(n2081), .B(n2082), .Z(n2067) );
  AND U2021 ( .A(n140), .B(n2083), .Z(n2082) );
  IV U2022 ( .A(n2078), .Z(n2080) );
  XOR U2023 ( .A(n2084), .B(n2085), .Z(n2078) );
  AND U2024 ( .A(n124), .B(n2077), .Z(n2085) );
  XNOR U2025 ( .A(n2075), .B(n2084), .Z(n2077) );
  XNOR U2026 ( .A(n2086), .B(n2087), .Z(n2075) );
  AND U2027 ( .A(n128), .B(n2088), .Z(n2087) );
  XOR U2028 ( .A(p_input[62]), .B(n2086), .Z(n2088) );
  XNOR U2029 ( .A(n2089), .B(n2090), .Z(n2086) );
  AND U2030 ( .A(n132), .B(n2091), .Z(n2090) );
  XOR U2031 ( .A(n2092), .B(n2093), .Z(n2084) );
  AND U2032 ( .A(n136), .B(n2083), .Z(n2093) );
  XNOR U2033 ( .A(n2094), .B(n2081), .Z(n2083) );
  XOR U2034 ( .A(n2095), .B(n2096), .Z(n2081) );
  AND U2035 ( .A(n159), .B(n2097), .Z(n2096) );
  IV U2036 ( .A(n2092), .Z(n2094) );
  XOR U2037 ( .A(n2098), .B(n2099), .Z(n2092) );
  AND U2038 ( .A(n143), .B(n2091), .Z(n2099) );
  XNOR U2039 ( .A(n2089), .B(n2098), .Z(n2091) );
  XNOR U2040 ( .A(n2100), .B(n2101), .Z(n2089) );
  AND U2041 ( .A(n147), .B(n2102), .Z(n2101) );
  XOR U2042 ( .A(p_input[78]), .B(n2100), .Z(n2102) );
  XNOR U2043 ( .A(n2103), .B(n2104), .Z(n2100) );
  AND U2044 ( .A(n151), .B(n2105), .Z(n2104) );
  XOR U2045 ( .A(n2106), .B(n2107), .Z(n2098) );
  AND U2046 ( .A(n155), .B(n2097), .Z(n2107) );
  XNOR U2047 ( .A(n2108), .B(n2095), .Z(n2097) );
  XOR U2048 ( .A(n2109), .B(n2110), .Z(n2095) );
  AND U2049 ( .A(n178), .B(n2111), .Z(n2110) );
  IV U2050 ( .A(n2106), .Z(n2108) );
  XOR U2051 ( .A(n2112), .B(n2113), .Z(n2106) );
  AND U2052 ( .A(n162), .B(n2105), .Z(n2113) );
  XNOR U2053 ( .A(n2103), .B(n2112), .Z(n2105) );
  XNOR U2054 ( .A(n2114), .B(n2115), .Z(n2103) );
  AND U2055 ( .A(n166), .B(n2116), .Z(n2115) );
  XOR U2056 ( .A(p_input[94]), .B(n2114), .Z(n2116) );
  XNOR U2057 ( .A(n2117), .B(n2118), .Z(n2114) );
  AND U2058 ( .A(n170), .B(n2119), .Z(n2118) );
  XOR U2059 ( .A(n2120), .B(n2121), .Z(n2112) );
  AND U2060 ( .A(n174), .B(n2111), .Z(n2121) );
  XNOR U2061 ( .A(n2122), .B(n2109), .Z(n2111) );
  XOR U2062 ( .A(n2123), .B(n2124), .Z(n2109) );
  AND U2063 ( .A(n197), .B(n2125), .Z(n2124) );
  IV U2064 ( .A(n2120), .Z(n2122) );
  XOR U2065 ( .A(n2126), .B(n2127), .Z(n2120) );
  AND U2066 ( .A(n181), .B(n2119), .Z(n2127) );
  XNOR U2067 ( .A(n2117), .B(n2126), .Z(n2119) );
  XNOR U2068 ( .A(n2128), .B(n2129), .Z(n2117) );
  AND U2069 ( .A(n185), .B(n2130), .Z(n2129) );
  XOR U2070 ( .A(p_input[110]), .B(n2128), .Z(n2130) );
  XNOR U2071 ( .A(n2131), .B(n2132), .Z(n2128) );
  AND U2072 ( .A(n189), .B(n2133), .Z(n2132) );
  XOR U2073 ( .A(n2134), .B(n2135), .Z(n2126) );
  AND U2074 ( .A(n193), .B(n2125), .Z(n2135) );
  XNOR U2075 ( .A(n2136), .B(n2123), .Z(n2125) );
  XOR U2076 ( .A(n2137), .B(n2138), .Z(n2123) );
  AND U2077 ( .A(n216), .B(n2139), .Z(n2138) );
  IV U2078 ( .A(n2134), .Z(n2136) );
  XOR U2079 ( .A(n2140), .B(n2141), .Z(n2134) );
  AND U2080 ( .A(n200), .B(n2133), .Z(n2141) );
  XNOR U2081 ( .A(n2131), .B(n2140), .Z(n2133) );
  XNOR U2082 ( .A(n2142), .B(n2143), .Z(n2131) );
  AND U2083 ( .A(n204), .B(n2144), .Z(n2143) );
  XOR U2084 ( .A(p_input[126]), .B(n2142), .Z(n2144) );
  XNOR U2085 ( .A(n2145), .B(n2146), .Z(n2142) );
  AND U2086 ( .A(n208), .B(n2147), .Z(n2146) );
  XOR U2087 ( .A(n2148), .B(n2149), .Z(n2140) );
  AND U2088 ( .A(n212), .B(n2139), .Z(n2149) );
  XNOR U2089 ( .A(n2150), .B(n2137), .Z(n2139) );
  XOR U2090 ( .A(n2151), .B(n2152), .Z(n2137) );
  AND U2091 ( .A(n235), .B(n2153), .Z(n2152) );
  IV U2092 ( .A(n2148), .Z(n2150) );
  XOR U2093 ( .A(n2154), .B(n2155), .Z(n2148) );
  AND U2094 ( .A(n219), .B(n2147), .Z(n2155) );
  XNOR U2095 ( .A(n2145), .B(n2154), .Z(n2147) );
  XNOR U2096 ( .A(n2156), .B(n2157), .Z(n2145) );
  AND U2097 ( .A(n223), .B(n2158), .Z(n2157) );
  XOR U2098 ( .A(p_input[142]), .B(n2156), .Z(n2158) );
  XNOR U2099 ( .A(n2159), .B(n2160), .Z(n2156) );
  AND U2100 ( .A(n227), .B(n2161), .Z(n2160) );
  XOR U2101 ( .A(n2162), .B(n2163), .Z(n2154) );
  AND U2102 ( .A(n231), .B(n2153), .Z(n2163) );
  XNOR U2103 ( .A(n2164), .B(n2151), .Z(n2153) );
  XOR U2104 ( .A(n2165), .B(n2166), .Z(n2151) );
  AND U2105 ( .A(n254), .B(n2167), .Z(n2166) );
  IV U2106 ( .A(n2162), .Z(n2164) );
  XOR U2107 ( .A(n2168), .B(n2169), .Z(n2162) );
  AND U2108 ( .A(n238), .B(n2161), .Z(n2169) );
  XNOR U2109 ( .A(n2159), .B(n2168), .Z(n2161) );
  XNOR U2110 ( .A(n2170), .B(n2171), .Z(n2159) );
  AND U2111 ( .A(n242), .B(n2172), .Z(n2171) );
  XOR U2112 ( .A(p_input[158]), .B(n2170), .Z(n2172) );
  XNOR U2113 ( .A(n2173), .B(n2174), .Z(n2170) );
  AND U2114 ( .A(n246), .B(n2175), .Z(n2174) );
  XOR U2115 ( .A(n2176), .B(n2177), .Z(n2168) );
  AND U2116 ( .A(n250), .B(n2167), .Z(n2177) );
  XNOR U2117 ( .A(n2178), .B(n2165), .Z(n2167) );
  XOR U2118 ( .A(n2179), .B(n2180), .Z(n2165) );
  AND U2119 ( .A(n273), .B(n2181), .Z(n2180) );
  IV U2120 ( .A(n2176), .Z(n2178) );
  XOR U2121 ( .A(n2182), .B(n2183), .Z(n2176) );
  AND U2122 ( .A(n257), .B(n2175), .Z(n2183) );
  XNOR U2123 ( .A(n2173), .B(n2182), .Z(n2175) );
  XNOR U2124 ( .A(n2184), .B(n2185), .Z(n2173) );
  AND U2125 ( .A(n261), .B(n2186), .Z(n2185) );
  XOR U2126 ( .A(p_input[174]), .B(n2184), .Z(n2186) );
  XNOR U2127 ( .A(n2187), .B(n2188), .Z(n2184) );
  AND U2128 ( .A(n265), .B(n2189), .Z(n2188) );
  XOR U2129 ( .A(n2190), .B(n2191), .Z(n2182) );
  AND U2130 ( .A(n269), .B(n2181), .Z(n2191) );
  XNOR U2131 ( .A(n2192), .B(n2179), .Z(n2181) );
  XOR U2132 ( .A(n2193), .B(n2194), .Z(n2179) );
  AND U2133 ( .A(n292), .B(n2195), .Z(n2194) );
  IV U2134 ( .A(n2190), .Z(n2192) );
  XOR U2135 ( .A(n2196), .B(n2197), .Z(n2190) );
  AND U2136 ( .A(n276), .B(n2189), .Z(n2197) );
  XNOR U2137 ( .A(n2187), .B(n2196), .Z(n2189) );
  XNOR U2138 ( .A(n2198), .B(n2199), .Z(n2187) );
  AND U2139 ( .A(n280), .B(n2200), .Z(n2199) );
  XOR U2140 ( .A(p_input[190]), .B(n2198), .Z(n2200) );
  XNOR U2141 ( .A(n2201), .B(n2202), .Z(n2198) );
  AND U2142 ( .A(n284), .B(n2203), .Z(n2202) );
  XOR U2143 ( .A(n2204), .B(n2205), .Z(n2196) );
  AND U2144 ( .A(n288), .B(n2195), .Z(n2205) );
  XNOR U2145 ( .A(n2206), .B(n2193), .Z(n2195) );
  XOR U2146 ( .A(n2207), .B(n2208), .Z(n2193) );
  AND U2147 ( .A(n310), .B(n2209), .Z(n2208) );
  IV U2148 ( .A(n2204), .Z(n2206) );
  XOR U2149 ( .A(n2210), .B(n2211), .Z(n2204) );
  AND U2150 ( .A(n295), .B(n2203), .Z(n2211) );
  XNOR U2151 ( .A(n2201), .B(n2210), .Z(n2203) );
  XNOR U2152 ( .A(n2212), .B(n2213), .Z(n2201) );
  AND U2153 ( .A(n299), .B(n2214), .Z(n2213) );
  XOR U2154 ( .A(p_input[206]), .B(n2212), .Z(n2214) );
  XOR U2155 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n2215), 
        .Z(n2212) );
  AND U2156 ( .A(n302), .B(n2216), .Z(n2215) );
  XOR U2157 ( .A(n2217), .B(n2218), .Z(n2210) );
  AND U2158 ( .A(n306), .B(n2209), .Z(n2218) );
  XNOR U2159 ( .A(n2219), .B(n2207), .Z(n2209) );
  XOR U2160 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n2220), .Z(n2207) );
  AND U2161 ( .A(n318), .B(n2221), .Z(n2220) );
  IV U2162 ( .A(n2217), .Z(n2219) );
  XOR U2163 ( .A(n2222), .B(n2223), .Z(n2217) );
  AND U2164 ( .A(n313), .B(n2216), .Z(n2223) );
  XOR U2165 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n2222), 
        .Z(n2216) );
  XOR U2166 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(n2224), 
        .Z(n2222) );
  AND U2167 ( .A(n315), .B(n2221), .Z(n2224) );
  XOR U2168 ( .A(n2225), .B(n2226), .Z(n2221) );
  IV U2169 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n2226) );
  IV U2170 ( .A(\knn_comb_/min_val_out[0][14] ), .Z(n2225) );
  XOR U2171 ( .A(n53), .B(n2227), .Z(o[13]) );
  AND U2172 ( .A(n62), .B(n2228), .Z(n53) );
  XOR U2173 ( .A(n54), .B(n2227), .Z(n2228) );
  XOR U2174 ( .A(n2229), .B(n2230), .Z(n2227) );
  AND U2175 ( .A(n82), .B(n2231), .Z(n2230) );
  XOR U2176 ( .A(n2232), .B(n17), .Z(n54) );
  AND U2177 ( .A(n65), .B(n2233), .Z(n17) );
  XOR U2178 ( .A(n18), .B(n2232), .Z(n2233) );
  XOR U2179 ( .A(n2234), .B(n2235), .Z(n18) );
  AND U2180 ( .A(n70), .B(n2236), .Z(n2235) );
  XOR U2181 ( .A(p_input[13]), .B(n2234), .Z(n2236) );
  XNOR U2182 ( .A(n2237), .B(n2238), .Z(n2234) );
  AND U2183 ( .A(n74), .B(n2239), .Z(n2238) );
  XOR U2184 ( .A(n2240), .B(n2241), .Z(n2232) );
  AND U2185 ( .A(n78), .B(n2231), .Z(n2241) );
  XNOR U2186 ( .A(n2242), .B(n2229), .Z(n2231) );
  XOR U2187 ( .A(n2243), .B(n2244), .Z(n2229) );
  AND U2188 ( .A(n102), .B(n2245), .Z(n2244) );
  IV U2189 ( .A(n2240), .Z(n2242) );
  XOR U2190 ( .A(n2246), .B(n2247), .Z(n2240) );
  AND U2191 ( .A(n86), .B(n2239), .Z(n2247) );
  XNOR U2192 ( .A(n2237), .B(n2246), .Z(n2239) );
  XNOR U2193 ( .A(n2248), .B(n2249), .Z(n2237) );
  AND U2194 ( .A(n90), .B(n2250), .Z(n2249) );
  XOR U2195 ( .A(p_input[29]), .B(n2248), .Z(n2250) );
  XNOR U2196 ( .A(n2251), .B(n2252), .Z(n2248) );
  AND U2197 ( .A(n94), .B(n2253), .Z(n2252) );
  XOR U2198 ( .A(n2254), .B(n2255), .Z(n2246) );
  AND U2199 ( .A(n98), .B(n2245), .Z(n2255) );
  XNOR U2200 ( .A(n2256), .B(n2243), .Z(n2245) );
  XOR U2201 ( .A(n2257), .B(n2258), .Z(n2243) );
  AND U2202 ( .A(n121), .B(n2259), .Z(n2258) );
  IV U2203 ( .A(n2254), .Z(n2256) );
  XOR U2204 ( .A(n2260), .B(n2261), .Z(n2254) );
  AND U2205 ( .A(n105), .B(n2253), .Z(n2261) );
  XNOR U2206 ( .A(n2251), .B(n2260), .Z(n2253) );
  XNOR U2207 ( .A(n2262), .B(n2263), .Z(n2251) );
  AND U2208 ( .A(n109), .B(n2264), .Z(n2263) );
  XOR U2209 ( .A(p_input[45]), .B(n2262), .Z(n2264) );
  XNOR U2210 ( .A(n2265), .B(n2266), .Z(n2262) );
  AND U2211 ( .A(n113), .B(n2267), .Z(n2266) );
  XOR U2212 ( .A(n2268), .B(n2269), .Z(n2260) );
  AND U2213 ( .A(n117), .B(n2259), .Z(n2269) );
  XNOR U2214 ( .A(n2270), .B(n2257), .Z(n2259) );
  XOR U2215 ( .A(n2271), .B(n2272), .Z(n2257) );
  AND U2216 ( .A(n140), .B(n2273), .Z(n2272) );
  IV U2217 ( .A(n2268), .Z(n2270) );
  XOR U2218 ( .A(n2274), .B(n2275), .Z(n2268) );
  AND U2219 ( .A(n124), .B(n2267), .Z(n2275) );
  XNOR U2220 ( .A(n2265), .B(n2274), .Z(n2267) );
  XNOR U2221 ( .A(n2276), .B(n2277), .Z(n2265) );
  AND U2222 ( .A(n128), .B(n2278), .Z(n2277) );
  XOR U2223 ( .A(p_input[61]), .B(n2276), .Z(n2278) );
  XNOR U2224 ( .A(n2279), .B(n2280), .Z(n2276) );
  AND U2225 ( .A(n132), .B(n2281), .Z(n2280) );
  XOR U2226 ( .A(n2282), .B(n2283), .Z(n2274) );
  AND U2227 ( .A(n136), .B(n2273), .Z(n2283) );
  XNOR U2228 ( .A(n2284), .B(n2271), .Z(n2273) );
  XOR U2229 ( .A(n2285), .B(n2286), .Z(n2271) );
  AND U2230 ( .A(n159), .B(n2287), .Z(n2286) );
  IV U2231 ( .A(n2282), .Z(n2284) );
  XOR U2232 ( .A(n2288), .B(n2289), .Z(n2282) );
  AND U2233 ( .A(n143), .B(n2281), .Z(n2289) );
  XNOR U2234 ( .A(n2279), .B(n2288), .Z(n2281) );
  XNOR U2235 ( .A(n2290), .B(n2291), .Z(n2279) );
  AND U2236 ( .A(n147), .B(n2292), .Z(n2291) );
  XOR U2237 ( .A(p_input[77]), .B(n2290), .Z(n2292) );
  XNOR U2238 ( .A(n2293), .B(n2294), .Z(n2290) );
  AND U2239 ( .A(n151), .B(n2295), .Z(n2294) );
  XOR U2240 ( .A(n2296), .B(n2297), .Z(n2288) );
  AND U2241 ( .A(n155), .B(n2287), .Z(n2297) );
  XNOR U2242 ( .A(n2298), .B(n2285), .Z(n2287) );
  XOR U2243 ( .A(n2299), .B(n2300), .Z(n2285) );
  AND U2244 ( .A(n178), .B(n2301), .Z(n2300) );
  IV U2245 ( .A(n2296), .Z(n2298) );
  XOR U2246 ( .A(n2302), .B(n2303), .Z(n2296) );
  AND U2247 ( .A(n162), .B(n2295), .Z(n2303) );
  XNOR U2248 ( .A(n2293), .B(n2302), .Z(n2295) );
  XNOR U2249 ( .A(n2304), .B(n2305), .Z(n2293) );
  AND U2250 ( .A(n166), .B(n2306), .Z(n2305) );
  XOR U2251 ( .A(p_input[93]), .B(n2304), .Z(n2306) );
  XNOR U2252 ( .A(n2307), .B(n2308), .Z(n2304) );
  AND U2253 ( .A(n170), .B(n2309), .Z(n2308) );
  XOR U2254 ( .A(n2310), .B(n2311), .Z(n2302) );
  AND U2255 ( .A(n174), .B(n2301), .Z(n2311) );
  XNOR U2256 ( .A(n2312), .B(n2299), .Z(n2301) );
  XOR U2257 ( .A(n2313), .B(n2314), .Z(n2299) );
  AND U2258 ( .A(n197), .B(n2315), .Z(n2314) );
  IV U2259 ( .A(n2310), .Z(n2312) );
  XOR U2260 ( .A(n2316), .B(n2317), .Z(n2310) );
  AND U2261 ( .A(n181), .B(n2309), .Z(n2317) );
  XNOR U2262 ( .A(n2307), .B(n2316), .Z(n2309) );
  XNOR U2263 ( .A(n2318), .B(n2319), .Z(n2307) );
  AND U2264 ( .A(n185), .B(n2320), .Z(n2319) );
  XOR U2265 ( .A(p_input[109]), .B(n2318), .Z(n2320) );
  XNOR U2266 ( .A(n2321), .B(n2322), .Z(n2318) );
  AND U2267 ( .A(n189), .B(n2323), .Z(n2322) );
  XOR U2268 ( .A(n2324), .B(n2325), .Z(n2316) );
  AND U2269 ( .A(n193), .B(n2315), .Z(n2325) );
  XNOR U2270 ( .A(n2326), .B(n2313), .Z(n2315) );
  XOR U2271 ( .A(n2327), .B(n2328), .Z(n2313) );
  AND U2272 ( .A(n216), .B(n2329), .Z(n2328) );
  IV U2273 ( .A(n2324), .Z(n2326) );
  XOR U2274 ( .A(n2330), .B(n2331), .Z(n2324) );
  AND U2275 ( .A(n200), .B(n2323), .Z(n2331) );
  XNOR U2276 ( .A(n2321), .B(n2330), .Z(n2323) );
  XNOR U2277 ( .A(n2332), .B(n2333), .Z(n2321) );
  AND U2278 ( .A(n204), .B(n2334), .Z(n2333) );
  XOR U2279 ( .A(p_input[125]), .B(n2332), .Z(n2334) );
  XNOR U2280 ( .A(n2335), .B(n2336), .Z(n2332) );
  AND U2281 ( .A(n208), .B(n2337), .Z(n2336) );
  XOR U2282 ( .A(n2338), .B(n2339), .Z(n2330) );
  AND U2283 ( .A(n212), .B(n2329), .Z(n2339) );
  XNOR U2284 ( .A(n2340), .B(n2327), .Z(n2329) );
  XOR U2285 ( .A(n2341), .B(n2342), .Z(n2327) );
  AND U2286 ( .A(n235), .B(n2343), .Z(n2342) );
  IV U2287 ( .A(n2338), .Z(n2340) );
  XOR U2288 ( .A(n2344), .B(n2345), .Z(n2338) );
  AND U2289 ( .A(n219), .B(n2337), .Z(n2345) );
  XNOR U2290 ( .A(n2335), .B(n2344), .Z(n2337) );
  XNOR U2291 ( .A(n2346), .B(n2347), .Z(n2335) );
  AND U2292 ( .A(n223), .B(n2348), .Z(n2347) );
  XOR U2293 ( .A(p_input[141]), .B(n2346), .Z(n2348) );
  XNOR U2294 ( .A(n2349), .B(n2350), .Z(n2346) );
  AND U2295 ( .A(n227), .B(n2351), .Z(n2350) );
  XOR U2296 ( .A(n2352), .B(n2353), .Z(n2344) );
  AND U2297 ( .A(n231), .B(n2343), .Z(n2353) );
  XNOR U2298 ( .A(n2354), .B(n2341), .Z(n2343) );
  XOR U2299 ( .A(n2355), .B(n2356), .Z(n2341) );
  AND U2300 ( .A(n254), .B(n2357), .Z(n2356) );
  IV U2301 ( .A(n2352), .Z(n2354) );
  XOR U2302 ( .A(n2358), .B(n2359), .Z(n2352) );
  AND U2303 ( .A(n238), .B(n2351), .Z(n2359) );
  XNOR U2304 ( .A(n2349), .B(n2358), .Z(n2351) );
  XNOR U2305 ( .A(n2360), .B(n2361), .Z(n2349) );
  AND U2306 ( .A(n242), .B(n2362), .Z(n2361) );
  XOR U2307 ( .A(p_input[157]), .B(n2360), .Z(n2362) );
  XNOR U2308 ( .A(n2363), .B(n2364), .Z(n2360) );
  AND U2309 ( .A(n246), .B(n2365), .Z(n2364) );
  XOR U2310 ( .A(n2366), .B(n2367), .Z(n2358) );
  AND U2311 ( .A(n250), .B(n2357), .Z(n2367) );
  XNOR U2312 ( .A(n2368), .B(n2355), .Z(n2357) );
  XOR U2313 ( .A(n2369), .B(n2370), .Z(n2355) );
  AND U2314 ( .A(n273), .B(n2371), .Z(n2370) );
  IV U2315 ( .A(n2366), .Z(n2368) );
  XOR U2316 ( .A(n2372), .B(n2373), .Z(n2366) );
  AND U2317 ( .A(n257), .B(n2365), .Z(n2373) );
  XNOR U2318 ( .A(n2363), .B(n2372), .Z(n2365) );
  XNOR U2319 ( .A(n2374), .B(n2375), .Z(n2363) );
  AND U2320 ( .A(n261), .B(n2376), .Z(n2375) );
  XOR U2321 ( .A(p_input[173]), .B(n2374), .Z(n2376) );
  XNOR U2322 ( .A(n2377), .B(n2378), .Z(n2374) );
  AND U2323 ( .A(n265), .B(n2379), .Z(n2378) );
  XOR U2324 ( .A(n2380), .B(n2381), .Z(n2372) );
  AND U2325 ( .A(n269), .B(n2371), .Z(n2381) );
  XNOR U2326 ( .A(n2382), .B(n2369), .Z(n2371) );
  XOR U2327 ( .A(n2383), .B(n2384), .Z(n2369) );
  AND U2328 ( .A(n292), .B(n2385), .Z(n2384) );
  IV U2329 ( .A(n2380), .Z(n2382) );
  XOR U2330 ( .A(n2386), .B(n2387), .Z(n2380) );
  AND U2331 ( .A(n276), .B(n2379), .Z(n2387) );
  XNOR U2332 ( .A(n2377), .B(n2386), .Z(n2379) );
  XNOR U2333 ( .A(n2388), .B(n2389), .Z(n2377) );
  AND U2334 ( .A(n280), .B(n2390), .Z(n2389) );
  XOR U2335 ( .A(p_input[189]), .B(n2388), .Z(n2390) );
  XNOR U2336 ( .A(n2391), .B(n2392), .Z(n2388) );
  AND U2337 ( .A(n284), .B(n2393), .Z(n2392) );
  XOR U2338 ( .A(n2394), .B(n2395), .Z(n2386) );
  AND U2339 ( .A(n288), .B(n2385), .Z(n2395) );
  XNOR U2340 ( .A(n2396), .B(n2383), .Z(n2385) );
  XOR U2341 ( .A(n2397), .B(n2398), .Z(n2383) );
  AND U2342 ( .A(n310), .B(n2399), .Z(n2398) );
  IV U2343 ( .A(n2394), .Z(n2396) );
  XOR U2344 ( .A(n2400), .B(n2401), .Z(n2394) );
  AND U2345 ( .A(n295), .B(n2393), .Z(n2401) );
  XNOR U2346 ( .A(n2391), .B(n2400), .Z(n2393) );
  XNOR U2347 ( .A(n2402), .B(n2403), .Z(n2391) );
  AND U2348 ( .A(n299), .B(n2404), .Z(n2403) );
  XOR U2349 ( .A(p_input[205]), .B(n2402), .Z(n2404) );
  XOR U2350 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(n2405), 
        .Z(n2402) );
  AND U2351 ( .A(n302), .B(n2406), .Z(n2405) );
  XOR U2352 ( .A(n2407), .B(n2408), .Z(n2400) );
  AND U2353 ( .A(n306), .B(n2399), .Z(n2408) );
  XNOR U2354 ( .A(n2409), .B(n2397), .Z(n2399) );
  XOR U2355 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n2410), .Z(n2397) );
  AND U2356 ( .A(n318), .B(n2411), .Z(n2410) );
  IV U2357 ( .A(n2407), .Z(n2409) );
  XOR U2358 ( .A(n2412), .B(n2413), .Z(n2407) );
  AND U2359 ( .A(n313), .B(n2406), .Z(n2413) );
  XOR U2360 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(n2412), 
        .Z(n2406) );
  XOR U2361 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(n2414), 
        .Z(n2412) );
  AND U2362 ( .A(n315), .B(n2411), .Z(n2414) );
  XOR U2363 ( .A(\knn_comb_/min_val_out[0][13] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n2411) );
  XOR U2364 ( .A(n55), .B(n2415), .Z(o[12]) );
  AND U2365 ( .A(n62), .B(n2416), .Z(n55) );
  XOR U2366 ( .A(n56), .B(n2415), .Z(n2416) );
  XOR U2367 ( .A(n2417), .B(n2418), .Z(n2415) );
  AND U2368 ( .A(n82), .B(n2419), .Z(n2418) );
  XOR U2369 ( .A(n2420), .B(n19), .Z(n56) );
  AND U2370 ( .A(n65), .B(n2421), .Z(n19) );
  XOR U2371 ( .A(n20), .B(n2420), .Z(n2421) );
  XOR U2372 ( .A(n2422), .B(n2423), .Z(n20) );
  AND U2373 ( .A(n70), .B(n2424), .Z(n2423) );
  XOR U2374 ( .A(p_input[12]), .B(n2422), .Z(n2424) );
  XNOR U2375 ( .A(n2425), .B(n2426), .Z(n2422) );
  AND U2376 ( .A(n74), .B(n2427), .Z(n2426) );
  XOR U2377 ( .A(n2428), .B(n2429), .Z(n2420) );
  AND U2378 ( .A(n78), .B(n2419), .Z(n2429) );
  XNOR U2379 ( .A(n2430), .B(n2417), .Z(n2419) );
  XOR U2380 ( .A(n2431), .B(n2432), .Z(n2417) );
  AND U2381 ( .A(n102), .B(n2433), .Z(n2432) );
  IV U2382 ( .A(n2428), .Z(n2430) );
  XOR U2383 ( .A(n2434), .B(n2435), .Z(n2428) );
  AND U2384 ( .A(n86), .B(n2427), .Z(n2435) );
  XNOR U2385 ( .A(n2425), .B(n2434), .Z(n2427) );
  XNOR U2386 ( .A(n2436), .B(n2437), .Z(n2425) );
  AND U2387 ( .A(n90), .B(n2438), .Z(n2437) );
  XOR U2388 ( .A(p_input[28]), .B(n2436), .Z(n2438) );
  XNOR U2389 ( .A(n2439), .B(n2440), .Z(n2436) );
  AND U2390 ( .A(n94), .B(n2441), .Z(n2440) );
  XOR U2391 ( .A(n2442), .B(n2443), .Z(n2434) );
  AND U2392 ( .A(n98), .B(n2433), .Z(n2443) );
  XNOR U2393 ( .A(n2444), .B(n2431), .Z(n2433) );
  XOR U2394 ( .A(n2445), .B(n2446), .Z(n2431) );
  AND U2395 ( .A(n121), .B(n2447), .Z(n2446) );
  IV U2396 ( .A(n2442), .Z(n2444) );
  XOR U2397 ( .A(n2448), .B(n2449), .Z(n2442) );
  AND U2398 ( .A(n105), .B(n2441), .Z(n2449) );
  XNOR U2399 ( .A(n2439), .B(n2448), .Z(n2441) );
  XNOR U2400 ( .A(n2450), .B(n2451), .Z(n2439) );
  AND U2401 ( .A(n109), .B(n2452), .Z(n2451) );
  XOR U2402 ( .A(p_input[44]), .B(n2450), .Z(n2452) );
  XNOR U2403 ( .A(n2453), .B(n2454), .Z(n2450) );
  AND U2404 ( .A(n113), .B(n2455), .Z(n2454) );
  XOR U2405 ( .A(n2456), .B(n2457), .Z(n2448) );
  AND U2406 ( .A(n117), .B(n2447), .Z(n2457) );
  XNOR U2407 ( .A(n2458), .B(n2445), .Z(n2447) );
  XOR U2408 ( .A(n2459), .B(n2460), .Z(n2445) );
  AND U2409 ( .A(n140), .B(n2461), .Z(n2460) );
  IV U2410 ( .A(n2456), .Z(n2458) );
  XOR U2411 ( .A(n2462), .B(n2463), .Z(n2456) );
  AND U2412 ( .A(n124), .B(n2455), .Z(n2463) );
  XNOR U2413 ( .A(n2453), .B(n2462), .Z(n2455) );
  XNOR U2414 ( .A(n2464), .B(n2465), .Z(n2453) );
  AND U2415 ( .A(n128), .B(n2466), .Z(n2465) );
  XOR U2416 ( .A(p_input[60]), .B(n2464), .Z(n2466) );
  XNOR U2417 ( .A(n2467), .B(n2468), .Z(n2464) );
  AND U2418 ( .A(n132), .B(n2469), .Z(n2468) );
  XOR U2419 ( .A(n2470), .B(n2471), .Z(n2462) );
  AND U2420 ( .A(n136), .B(n2461), .Z(n2471) );
  XNOR U2421 ( .A(n2472), .B(n2459), .Z(n2461) );
  XOR U2422 ( .A(n2473), .B(n2474), .Z(n2459) );
  AND U2423 ( .A(n159), .B(n2475), .Z(n2474) );
  IV U2424 ( .A(n2470), .Z(n2472) );
  XOR U2425 ( .A(n2476), .B(n2477), .Z(n2470) );
  AND U2426 ( .A(n143), .B(n2469), .Z(n2477) );
  XNOR U2427 ( .A(n2467), .B(n2476), .Z(n2469) );
  XNOR U2428 ( .A(n2478), .B(n2479), .Z(n2467) );
  AND U2429 ( .A(n147), .B(n2480), .Z(n2479) );
  XOR U2430 ( .A(p_input[76]), .B(n2478), .Z(n2480) );
  XNOR U2431 ( .A(n2481), .B(n2482), .Z(n2478) );
  AND U2432 ( .A(n151), .B(n2483), .Z(n2482) );
  XOR U2433 ( .A(n2484), .B(n2485), .Z(n2476) );
  AND U2434 ( .A(n155), .B(n2475), .Z(n2485) );
  XNOR U2435 ( .A(n2486), .B(n2473), .Z(n2475) );
  XOR U2436 ( .A(n2487), .B(n2488), .Z(n2473) );
  AND U2437 ( .A(n178), .B(n2489), .Z(n2488) );
  IV U2438 ( .A(n2484), .Z(n2486) );
  XOR U2439 ( .A(n2490), .B(n2491), .Z(n2484) );
  AND U2440 ( .A(n162), .B(n2483), .Z(n2491) );
  XNOR U2441 ( .A(n2481), .B(n2490), .Z(n2483) );
  XNOR U2442 ( .A(n2492), .B(n2493), .Z(n2481) );
  AND U2443 ( .A(n166), .B(n2494), .Z(n2493) );
  XOR U2444 ( .A(p_input[92]), .B(n2492), .Z(n2494) );
  XNOR U2445 ( .A(n2495), .B(n2496), .Z(n2492) );
  AND U2446 ( .A(n170), .B(n2497), .Z(n2496) );
  XOR U2447 ( .A(n2498), .B(n2499), .Z(n2490) );
  AND U2448 ( .A(n174), .B(n2489), .Z(n2499) );
  XNOR U2449 ( .A(n2500), .B(n2487), .Z(n2489) );
  XOR U2450 ( .A(n2501), .B(n2502), .Z(n2487) );
  AND U2451 ( .A(n197), .B(n2503), .Z(n2502) );
  IV U2452 ( .A(n2498), .Z(n2500) );
  XOR U2453 ( .A(n2504), .B(n2505), .Z(n2498) );
  AND U2454 ( .A(n181), .B(n2497), .Z(n2505) );
  XNOR U2455 ( .A(n2495), .B(n2504), .Z(n2497) );
  XNOR U2456 ( .A(n2506), .B(n2507), .Z(n2495) );
  AND U2457 ( .A(n185), .B(n2508), .Z(n2507) );
  XOR U2458 ( .A(p_input[108]), .B(n2506), .Z(n2508) );
  XNOR U2459 ( .A(n2509), .B(n2510), .Z(n2506) );
  AND U2460 ( .A(n189), .B(n2511), .Z(n2510) );
  XOR U2461 ( .A(n2512), .B(n2513), .Z(n2504) );
  AND U2462 ( .A(n193), .B(n2503), .Z(n2513) );
  XNOR U2463 ( .A(n2514), .B(n2501), .Z(n2503) );
  XOR U2464 ( .A(n2515), .B(n2516), .Z(n2501) );
  AND U2465 ( .A(n216), .B(n2517), .Z(n2516) );
  IV U2466 ( .A(n2512), .Z(n2514) );
  XOR U2467 ( .A(n2518), .B(n2519), .Z(n2512) );
  AND U2468 ( .A(n200), .B(n2511), .Z(n2519) );
  XNOR U2469 ( .A(n2509), .B(n2518), .Z(n2511) );
  XNOR U2470 ( .A(n2520), .B(n2521), .Z(n2509) );
  AND U2471 ( .A(n204), .B(n2522), .Z(n2521) );
  XOR U2472 ( .A(p_input[124]), .B(n2520), .Z(n2522) );
  XNOR U2473 ( .A(n2523), .B(n2524), .Z(n2520) );
  AND U2474 ( .A(n208), .B(n2525), .Z(n2524) );
  XOR U2475 ( .A(n2526), .B(n2527), .Z(n2518) );
  AND U2476 ( .A(n212), .B(n2517), .Z(n2527) );
  XNOR U2477 ( .A(n2528), .B(n2515), .Z(n2517) );
  XOR U2478 ( .A(n2529), .B(n2530), .Z(n2515) );
  AND U2479 ( .A(n235), .B(n2531), .Z(n2530) );
  IV U2480 ( .A(n2526), .Z(n2528) );
  XOR U2481 ( .A(n2532), .B(n2533), .Z(n2526) );
  AND U2482 ( .A(n219), .B(n2525), .Z(n2533) );
  XNOR U2483 ( .A(n2523), .B(n2532), .Z(n2525) );
  XNOR U2484 ( .A(n2534), .B(n2535), .Z(n2523) );
  AND U2485 ( .A(n223), .B(n2536), .Z(n2535) );
  XOR U2486 ( .A(p_input[140]), .B(n2534), .Z(n2536) );
  XNOR U2487 ( .A(n2537), .B(n2538), .Z(n2534) );
  AND U2488 ( .A(n227), .B(n2539), .Z(n2538) );
  XOR U2489 ( .A(n2540), .B(n2541), .Z(n2532) );
  AND U2490 ( .A(n231), .B(n2531), .Z(n2541) );
  XNOR U2491 ( .A(n2542), .B(n2529), .Z(n2531) );
  XOR U2492 ( .A(n2543), .B(n2544), .Z(n2529) );
  AND U2493 ( .A(n254), .B(n2545), .Z(n2544) );
  IV U2494 ( .A(n2540), .Z(n2542) );
  XOR U2495 ( .A(n2546), .B(n2547), .Z(n2540) );
  AND U2496 ( .A(n238), .B(n2539), .Z(n2547) );
  XNOR U2497 ( .A(n2537), .B(n2546), .Z(n2539) );
  XNOR U2498 ( .A(n2548), .B(n2549), .Z(n2537) );
  AND U2499 ( .A(n242), .B(n2550), .Z(n2549) );
  XOR U2500 ( .A(p_input[156]), .B(n2548), .Z(n2550) );
  XNOR U2501 ( .A(n2551), .B(n2552), .Z(n2548) );
  AND U2502 ( .A(n246), .B(n2553), .Z(n2552) );
  XOR U2503 ( .A(n2554), .B(n2555), .Z(n2546) );
  AND U2504 ( .A(n250), .B(n2545), .Z(n2555) );
  XNOR U2505 ( .A(n2556), .B(n2543), .Z(n2545) );
  XOR U2506 ( .A(n2557), .B(n2558), .Z(n2543) );
  AND U2507 ( .A(n273), .B(n2559), .Z(n2558) );
  IV U2508 ( .A(n2554), .Z(n2556) );
  XOR U2509 ( .A(n2560), .B(n2561), .Z(n2554) );
  AND U2510 ( .A(n257), .B(n2553), .Z(n2561) );
  XNOR U2511 ( .A(n2551), .B(n2560), .Z(n2553) );
  XNOR U2512 ( .A(n2562), .B(n2563), .Z(n2551) );
  AND U2513 ( .A(n261), .B(n2564), .Z(n2563) );
  XOR U2514 ( .A(p_input[172]), .B(n2562), .Z(n2564) );
  XNOR U2515 ( .A(n2565), .B(n2566), .Z(n2562) );
  AND U2516 ( .A(n265), .B(n2567), .Z(n2566) );
  XOR U2517 ( .A(n2568), .B(n2569), .Z(n2560) );
  AND U2518 ( .A(n269), .B(n2559), .Z(n2569) );
  XNOR U2519 ( .A(n2570), .B(n2557), .Z(n2559) );
  XOR U2520 ( .A(n2571), .B(n2572), .Z(n2557) );
  AND U2521 ( .A(n292), .B(n2573), .Z(n2572) );
  IV U2522 ( .A(n2568), .Z(n2570) );
  XOR U2523 ( .A(n2574), .B(n2575), .Z(n2568) );
  AND U2524 ( .A(n276), .B(n2567), .Z(n2575) );
  XNOR U2525 ( .A(n2565), .B(n2574), .Z(n2567) );
  XNOR U2526 ( .A(n2576), .B(n2577), .Z(n2565) );
  AND U2527 ( .A(n280), .B(n2578), .Z(n2577) );
  XOR U2528 ( .A(p_input[188]), .B(n2576), .Z(n2578) );
  XNOR U2529 ( .A(n2579), .B(n2580), .Z(n2576) );
  AND U2530 ( .A(n284), .B(n2581), .Z(n2580) );
  XOR U2531 ( .A(n2582), .B(n2583), .Z(n2574) );
  AND U2532 ( .A(n288), .B(n2573), .Z(n2583) );
  XNOR U2533 ( .A(n2584), .B(n2571), .Z(n2573) );
  XOR U2534 ( .A(n2585), .B(n2586), .Z(n2571) );
  AND U2535 ( .A(n310), .B(n2587), .Z(n2586) );
  IV U2536 ( .A(n2582), .Z(n2584) );
  XOR U2537 ( .A(n2588), .B(n2589), .Z(n2582) );
  AND U2538 ( .A(n295), .B(n2581), .Z(n2589) );
  XNOR U2539 ( .A(n2579), .B(n2588), .Z(n2581) );
  XNOR U2540 ( .A(n2590), .B(n2591), .Z(n2579) );
  AND U2541 ( .A(n299), .B(n2592), .Z(n2591) );
  XOR U2542 ( .A(p_input[204]), .B(n2590), .Z(n2592) );
  XOR U2543 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n2593), 
        .Z(n2590) );
  AND U2544 ( .A(n302), .B(n2594), .Z(n2593) );
  XOR U2545 ( .A(n2595), .B(n2596), .Z(n2588) );
  AND U2546 ( .A(n306), .B(n2587), .Z(n2596) );
  XNOR U2547 ( .A(n2597), .B(n2585), .Z(n2587) );
  XOR U2548 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n2598), .Z(n2585) );
  AND U2549 ( .A(n318), .B(n2599), .Z(n2598) );
  IV U2550 ( .A(n2595), .Z(n2597) );
  XOR U2551 ( .A(n2600), .B(n2601), .Z(n2595) );
  AND U2552 ( .A(n313), .B(n2594), .Z(n2601) );
  XOR U2553 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n2600), 
        .Z(n2594) );
  XOR U2554 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(n2602), 
        .Z(n2600) );
  AND U2555 ( .A(n315), .B(n2599), .Z(n2602) );
  XOR U2556 ( .A(\knn_comb_/min_val_out[0][12] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n2599) );
  XOR U2557 ( .A(n57), .B(n2603), .Z(o[11]) );
  AND U2558 ( .A(n62), .B(n2604), .Z(n57) );
  XOR U2559 ( .A(n58), .B(n2603), .Z(n2604) );
  XOR U2560 ( .A(n2605), .B(n2606), .Z(n2603) );
  AND U2561 ( .A(n82), .B(n2607), .Z(n2606) );
  XOR U2562 ( .A(n2608), .B(n21), .Z(n58) );
  AND U2563 ( .A(n65), .B(n2609), .Z(n21) );
  XOR U2564 ( .A(n22), .B(n2608), .Z(n2609) );
  XOR U2565 ( .A(n2610), .B(n2611), .Z(n22) );
  AND U2566 ( .A(n70), .B(n2612), .Z(n2611) );
  XOR U2567 ( .A(p_input[11]), .B(n2610), .Z(n2612) );
  XNOR U2568 ( .A(n2613), .B(n2614), .Z(n2610) );
  AND U2569 ( .A(n74), .B(n2615), .Z(n2614) );
  XOR U2570 ( .A(n2616), .B(n2617), .Z(n2608) );
  AND U2571 ( .A(n78), .B(n2607), .Z(n2617) );
  XNOR U2572 ( .A(n2618), .B(n2605), .Z(n2607) );
  XOR U2573 ( .A(n2619), .B(n2620), .Z(n2605) );
  AND U2574 ( .A(n102), .B(n2621), .Z(n2620) );
  IV U2575 ( .A(n2616), .Z(n2618) );
  XOR U2576 ( .A(n2622), .B(n2623), .Z(n2616) );
  AND U2577 ( .A(n86), .B(n2615), .Z(n2623) );
  XNOR U2578 ( .A(n2613), .B(n2622), .Z(n2615) );
  XNOR U2579 ( .A(n2624), .B(n2625), .Z(n2613) );
  AND U2580 ( .A(n90), .B(n2626), .Z(n2625) );
  XOR U2581 ( .A(p_input[27]), .B(n2624), .Z(n2626) );
  XNOR U2582 ( .A(n2627), .B(n2628), .Z(n2624) );
  AND U2583 ( .A(n94), .B(n2629), .Z(n2628) );
  XOR U2584 ( .A(n2630), .B(n2631), .Z(n2622) );
  AND U2585 ( .A(n98), .B(n2621), .Z(n2631) );
  XNOR U2586 ( .A(n2632), .B(n2619), .Z(n2621) );
  XOR U2587 ( .A(n2633), .B(n2634), .Z(n2619) );
  AND U2588 ( .A(n121), .B(n2635), .Z(n2634) );
  IV U2589 ( .A(n2630), .Z(n2632) );
  XOR U2590 ( .A(n2636), .B(n2637), .Z(n2630) );
  AND U2591 ( .A(n105), .B(n2629), .Z(n2637) );
  XNOR U2592 ( .A(n2627), .B(n2636), .Z(n2629) );
  XNOR U2593 ( .A(n2638), .B(n2639), .Z(n2627) );
  AND U2594 ( .A(n109), .B(n2640), .Z(n2639) );
  XOR U2595 ( .A(p_input[43]), .B(n2638), .Z(n2640) );
  XNOR U2596 ( .A(n2641), .B(n2642), .Z(n2638) );
  AND U2597 ( .A(n113), .B(n2643), .Z(n2642) );
  XOR U2598 ( .A(n2644), .B(n2645), .Z(n2636) );
  AND U2599 ( .A(n117), .B(n2635), .Z(n2645) );
  XNOR U2600 ( .A(n2646), .B(n2633), .Z(n2635) );
  XOR U2601 ( .A(n2647), .B(n2648), .Z(n2633) );
  AND U2602 ( .A(n140), .B(n2649), .Z(n2648) );
  IV U2603 ( .A(n2644), .Z(n2646) );
  XOR U2604 ( .A(n2650), .B(n2651), .Z(n2644) );
  AND U2605 ( .A(n124), .B(n2643), .Z(n2651) );
  XNOR U2606 ( .A(n2641), .B(n2650), .Z(n2643) );
  XNOR U2607 ( .A(n2652), .B(n2653), .Z(n2641) );
  AND U2608 ( .A(n128), .B(n2654), .Z(n2653) );
  XOR U2609 ( .A(p_input[59]), .B(n2652), .Z(n2654) );
  XNOR U2610 ( .A(n2655), .B(n2656), .Z(n2652) );
  AND U2611 ( .A(n132), .B(n2657), .Z(n2656) );
  XOR U2612 ( .A(n2658), .B(n2659), .Z(n2650) );
  AND U2613 ( .A(n136), .B(n2649), .Z(n2659) );
  XNOR U2614 ( .A(n2660), .B(n2647), .Z(n2649) );
  XOR U2615 ( .A(n2661), .B(n2662), .Z(n2647) );
  AND U2616 ( .A(n159), .B(n2663), .Z(n2662) );
  IV U2617 ( .A(n2658), .Z(n2660) );
  XOR U2618 ( .A(n2664), .B(n2665), .Z(n2658) );
  AND U2619 ( .A(n143), .B(n2657), .Z(n2665) );
  XNOR U2620 ( .A(n2655), .B(n2664), .Z(n2657) );
  XNOR U2621 ( .A(n2666), .B(n2667), .Z(n2655) );
  AND U2622 ( .A(n147), .B(n2668), .Z(n2667) );
  XOR U2623 ( .A(p_input[75]), .B(n2666), .Z(n2668) );
  XNOR U2624 ( .A(n2669), .B(n2670), .Z(n2666) );
  AND U2625 ( .A(n151), .B(n2671), .Z(n2670) );
  XOR U2626 ( .A(n2672), .B(n2673), .Z(n2664) );
  AND U2627 ( .A(n155), .B(n2663), .Z(n2673) );
  XNOR U2628 ( .A(n2674), .B(n2661), .Z(n2663) );
  XOR U2629 ( .A(n2675), .B(n2676), .Z(n2661) );
  AND U2630 ( .A(n178), .B(n2677), .Z(n2676) );
  IV U2631 ( .A(n2672), .Z(n2674) );
  XOR U2632 ( .A(n2678), .B(n2679), .Z(n2672) );
  AND U2633 ( .A(n162), .B(n2671), .Z(n2679) );
  XNOR U2634 ( .A(n2669), .B(n2678), .Z(n2671) );
  XNOR U2635 ( .A(n2680), .B(n2681), .Z(n2669) );
  AND U2636 ( .A(n166), .B(n2682), .Z(n2681) );
  XOR U2637 ( .A(p_input[91]), .B(n2680), .Z(n2682) );
  XNOR U2638 ( .A(n2683), .B(n2684), .Z(n2680) );
  AND U2639 ( .A(n170), .B(n2685), .Z(n2684) );
  XOR U2640 ( .A(n2686), .B(n2687), .Z(n2678) );
  AND U2641 ( .A(n174), .B(n2677), .Z(n2687) );
  XNOR U2642 ( .A(n2688), .B(n2675), .Z(n2677) );
  XOR U2643 ( .A(n2689), .B(n2690), .Z(n2675) );
  AND U2644 ( .A(n197), .B(n2691), .Z(n2690) );
  IV U2645 ( .A(n2686), .Z(n2688) );
  XOR U2646 ( .A(n2692), .B(n2693), .Z(n2686) );
  AND U2647 ( .A(n181), .B(n2685), .Z(n2693) );
  XNOR U2648 ( .A(n2683), .B(n2692), .Z(n2685) );
  XNOR U2649 ( .A(n2694), .B(n2695), .Z(n2683) );
  AND U2650 ( .A(n185), .B(n2696), .Z(n2695) );
  XOR U2651 ( .A(p_input[107]), .B(n2694), .Z(n2696) );
  XNOR U2652 ( .A(n2697), .B(n2698), .Z(n2694) );
  AND U2653 ( .A(n189), .B(n2699), .Z(n2698) );
  XOR U2654 ( .A(n2700), .B(n2701), .Z(n2692) );
  AND U2655 ( .A(n193), .B(n2691), .Z(n2701) );
  XNOR U2656 ( .A(n2702), .B(n2689), .Z(n2691) );
  XOR U2657 ( .A(n2703), .B(n2704), .Z(n2689) );
  AND U2658 ( .A(n216), .B(n2705), .Z(n2704) );
  IV U2659 ( .A(n2700), .Z(n2702) );
  XOR U2660 ( .A(n2706), .B(n2707), .Z(n2700) );
  AND U2661 ( .A(n200), .B(n2699), .Z(n2707) );
  XNOR U2662 ( .A(n2697), .B(n2706), .Z(n2699) );
  XNOR U2663 ( .A(n2708), .B(n2709), .Z(n2697) );
  AND U2664 ( .A(n204), .B(n2710), .Z(n2709) );
  XOR U2665 ( .A(p_input[123]), .B(n2708), .Z(n2710) );
  XNOR U2666 ( .A(n2711), .B(n2712), .Z(n2708) );
  AND U2667 ( .A(n208), .B(n2713), .Z(n2712) );
  XOR U2668 ( .A(n2714), .B(n2715), .Z(n2706) );
  AND U2669 ( .A(n212), .B(n2705), .Z(n2715) );
  XNOR U2670 ( .A(n2716), .B(n2703), .Z(n2705) );
  XOR U2671 ( .A(n2717), .B(n2718), .Z(n2703) );
  AND U2672 ( .A(n235), .B(n2719), .Z(n2718) );
  IV U2673 ( .A(n2714), .Z(n2716) );
  XOR U2674 ( .A(n2720), .B(n2721), .Z(n2714) );
  AND U2675 ( .A(n219), .B(n2713), .Z(n2721) );
  XNOR U2676 ( .A(n2711), .B(n2720), .Z(n2713) );
  XNOR U2677 ( .A(n2722), .B(n2723), .Z(n2711) );
  AND U2678 ( .A(n223), .B(n2724), .Z(n2723) );
  XOR U2679 ( .A(p_input[139]), .B(n2722), .Z(n2724) );
  XNOR U2680 ( .A(n2725), .B(n2726), .Z(n2722) );
  AND U2681 ( .A(n227), .B(n2727), .Z(n2726) );
  XOR U2682 ( .A(n2728), .B(n2729), .Z(n2720) );
  AND U2683 ( .A(n231), .B(n2719), .Z(n2729) );
  XNOR U2684 ( .A(n2730), .B(n2717), .Z(n2719) );
  XOR U2685 ( .A(n2731), .B(n2732), .Z(n2717) );
  AND U2686 ( .A(n254), .B(n2733), .Z(n2732) );
  IV U2687 ( .A(n2728), .Z(n2730) );
  XOR U2688 ( .A(n2734), .B(n2735), .Z(n2728) );
  AND U2689 ( .A(n238), .B(n2727), .Z(n2735) );
  XNOR U2690 ( .A(n2725), .B(n2734), .Z(n2727) );
  XNOR U2691 ( .A(n2736), .B(n2737), .Z(n2725) );
  AND U2692 ( .A(n242), .B(n2738), .Z(n2737) );
  XOR U2693 ( .A(p_input[155]), .B(n2736), .Z(n2738) );
  XNOR U2694 ( .A(n2739), .B(n2740), .Z(n2736) );
  AND U2695 ( .A(n246), .B(n2741), .Z(n2740) );
  XOR U2696 ( .A(n2742), .B(n2743), .Z(n2734) );
  AND U2697 ( .A(n250), .B(n2733), .Z(n2743) );
  XNOR U2698 ( .A(n2744), .B(n2731), .Z(n2733) );
  XOR U2699 ( .A(n2745), .B(n2746), .Z(n2731) );
  AND U2700 ( .A(n273), .B(n2747), .Z(n2746) );
  IV U2701 ( .A(n2742), .Z(n2744) );
  XOR U2702 ( .A(n2748), .B(n2749), .Z(n2742) );
  AND U2703 ( .A(n257), .B(n2741), .Z(n2749) );
  XNOR U2704 ( .A(n2739), .B(n2748), .Z(n2741) );
  XNOR U2705 ( .A(n2750), .B(n2751), .Z(n2739) );
  AND U2706 ( .A(n261), .B(n2752), .Z(n2751) );
  XOR U2707 ( .A(p_input[171]), .B(n2750), .Z(n2752) );
  XNOR U2708 ( .A(n2753), .B(n2754), .Z(n2750) );
  AND U2709 ( .A(n265), .B(n2755), .Z(n2754) );
  XOR U2710 ( .A(n2756), .B(n2757), .Z(n2748) );
  AND U2711 ( .A(n269), .B(n2747), .Z(n2757) );
  XNOR U2712 ( .A(n2758), .B(n2745), .Z(n2747) );
  XOR U2713 ( .A(n2759), .B(n2760), .Z(n2745) );
  AND U2714 ( .A(n292), .B(n2761), .Z(n2760) );
  IV U2715 ( .A(n2756), .Z(n2758) );
  XOR U2716 ( .A(n2762), .B(n2763), .Z(n2756) );
  AND U2717 ( .A(n276), .B(n2755), .Z(n2763) );
  XNOR U2718 ( .A(n2753), .B(n2762), .Z(n2755) );
  XNOR U2719 ( .A(n2764), .B(n2765), .Z(n2753) );
  AND U2720 ( .A(n280), .B(n2766), .Z(n2765) );
  XOR U2721 ( .A(p_input[187]), .B(n2764), .Z(n2766) );
  XNOR U2722 ( .A(n2767), .B(n2768), .Z(n2764) );
  AND U2723 ( .A(n284), .B(n2769), .Z(n2768) );
  XOR U2724 ( .A(n2770), .B(n2771), .Z(n2762) );
  AND U2725 ( .A(n288), .B(n2761), .Z(n2771) );
  XNOR U2726 ( .A(n2772), .B(n2759), .Z(n2761) );
  XOR U2727 ( .A(n2773), .B(n2774), .Z(n2759) );
  AND U2728 ( .A(n310), .B(n2775), .Z(n2774) );
  IV U2729 ( .A(n2770), .Z(n2772) );
  XOR U2730 ( .A(n2776), .B(n2777), .Z(n2770) );
  AND U2731 ( .A(n295), .B(n2769), .Z(n2777) );
  XNOR U2732 ( .A(n2767), .B(n2776), .Z(n2769) );
  XNOR U2733 ( .A(n2778), .B(n2779), .Z(n2767) );
  AND U2734 ( .A(n299), .B(n2780), .Z(n2779) );
  XOR U2735 ( .A(p_input[203]), .B(n2778), .Z(n2780) );
  XOR U2736 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n2781), 
        .Z(n2778) );
  AND U2737 ( .A(n302), .B(n2782), .Z(n2781) );
  XOR U2738 ( .A(n2783), .B(n2784), .Z(n2776) );
  AND U2739 ( .A(n306), .B(n2775), .Z(n2784) );
  XNOR U2740 ( .A(n2785), .B(n2773), .Z(n2775) );
  XOR U2741 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n2786), .Z(n2773) );
  AND U2742 ( .A(n318), .B(n2787), .Z(n2786) );
  IV U2743 ( .A(n2783), .Z(n2785) );
  XOR U2744 ( .A(n2788), .B(n2789), .Z(n2783) );
  AND U2745 ( .A(n313), .B(n2782), .Z(n2789) );
  XOR U2746 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n2788), 
        .Z(n2782) );
  XOR U2747 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n2790), 
        .Z(n2788) );
  AND U2748 ( .A(n315), .B(n2787), .Z(n2790) );
  XOR U2749 ( .A(n2791), .B(n2792), .Z(n2787) );
  IV U2750 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n2792) );
  IV U2751 ( .A(\knn_comb_/min_val_out[0][11] ), .Z(n2791) );
  XOR U2752 ( .A(n59), .B(n2793), .Z(o[10]) );
  AND U2753 ( .A(n62), .B(n2794), .Z(n59) );
  XOR U2754 ( .A(n60), .B(n2793), .Z(n2794) );
  XOR U2755 ( .A(n2795), .B(n2796), .Z(n2793) );
  AND U2756 ( .A(n82), .B(n2797), .Z(n2796) );
  XOR U2757 ( .A(n2798), .B(n23), .Z(n60) );
  AND U2758 ( .A(n65), .B(n2799), .Z(n23) );
  XOR U2759 ( .A(n24), .B(n2798), .Z(n2799) );
  XOR U2760 ( .A(n2800), .B(n2801), .Z(n24) );
  AND U2761 ( .A(n70), .B(n2802), .Z(n2801) );
  XOR U2762 ( .A(p_input[10]), .B(n2800), .Z(n2802) );
  XNOR U2763 ( .A(n2803), .B(n2804), .Z(n2800) );
  AND U2764 ( .A(n74), .B(n2805), .Z(n2804) );
  XOR U2765 ( .A(n2806), .B(n2807), .Z(n2798) );
  AND U2766 ( .A(n78), .B(n2797), .Z(n2807) );
  XNOR U2767 ( .A(n2808), .B(n2795), .Z(n2797) );
  XOR U2768 ( .A(n2809), .B(n2810), .Z(n2795) );
  AND U2769 ( .A(n102), .B(n2811), .Z(n2810) );
  IV U2770 ( .A(n2806), .Z(n2808) );
  XOR U2771 ( .A(n2812), .B(n2813), .Z(n2806) );
  AND U2772 ( .A(n86), .B(n2805), .Z(n2813) );
  XNOR U2773 ( .A(n2803), .B(n2812), .Z(n2805) );
  XNOR U2774 ( .A(n2814), .B(n2815), .Z(n2803) );
  AND U2775 ( .A(n90), .B(n2816), .Z(n2815) );
  XOR U2776 ( .A(p_input[26]), .B(n2814), .Z(n2816) );
  XNOR U2777 ( .A(n2817), .B(n2818), .Z(n2814) );
  AND U2778 ( .A(n94), .B(n2819), .Z(n2818) );
  XOR U2779 ( .A(n2820), .B(n2821), .Z(n2812) );
  AND U2780 ( .A(n98), .B(n2811), .Z(n2821) );
  XNOR U2781 ( .A(n2822), .B(n2809), .Z(n2811) );
  XOR U2782 ( .A(n2823), .B(n2824), .Z(n2809) );
  AND U2783 ( .A(n121), .B(n2825), .Z(n2824) );
  IV U2784 ( .A(n2820), .Z(n2822) );
  XOR U2785 ( .A(n2826), .B(n2827), .Z(n2820) );
  AND U2786 ( .A(n105), .B(n2819), .Z(n2827) );
  XNOR U2787 ( .A(n2817), .B(n2826), .Z(n2819) );
  XNOR U2788 ( .A(n2828), .B(n2829), .Z(n2817) );
  AND U2789 ( .A(n109), .B(n2830), .Z(n2829) );
  XOR U2790 ( .A(p_input[42]), .B(n2828), .Z(n2830) );
  XNOR U2791 ( .A(n2831), .B(n2832), .Z(n2828) );
  AND U2792 ( .A(n113), .B(n2833), .Z(n2832) );
  XOR U2793 ( .A(n2834), .B(n2835), .Z(n2826) );
  AND U2794 ( .A(n117), .B(n2825), .Z(n2835) );
  XNOR U2795 ( .A(n2836), .B(n2823), .Z(n2825) );
  XOR U2796 ( .A(n2837), .B(n2838), .Z(n2823) );
  AND U2797 ( .A(n140), .B(n2839), .Z(n2838) );
  IV U2798 ( .A(n2834), .Z(n2836) );
  XOR U2799 ( .A(n2840), .B(n2841), .Z(n2834) );
  AND U2800 ( .A(n124), .B(n2833), .Z(n2841) );
  XNOR U2801 ( .A(n2831), .B(n2840), .Z(n2833) );
  XNOR U2802 ( .A(n2842), .B(n2843), .Z(n2831) );
  AND U2803 ( .A(n128), .B(n2844), .Z(n2843) );
  XOR U2804 ( .A(p_input[58]), .B(n2842), .Z(n2844) );
  XNOR U2805 ( .A(n2845), .B(n2846), .Z(n2842) );
  AND U2806 ( .A(n132), .B(n2847), .Z(n2846) );
  XOR U2807 ( .A(n2848), .B(n2849), .Z(n2840) );
  AND U2808 ( .A(n136), .B(n2839), .Z(n2849) );
  XNOR U2809 ( .A(n2850), .B(n2837), .Z(n2839) );
  XOR U2810 ( .A(n2851), .B(n2852), .Z(n2837) );
  AND U2811 ( .A(n159), .B(n2853), .Z(n2852) );
  IV U2812 ( .A(n2848), .Z(n2850) );
  XOR U2813 ( .A(n2854), .B(n2855), .Z(n2848) );
  AND U2814 ( .A(n143), .B(n2847), .Z(n2855) );
  XNOR U2815 ( .A(n2845), .B(n2854), .Z(n2847) );
  XNOR U2816 ( .A(n2856), .B(n2857), .Z(n2845) );
  AND U2817 ( .A(n147), .B(n2858), .Z(n2857) );
  XOR U2818 ( .A(p_input[74]), .B(n2856), .Z(n2858) );
  XNOR U2819 ( .A(n2859), .B(n2860), .Z(n2856) );
  AND U2820 ( .A(n151), .B(n2861), .Z(n2860) );
  XOR U2821 ( .A(n2862), .B(n2863), .Z(n2854) );
  AND U2822 ( .A(n155), .B(n2853), .Z(n2863) );
  XNOR U2823 ( .A(n2864), .B(n2851), .Z(n2853) );
  XOR U2824 ( .A(n2865), .B(n2866), .Z(n2851) );
  AND U2825 ( .A(n178), .B(n2867), .Z(n2866) );
  IV U2826 ( .A(n2862), .Z(n2864) );
  XOR U2827 ( .A(n2868), .B(n2869), .Z(n2862) );
  AND U2828 ( .A(n162), .B(n2861), .Z(n2869) );
  XNOR U2829 ( .A(n2859), .B(n2868), .Z(n2861) );
  XNOR U2830 ( .A(n2870), .B(n2871), .Z(n2859) );
  AND U2831 ( .A(n166), .B(n2872), .Z(n2871) );
  XOR U2832 ( .A(p_input[90]), .B(n2870), .Z(n2872) );
  XNOR U2833 ( .A(n2873), .B(n2874), .Z(n2870) );
  AND U2834 ( .A(n170), .B(n2875), .Z(n2874) );
  XOR U2835 ( .A(n2876), .B(n2877), .Z(n2868) );
  AND U2836 ( .A(n174), .B(n2867), .Z(n2877) );
  XNOR U2837 ( .A(n2878), .B(n2865), .Z(n2867) );
  XOR U2838 ( .A(n2879), .B(n2880), .Z(n2865) );
  AND U2839 ( .A(n197), .B(n2881), .Z(n2880) );
  IV U2840 ( .A(n2876), .Z(n2878) );
  XOR U2841 ( .A(n2882), .B(n2883), .Z(n2876) );
  AND U2842 ( .A(n181), .B(n2875), .Z(n2883) );
  XNOR U2843 ( .A(n2873), .B(n2882), .Z(n2875) );
  XNOR U2844 ( .A(n2884), .B(n2885), .Z(n2873) );
  AND U2845 ( .A(n185), .B(n2886), .Z(n2885) );
  XOR U2846 ( .A(p_input[106]), .B(n2884), .Z(n2886) );
  XNOR U2847 ( .A(n2887), .B(n2888), .Z(n2884) );
  AND U2848 ( .A(n189), .B(n2889), .Z(n2888) );
  XOR U2849 ( .A(n2890), .B(n2891), .Z(n2882) );
  AND U2850 ( .A(n193), .B(n2881), .Z(n2891) );
  XNOR U2851 ( .A(n2892), .B(n2879), .Z(n2881) );
  XOR U2852 ( .A(n2893), .B(n2894), .Z(n2879) );
  AND U2853 ( .A(n216), .B(n2895), .Z(n2894) );
  IV U2854 ( .A(n2890), .Z(n2892) );
  XOR U2855 ( .A(n2896), .B(n2897), .Z(n2890) );
  AND U2856 ( .A(n200), .B(n2889), .Z(n2897) );
  XNOR U2857 ( .A(n2887), .B(n2896), .Z(n2889) );
  XNOR U2858 ( .A(n2898), .B(n2899), .Z(n2887) );
  AND U2859 ( .A(n204), .B(n2900), .Z(n2899) );
  XOR U2860 ( .A(p_input[122]), .B(n2898), .Z(n2900) );
  XNOR U2861 ( .A(n2901), .B(n2902), .Z(n2898) );
  AND U2862 ( .A(n208), .B(n2903), .Z(n2902) );
  XOR U2863 ( .A(n2904), .B(n2905), .Z(n2896) );
  AND U2864 ( .A(n212), .B(n2895), .Z(n2905) );
  XNOR U2865 ( .A(n2906), .B(n2893), .Z(n2895) );
  XOR U2866 ( .A(n2907), .B(n2908), .Z(n2893) );
  AND U2867 ( .A(n235), .B(n2909), .Z(n2908) );
  IV U2868 ( .A(n2904), .Z(n2906) );
  XOR U2869 ( .A(n2910), .B(n2911), .Z(n2904) );
  AND U2870 ( .A(n219), .B(n2903), .Z(n2911) );
  XNOR U2871 ( .A(n2901), .B(n2910), .Z(n2903) );
  XNOR U2872 ( .A(n2912), .B(n2913), .Z(n2901) );
  AND U2873 ( .A(n223), .B(n2914), .Z(n2913) );
  XOR U2874 ( .A(p_input[138]), .B(n2912), .Z(n2914) );
  XNOR U2875 ( .A(n2915), .B(n2916), .Z(n2912) );
  AND U2876 ( .A(n227), .B(n2917), .Z(n2916) );
  XOR U2877 ( .A(n2918), .B(n2919), .Z(n2910) );
  AND U2878 ( .A(n231), .B(n2909), .Z(n2919) );
  XNOR U2879 ( .A(n2920), .B(n2907), .Z(n2909) );
  XOR U2880 ( .A(n2921), .B(n2922), .Z(n2907) );
  AND U2881 ( .A(n254), .B(n2923), .Z(n2922) );
  IV U2882 ( .A(n2918), .Z(n2920) );
  XOR U2883 ( .A(n2924), .B(n2925), .Z(n2918) );
  AND U2884 ( .A(n238), .B(n2917), .Z(n2925) );
  XNOR U2885 ( .A(n2915), .B(n2924), .Z(n2917) );
  XNOR U2886 ( .A(n2926), .B(n2927), .Z(n2915) );
  AND U2887 ( .A(n242), .B(n2928), .Z(n2927) );
  XOR U2888 ( .A(p_input[154]), .B(n2926), .Z(n2928) );
  XNOR U2889 ( .A(n2929), .B(n2930), .Z(n2926) );
  AND U2890 ( .A(n246), .B(n2931), .Z(n2930) );
  XOR U2891 ( .A(n2932), .B(n2933), .Z(n2924) );
  AND U2892 ( .A(n250), .B(n2923), .Z(n2933) );
  XNOR U2893 ( .A(n2934), .B(n2921), .Z(n2923) );
  XOR U2894 ( .A(n2935), .B(n2936), .Z(n2921) );
  AND U2895 ( .A(n273), .B(n2937), .Z(n2936) );
  IV U2896 ( .A(n2932), .Z(n2934) );
  XOR U2897 ( .A(n2938), .B(n2939), .Z(n2932) );
  AND U2898 ( .A(n257), .B(n2931), .Z(n2939) );
  XNOR U2899 ( .A(n2929), .B(n2938), .Z(n2931) );
  XNOR U2900 ( .A(n2940), .B(n2941), .Z(n2929) );
  AND U2901 ( .A(n261), .B(n2942), .Z(n2941) );
  XOR U2902 ( .A(p_input[170]), .B(n2940), .Z(n2942) );
  XNOR U2903 ( .A(n2943), .B(n2944), .Z(n2940) );
  AND U2904 ( .A(n265), .B(n2945), .Z(n2944) );
  XOR U2905 ( .A(n2946), .B(n2947), .Z(n2938) );
  AND U2906 ( .A(n269), .B(n2937), .Z(n2947) );
  XNOR U2907 ( .A(n2948), .B(n2935), .Z(n2937) );
  XOR U2908 ( .A(n2949), .B(n2950), .Z(n2935) );
  AND U2909 ( .A(n292), .B(n2951), .Z(n2950) );
  IV U2910 ( .A(n2946), .Z(n2948) );
  XOR U2911 ( .A(n2952), .B(n2953), .Z(n2946) );
  AND U2912 ( .A(n276), .B(n2945), .Z(n2953) );
  XNOR U2913 ( .A(n2943), .B(n2952), .Z(n2945) );
  XNOR U2914 ( .A(n2954), .B(n2955), .Z(n2943) );
  AND U2915 ( .A(n280), .B(n2956), .Z(n2955) );
  XOR U2916 ( .A(p_input[186]), .B(n2954), .Z(n2956) );
  XNOR U2917 ( .A(n2957), .B(n2958), .Z(n2954) );
  AND U2918 ( .A(n284), .B(n2959), .Z(n2958) );
  XOR U2919 ( .A(n2960), .B(n2961), .Z(n2952) );
  AND U2920 ( .A(n288), .B(n2951), .Z(n2961) );
  XNOR U2921 ( .A(n2962), .B(n2949), .Z(n2951) );
  XOR U2922 ( .A(n2963), .B(n2964), .Z(n2949) );
  AND U2923 ( .A(n310), .B(n2965), .Z(n2964) );
  IV U2924 ( .A(n2960), .Z(n2962) );
  XOR U2925 ( .A(n2966), .B(n2967), .Z(n2960) );
  AND U2926 ( .A(n295), .B(n2959), .Z(n2967) );
  XNOR U2927 ( .A(n2957), .B(n2966), .Z(n2959) );
  XNOR U2928 ( .A(n2968), .B(n2969), .Z(n2957) );
  AND U2929 ( .A(n299), .B(n2970), .Z(n2969) );
  XOR U2930 ( .A(p_input[202]), .B(n2968), .Z(n2970) );
  XOR U2931 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n2971), 
        .Z(n2968) );
  AND U2932 ( .A(n302), .B(n2972), .Z(n2971) );
  XOR U2933 ( .A(n2973), .B(n2974), .Z(n2966) );
  AND U2934 ( .A(n306), .B(n2965), .Z(n2974) );
  XNOR U2935 ( .A(n2975), .B(n2963), .Z(n2965) );
  XOR U2936 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n2976), .Z(n2963) );
  AND U2937 ( .A(n318), .B(n2977), .Z(n2976) );
  IV U2938 ( .A(n2973), .Z(n2975) );
  XOR U2939 ( .A(n2978), .B(n2979), .Z(n2973) );
  AND U2940 ( .A(n313), .B(n2972), .Z(n2979) );
  XOR U2941 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n2978), 
        .Z(n2972) );
  XOR U2942 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(n2980), 
        .Z(n2978) );
  AND U2943 ( .A(n315), .B(n2977), .Z(n2980) );
  XOR U2944 ( .A(\knn_comb_/min_val_out[0][10] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n2977) );
  XOR U2945 ( .A(n1845), .B(n2981), .Z(o[0]) );
  AND U2946 ( .A(n62), .B(n2982), .Z(n1845) );
  XOR U2947 ( .A(n1846), .B(n2981), .Z(n2982) );
  XOR U2948 ( .A(n2983), .B(n2984), .Z(n2981) );
  AND U2949 ( .A(n82), .B(n2985), .Z(n2984) );
  XOR U2950 ( .A(n2986), .B(n45), .Z(n1846) );
  AND U2951 ( .A(n65), .B(n2987), .Z(n45) );
  XOR U2952 ( .A(n46), .B(n2986), .Z(n2987) );
  XOR U2953 ( .A(n2988), .B(n2989), .Z(n46) );
  AND U2954 ( .A(n70), .B(n2990), .Z(n2989) );
  XOR U2955 ( .A(p_input[0]), .B(n2988), .Z(n2990) );
  XNOR U2956 ( .A(n2991), .B(n2992), .Z(n2988) );
  AND U2957 ( .A(n74), .B(n2993), .Z(n2992) );
  XOR U2958 ( .A(n2994), .B(n2995), .Z(n2986) );
  AND U2959 ( .A(n78), .B(n2985), .Z(n2995) );
  XNOR U2960 ( .A(n2996), .B(n2983), .Z(n2985) );
  XOR U2961 ( .A(n2997), .B(n2998), .Z(n2983) );
  AND U2962 ( .A(n102), .B(n2999), .Z(n2998) );
  IV U2963 ( .A(n2994), .Z(n2996) );
  XOR U2964 ( .A(n3000), .B(n3001), .Z(n2994) );
  AND U2965 ( .A(n86), .B(n2993), .Z(n3001) );
  XNOR U2966 ( .A(n2991), .B(n3000), .Z(n2993) );
  XNOR U2967 ( .A(n3002), .B(n3003), .Z(n2991) );
  AND U2968 ( .A(n90), .B(n3004), .Z(n3003) );
  XOR U2969 ( .A(p_input[16]), .B(n3002), .Z(n3004) );
  XNOR U2970 ( .A(n3005), .B(n3006), .Z(n3002) );
  AND U2971 ( .A(n94), .B(n3007), .Z(n3006) );
  XOR U2972 ( .A(n3008), .B(n3009), .Z(n3000) );
  AND U2973 ( .A(n98), .B(n2999), .Z(n3009) );
  XNOR U2974 ( .A(n3010), .B(n2997), .Z(n2999) );
  XOR U2975 ( .A(n3011), .B(n3012), .Z(n2997) );
  AND U2976 ( .A(n121), .B(n3013), .Z(n3012) );
  IV U2977 ( .A(n3008), .Z(n3010) );
  XOR U2978 ( .A(n3014), .B(n3015), .Z(n3008) );
  AND U2979 ( .A(n105), .B(n3007), .Z(n3015) );
  XNOR U2980 ( .A(n3005), .B(n3014), .Z(n3007) );
  XNOR U2981 ( .A(n3016), .B(n3017), .Z(n3005) );
  AND U2982 ( .A(n109), .B(n3018), .Z(n3017) );
  XOR U2983 ( .A(p_input[32]), .B(n3016), .Z(n3018) );
  XNOR U2984 ( .A(n3019), .B(n3020), .Z(n3016) );
  AND U2985 ( .A(n113), .B(n3021), .Z(n3020) );
  XOR U2986 ( .A(n3022), .B(n3023), .Z(n3014) );
  AND U2987 ( .A(n117), .B(n3013), .Z(n3023) );
  XNOR U2988 ( .A(n3024), .B(n3011), .Z(n3013) );
  XOR U2989 ( .A(n3025), .B(n3026), .Z(n3011) );
  AND U2990 ( .A(n140), .B(n3027), .Z(n3026) );
  IV U2991 ( .A(n3022), .Z(n3024) );
  XOR U2992 ( .A(n3028), .B(n3029), .Z(n3022) );
  AND U2993 ( .A(n124), .B(n3021), .Z(n3029) );
  XNOR U2994 ( .A(n3019), .B(n3028), .Z(n3021) );
  XNOR U2995 ( .A(n3030), .B(n3031), .Z(n3019) );
  AND U2996 ( .A(n128), .B(n3032), .Z(n3031) );
  XOR U2997 ( .A(p_input[48]), .B(n3030), .Z(n3032) );
  XNOR U2998 ( .A(n3033), .B(n3034), .Z(n3030) );
  AND U2999 ( .A(n132), .B(n3035), .Z(n3034) );
  XOR U3000 ( .A(n3036), .B(n3037), .Z(n3028) );
  AND U3001 ( .A(n136), .B(n3027), .Z(n3037) );
  XNOR U3002 ( .A(n3038), .B(n3025), .Z(n3027) );
  XOR U3003 ( .A(n3039), .B(n3040), .Z(n3025) );
  AND U3004 ( .A(n159), .B(n3041), .Z(n3040) );
  IV U3005 ( .A(n3036), .Z(n3038) );
  XOR U3006 ( .A(n3042), .B(n3043), .Z(n3036) );
  AND U3007 ( .A(n143), .B(n3035), .Z(n3043) );
  XNOR U3008 ( .A(n3033), .B(n3042), .Z(n3035) );
  XNOR U3009 ( .A(n3044), .B(n3045), .Z(n3033) );
  AND U3010 ( .A(n147), .B(n3046), .Z(n3045) );
  XOR U3011 ( .A(p_input[64]), .B(n3044), .Z(n3046) );
  XNOR U3012 ( .A(n3047), .B(n3048), .Z(n3044) );
  AND U3013 ( .A(n151), .B(n3049), .Z(n3048) );
  XOR U3014 ( .A(n3050), .B(n3051), .Z(n3042) );
  AND U3015 ( .A(n155), .B(n3041), .Z(n3051) );
  XNOR U3016 ( .A(n3052), .B(n3039), .Z(n3041) );
  XOR U3017 ( .A(n3053), .B(n3054), .Z(n3039) );
  AND U3018 ( .A(n178), .B(n3055), .Z(n3054) );
  IV U3019 ( .A(n3050), .Z(n3052) );
  XOR U3020 ( .A(n3056), .B(n3057), .Z(n3050) );
  AND U3021 ( .A(n162), .B(n3049), .Z(n3057) );
  XNOR U3022 ( .A(n3047), .B(n3056), .Z(n3049) );
  XNOR U3023 ( .A(n3058), .B(n3059), .Z(n3047) );
  AND U3024 ( .A(n166), .B(n3060), .Z(n3059) );
  XOR U3025 ( .A(p_input[80]), .B(n3058), .Z(n3060) );
  XNOR U3026 ( .A(n3061), .B(n3062), .Z(n3058) );
  AND U3027 ( .A(n170), .B(n3063), .Z(n3062) );
  XOR U3028 ( .A(n3064), .B(n3065), .Z(n3056) );
  AND U3029 ( .A(n174), .B(n3055), .Z(n3065) );
  XNOR U3030 ( .A(n3066), .B(n3053), .Z(n3055) );
  XOR U3031 ( .A(n3067), .B(n3068), .Z(n3053) );
  AND U3032 ( .A(n197), .B(n3069), .Z(n3068) );
  IV U3033 ( .A(n3064), .Z(n3066) );
  XOR U3034 ( .A(n3070), .B(n3071), .Z(n3064) );
  AND U3035 ( .A(n181), .B(n3063), .Z(n3071) );
  XNOR U3036 ( .A(n3061), .B(n3070), .Z(n3063) );
  XNOR U3037 ( .A(n3072), .B(n3073), .Z(n3061) );
  AND U3038 ( .A(n185), .B(n3074), .Z(n3073) );
  XOR U3039 ( .A(p_input[96]), .B(n3072), .Z(n3074) );
  XNOR U3040 ( .A(n3075), .B(n3076), .Z(n3072) );
  AND U3041 ( .A(n189), .B(n3077), .Z(n3076) );
  XOR U3042 ( .A(n3078), .B(n3079), .Z(n3070) );
  AND U3043 ( .A(n193), .B(n3069), .Z(n3079) );
  XNOR U3044 ( .A(n3080), .B(n3067), .Z(n3069) );
  XOR U3045 ( .A(n3081), .B(n3082), .Z(n3067) );
  AND U3046 ( .A(n216), .B(n3083), .Z(n3082) );
  IV U3047 ( .A(n3078), .Z(n3080) );
  XOR U3048 ( .A(n3084), .B(n3085), .Z(n3078) );
  AND U3049 ( .A(n200), .B(n3077), .Z(n3085) );
  XNOR U3050 ( .A(n3075), .B(n3084), .Z(n3077) );
  XNOR U3051 ( .A(n3086), .B(n3087), .Z(n3075) );
  AND U3052 ( .A(n204), .B(n3088), .Z(n3087) );
  XOR U3053 ( .A(p_input[112]), .B(n3086), .Z(n3088) );
  XNOR U3054 ( .A(n3089), .B(n3090), .Z(n3086) );
  AND U3055 ( .A(n208), .B(n3091), .Z(n3090) );
  XOR U3056 ( .A(n3092), .B(n3093), .Z(n3084) );
  AND U3057 ( .A(n212), .B(n3083), .Z(n3093) );
  XNOR U3058 ( .A(n3094), .B(n3081), .Z(n3083) );
  XOR U3059 ( .A(n3095), .B(n3096), .Z(n3081) );
  AND U3060 ( .A(n235), .B(n3097), .Z(n3096) );
  IV U3061 ( .A(n3092), .Z(n3094) );
  XOR U3062 ( .A(n3098), .B(n3099), .Z(n3092) );
  AND U3063 ( .A(n219), .B(n3091), .Z(n3099) );
  XNOR U3064 ( .A(n3089), .B(n3098), .Z(n3091) );
  XNOR U3065 ( .A(n3100), .B(n3101), .Z(n3089) );
  AND U3066 ( .A(n223), .B(n3102), .Z(n3101) );
  XOR U3067 ( .A(p_input[128]), .B(n3100), .Z(n3102) );
  XNOR U3068 ( .A(n3103), .B(n3104), .Z(n3100) );
  AND U3069 ( .A(n227), .B(n3105), .Z(n3104) );
  XOR U3070 ( .A(n3106), .B(n3107), .Z(n3098) );
  AND U3071 ( .A(n231), .B(n3097), .Z(n3107) );
  XNOR U3072 ( .A(n3108), .B(n3095), .Z(n3097) );
  XOR U3073 ( .A(n3109), .B(n3110), .Z(n3095) );
  AND U3074 ( .A(n254), .B(n3111), .Z(n3110) );
  IV U3075 ( .A(n3106), .Z(n3108) );
  XOR U3076 ( .A(n3112), .B(n3113), .Z(n3106) );
  AND U3077 ( .A(n238), .B(n3105), .Z(n3113) );
  XNOR U3078 ( .A(n3103), .B(n3112), .Z(n3105) );
  XNOR U3079 ( .A(n3114), .B(n3115), .Z(n3103) );
  AND U3080 ( .A(n242), .B(n3116), .Z(n3115) );
  XOR U3081 ( .A(p_input[144]), .B(n3114), .Z(n3116) );
  XNOR U3082 ( .A(n3117), .B(n3118), .Z(n3114) );
  AND U3083 ( .A(n246), .B(n3119), .Z(n3118) );
  XOR U3084 ( .A(n3120), .B(n3121), .Z(n3112) );
  AND U3085 ( .A(n250), .B(n3111), .Z(n3121) );
  XNOR U3086 ( .A(n3122), .B(n3109), .Z(n3111) );
  XOR U3087 ( .A(n3123), .B(n3124), .Z(n3109) );
  AND U3088 ( .A(n273), .B(n3125), .Z(n3124) );
  IV U3089 ( .A(n3120), .Z(n3122) );
  XOR U3090 ( .A(n3126), .B(n3127), .Z(n3120) );
  AND U3091 ( .A(n257), .B(n3119), .Z(n3127) );
  XNOR U3092 ( .A(n3117), .B(n3126), .Z(n3119) );
  XNOR U3093 ( .A(n3128), .B(n3129), .Z(n3117) );
  AND U3094 ( .A(n261), .B(n3130), .Z(n3129) );
  XOR U3095 ( .A(p_input[160]), .B(n3128), .Z(n3130) );
  XNOR U3096 ( .A(n3131), .B(n3132), .Z(n3128) );
  AND U3097 ( .A(n265), .B(n3133), .Z(n3132) );
  XOR U3098 ( .A(n3134), .B(n3135), .Z(n3126) );
  AND U3099 ( .A(n269), .B(n3125), .Z(n3135) );
  XNOR U3100 ( .A(n3136), .B(n3123), .Z(n3125) );
  XOR U3101 ( .A(n3137), .B(n3138), .Z(n3123) );
  AND U3102 ( .A(n292), .B(n3139), .Z(n3138) );
  IV U3103 ( .A(n3134), .Z(n3136) );
  XOR U3104 ( .A(n3140), .B(n3141), .Z(n3134) );
  AND U3105 ( .A(n276), .B(n3133), .Z(n3141) );
  XNOR U3106 ( .A(n3131), .B(n3140), .Z(n3133) );
  XNOR U3107 ( .A(n3142), .B(n3143), .Z(n3131) );
  AND U3108 ( .A(n280), .B(n3144), .Z(n3143) );
  XOR U3109 ( .A(p_input[176]), .B(n3142), .Z(n3144) );
  XNOR U3110 ( .A(n3145), .B(n3146), .Z(n3142) );
  AND U3111 ( .A(n284), .B(n3147), .Z(n3146) );
  XOR U3112 ( .A(n3148), .B(n3149), .Z(n3140) );
  AND U3113 ( .A(n288), .B(n3139), .Z(n3149) );
  XNOR U3114 ( .A(n3150), .B(n3137), .Z(n3139) );
  XOR U3115 ( .A(n3151), .B(n3152), .Z(n3137) );
  AND U3116 ( .A(n310), .B(n3153), .Z(n3152) );
  IV U3117 ( .A(n3148), .Z(n3150) );
  XOR U3118 ( .A(n3154), .B(n3155), .Z(n3148) );
  AND U3119 ( .A(n295), .B(n3147), .Z(n3155) );
  XNOR U3120 ( .A(n3145), .B(n3154), .Z(n3147) );
  XNOR U3121 ( .A(n3156), .B(n3157), .Z(n3145) );
  AND U3122 ( .A(n299), .B(n3158), .Z(n3157) );
  XOR U3123 ( .A(p_input[192]), .B(n3156), .Z(n3158) );
  XOR U3124 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(n3159), 
        .Z(n3156) );
  AND U3125 ( .A(n302), .B(n3160), .Z(n3159) );
  XOR U3126 ( .A(n3161), .B(n3162), .Z(n3154) );
  AND U3127 ( .A(n306), .B(n3153), .Z(n3162) );
  XNOR U3128 ( .A(n3163), .B(n3151), .Z(n3153) );
  XOR U3129 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n3164), .Z(n3151) );
  AND U3130 ( .A(n318), .B(n3165), .Z(n3164) );
  IV U3131 ( .A(n3161), .Z(n3163) );
  XOR U3132 ( .A(n3166), .B(n3167), .Z(n3161) );
  AND U3133 ( .A(n313), .B(n3160), .Z(n3167) );
  XOR U3134 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(n3166), 
        .Z(n3160) );
  XOR U3135 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(n3168), 
        .Z(n3166) );
  AND U3136 ( .A(n315), .B(n3165), .Z(n3168) );
  XOR U3137 ( .A(\knn_comb_/min_val_out[0][0] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n3165) );
  XNOR U3138 ( .A(n3169), .B(n3170), .Z(n62) );
  AND U3139 ( .A(n3171), .B(n3172), .Z(n3170) );
  XNOR U3140 ( .A(n3169), .B(n3173), .Z(n3172) );
  XOR U3141 ( .A(n3174), .B(n3175), .Z(n3173) );
  AND U3142 ( .A(n65), .B(n3176), .Z(n3175) );
  XNOR U3143 ( .A(n3174), .B(n3177), .Z(n3176) );
  IV U3144 ( .A(n3178), .Z(n3174) );
  XNOR U3145 ( .A(n3169), .B(n3179), .Z(n3171) );
  XOR U3146 ( .A(n3180), .B(n3181), .Z(n3179) );
  AND U3147 ( .A(n82), .B(n3182), .Z(n3181) );
  XOR U3148 ( .A(n3183), .B(n3184), .Z(n3169) );
  AND U3149 ( .A(n3185), .B(n3186), .Z(n3184) );
  XOR U3150 ( .A(n3187), .B(n3183), .Z(n3186) );
  XNOR U3151 ( .A(n3188), .B(n3189), .Z(n3187) );
  AND U3152 ( .A(n65), .B(n3190), .Z(n3189) );
  XNOR U3153 ( .A(n3191), .B(n3188), .Z(n3190) );
  XNOR U3154 ( .A(n3183), .B(n3192), .Z(n3185) );
  XOR U3155 ( .A(n3193), .B(n3194), .Z(n3192) );
  AND U3156 ( .A(n82), .B(n3195), .Z(n3194) );
  XOR U3157 ( .A(n3196), .B(n3197), .Z(n3183) );
  AND U3158 ( .A(n3198), .B(n3199), .Z(n3197) );
  XOR U3159 ( .A(n3200), .B(n3196), .Z(n3199) );
  XNOR U3160 ( .A(n3201), .B(n3202), .Z(n3200) );
  AND U3161 ( .A(n65), .B(n3203), .Z(n3202) );
  XNOR U3162 ( .A(n3204), .B(n3201), .Z(n3203) );
  XNOR U3163 ( .A(n3196), .B(n3205), .Z(n3198) );
  XOR U3164 ( .A(n3206), .B(n3207), .Z(n3205) );
  AND U3165 ( .A(n82), .B(n3208), .Z(n3207) );
  XOR U3166 ( .A(n3209), .B(n3210), .Z(n3196) );
  AND U3167 ( .A(n3211), .B(n3212), .Z(n3210) );
  XOR U3168 ( .A(n3209), .B(n3213), .Z(n3212) );
  XOR U3169 ( .A(n3214), .B(n3215), .Z(n3213) );
  AND U3170 ( .A(n65), .B(n3216), .Z(n3215) );
  XOR U3171 ( .A(n3217), .B(n3214), .Z(n3216) );
  XNOR U3172 ( .A(n3218), .B(n3209), .Z(n3211) );
  XNOR U3173 ( .A(n3219), .B(n3220), .Z(n3218) );
  AND U3174 ( .A(n82), .B(n3221), .Z(n3220) );
  AND U3175 ( .A(n3222), .B(n3223), .Z(n3209) );
  XNOR U3176 ( .A(n3224), .B(n3225), .Z(n3223) );
  AND U3177 ( .A(n65), .B(n3226), .Z(n3225) );
  XNOR U3178 ( .A(n3227), .B(n3224), .Z(n3226) );
  XNOR U3179 ( .A(n3228), .B(n3229), .Z(n65) );
  AND U3180 ( .A(n3230), .B(n3231), .Z(n3229) );
  XOR U3181 ( .A(n3177), .B(n3228), .Z(n3231) );
  XOR U3182 ( .A(n3232), .B(n3233), .Z(n3177) );
  AND U3183 ( .A(n70), .B(n3234), .Z(n3233) );
  XOR U3184 ( .A(n3235), .B(n3232), .Z(n3234) );
  XNOR U3185 ( .A(n3178), .B(n3228), .Z(n3230) );
  XOR U3186 ( .A(n3236), .B(n3237), .Z(n3178) );
  AND U3187 ( .A(n78), .B(n3182), .Z(n3237) );
  XOR U3188 ( .A(n3180), .B(n3236), .Z(n3182) );
  XOR U3189 ( .A(n3238), .B(n3239), .Z(n3228) );
  AND U3190 ( .A(n3240), .B(n3241), .Z(n3239) );
  XOR U3191 ( .A(n3191), .B(n3238), .Z(n3241) );
  XOR U3192 ( .A(n3242), .B(n3243), .Z(n3191) );
  AND U3193 ( .A(n70), .B(n3244), .Z(n3243) );
  XOR U3194 ( .A(n3245), .B(n3242), .Z(n3244) );
  XOR U3195 ( .A(n3238), .B(n3188), .Z(n3240) );
  XOR U3196 ( .A(n3246), .B(n3247), .Z(n3188) );
  AND U3197 ( .A(n78), .B(n3195), .Z(n3247) );
  XOR U3198 ( .A(n3246), .B(n3248), .Z(n3195) );
  XOR U3199 ( .A(n3249), .B(n3250), .Z(n3238) );
  AND U3200 ( .A(n3251), .B(n3252), .Z(n3250) );
  XOR U3201 ( .A(n3204), .B(n3249), .Z(n3252) );
  XOR U3202 ( .A(n3253), .B(n3254), .Z(n3204) );
  AND U3203 ( .A(n70), .B(n3255), .Z(n3254) );
  XNOR U3204 ( .A(n3256), .B(n3253), .Z(n3255) );
  XOR U3205 ( .A(n3249), .B(n3201), .Z(n3251) );
  XOR U3206 ( .A(n3257), .B(n3258), .Z(n3201) );
  AND U3207 ( .A(n78), .B(n3208), .Z(n3258) );
  XOR U3208 ( .A(n3257), .B(n3259), .Z(n3208) );
  XOR U3209 ( .A(n3260), .B(n3261), .Z(n3249) );
  AND U3210 ( .A(n3262), .B(n3263), .Z(n3261) );
  XOR U3211 ( .A(n3260), .B(n3217), .Z(n3263) );
  XOR U3212 ( .A(n3264), .B(n3265), .Z(n3217) );
  AND U3213 ( .A(n70), .B(n3266), .Z(n3265) );
  XOR U3214 ( .A(n3267), .B(n3264), .Z(n3266) );
  XNOR U3215 ( .A(n3214), .B(n3260), .Z(n3262) );
  XNOR U3216 ( .A(n3268), .B(n3269), .Z(n3214) );
  AND U3217 ( .A(n78), .B(n3221), .Z(n3269) );
  XOR U3218 ( .A(n3268), .B(n3219), .Z(n3221) );
  AND U3219 ( .A(n3224), .B(n3227), .Z(n3260) );
  XOR U3220 ( .A(n3270), .B(n3271), .Z(n3227) );
  AND U3221 ( .A(n70), .B(n3272), .Z(n3271) );
  XNOR U3222 ( .A(n3273), .B(n3274), .Z(n3272) );
  XNOR U3223 ( .A(n3275), .B(n3276), .Z(n70) );
  AND U3224 ( .A(n3277), .B(n3278), .Z(n3276) );
  XOR U3225 ( .A(n3235), .B(n3275), .Z(n3278) );
  AND U3226 ( .A(n3279), .B(n3280), .Z(n3235) );
  XNOR U3227 ( .A(n3232), .B(n3275), .Z(n3277) );
  XNOR U3228 ( .A(n3281), .B(n3282), .Z(n3232) );
  AND U3229 ( .A(n74), .B(n3283), .Z(n3282) );
  XNOR U3230 ( .A(n3284), .B(n3285), .Z(n3283) );
  XOR U3231 ( .A(n3286), .B(n3287), .Z(n3275) );
  AND U3232 ( .A(n3288), .B(n3289), .Z(n3287) );
  XNOR U3233 ( .A(n3286), .B(n3279), .Z(n3289) );
  IV U3234 ( .A(n3245), .Z(n3279) );
  XOR U3235 ( .A(n3290), .B(n3291), .Z(n3245) );
  XOR U3236 ( .A(n3292), .B(n3280), .Z(n3291) );
  AND U3237 ( .A(n3256), .B(n3293), .Z(n3280) );
  AND U3238 ( .A(n3294), .B(n3295), .Z(n3292) );
  XOR U3239 ( .A(n3296), .B(n3290), .Z(n3294) );
  XNOR U3240 ( .A(n3242), .B(n3286), .Z(n3288) );
  XNOR U3241 ( .A(n3297), .B(n3298), .Z(n3242) );
  AND U3242 ( .A(n74), .B(n3299), .Z(n3298) );
  XNOR U3243 ( .A(n3300), .B(n3301), .Z(n3299) );
  XOR U3244 ( .A(n3302), .B(n3303), .Z(n3286) );
  AND U3245 ( .A(n3304), .B(n3305), .Z(n3303) );
  XNOR U3246 ( .A(n3302), .B(n3256), .Z(n3305) );
  XOR U3247 ( .A(n3306), .B(n3295), .Z(n3256) );
  XNOR U3248 ( .A(n3307), .B(n3290), .Z(n3295) );
  XOR U3249 ( .A(n3308), .B(n3309), .Z(n3290) );
  AND U3250 ( .A(n3310), .B(n3311), .Z(n3309) );
  XOR U3251 ( .A(n3312), .B(n3308), .Z(n3310) );
  XNOR U3252 ( .A(n3313), .B(n3314), .Z(n3307) );
  AND U3253 ( .A(n3315), .B(n3316), .Z(n3314) );
  XOR U3254 ( .A(n3313), .B(n3317), .Z(n3315) );
  XNOR U3255 ( .A(n3296), .B(n3293), .Z(n3306) );
  AND U3256 ( .A(n3318), .B(n3319), .Z(n3293) );
  XOR U3257 ( .A(n3320), .B(n3321), .Z(n3296) );
  AND U3258 ( .A(n3322), .B(n3323), .Z(n3321) );
  XOR U3259 ( .A(n3320), .B(n3324), .Z(n3322) );
  XNOR U3260 ( .A(n3253), .B(n3302), .Z(n3304) );
  XNOR U3261 ( .A(n3325), .B(n3326), .Z(n3253) );
  AND U3262 ( .A(n74), .B(n3327), .Z(n3326) );
  XNOR U3263 ( .A(n3328), .B(n3329), .Z(n3327) );
  XOR U3264 ( .A(n3330), .B(n3331), .Z(n3302) );
  AND U3265 ( .A(n3332), .B(n3333), .Z(n3331) );
  XNOR U3266 ( .A(n3330), .B(n3318), .Z(n3333) );
  IV U3267 ( .A(n3267), .Z(n3318) );
  XNOR U3268 ( .A(n3334), .B(n3311), .Z(n3267) );
  XNOR U3269 ( .A(n3335), .B(n3317), .Z(n3311) );
  XNOR U3270 ( .A(n3336), .B(n3337), .Z(n3317) );
  NOR U3271 ( .A(n3338), .B(n3339), .Z(n3337) );
  XOR U3272 ( .A(n3336), .B(n3340), .Z(n3338) );
  XNOR U3273 ( .A(n3316), .B(n3308), .Z(n3335) );
  XOR U3274 ( .A(n3341), .B(n3342), .Z(n3308) );
  AND U3275 ( .A(n3343), .B(n3344), .Z(n3342) );
  XNOR U3276 ( .A(n3341), .B(n3345), .Z(n3343) );
  XNOR U3277 ( .A(n3346), .B(n3313), .Z(n3316) );
  XOR U3278 ( .A(n3347), .B(n3348), .Z(n3313) );
  AND U3279 ( .A(n3349), .B(n3350), .Z(n3348) );
  XOR U3280 ( .A(n3347), .B(n3351), .Z(n3349) );
  XNOR U3281 ( .A(n3352), .B(n3353), .Z(n3346) );
  NOR U3282 ( .A(n3354), .B(n3355), .Z(n3353) );
  XNOR U3283 ( .A(n3352), .B(n3356), .Z(n3354) );
  XNOR U3284 ( .A(n3312), .B(n3319), .Z(n3334) );
  NOR U3285 ( .A(n3273), .B(n3357), .Z(n3319) );
  XOR U3286 ( .A(n3324), .B(n3323), .Z(n3312) );
  XNOR U3287 ( .A(n3358), .B(n3320), .Z(n3323) );
  XOR U3288 ( .A(n3359), .B(n3360), .Z(n3320) );
  AND U3289 ( .A(n3361), .B(n3362), .Z(n3360) );
  XOR U3290 ( .A(n3359), .B(n3363), .Z(n3361) );
  XNOR U3291 ( .A(n3364), .B(n3365), .Z(n3358) );
  NOR U3292 ( .A(n3366), .B(n3367), .Z(n3365) );
  XNOR U3293 ( .A(n3364), .B(n3368), .Z(n3366) );
  XOR U3294 ( .A(n3369), .B(n3370), .Z(n3324) );
  NOR U3295 ( .A(n3371), .B(n3372), .Z(n3370) );
  XNOR U3296 ( .A(n3369), .B(n3373), .Z(n3371) );
  XNOR U3297 ( .A(n3264), .B(n3330), .Z(n3332) );
  XNOR U3298 ( .A(n3374), .B(n3375), .Z(n3264) );
  AND U3299 ( .A(n74), .B(n3376), .Z(n3375) );
  XNOR U3300 ( .A(n3377), .B(n3378), .Z(n3376) );
  AND U3301 ( .A(n3274), .B(n3273), .Z(n3330) );
  XOR U3302 ( .A(n3379), .B(n3357), .Z(n3273) );
  XNOR U3303 ( .A(p_input[0]), .B(p_input[256]), .Z(n3357) );
  XOR U3304 ( .A(n3345), .B(n3344), .Z(n3379) );
  XNOR U3305 ( .A(n3380), .B(n3351), .Z(n3344) );
  XNOR U3306 ( .A(n3340), .B(n3339), .Z(n3351) );
  XNOR U3307 ( .A(n3381), .B(n3336), .Z(n3339) );
  XNOR U3308 ( .A(p_input[10]), .B(p_input[266]), .Z(n3336) );
  XOR U3309 ( .A(p_input[11]), .B(n3382), .Z(n3381) );
  XOR U3310 ( .A(p_input[12]), .B(p_input[268]), .Z(n3340) );
  XOR U3311 ( .A(n3350), .B(n3383), .Z(n3380) );
  IV U3312 ( .A(n3341), .Z(n3383) );
  XOR U3313 ( .A(p_input[1]), .B(p_input[257]), .Z(n3341) );
  XNOR U3314 ( .A(n3384), .B(n3356), .Z(n3350) );
  XNOR U3315 ( .A(p_input[15]), .B(n3385), .Z(n3356) );
  XOR U3316 ( .A(n3347), .B(n3355), .Z(n3384) );
  XOR U3317 ( .A(n3386), .B(n3352), .Z(n3355) );
  XOR U3318 ( .A(p_input[13]), .B(p_input[269]), .Z(n3352) );
  XOR U3319 ( .A(p_input[14]), .B(n3387), .Z(n3386) );
  XNOR U3320 ( .A(n3388), .B(p_input[9]), .Z(n3347) );
  XNOR U3321 ( .A(n3363), .B(n3362), .Z(n3345) );
  XNOR U3322 ( .A(n3389), .B(n3368), .Z(n3362) );
  XOR U3323 ( .A(p_input[264]), .B(p_input[8]), .Z(n3368) );
  XOR U3324 ( .A(n3359), .B(n3367), .Z(n3389) );
  XOR U3325 ( .A(n3390), .B(n3364), .Z(n3367) );
  XOR U3326 ( .A(p_input[262]), .B(p_input[6]), .Z(n3364) );
  XNOR U3327 ( .A(p_input[263]), .B(p_input[7]), .Z(n3390) );
  XNOR U3328 ( .A(n3391), .B(p_input[2]), .Z(n3359) );
  XNOR U3329 ( .A(n3373), .B(n3372), .Z(n3363) );
  XOR U3330 ( .A(n3392), .B(n3369), .Z(n3372) );
  XOR U3331 ( .A(p_input[259]), .B(p_input[3]), .Z(n3369) );
  XNOR U3332 ( .A(p_input[260]), .B(p_input[4]), .Z(n3392) );
  XOR U3333 ( .A(p_input[261]), .B(p_input[5]), .Z(n3373) );
  IV U3334 ( .A(n3270), .Z(n3274) );
  XOR U3335 ( .A(n3393), .B(n3394), .Z(n3270) );
  AND U3336 ( .A(n74), .B(n3395), .Z(n3394) );
  XNOR U3337 ( .A(n3396), .B(n3397), .Z(n74) );
  AND U3338 ( .A(n3398), .B(n3399), .Z(n3397) );
  XOR U3339 ( .A(n3285), .B(n3396), .Z(n3399) );
  XNOR U3340 ( .A(n3400), .B(n3396), .Z(n3398) );
  XOR U3341 ( .A(n3401), .B(n3402), .Z(n3396) );
  AND U3342 ( .A(n3403), .B(n3404), .Z(n3402) );
  XOR U3343 ( .A(n3300), .B(n3401), .Z(n3404) );
  XOR U3344 ( .A(n3401), .B(n3301), .Z(n3403) );
  XOR U3345 ( .A(n3405), .B(n3406), .Z(n3401) );
  AND U3346 ( .A(n3407), .B(n3408), .Z(n3406) );
  XOR U3347 ( .A(n3328), .B(n3405), .Z(n3408) );
  XOR U3348 ( .A(n3405), .B(n3329), .Z(n3407) );
  XOR U3349 ( .A(n3409), .B(n3410), .Z(n3405) );
  AND U3350 ( .A(n3411), .B(n3412), .Z(n3410) );
  XOR U3351 ( .A(n3409), .B(n3377), .Z(n3412) );
  XNOR U3352 ( .A(n3413), .B(n3414), .Z(n3224) );
  AND U3353 ( .A(n78), .B(n3415), .Z(n3414) );
  XNOR U3354 ( .A(n3416), .B(n3417), .Z(n78) );
  AND U3355 ( .A(n3418), .B(n3419), .Z(n3417) );
  XOR U3356 ( .A(n3416), .B(n3236), .Z(n3419) );
  XNOR U3357 ( .A(n3416), .B(n3180), .Z(n3418) );
  XOR U3358 ( .A(n3420), .B(n3421), .Z(n3416) );
  AND U3359 ( .A(n3422), .B(n3423), .Z(n3421) );
  XNOR U3360 ( .A(n3246), .B(n3420), .Z(n3423) );
  XOR U3361 ( .A(n3420), .B(n3248), .Z(n3422) );
  XOR U3362 ( .A(n3424), .B(n3425), .Z(n3420) );
  AND U3363 ( .A(n3426), .B(n3427), .Z(n3425) );
  XOR U3364 ( .A(n3424), .B(n3259), .Z(n3426) );
  IV U3365 ( .A(n3206), .Z(n3259) );
  XOR U3366 ( .A(n3428), .B(n3429), .Z(n3222) );
  AND U3367 ( .A(n82), .B(n3415), .Z(n3429) );
  XNOR U3368 ( .A(n3413), .B(n3428), .Z(n3415) );
  XNOR U3369 ( .A(n3430), .B(n3431), .Z(n82) );
  AND U3370 ( .A(n3432), .B(n3433), .Z(n3431) );
  XNOR U3371 ( .A(n3434), .B(n3430), .Z(n3433) );
  IV U3372 ( .A(n3236), .Z(n3434) );
  XOR U3373 ( .A(n3400), .B(n3435), .Z(n3236) );
  AND U3374 ( .A(n86), .B(n3436), .Z(n3435) );
  XOR U3375 ( .A(n3284), .B(n3281), .Z(n3436) );
  IV U3376 ( .A(n3400), .Z(n3284) );
  XNOR U3377 ( .A(n3180), .B(n3430), .Z(n3432) );
  XOR U3378 ( .A(n3437), .B(n3438), .Z(n3180) );
  AND U3379 ( .A(n102), .B(n3439), .Z(n3438) );
  XOR U3380 ( .A(n3440), .B(n3441), .Z(n3430) );
  AND U3381 ( .A(n3442), .B(n3443), .Z(n3441) );
  XNOR U3382 ( .A(n3440), .B(n3246), .Z(n3443) );
  XOR U3383 ( .A(n3301), .B(n3444), .Z(n3246) );
  AND U3384 ( .A(n86), .B(n3445), .Z(n3444) );
  XOR U3385 ( .A(n3297), .B(n3301), .Z(n3445) );
  XNOR U3386 ( .A(n3193), .B(n3440), .Z(n3442) );
  IV U3387 ( .A(n3248), .Z(n3193) );
  XOR U3388 ( .A(n3446), .B(n3447), .Z(n3248) );
  AND U3389 ( .A(n102), .B(n3448), .Z(n3447) );
  XOR U3390 ( .A(n3424), .B(n3449), .Z(n3440) );
  AND U3391 ( .A(n3450), .B(n3427), .Z(n3449) );
  XNOR U3392 ( .A(n3257), .B(n3424), .Z(n3427) );
  XOR U3393 ( .A(n3329), .B(n3451), .Z(n3257) );
  AND U3394 ( .A(n86), .B(n3452), .Z(n3451) );
  XOR U3395 ( .A(n3325), .B(n3329), .Z(n3452) );
  XNOR U3396 ( .A(n3206), .B(n3424), .Z(n3450) );
  XNOR U3397 ( .A(n3453), .B(n3454), .Z(n3206) );
  AND U3398 ( .A(n102), .B(n3455), .Z(n3454) );
  XOR U3399 ( .A(n3456), .B(n3457), .Z(n3424) );
  AND U3400 ( .A(n3458), .B(n3459), .Z(n3457) );
  XNOR U3401 ( .A(n3456), .B(n3268), .Z(n3459) );
  XOR U3402 ( .A(n3378), .B(n3460), .Z(n3268) );
  AND U3403 ( .A(n86), .B(n3461), .Z(n3460) );
  XOR U3404 ( .A(n3374), .B(n3378), .Z(n3461) );
  XNOR U3405 ( .A(n3462), .B(n3456), .Z(n3458) );
  IV U3406 ( .A(n3219), .Z(n3462) );
  XOR U3407 ( .A(n3463), .B(n3464), .Z(n3219) );
  AND U3408 ( .A(n102), .B(n3465), .Z(n3464) );
  AND U3409 ( .A(n3428), .B(n3413), .Z(n3456) );
  XNOR U3410 ( .A(n3466), .B(n3467), .Z(n3413) );
  AND U3411 ( .A(n86), .B(n3395), .Z(n3467) );
  XNOR U3412 ( .A(n3393), .B(n3466), .Z(n3395) );
  XNOR U3413 ( .A(n3468), .B(n3469), .Z(n86) );
  AND U3414 ( .A(n3470), .B(n3471), .Z(n3469) );
  XNOR U3415 ( .A(n3468), .B(n3281), .Z(n3471) );
  IV U3416 ( .A(n3285), .Z(n3281) );
  XOR U3417 ( .A(n3472), .B(n3473), .Z(n3285) );
  AND U3418 ( .A(n90), .B(n3474), .Z(n3473) );
  XOR U3419 ( .A(n3475), .B(n3472), .Z(n3474) );
  XNOR U3420 ( .A(n3468), .B(n3400), .Z(n3470) );
  XOR U3421 ( .A(n3476), .B(n3477), .Z(n3400) );
  AND U3422 ( .A(n98), .B(n3439), .Z(n3477) );
  XOR U3423 ( .A(n3437), .B(n3476), .Z(n3439) );
  XOR U3424 ( .A(n3478), .B(n3479), .Z(n3468) );
  AND U3425 ( .A(n3480), .B(n3481), .Z(n3479) );
  XNOR U3426 ( .A(n3478), .B(n3297), .Z(n3481) );
  IV U3427 ( .A(n3300), .Z(n3297) );
  XOR U3428 ( .A(n3482), .B(n3483), .Z(n3300) );
  AND U3429 ( .A(n90), .B(n3484), .Z(n3483) );
  XOR U3430 ( .A(n3485), .B(n3482), .Z(n3484) );
  XOR U3431 ( .A(n3301), .B(n3478), .Z(n3480) );
  XOR U3432 ( .A(n3486), .B(n3487), .Z(n3301) );
  AND U3433 ( .A(n98), .B(n3448), .Z(n3487) );
  XOR U3434 ( .A(n3486), .B(n3446), .Z(n3448) );
  XOR U3435 ( .A(n3488), .B(n3489), .Z(n3478) );
  AND U3436 ( .A(n3490), .B(n3491), .Z(n3489) );
  XNOR U3437 ( .A(n3488), .B(n3325), .Z(n3491) );
  IV U3438 ( .A(n3328), .Z(n3325) );
  XOR U3439 ( .A(n3492), .B(n3493), .Z(n3328) );
  AND U3440 ( .A(n90), .B(n3494), .Z(n3493) );
  XNOR U3441 ( .A(n3495), .B(n3492), .Z(n3494) );
  XOR U3442 ( .A(n3329), .B(n3488), .Z(n3490) );
  XOR U3443 ( .A(n3496), .B(n3497), .Z(n3329) );
  AND U3444 ( .A(n98), .B(n3455), .Z(n3497) );
  XOR U3445 ( .A(n3496), .B(n3453), .Z(n3455) );
  XOR U3446 ( .A(n3409), .B(n3498), .Z(n3488) );
  AND U3447 ( .A(n3411), .B(n3499), .Z(n3498) );
  XNOR U3448 ( .A(n3409), .B(n3374), .Z(n3499) );
  IV U3449 ( .A(n3377), .Z(n3374) );
  XOR U3450 ( .A(n3500), .B(n3501), .Z(n3377) );
  AND U3451 ( .A(n90), .B(n3502), .Z(n3501) );
  XOR U3452 ( .A(n3503), .B(n3500), .Z(n3502) );
  XOR U3453 ( .A(n3378), .B(n3409), .Z(n3411) );
  XOR U3454 ( .A(n3504), .B(n3505), .Z(n3378) );
  AND U3455 ( .A(n98), .B(n3465), .Z(n3505) );
  XOR U3456 ( .A(n3504), .B(n3463), .Z(n3465) );
  AND U3457 ( .A(n3466), .B(n3393), .Z(n3409) );
  XNOR U3458 ( .A(n3506), .B(n3507), .Z(n3393) );
  AND U3459 ( .A(n90), .B(n3508), .Z(n3507) );
  XNOR U3460 ( .A(n3509), .B(n3506), .Z(n3508) );
  XNOR U3461 ( .A(n3510), .B(n3511), .Z(n90) );
  AND U3462 ( .A(n3512), .B(n3513), .Z(n3511) );
  XOR U3463 ( .A(n3475), .B(n3510), .Z(n3513) );
  AND U3464 ( .A(n3514), .B(n3515), .Z(n3475) );
  XNOR U3465 ( .A(n3472), .B(n3510), .Z(n3512) );
  XNOR U3466 ( .A(n3516), .B(n3517), .Z(n3472) );
  AND U3467 ( .A(n94), .B(n3518), .Z(n3517) );
  XNOR U3468 ( .A(n3519), .B(n3520), .Z(n3518) );
  XOR U3469 ( .A(n3521), .B(n3522), .Z(n3510) );
  AND U3470 ( .A(n3523), .B(n3524), .Z(n3522) );
  XNOR U3471 ( .A(n3521), .B(n3514), .Z(n3524) );
  IV U3472 ( .A(n3485), .Z(n3514) );
  XOR U3473 ( .A(n3525), .B(n3526), .Z(n3485) );
  XOR U3474 ( .A(n3527), .B(n3515), .Z(n3526) );
  AND U3475 ( .A(n3495), .B(n3528), .Z(n3515) );
  AND U3476 ( .A(n3529), .B(n3530), .Z(n3527) );
  XOR U3477 ( .A(n3531), .B(n3525), .Z(n3529) );
  XNOR U3478 ( .A(n3482), .B(n3521), .Z(n3523) );
  XNOR U3479 ( .A(n3532), .B(n3533), .Z(n3482) );
  AND U3480 ( .A(n94), .B(n3534), .Z(n3533) );
  XNOR U3481 ( .A(n3535), .B(n3536), .Z(n3534) );
  XOR U3482 ( .A(n3537), .B(n3538), .Z(n3521) );
  AND U3483 ( .A(n3539), .B(n3540), .Z(n3538) );
  XNOR U3484 ( .A(n3537), .B(n3495), .Z(n3540) );
  XOR U3485 ( .A(n3541), .B(n3530), .Z(n3495) );
  XNOR U3486 ( .A(n3542), .B(n3525), .Z(n3530) );
  XOR U3487 ( .A(n3543), .B(n3544), .Z(n3525) );
  AND U3488 ( .A(n3545), .B(n3546), .Z(n3544) );
  XOR U3489 ( .A(n3547), .B(n3543), .Z(n3545) );
  XNOR U3490 ( .A(n3548), .B(n3549), .Z(n3542) );
  AND U3491 ( .A(n3550), .B(n3551), .Z(n3549) );
  XOR U3492 ( .A(n3548), .B(n3552), .Z(n3550) );
  XNOR U3493 ( .A(n3531), .B(n3528), .Z(n3541) );
  AND U3494 ( .A(n3553), .B(n3554), .Z(n3528) );
  XOR U3495 ( .A(n3555), .B(n3556), .Z(n3531) );
  AND U3496 ( .A(n3557), .B(n3558), .Z(n3556) );
  XOR U3497 ( .A(n3555), .B(n3559), .Z(n3557) );
  XNOR U3498 ( .A(n3492), .B(n3537), .Z(n3539) );
  XNOR U3499 ( .A(n3560), .B(n3561), .Z(n3492) );
  AND U3500 ( .A(n94), .B(n3562), .Z(n3561) );
  XNOR U3501 ( .A(n3563), .B(n3564), .Z(n3562) );
  XOR U3502 ( .A(n3565), .B(n3566), .Z(n3537) );
  AND U3503 ( .A(n3567), .B(n3568), .Z(n3566) );
  XNOR U3504 ( .A(n3565), .B(n3553), .Z(n3568) );
  IV U3505 ( .A(n3503), .Z(n3553) );
  XNOR U3506 ( .A(n3569), .B(n3546), .Z(n3503) );
  XNOR U3507 ( .A(n3570), .B(n3552), .Z(n3546) );
  XOR U3508 ( .A(n3571), .B(n3572), .Z(n3552) );
  NOR U3509 ( .A(n3573), .B(n3574), .Z(n3572) );
  XNOR U3510 ( .A(n3571), .B(n3575), .Z(n3573) );
  XNOR U3511 ( .A(n3551), .B(n3543), .Z(n3570) );
  XOR U3512 ( .A(n3576), .B(n3577), .Z(n3543) );
  AND U3513 ( .A(n3578), .B(n3579), .Z(n3577) );
  XOR U3514 ( .A(n3576), .B(n3580), .Z(n3578) );
  XNOR U3515 ( .A(n3581), .B(n3548), .Z(n3551) );
  XOR U3516 ( .A(n3582), .B(n3583), .Z(n3548) );
  AND U3517 ( .A(n3584), .B(n3585), .Z(n3583) );
  XNOR U3518 ( .A(n3586), .B(n3587), .Z(n3584) );
  IV U3519 ( .A(n3582), .Z(n3586) );
  XNOR U3520 ( .A(n3588), .B(n3589), .Z(n3581) );
  NOR U3521 ( .A(n3590), .B(n3591), .Z(n3589) );
  XOR U3522 ( .A(n3588), .B(n3592), .Z(n3590) );
  XNOR U3523 ( .A(n3547), .B(n3554), .Z(n3569) );
  NOR U3524 ( .A(n3509), .B(n3593), .Z(n3554) );
  XOR U3525 ( .A(n3559), .B(n3558), .Z(n3547) );
  XNOR U3526 ( .A(n3594), .B(n3555), .Z(n3558) );
  XOR U3527 ( .A(n3595), .B(n3596), .Z(n3555) );
  AND U3528 ( .A(n3597), .B(n3598), .Z(n3596) );
  XNOR U3529 ( .A(n3599), .B(n3600), .Z(n3597) );
  IV U3530 ( .A(n3595), .Z(n3599) );
  XNOR U3531 ( .A(n3601), .B(n3602), .Z(n3594) );
  NOR U3532 ( .A(n3603), .B(n3604), .Z(n3602) );
  XNOR U3533 ( .A(n3601), .B(n3605), .Z(n3603) );
  XOR U3534 ( .A(n3606), .B(n3607), .Z(n3559) );
  NOR U3535 ( .A(n3608), .B(n3609), .Z(n3607) );
  XNOR U3536 ( .A(n3606), .B(n3610), .Z(n3608) );
  XNOR U3537 ( .A(n3500), .B(n3565), .Z(n3567) );
  XNOR U3538 ( .A(n3611), .B(n3612), .Z(n3500) );
  AND U3539 ( .A(n94), .B(n3613), .Z(n3612) );
  XNOR U3540 ( .A(n3614), .B(n3615), .Z(n3613) );
  AND U3541 ( .A(n3506), .B(n3509), .Z(n3565) );
  XOR U3542 ( .A(n3616), .B(n3593), .Z(n3509) );
  XNOR U3543 ( .A(p_input[16]), .B(p_input[256]), .Z(n3593) );
  XNOR U3544 ( .A(n3580), .B(n3579), .Z(n3616) );
  XNOR U3545 ( .A(n3617), .B(n3587), .Z(n3579) );
  XNOR U3546 ( .A(n3575), .B(n3574), .Z(n3587) );
  XOR U3547 ( .A(n3618), .B(n3571), .Z(n3574) );
  XNOR U3548 ( .A(n3619), .B(p_input[26]), .Z(n3571) );
  XNOR U3549 ( .A(p_input[267]), .B(p_input[27]), .Z(n3618) );
  XOR U3550 ( .A(p_input[268]), .B(p_input[28]), .Z(n3575) );
  XOR U3551 ( .A(n3585), .B(n3620), .Z(n3617) );
  IV U3552 ( .A(n3576), .Z(n3620) );
  XOR U3553 ( .A(p_input[17]), .B(p_input[257]), .Z(n3576) );
  XOR U3554 ( .A(n3621), .B(n3592), .Z(n3585) );
  XNOR U3555 ( .A(p_input[271]), .B(p_input[31]), .Z(n3592) );
  XOR U3556 ( .A(n3582), .B(n3591), .Z(n3621) );
  XOR U3557 ( .A(n3622), .B(n3588), .Z(n3591) );
  XOR U3558 ( .A(p_input[269]), .B(p_input[29]), .Z(n3588) );
  XNOR U3559 ( .A(p_input[270]), .B(p_input[30]), .Z(n3622) );
  XOR U3560 ( .A(p_input[25]), .B(p_input[265]), .Z(n3582) );
  XOR U3561 ( .A(n3600), .B(n3598), .Z(n3580) );
  XNOR U3562 ( .A(n3623), .B(n3605), .Z(n3598) );
  XOR U3563 ( .A(p_input[24]), .B(p_input[264]), .Z(n3605) );
  XOR U3564 ( .A(n3595), .B(n3604), .Z(n3623) );
  XOR U3565 ( .A(n3624), .B(n3601), .Z(n3604) );
  XOR U3566 ( .A(p_input[22]), .B(p_input[262]), .Z(n3601) );
  XOR U3567 ( .A(p_input[23]), .B(n3625), .Z(n3624) );
  XOR U3568 ( .A(p_input[18]), .B(p_input[258]), .Z(n3595) );
  XNOR U3569 ( .A(n3610), .B(n3609), .Z(n3600) );
  XOR U3570 ( .A(n3626), .B(n3606), .Z(n3609) );
  XOR U3571 ( .A(p_input[19]), .B(p_input[259]), .Z(n3606) );
  XOR U3572 ( .A(p_input[20]), .B(n3627), .Z(n3626) );
  XOR U3573 ( .A(p_input[21]), .B(p_input[261]), .Z(n3610) );
  XNOR U3574 ( .A(n3628), .B(n3629), .Z(n3506) );
  AND U3575 ( .A(n94), .B(n3630), .Z(n3629) );
  XNOR U3576 ( .A(n3631), .B(n3632), .Z(n94) );
  AND U3577 ( .A(n3633), .B(n3634), .Z(n3632) );
  XOR U3578 ( .A(n3520), .B(n3631), .Z(n3634) );
  XNOR U3579 ( .A(n3635), .B(n3631), .Z(n3633) );
  XOR U3580 ( .A(n3636), .B(n3637), .Z(n3631) );
  AND U3581 ( .A(n3638), .B(n3639), .Z(n3637) );
  XOR U3582 ( .A(n3535), .B(n3636), .Z(n3639) );
  XOR U3583 ( .A(n3636), .B(n3536), .Z(n3638) );
  XOR U3584 ( .A(n3640), .B(n3641), .Z(n3636) );
  AND U3585 ( .A(n3642), .B(n3643), .Z(n3641) );
  XOR U3586 ( .A(n3563), .B(n3640), .Z(n3643) );
  XOR U3587 ( .A(n3640), .B(n3564), .Z(n3642) );
  XOR U3588 ( .A(n3644), .B(n3645), .Z(n3640) );
  AND U3589 ( .A(n3646), .B(n3647), .Z(n3645) );
  XOR U3590 ( .A(n3644), .B(n3614), .Z(n3647) );
  XNOR U3591 ( .A(n3648), .B(n3649), .Z(n3466) );
  AND U3592 ( .A(n98), .B(n3650), .Z(n3649) );
  XNOR U3593 ( .A(n3651), .B(n3652), .Z(n98) );
  AND U3594 ( .A(n3653), .B(n3654), .Z(n3652) );
  XOR U3595 ( .A(n3651), .B(n3476), .Z(n3654) );
  XNOR U3596 ( .A(n3651), .B(n3437), .Z(n3653) );
  XOR U3597 ( .A(n3655), .B(n3656), .Z(n3651) );
  AND U3598 ( .A(n3657), .B(n3658), .Z(n3656) );
  XOR U3599 ( .A(n3655), .B(n3446), .Z(n3657) );
  XOR U3600 ( .A(n3659), .B(n3660), .Z(n3428) );
  AND U3601 ( .A(n102), .B(n3650), .Z(n3660) );
  XNOR U3602 ( .A(n3648), .B(n3659), .Z(n3650) );
  XNOR U3603 ( .A(n3661), .B(n3662), .Z(n102) );
  AND U3604 ( .A(n3663), .B(n3664), .Z(n3662) );
  XNOR U3605 ( .A(n3665), .B(n3661), .Z(n3664) );
  IV U3606 ( .A(n3476), .Z(n3665) );
  XOR U3607 ( .A(n3635), .B(n3666), .Z(n3476) );
  AND U3608 ( .A(n105), .B(n3667), .Z(n3666) );
  XOR U3609 ( .A(n3519), .B(n3516), .Z(n3667) );
  IV U3610 ( .A(n3635), .Z(n3519) );
  XNOR U3611 ( .A(n3437), .B(n3661), .Z(n3663) );
  XOR U3612 ( .A(n3668), .B(n3669), .Z(n3437) );
  AND U3613 ( .A(n121), .B(n3670), .Z(n3669) );
  XOR U3614 ( .A(n3655), .B(n3671), .Z(n3661) );
  AND U3615 ( .A(n3672), .B(n3658), .Z(n3671) );
  XNOR U3616 ( .A(n3486), .B(n3655), .Z(n3658) );
  XOR U3617 ( .A(n3536), .B(n3673), .Z(n3486) );
  AND U3618 ( .A(n105), .B(n3674), .Z(n3673) );
  XOR U3619 ( .A(n3532), .B(n3536), .Z(n3674) );
  XNOR U3620 ( .A(n3675), .B(n3655), .Z(n3672) );
  IV U3621 ( .A(n3446), .Z(n3675) );
  XOR U3622 ( .A(n3676), .B(n3677), .Z(n3446) );
  AND U3623 ( .A(n121), .B(n3678), .Z(n3677) );
  XOR U3624 ( .A(n3679), .B(n3680), .Z(n3655) );
  AND U3625 ( .A(n3681), .B(n3682), .Z(n3680) );
  XNOR U3626 ( .A(n3496), .B(n3679), .Z(n3682) );
  XOR U3627 ( .A(n3564), .B(n3683), .Z(n3496) );
  AND U3628 ( .A(n105), .B(n3684), .Z(n3683) );
  XOR U3629 ( .A(n3560), .B(n3564), .Z(n3684) );
  XOR U3630 ( .A(n3679), .B(n3453), .Z(n3681) );
  XOR U3631 ( .A(n3685), .B(n3686), .Z(n3453) );
  AND U3632 ( .A(n121), .B(n3687), .Z(n3686) );
  XOR U3633 ( .A(n3688), .B(n3689), .Z(n3679) );
  AND U3634 ( .A(n3690), .B(n3691), .Z(n3689) );
  XNOR U3635 ( .A(n3688), .B(n3504), .Z(n3691) );
  XOR U3636 ( .A(n3615), .B(n3692), .Z(n3504) );
  AND U3637 ( .A(n105), .B(n3693), .Z(n3692) );
  XOR U3638 ( .A(n3611), .B(n3615), .Z(n3693) );
  XNOR U3639 ( .A(n3694), .B(n3688), .Z(n3690) );
  IV U3640 ( .A(n3463), .Z(n3694) );
  XOR U3641 ( .A(n3695), .B(n3696), .Z(n3463) );
  AND U3642 ( .A(n121), .B(n3697), .Z(n3696) );
  AND U3643 ( .A(n3659), .B(n3648), .Z(n3688) );
  XNOR U3644 ( .A(n3698), .B(n3699), .Z(n3648) );
  AND U3645 ( .A(n105), .B(n3630), .Z(n3699) );
  XNOR U3646 ( .A(n3628), .B(n3698), .Z(n3630) );
  XNOR U3647 ( .A(n3700), .B(n3701), .Z(n105) );
  AND U3648 ( .A(n3702), .B(n3703), .Z(n3701) );
  XNOR U3649 ( .A(n3700), .B(n3516), .Z(n3703) );
  IV U3650 ( .A(n3520), .Z(n3516) );
  XOR U3651 ( .A(n3704), .B(n3705), .Z(n3520) );
  AND U3652 ( .A(n109), .B(n3706), .Z(n3705) );
  XOR U3653 ( .A(n3707), .B(n3704), .Z(n3706) );
  XNOR U3654 ( .A(n3700), .B(n3635), .Z(n3702) );
  XOR U3655 ( .A(n3708), .B(n3709), .Z(n3635) );
  AND U3656 ( .A(n117), .B(n3670), .Z(n3709) );
  XOR U3657 ( .A(n3668), .B(n3708), .Z(n3670) );
  XOR U3658 ( .A(n3710), .B(n3711), .Z(n3700) );
  AND U3659 ( .A(n3712), .B(n3713), .Z(n3711) );
  XNOR U3660 ( .A(n3710), .B(n3532), .Z(n3713) );
  IV U3661 ( .A(n3535), .Z(n3532) );
  XOR U3662 ( .A(n3714), .B(n3715), .Z(n3535) );
  AND U3663 ( .A(n109), .B(n3716), .Z(n3715) );
  XOR U3664 ( .A(n3717), .B(n3714), .Z(n3716) );
  XOR U3665 ( .A(n3536), .B(n3710), .Z(n3712) );
  XOR U3666 ( .A(n3718), .B(n3719), .Z(n3536) );
  AND U3667 ( .A(n117), .B(n3678), .Z(n3719) );
  XOR U3668 ( .A(n3718), .B(n3676), .Z(n3678) );
  XOR U3669 ( .A(n3720), .B(n3721), .Z(n3710) );
  AND U3670 ( .A(n3722), .B(n3723), .Z(n3721) );
  XNOR U3671 ( .A(n3720), .B(n3560), .Z(n3723) );
  IV U3672 ( .A(n3563), .Z(n3560) );
  XOR U3673 ( .A(n3724), .B(n3725), .Z(n3563) );
  AND U3674 ( .A(n109), .B(n3726), .Z(n3725) );
  XNOR U3675 ( .A(n3727), .B(n3724), .Z(n3726) );
  XOR U3676 ( .A(n3564), .B(n3720), .Z(n3722) );
  XOR U3677 ( .A(n3728), .B(n3729), .Z(n3564) );
  AND U3678 ( .A(n117), .B(n3687), .Z(n3729) );
  XOR U3679 ( .A(n3728), .B(n3685), .Z(n3687) );
  XOR U3680 ( .A(n3644), .B(n3730), .Z(n3720) );
  AND U3681 ( .A(n3646), .B(n3731), .Z(n3730) );
  XNOR U3682 ( .A(n3644), .B(n3611), .Z(n3731) );
  IV U3683 ( .A(n3614), .Z(n3611) );
  XOR U3684 ( .A(n3732), .B(n3733), .Z(n3614) );
  AND U3685 ( .A(n109), .B(n3734), .Z(n3733) );
  XOR U3686 ( .A(n3735), .B(n3732), .Z(n3734) );
  XOR U3687 ( .A(n3615), .B(n3644), .Z(n3646) );
  XOR U3688 ( .A(n3736), .B(n3737), .Z(n3615) );
  AND U3689 ( .A(n117), .B(n3697), .Z(n3737) );
  XOR U3690 ( .A(n3736), .B(n3695), .Z(n3697) );
  AND U3691 ( .A(n3698), .B(n3628), .Z(n3644) );
  XNOR U3692 ( .A(n3738), .B(n3739), .Z(n3628) );
  AND U3693 ( .A(n109), .B(n3740), .Z(n3739) );
  XNOR U3694 ( .A(n3741), .B(n3738), .Z(n3740) );
  XNOR U3695 ( .A(n3742), .B(n3743), .Z(n109) );
  AND U3696 ( .A(n3744), .B(n3745), .Z(n3743) );
  XOR U3697 ( .A(n3707), .B(n3742), .Z(n3745) );
  AND U3698 ( .A(n3746), .B(n3747), .Z(n3707) );
  XNOR U3699 ( .A(n3704), .B(n3742), .Z(n3744) );
  XNOR U3700 ( .A(n3748), .B(n3749), .Z(n3704) );
  AND U3701 ( .A(n113), .B(n3750), .Z(n3749) );
  XNOR U3702 ( .A(n3751), .B(n3752), .Z(n3750) );
  XOR U3703 ( .A(n3753), .B(n3754), .Z(n3742) );
  AND U3704 ( .A(n3755), .B(n3756), .Z(n3754) );
  XNOR U3705 ( .A(n3753), .B(n3746), .Z(n3756) );
  IV U3706 ( .A(n3717), .Z(n3746) );
  XOR U3707 ( .A(n3757), .B(n3758), .Z(n3717) );
  XOR U3708 ( .A(n3759), .B(n3747), .Z(n3758) );
  AND U3709 ( .A(n3727), .B(n3760), .Z(n3747) );
  AND U3710 ( .A(n3761), .B(n3762), .Z(n3759) );
  XOR U3711 ( .A(n3763), .B(n3757), .Z(n3761) );
  XNOR U3712 ( .A(n3714), .B(n3753), .Z(n3755) );
  XNOR U3713 ( .A(n3764), .B(n3765), .Z(n3714) );
  AND U3714 ( .A(n113), .B(n3766), .Z(n3765) );
  XNOR U3715 ( .A(n3767), .B(n3768), .Z(n3766) );
  XOR U3716 ( .A(n3769), .B(n3770), .Z(n3753) );
  AND U3717 ( .A(n3771), .B(n3772), .Z(n3770) );
  XNOR U3718 ( .A(n3769), .B(n3727), .Z(n3772) );
  XOR U3719 ( .A(n3773), .B(n3762), .Z(n3727) );
  XNOR U3720 ( .A(n3774), .B(n3757), .Z(n3762) );
  XOR U3721 ( .A(n3775), .B(n3776), .Z(n3757) );
  AND U3722 ( .A(n3777), .B(n3778), .Z(n3776) );
  XOR U3723 ( .A(n3779), .B(n3775), .Z(n3777) );
  XNOR U3724 ( .A(n3780), .B(n3781), .Z(n3774) );
  AND U3725 ( .A(n3782), .B(n3783), .Z(n3781) );
  XOR U3726 ( .A(n3780), .B(n3784), .Z(n3782) );
  XNOR U3727 ( .A(n3763), .B(n3760), .Z(n3773) );
  AND U3728 ( .A(n3785), .B(n3786), .Z(n3760) );
  XOR U3729 ( .A(n3787), .B(n3788), .Z(n3763) );
  AND U3730 ( .A(n3789), .B(n3790), .Z(n3788) );
  XOR U3731 ( .A(n3787), .B(n3791), .Z(n3789) );
  XNOR U3732 ( .A(n3724), .B(n3769), .Z(n3771) );
  XNOR U3733 ( .A(n3792), .B(n3793), .Z(n3724) );
  AND U3734 ( .A(n113), .B(n3794), .Z(n3793) );
  XNOR U3735 ( .A(n3795), .B(n3796), .Z(n3794) );
  XOR U3736 ( .A(n3797), .B(n3798), .Z(n3769) );
  AND U3737 ( .A(n3799), .B(n3800), .Z(n3798) );
  XNOR U3738 ( .A(n3797), .B(n3785), .Z(n3800) );
  IV U3739 ( .A(n3735), .Z(n3785) );
  XNOR U3740 ( .A(n3801), .B(n3778), .Z(n3735) );
  XNOR U3741 ( .A(n3802), .B(n3784), .Z(n3778) );
  XOR U3742 ( .A(n3803), .B(n3804), .Z(n3784) );
  NOR U3743 ( .A(n3805), .B(n3806), .Z(n3804) );
  XNOR U3744 ( .A(n3803), .B(n3807), .Z(n3805) );
  XNOR U3745 ( .A(n3783), .B(n3775), .Z(n3802) );
  XOR U3746 ( .A(n3808), .B(n3809), .Z(n3775) );
  AND U3747 ( .A(n3810), .B(n3811), .Z(n3809) );
  XNOR U3748 ( .A(n3808), .B(n3812), .Z(n3810) );
  XNOR U3749 ( .A(n3813), .B(n3780), .Z(n3783) );
  XOR U3750 ( .A(n3814), .B(n3815), .Z(n3780) );
  AND U3751 ( .A(n3816), .B(n3817), .Z(n3815) );
  XOR U3752 ( .A(n3814), .B(n3818), .Z(n3816) );
  XNOR U3753 ( .A(n3819), .B(n3820), .Z(n3813) );
  NOR U3754 ( .A(n3821), .B(n3822), .Z(n3820) );
  XOR U3755 ( .A(n3819), .B(n3823), .Z(n3821) );
  XNOR U3756 ( .A(n3779), .B(n3786), .Z(n3801) );
  NOR U3757 ( .A(n3741), .B(n3824), .Z(n3786) );
  XOR U3758 ( .A(n3791), .B(n3790), .Z(n3779) );
  XNOR U3759 ( .A(n3825), .B(n3787), .Z(n3790) );
  XOR U3760 ( .A(n3826), .B(n3827), .Z(n3787) );
  AND U3761 ( .A(n3828), .B(n3829), .Z(n3827) );
  XOR U3762 ( .A(n3826), .B(n3830), .Z(n3828) );
  XNOR U3763 ( .A(n3831), .B(n3832), .Z(n3825) );
  NOR U3764 ( .A(n3833), .B(n3834), .Z(n3832) );
  XNOR U3765 ( .A(n3831), .B(n3835), .Z(n3833) );
  XOR U3766 ( .A(n3836), .B(n3837), .Z(n3791) );
  NOR U3767 ( .A(n3838), .B(n3839), .Z(n3837) );
  XNOR U3768 ( .A(n3836), .B(n3840), .Z(n3838) );
  XNOR U3769 ( .A(n3732), .B(n3797), .Z(n3799) );
  XNOR U3770 ( .A(n3841), .B(n3842), .Z(n3732) );
  AND U3771 ( .A(n113), .B(n3843), .Z(n3842) );
  XNOR U3772 ( .A(n3844), .B(n3845), .Z(n3843) );
  AND U3773 ( .A(n3738), .B(n3741), .Z(n3797) );
  XOR U3774 ( .A(n3846), .B(n3824), .Z(n3741) );
  XNOR U3775 ( .A(p_input[256]), .B(p_input[32]), .Z(n3824) );
  XOR U3776 ( .A(n3812), .B(n3811), .Z(n3846) );
  XNOR U3777 ( .A(n3847), .B(n3818), .Z(n3811) );
  XNOR U3778 ( .A(n3807), .B(n3806), .Z(n3818) );
  XOR U3779 ( .A(n3848), .B(n3803), .Z(n3806) );
  XNOR U3780 ( .A(n3619), .B(p_input[42]), .Z(n3803) );
  XNOR U3781 ( .A(p_input[267]), .B(p_input[43]), .Z(n3848) );
  XOR U3782 ( .A(p_input[268]), .B(p_input[44]), .Z(n3807) );
  XNOR U3783 ( .A(n3817), .B(n3808), .Z(n3847) );
  XNOR U3784 ( .A(n3849), .B(p_input[33]), .Z(n3808) );
  XOR U3785 ( .A(n3850), .B(n3823), .Z(n3817) );
  XNOR U3786 ( .A(p_input[271]), .B(p_input[47]), .Z(n3823) );
  XOR U3787 ( .A(n3814), .B(n3822), .Z(n3850) );
  XOR U3788 ( .A(n3851), .B(n3819), .Z(n3822) );
  XOR U3789 ( .A(p_input[269]), .B(p_input[45]), .Z(n3819) );
  XNOR U3790 ( .A(p_input[270]), .B(p_input[46]), .Z(n3851) );
  XNOR U3791 ( .A(n3388), .B(p_input[41]), .Z(n3814) );
  XNOR U3792 ( .A(n3830), .B(n3829), .Z(n3812) );
  XNOR U3793 ( .A(n3852), .B(n3835), .Z(n3829) );
  XOR U3794 ( .A(p_input[264]), .B(p_input[40]), .Z(n3835) );
  XOR U3795 ( .A(n3826), .B(n3834), .Z(n3852) );
  XOR U3796 ( .A(n3853), .B(n3831), .Z(n3834) );
  XOR U3797 ( .A(p_input[262]), .B(p_input[38]), .Z(n3831) );
  XNOR U3798 ( .A(p_input[263]), .B(p_input[39]), .Z(n3853) );
  XNOR U3799 ( .A(n3391), .B(p_input[34]), .Z(n3826) );
  XNOR U3800 ( .A(n3840), .B(n3839), .Z(n3830) );
  XOR U3801 ( .A(n3854), .B(n3836), .Z(n3839) );
  XOR U3802 ( .A(p_input[259]), .B(p_input[35]), .Z(n3836) );
  XNOR U3803 ( .A(p_input[260]), .B(p_input[36]), .Z(n3854) );
  XOR U3804 ( .A(p_input[261]), .B(p_input[37]), .Z(n3840) );
  XNOR U3805 ( .A(n3855), .B(n3856), .Z(n3738) );
  AND U3806 ( .A(n113), .B(n3857), .Z(n3856) );
  XNOR U3807 ( .A(n3858), .B(n3859), .Z(n113) );
  AND U3808 ( .A(n3860), .B(n3861), .Z(n3859) );
  XOR U3809 ( .A(n3752), .B(n3858), .Z(n3861) );
  XNOR U3810 ( .A(n3862), .B(n3858), .Z(n3860) );
  XOR U3811 ( .A(n3863), .B(n3864), .Z(n3858) );
  AND U3812 ( .A(n3865), .B(n3866), .Z(n3864) );
  XOR U3813 ( .A(n3767), .B(n3863), .Z(n3866) );
  XOR U3814 ( .A(n3863), .B(n3768), .Z(n3865) );
  XOR U3815 ( .A(n3867), .B(n3868), .Z(n3863) );
  AND U3816 ( .A(n3869), .B(n3870), .Z(n3868) );
  XOR U3817 ( .A(n3795), .B(n3867), .Z(n3870) );
  XOR U3818 ( .A(n3867), .B(n3796), .Z(n3869) );
  XOR U3819 ( .A(n3871), .B(n3872), .Z(n3867) );
  AND U3820 ( .A(n3873), .B(n3874), .Z(n3872) );
  XOR U3821 ( .A(n3871), .B(n3844), .Z(n3874) );
  XNOR U3822 ( .A(n3875), .B(n3876), .Z(n3698) );
  AND U3823 ( .A(n117), .B(n3877), .Z(n3876) );
  XNOR U3824 ( .A(n3878), .B(n3879), .Z(n117) );
  AND U3825 ( .A(n3880), .B(n3881), .Z(n3879) );
  XOR U3826 ( .A(n3878), .B(n3708), .Z(n3881) );
  XNOR U3827 ( .A(n3878), .B(n3668), .Z(n3880) );
  XOR U3828 ( .A(n3882), .B(n3883), .Z(n3878) );
  AND U3829 ( .A(n3884), .B(n3885), .Z(n3883) );
  XOR U3830 ( .A(n3882), .B(n3676), .Z(n3884) );
  XOR U3831 ( .A(n3886), .B(n3887), .Z(n3659) );
  AND U3832 ( .A(n121), .B(n3877), .Z(n3887) );
  XNOR U3833 ( .A(n3875), .B(n3886), .Z(n3877) );
  XNOR U3834 ( .A(n3888), .B(n3889), .Z(n121) );
  AND U3835 ( .A(n3890), .B(n3891), .Z(n3889) );
  XNOR U3836 ( .A(n3892), .B(n3888), .Z(n3891) );
  IV U3837 ( .A(n3708), .Z(n3892) );
  XOR U3838 ( .A(n3862), .B(n3893), .Z(n3708) );
  AND U3839 ( .A(n124), .B(n3894), .Z(n3893) );
  XOR U3840 ( .A(n3751), .B(n3748), .Z(n3894) );
  IV U3841 ( .A(n3862), .Z(n3751) );
  XNOR U3842 ( .A(n3668), .B(n3888), .Z(n3890) );
  XOR U3843 ( .A(n3895), .B(n3896), .Z(n3668) );
  AND U3844 ( .A(n140), .B(n3897), .Z(n3896) );
  XOR U3845 ( .A(n3882), .B(n3898), .Z(n3888) );
  AND U3846 ( .A(n3899), .B(n3885), .Z(n3898) );
  XNOR U3847 ( .A(n3718), .B(n3882), .Z(n3885) );
  XOR U3848 ( .A(n3768), .B(n3900), .Z(n3718) );
  AND U3849 ( .A(n124), .B(n3901), .Z(n3900) );
  XOR U3850 ( .A(n3764), .B(n3768), .Z(n3901) );
  XNOR U3851 ( .A(n3902), .B(n3882), .Z(n3899) );
  IV U3852 ( .A(n3676), .Z(n3902) );
  XOR U3853 ( .A(n3903), .B(n3904), .Z(n3676) );
  AND U3854 ( .A(n140), .B(n3905), .Z(n3904) );
  XOR U3855 ( .A(n3906), .B(n3907), .Z(n3882) );
  AND U3856 ( .A(n3908), .B(n3909), .Z(n3907) );
  XNOR U3857 ( .A(n3728), .B(n3906), .Z(n3909) );
  XOR U3858 ( .A(n3796), .B(n3910), .Z(n3728) );
  AND U3859 ( .A(n124), .B(n3911), .Z(n3910) );
  XOR U3860 ( .A(n3792), .B(n3796), .Z(n3911) );
  XOR U3861 ( .A(n3906), .B(n3685), .Z(n3908) );
  XOR U3862 ( .A(n3912), .B(n3913), .Z(n3685) );
  AND U3863 ( .A(n140), .B(n3914), .Z(n3913) );
  XOR U3864 ( .A(n3915), .B(n3916), .Z(n3906) );
  AND U3865 ( .A(n3917), .B(n3918), .Z(n3916) );
  XNOR U3866 ( .A(n3915), .B(n3736), .Z(n3918) );
  XOR U3867 ( .A(n3845), .B(n3919), .Z(n3736) );
  AND U3868 ( .A(n124), .B(n3920), .Z(n3919) );
  XOR U3869 ( .A(n3841), .B(n3845), .Z(n3920) );
  XNOR U3870 ( .A(n3921), .B(n3915), .Z(n3917) );
  IV U3871 ( .A(n3695), .Z(n3921) );
  XOR U3872 ( .A(n3922), .B(n3923), .Z(n3695) );
  AND U3873 ( .A(n140), .B(n3924), .Z(n3923) );
  AND U3874 ( .A(n3886), .B(n3875), .Z(n3915) );
  XNOR U3875 ( .A(n3925), .B(n3926), .Z(n3875) );
  AND U3876 ( .A(n124), .B(n3857), .Z(n3926) );
  XNOR U3877 ( .A(n3855), .B(n3925), .Z(n3857) );
  XNOR U3878 ( .A(n3927), .B(n3928), .Z(n124) );
  AND U3879 ( .A(n3929), .B(n3930), .Z(n3928) );
  XNOR U3880 ( .A(n3927), .B(n3748), .Z(n3930) );
  IV U3881 ( .A(n3752), .Z(n3748) );
  XOR U3882 ( .A(n3931), .B(n3932), .Z(n3752) );
  AND U3883 ( .A(n128), .B(n3933), .Z(n3932) );
  XOR U3884 ( .A(n3934), .B(n3931), .Z(n3933) );
  XNOR U3885 ( .A(n3927), .B(n3862), .Z(n3929) );
  XOR U3886 ( .A(n3935), .B(n3936), .Z(n3862) );
  AND U3887 ( .A(n136), .B(n3897), .Z(n3936) );
  XOR U3888 ( .A(n3895), .B(n3935), .Z(n3897) );
  XOR U3889 ( .A(n3937), .B(n3938), .Z(n3927) );
  AND U3890 ( .A(n3939), .B(n3940), .Z(n3938) );
  XNOR U3891 ( .A(n3937), .B(n3764), .Z(n3940) );
  IV U3892 ( .A(n3767), .Z(n3764) );
  XOR U3893 ( .A(n3941), .B(n3942), .Z(n3767) );
  AND U3894 ( .A(n128), .B(n3943), .Z(n3942) );
  XOR U3895 ( .A(n3944), .B(n3941), .Z(n3943) );
  XOR U3896 ( .A(n3768), .B(n3937), .Z(n3939) );
  XOR U3897 ( .A(n3945), .B(n3946), .Z(n3768) );
  AND U3898 ( .A(n136), .B(n3905), .Z(n3946) );
  XOR U3899 ( .A(n3945), .B(n3903), .Z(n3905) );
  XOR U3900 ( .A(n3947), .B(n3948), .Z(n3937) );
  AND U3901 ( .A(n3949), .B(n3950), .Z(n3948) );
  XNOR U3902 ( .A(n3947), .B(n3792), .Z(n3950) );
  IV U3903 ( .A(n3795), .Z(n3792) );
  XOR U3904 ( .A(n3951), .B(n3952), .Z(n3795) );
  AND U3905 ( .A(n128), .B(n3953), .Z(n3952) );
  XNOR U3906 ( .A(n3954), .B(n3951), .Z(n3953) );
  XOR U3907 ( .A(n3796), .B(n3947), .Z(n3949) );
  XOR U3908 ( .A(n3955), .B(n3956), .Z(n3796) );
  AND U3909 ( .A(n136), .B(n3914), .Z(n3956) );
  XOR U3910 ( .A(n3955), .B(n3912), .Z(n3914) );
  XOR U3911 ( .A(n3871), .B(n3957), .Z(n3947) );
  AND U3912 ( .A(n3873), .B(n3958), .Z(n3957) );
  XNOR U3913 ( .A(n3871), .B(n3841), .Z(n3958) );
  IV U3914 ( .A(n3844), .Z(n3841) );
  XOR U3915 ( .A(n3959), .B(n3960), .Z(n3844) );
  AND U3916 ( .A(n128), .B(n3961), .Z(n3960) );
  XOR U3917 ( .A(n3962), .B(n3959), .Z(n3961) );
  XOR U3918 ( .A(n3845), .B(n3871), .Z(n3873) );
  XOR U3919 ( .A(n3963), .B(n3964), .Z(n3845) );
  AND U3920 ( .A(n136), .B(n3924), .Z(n3964) );
  XOR U3921 ( .A(n3963), .B(n3922), .Z(n3924) );
  AND U3922 ( .A(n3925), .B(n3855), .Z(n3871) );
  XNOR U3923 ( .A(n3965), .B(n3966), .Z(n3855) );
  AND U3924 ( .A(n128), .B(n3967), .Z(n3966) );
  XNOR U3925 ( .A(n3968), .B(n3965), .Z(n3967) );
  XNOR U3926 ( .A(n3969), .B(n3970), .Z(n128) );
  AND U3927 ( .A(n3971), .B(n3972), .Z(n3970) );
  XOR U3928 ( .A(n3934), .B(n3969), .Z(n3972) );
  AND U3929 ( .A(n3973), .B(n3974), .Z(n3934) );
  XNOR U3930 ( .A(n3931), .B(n3969), .Z(n3971) );
  XNOR U3931 ( .A(n3975), .B(n3976), .Z(n3931) );
  AND U3932 ( .A(n132), .B(n3977), .Z(n3976) );
  XNOR U3933 ( .A(n3978), .B(n3979), .Z(n3977) );
  XOR U3934 ( .A(n3980), .B(n3981), .Z(n3969) );
  AND U3935 ( .A(n3982), .B(n3983), .Z(n3981) );
  XNOR U3936 ( .A(n3980), .B(n3973), .Z(n3983) );
  IV U3937 ( .A(n3944), .Z(n3973) );
  XOR U3938 ( .A(n3984), .B(n3985), .Z(n3944) );
  XOR U3939 ( .A(n3986), .B(n3974), .Z(n3985) );
  AND U3940 ( .A(n3954), .B(n3987), .Z(n3974) );
  AND U3941 ( .A(n3988), .B(n3989), .Z(n3986) );
  XOR U3942 ( .A(n3990), .B(n3984), .Z(n3988) );
  XNOR U3943 ( .A(n3941), .B(n3980), .Z(n3982) );
  XNOR U3944 ( .A(n3991), .B(n3992), .Z(n3941) );
  AND U3945 ( .A(n132), .B(n3993), .Z(n3992) );
  XNOR U3946 ( .A(n3994), .B(n3995), .Z(n3993) );
  XOR U3947 ( .A(n3996), .B(n3997), .Z(n3980) );
  AND U3948 ( .A(n3998), .B(n3999), .Z(n3997) );
  XNOR U3949 ( .A(n3996), .B(n3954), .Z(n3999) );
  XOR U3950 ( .A(n4000), .B(n3989), .Z(n3954) );
  XNOR U3951 ( .A(n4001), .B(n3984), .Z(n3989) );
  XOR U3952 ( .A(n4002), .B(n4003), .Z(n3984) );
  AND U3953 ( .A(n4004), .B(n4005), .Z(n4003) );
  XOR U3954 ( .A(n4006), .B(n4002), .Z(n4004) );
  XNOR U3955 ( .A(n4007), .B(n4008), .Z(n4001) );
  AND U3956 ( .A(n4009), .B(n4010), .Z(n4008) );
  XOR U3957 ( .A(n4007), .B(n4011), .Z(n4009) );
  XNOR U3958 ( .A(n3990), .B(n3987), .Z(n4000) );
  AND U3959 ( .A(n4012), .B(n4013), .Z(n3987) );
  XOR U3960 ( .A(n4014), .B(n4015), .Z(n3990) );
  AND U3961 ( .A(n4016), .B(n4017), .Z(n4015) );
  XOR U3962 ( .A(n4014), .B(n4018), .Z(n4016) );
  XNOR U3963 ( .A(n3951), .B(n3996), .Z(n3998) );
  XNOR U3964 ( .A(n4019), .B(n4020), .Z(n3951) );
  AND U3965 ( .A(n132), .B(n4021), .Z(n4020) );
  XNOR U3966 ( .A(n4022), .B(n4023), .Z(n4021) );
  XOR U3967 ( .A(n4024), .B(n4025), .Z(n3996) );
  AND U3968 ( .A(n4026), .B(n4027), .Z(n4025) );
  XNOR U3969 ( .A(n4024), .B(n4012), .Z(n4027) );
  IV U3970 ( .A(n3962), .Z(n4012) );
  XNOR U3971 ( .A(n4028), .B(n4005), .Z(n3962) );
  XNOR U3972 ( .A(n4029), .B(n4011), .Z(n4005) );
  XOR U3973 ( .A(n4030), .B(n4031), .Z(n4011) );
  NOR U3974 ( .A(n4032), .B(n4033), .Z(n4031) );
  XNOR U3975 ( .A(n4030), .B(n4034), .Z(n4032) );
  XNOR U3976 ( .A(n4010), .B(n4002), .Z(n4029) );
  XOR U3977 ( .A(n4035), .B(n4036), .Z(n4002) );
  AND U3978 ( .A(n4037), .B(n4038), .Z(n4036) );
  XNOR U3979 ( .A(n4035), .B(n4039), .Z(n4037) );
  XNOR U3980 ( .A(n4040), .B(n4007), .Z(n4010) );
  XOR U3981 ( .A(n4041), .B(n4042), .Z(n4007) );
  AND U3982 ( .A(n4043), .B(n4044), .Z(n4042) );
  XOR U3983 ( .A(n4041), .B(n4045), .Z(n4043) );
  XNOR U3984 ( .A(n4046), .B(n4047), .Z(n4040) );
  NOR U3985 ( .A(n4048), .B(n4049), .Z(n4047) );
  XOR U3986 ( .A(n4046), .B(n4050), .Z(n4048) );
  XNOR U3987 ( .A(n4006), .B(n4013), .Z(n4028) );
  NOR U3988 ( .A(n3968), .B(n4051), .Z(n4013) );
  XOR U3989 ( .A(n4018), .B(n4017), .Z(n4006) );
  XNOR U3990 ( .A(n4052), .B(n4014), .Z(n4017) );
  XOR U3991 ( .A(n4053), .B(n4054), .Z(n4014) );
  AND U3992 ( .A(n4055), .B(n4056), .Z(n4054) );
  XOR U3993 ( .A(n4053), .B(n4057), .Z(n4055) );
  XNOR U3994 ( .A(n4058), .B(n4059), .Z(n4052) );
  NOR U3995 ( .A(n4060), .B(n4061), .Z(n4059) );
  XNOR U3996 ( .A(n4058), .B(n4062), .Z(n4060) );
  XOR U3997 ( .A(n4063), .B(n4064), .Z(n4018) );
  NOR U3998 ( .A(n4065), .B(n4066), .Z(n4064) );
  XNOR U3999 ( .A(n4063), .B(n4067), .Z(n4065) );
  XNOR U4000 ( .A(n3959), .B(n4024), .Z(n4026) );
  XNOR U4001 ( .A(n4068), .B(n4069), .Z(n3959) );
  AND U4002 ( .A(n132), .B(n4070), .Z(n4069) );
  XNOR U4003 ( .A(n4071), .B(n4072), .Z(n4070) );
  AND U4004 ( .A(n3965), .B(n3968), .Z(n4024) );
  XOR U4005 ( .A(n4073), .B(n4051), .Z(n3968) );
  XNOR U4006 ( .A(p_input[256]), .B(p_input[48]), .Z(n4051) );
  XOR U4007 ( .A(n4039), .B(n4038), .Z(n4073) );
  XNOR U4008 ( .A(n4074), .B(n4045), .Z(n4038) );
  XNOR U4009 ( .A(n4034), .B(n4033), .Z(n4045) );
  XOR U4010 ( .A(n4075), .B(n4030), .Z(n4033) );
  XNOR U4011 ( .A(n3619), .B(p_input[58]), .Z(n4030) );
  XNOR U4012 ( .A(p_input[267]), .B(p_input[59]), .Z(n4075) );
  XOR U4013 ( .A(p_input[268]), .B(p_input[60]), .Z(n4034) );
  XNOR U4014 ( .A(n4044), .B(n4035), .Z(n4074) );
  XNOR U4015 ( .A(n3849), .B(p_input[49]), .Z(n4035) );
  XOR U4016 ( .A(n4076), .B(n4050), .Z(n4044) );
  XNOR U4017 ( .A(p_input[271]), .B(p_input[63]), .Z(n4050) );
  XOR U4018 ( .A(n4041), .B(n4049), .Z(n4076) );
  XOR U4019 ( .A(n4077), .B(n4046), .Z(n4049) );
  XOR U4020 ( .A(p_input[269]), .B(p_input[61]), .Z(n4046) );
  XNOR U4021 ( .A(p_input[270]), .B(p_input[62]), .Z(n4077) );
  XNOR U4022 ( .A(n3388), .B(p_input[57]), .Z(n4041) );
  XNOR U4023 ( .A(n4057), .B(n4056), .Z(n4039) );
  XNOR U4024 ( .A(n4078), .B(n4062), .Z(n4056) );
  XOR U4025 ( .A(p_input[264]), .B(p_input[56]), .Z(n4062) );
  XOR U4026 ( .A(n4053), .B(n4061), .Z(n4078) );
  XOR U4027 ( .A(n4079), .B(n4058), .Z(n4061) );
  XOR U4028 ( .A(p_input[262]), .B(p_input[54]), .Z(n4058) );
  XNOR U4029 ( .A(p_input[263]), .B(p_input[55]), .Z(n4079) );
  XNOR U4030 ( .A(n3391), .B(p_input[50]), .Z(n4053) );
  XNOR U4031 ( .A(n4067), .B(n4066), .Z(n4057) );
  XOR U4032 ( .A(n4080), .B(n4063), .Z(n4066) );
  XOR U4033 ( .A(p_input[259]), .B(p_input[51]), .Z(n4063) );
  XNOR U4034 ( .A(p_input[260]), .B(p_input[52]), .Z(n4080) );
  XOR U4035 ( .A(p_input[261]), .B(p_input[53]), .Z(n4067) );
  XNOR U4036 ( .A(n4081), .B(n4082), .Z(n3965) );
  AND U4037 ( .A(n132), .B(n4083), .Z(n4082) );
  XNOR U4038 ( .A(n4084), .B(n4085), .Z(n132) );
  AND U4039 ( .A(n4086), .B(n4087), .Z(n4085) );
  XOR U4040 ( .A(n3979), .B(n4084), .Z(n4087) );
  XNOR U4041 ( .A(n4088), .B(n4084), .Z(n4086) );
  XOR U4042 ( .A(n4089), .B(n4090), .Z(n4084) );
  AND U4043 ( .A(n4091), .B(n4092), .Z(n4090) );
  XOR U4044 ( .A(n3994), .B(n4089), .Z(n4092) );
  XOR U4045 ( .A(n4089), .B(n3995), .Z(n4091) );
  XOR U4046 ( .A(n4093), .B(n4094), .Z(n4089) );
  AND U4047 ( .A(n4095), .B(n4096), .Z(n4094) );
  XOR U4048 ( .A(n4022), .B(n4093), .Z(n4096) );
  XOR U4049 ( .A(n4093), .B(n4023), .Z(n4095) );
  XOR U4050 ( .A(n4097), .B(n4098), .Z(n4093) );
  AND U4051 ( .A(n4099), .B(n4100), .Z(n4098) );
  XOR U4052 ( .A(n4097), .B(n4071), .Z(n4100) );
  XNOR U4053 ( .A(n4101), .B(n4102), .Z(n3925) );
  AND U4054 ( .A(n136), .B(n4103), .Z(n4102) );
  XNOR U4055 ( .A(n4104), .B(n4105), .Z(n136) );
  AND U4056 ( .A(n4106), .B(n4107), .Z(n4105) );
  XOR U4057 ( .A(n4104), .B(n3935), .Z(n4107) );
  XNOR U4058 ( .A(n4104), .B(n3895), .Z(n4106) );
  XOR U4059 ( .A(n4108), .B(n4109), .Z(n4104) );
  AND U4060 ( .A(n4110), .B(n4111), .Z(n4109) );
  XOR U4061 ( .A(n4108), .B(n3903), .Z(n4110) );
  XOR U4062 ( .A(n4112), .B(n4113), .Z(n3886) );
  AND U4063 ( .A(n140), .B(n4103), .Z(n4113) );
  XNOR U4064 ( .A(n4101), .B(n4112), .Z(n4103) );
  XNOR U4065 ( .A(n4114), .B(n4115), .Z(n140) );
  AND U4066 ( .A(n4116), .B(n4117), .Z(n4115) );
  XNOR U4067 ( .A(n4118), .B(n4114), .Z(n4117) );
  IV U4068 ( .A(n3935), .Z(n4118) );
  XOR U4069 ( .A(n4088), .B(n4119), .Z(n3935) );
  AND U4070 ( .A(n143), .B(n4120), .Z(n4119) );
  XOR U4071 ( .A(n3978), .B(n3975), .Z(n4120) );
  IV U4072 ( .A(n4088), .Z(n3978) );
  XNOR U4073 ( .A(n3895), .B(n4114), .Z(n4116) );
  XOR U4074 ( .A(n4121), .B(n4122), .Z(n3895) );
  AND U4075 ( .A(n159), .B(n4123), .Z(n4122) );
  XOR U4076 ( .A(n4108), .B(n4124), .Z(n4114) );
  AND U4077 ( .A(n4125), .B(n4111), .Z(n4124) );
  XNOR U4078 ( .A(n3945), .B(n4108), .Z(n4111) );
  XOR U4079 ( .A(n3995), .B(n4126), .Z(n3945) );
  AND U4080 ( .A(n143), .B(n4127), .Z(n4126) );
  XOR U4081 ( .A(n3991), .B(n3995), .Z(n4127) );
  XNOR U4082 ( .A(n4128), .B(n4108), .Z(n4125) );
  IV U4083 ( .A(n3903), .Z(n4128) );
  XOR U4084 ( .A(n4129), .B(n4130), .Z(n3903) );
  AND U4085 ( .A(n159), .B(n4131), .Z(n4130) );
  XOR U4086 ( .A(n4132), .B(n4133), .Z(n4108) );
  AND U4087 ( .A(n4134), .B(n4135), .Z(n4133) );
  XNOR U4088 ( .A(n3955), .B(n4132), .Z(n4135) );
  XOR U4089 ( .A(n4023), .B(n4136), .Z(n3955) );
  AND U4090 ( .A(n143), .B(n4137), .Z(n4136) );
  XOR U4091 ( .A(n4019), .B(n4023), .Z(n4137) );
  XOR U4092 ( .A(n4132), .B(n3912), .Z(n4134) );
  XOR U4093 ( .A(n4138), .B(n4139), .Z(n3912) );
  AND U4094 ( .A(n159), .B(n4140), .Z(n4139) );
  XOR U4095 ( .A(n4141), .B(n4142), .Z(n4132) );
  AND U4096 ( .A(n4143), .B(n4144), .Z(n4142) );
  XNOR U4097 ( .A(n4141), .B(n3963), .Z(n4144) );
  XOR U4098 ( .A(n4072), .B(n4145), .Z(n3963) );
  AND U4099 ( .A(n143), .B(n4146), .Z(n4145) );
  XOR U4100 ( .A(n4068), .B(n4072), .Z(n4146) );
  XNOR U4101 ( .A(n4147), .B(n4141), .Z(n4143) );
  IV U4102 ( .A(n3922), .Z(n4147) );
  XOR U4103 ( .A(n4148), .B(n4149), .Z(n3922) );
  AND U4104 ( .A(n159), .B(n4150), .Z(n4149) );
  AND U4105 ( .A(n4112), .B(n4101), .Z(n4141) );
  XNOR U4106 ( .A(n4151), .B(n4152), .Z(n4101) );
  AND U4107 ( .A(n143), .B(n4083), .Z(n4152) );
  XNOR U4108 ( .A(n4081), .B(n4151), .Z(n4083) );
  XNOR U4109 ( .A(n4153), .B(n4154), .Z(n143) );
  AND U4110 ( .A(n4155), .B(n4156), .Z(n4154) );
  XNOR U4111 ( .A(n4153), .B(n3975), .Z(n4156) );
  IV U4112 ( .A(n3979), .Z(n3975) );
  XOR U4113 ( .A(n4157), .B(n4158), .Z(n3979) );
  AND U4114 ( .A(n147), .B(n4159), .Z(n4158) );
  XOR U4115 ( .A(n4160), .B(n4157), .Z(n4159) );
  XNOR U4116 ( .A(n4153), .B(n4088), .Z(n4155) );
  XOR U4117 ( .A(n4161), .B(n4162), .Z(n4088) );
  AND U4118 ( .A(n155), .B(n4123), .Z(n4162) );
  XOR U4119 ( .A(n4121), .B(n4161), .Z(n4123) );
  XOR U4120 ( .A(n4163), .B(n4164), .Z(n4153) );
  AND U4121 ( .A(n4165), .B(n4166), .Z(n4164) );
  XNOR U4122 ( .A(n4163), .B(n3991), .Z(n4166) );
  IV U4123 ( .A(n3994), .Z(n3991) );
  XOR U4124 ( .A(n4167), .B(n4168), .Z(n3994) );
  AND U4125 ( .A(n147), .B(n4169), .Z(n4168) );
  XOR U4126 ( .A(n4170), .B(n4167), .Z(n4169) );
  XOR U4127 ( .A(n3995), .B(n4163), .Z(n4165) );
  XOR U4128 ( .A(n4171), .B(n4172), .Z(n3995) );
  AND U4129 ( .A(n155), .B(n4131), .Z(n4172) );
  XOR U4130 ( .A(n4171), .B(n4129), .Z(n4131) );
  XOR U4131 ( .A(n4173), .B(n4174), .Z(n4163) );
  AND U4132 ( .A(n4175), .B(n4176), .Z(n4174) );
  XNOR U4133 ( .A(n4173), .B(n4019), .Z(n4176) );
  IV U4134 ( .A(n4022), .Z(n4019) );
  XOR U4135 ( .A(n4177), .B(n4178), .Z(n4022) );
  AND U4136 ( .A(n147), .B(n4179), .Z(n4178) );
  XNOR U4137 ( .A(n4180), .B(n4177), .Z(n4179) );
  XOR U4138 ( .A(n4023), .B(n4173), .Z(n4175) );
  XOR U4139 ( .A(n4181), .B(n4182), .Z(n4023) );
  AND U4140 ( .A(n155), .B(n4140), .Z(n4182) );
  XOR U4141 ( .A(n4181), .B(n4138), .Z(n4140) );
  XOR U4142 ( .A(n4097), .B(n4183), .Z(n4173) );
  AND U4143 ( .A(n4099), .B(n4184), .Z(n4183) );
  XNOR U4144 ( .A(n4097), .B(n4068), .Z(n4184) );
  IV U4145 ( .A(n4071), .Z(n4068) );
  XOR U4146 ( .A(n4185), .B(n4186), .Z(n4071) );
  AND U4147 ( .A(n147), .B(n4187), .Z(n4186) );
  XOR U4148 ( .A(n4188), .B(n4185), .Z(n4187) );
  XOR U4149 ( .A(n4072), .B(n4097), .Z(n4099) );
  XOR U4150 ( .A(n4189), .B(n4190), .Z(n4072) );
  AND U4151 ( .A(n155), .B(n4150), .Z(n4190) );
  XOR U4152 ( .A(n4189), .B(n4148), .Z(n4150) );
  AND U4153 ( .A(n4151), .B(n4081), .Z(n4097) );
  XNOR U4154 ( .A(n4191), .B(n4192), .Z(n4081) );
  AND U4155 ( .A(n147), .B(n4193), .Z(n4192) );
  XNOR U4156 ( .A(n4194), .B(n4191), .Z(n4193) );
  XNOR U4157 ( .A(n4195), .B(n4196), .Z(n147) );
  AND U4158 ( .A(n4197), .B(n4198), .Z(n4196) );
  XOR U4159 ( .A(n4160), .B(n4195), .Z(n4198) );
  AND U4160 ( .A(n4199), .B(n4200), .Z(n4160) );
  XNOR U4161 ( .A(n4157), .B(n4195), .Z(n4197) );
  XNOR U4162 ( .A(n4201), .B(n4202), .Z(n4157) );
  AND U4163 ( .A(n151), .B(n4203), .Z(n4202) );
  XNOR U4164 ( .A(n4204), .B(n4205), .Z(n4203) );
  XOR U4165 ( .A(n4206), .B(n4207), .Z(n4195) );
  AND U4166 ( .A(n4208), .B(n4209), .Z(n4207) );
  XNOR U4167 ( .A(n4206), .B(n4199), .Z(n4209) );
  IV U4168 ( .A(n4170), .Z(n4199) );
  XOR U4169 ( .A(n4210), .B(n4211), .Z(n4170) );
  XOR U4170 ( .A(n4212), .B(n4200), .Z(n4211) );
  AND U4171 ( .A(n4180), .B(n4213), .Z(n4200) );
  AND U4172 ( .A(n4214), .B(n4215), .Z(n4212) );
  XOR U4173 ( .A(n4216), .B(n4210), .Z(n4214) );
  XNOR U4174 ( .A(n4167), .B(n4206), .Z(n4208) );
  XNOR U4175 ( .A(n4217), .B(n4218), .Z(n4167) );
  AND U4176 ( .A(n151), .B(n4219), .Z(n4218) );
  XNOR U4177 ( .A(n4220), .B(n4221), .Z(n4219) );
  XOR U4178 ( .A(n4222), .B(n4223), .Z(n4206) );
  AND U4179 ( .A(n4224), .B(n4225), .Z(n4223) );
  XNOR U4180 ( .A(n4222), .B(n4180), .Z(n4225) );
  XOR U4181 ( .A(n4226), .B(n4215), .Z(n4180) );
  XNOR U4182 ( .A(n4227), .B(n4210), .Z(n4215) );
  XOR U4183 ( .A(n4228), .B(n4229), .Z(n4210) );
  AND U4184 ( .A(n4230), .B(n4231), .Z(n4229) );
  XOR U4185 ( .A(n4232), .B(n4228), .Z(n4230) );
  XNOR U4186 ( .A(n4233), .B(n4234), .Z(n4227) );
  AND U4187 ( .A(n4235), .B(n4236), .Z(n4234) );
  XOR U4188 ( .A(n4233), .B(n4237), .Z(n4235) );
  XNOR U4189 ( .A(n4216), .B(n4213), .Z(n4226) );
  AND U4190 ( .A(n4238), .B(n4239), .Z(n4213) );
  XOR U4191 ( .A(n4240), .B(n4241), .Z(n4216) );
  AND U4192 ( .A(n4242), .B(n4243), .Z(n4241) );
  XOR U4193 ( .A(n4240), .B(n4244), .Z(n4242) );
  XNOR U4194 ( .A(n4177), .B(n4222), .Z(n4224) );
  XNOR U4195 ( .A(n4245), .B(n4246), .Z(n4177) );
  AND U4196 ( .A(n151), .B(n4247), .Z(n4246) );
  XNOR U4197 ( .A(n4248), .B(n4249), .Z(n4247) );
  XOR U4198 ( .A(n4250), .B(n4251), .Z(n4222) );
  AND U4199 ( .A(n4252), .B(n4253), .Z(n4251) );
  XNOR U4200 ( .A(n4250), .B(n4238), .Z(n4253) );
  IV U4201 ( .A(n4188), .Z(n4238) );
  XNOR U4202 ( .A(n4254), .B(n4231), .Z(n4188) );
  XNOR U4203 ( .A(n4255), .B(n4237), .Z(n4231) );
  XOR U4204 ( .A(n4256), .B(n4257), .Z(n4237) );
  NOR U4205 ( .A(n4258), .B(n4259), .Z(n4257) );
  XNOR U4206 ( .A(n4256), .B(n4260), .Z(n4258) );
  XNOR U4207 ( .A(n4236), .B(n4228), .Z(n4255) );
  XOR U4208 ( .A(n4261), .B(n4262), .Z(n4228) );
  AND U4209 ( .A(n4263), .B(n4264), .Z(n4262) );
  XNOR U4210 ( .A(n4261), .B(n4265), .Z(n4263) );
  XNOR U4211 ( .A(n4266), .B(n4233), .Z(n4236) );
  XOR U4212 ( .A(n4267), .B(n4268), .Z(n4233) );
  AND U4213 ( .A(n4269), .B(n4270), .Z(n4268) );
  XOR U4214 ( .A(n4267), .B(n4271), .Z(n4269) );
  XNOR U4215 ( .A(n4272), .B(n4273), .Z(n4266) );
  NOR U4216 ( .A(n4274), .B(n4275), .Z(n4273) );
  XOR U4217 ( .A(n4272), .B(n4276), .Z(n4274) );
  XNOR U4218 ( .A(n4232), .B(n4239), .Z(n4254) );
  NOR U4219 ( .A(n4194), .B(n4277), .Z(n4239) );
  XOR U4220 ( .A(n4244), .B(n4243), .Z(n4232) );
  XNOR U4221 ( .A(n4278), .B(n4240), .Z(n4243) );
  XOR U4222 ( .A(n4279), .B(n4280), .Z(n4240) );
  AND U4223 ( .A(n4281), .B(n4282), .Z(n4280) );
  XOR U4224 ( .A(n4279), .B(n4283), .Z(n4281) );
  XNOR U4225 ( .A(n4284), .B(n4285), .Z(n4278) );
  NOR U4226 ( .A(n4286), .B(n4287), .Z(n4285) );
  XNOR U4227 ( .A(n4284), .B(n4288), .Z(n4286) );
  XOR U4228 ( .A(n4289), .B(n4290), .Z(n4244) );
  NOR U4229 ( .A(n4291), .B(n4292), .Z(n4290) );
  XNOR U4230 ( .A(n4289), .B(n4293), .Z(n4291) );
  XNOR U4231 ( .A(n4185), .B(n4250), .Z(n4252) );
  XNOR U4232 ( .A(n4294), .B(n4295), .Z(n4185) );
  AND U4233 ( .A(n151), .B(n4296), .Z(n4295) );
  XNOR U4234 ( .A(n4297), .B(n4298), .Z(n4296) );
  AND U4235 ( .A(n4191), .B(n4194), .Z(n4250) );
  XOR U4236 ( .A(n4299), .B(n4277), .Z(n4194) );
  XNOR U4237 ( .A(p_input[256]), .B(p_input[64]), .Z(n4277) );
  XOR U4238 ( .A(n4265), .B(n4264), .Z(n4299) );
  XNOR U4239 ( .A(n4300), .B(n4271), .Z(n4264) );
  XNOR U4240 ( .A(n4260), .B(n4259), .Z(n4271) );
  XOR U4241 ( .A(n4301), .B(n4256), .Z(n4259) );
  XNOR U4242 ( .A(n3619), .B(p_input[74]), .Z(n4256) );
  XNOR U4243 ( .A(p_input[267]), .B(p_input[75]), .Z(n4301) );
  XOR U4244 ( .A(p_input[268]), .B(p_input[76]), .Z(n4260) );
  XNOR U4245 ( .A(n4270), .B(n4261), .Z(n4300) );
  XNOR U4246 ( .A(n3849), .B(p_input[65]), .Z(n4261) );
  XOR U4247 ( .A(n4302), .B(n4276), .Z(n4270) );
  XNOR U4248 ( .A(p_input[271]), .B(p_input[79]), .Z(n4276) );
  XOR U4249 ( .A(n4267), .B(n4275), .Z(n4302) );
  XOR U4250 ( .A(n4303), .B(n4272), .Z(n4275) );
  XOR U4251 ( .A(p_input[269]), .B(p_input[77]), .Z(n4272) );
  XNOR U4252 ( .A(p_input[270]), .B(p_input[78]), .Z(n4303) );
  XNOR U4253 ( .A(n3388), .B(p_input[73]), .Z(n4267) );
  XNOR U4254 ( .A(n4283), .B(n4282), .Z(n4265) );
  XNOR U4255 ( .A(n4304), .B(n4288), .Z(n4282) );
  XOR U4256 ( .A(p_input[264]), .B(p_input[72]), .Z(n4288) );
  XOR U4257 ( .A(n4279), .B(n4287), .Z(n4304) );
  XOR U4258 ( .A(n4305), .B(n4284), .Z(n4287) );
  XOR U4259 ( .A(p_input[262]), .B(p_input[70]), .Z(n4284) );
  XNOR U4260 ( .A(p_input[263]), .B(p_input[71]), .Z(n4305) );
  XNOR U4261 ( .A(n3391), .B(p_input[66]), .Z(n4279) );
  XNOR U4262 ( .A(n4293), .B(n4292), .Z(n4283) );
  XOR U4263 ( .A(n4306), .B(n4289), .Z(n4292) );
  XOR U4264 ( .A(p_input[259]), .B(p_input[67]), .Z(n4289) );
  XNOR U4265 ( .A(p_input[260]), .B(p_input[68]), .Z(n4306) );
  XOR U4266 ( .A(p_input[261]), .B(p_input[69]), .Z(n4293) );
  XNOR U4267 ( .A(n4307), .B(n4308), .Z(n4191) );
  AND U4268 ( .A(n151), .B(n4309), .Z(n4308) );
  XNOR U4269 ( .A(n4310), .B(n4311), .Z(n151) );
  AND U4270 ( .A(n4312), .B(n4313), .Z(n4311) );
  XOR U4271 ( .A(n4205), .B(n4310), .Z(n4313) );
  XNOR U4272 ( .A(n4314), .B(n4310), .Z(n4312) );
  XOR U4273 ( .A(n4315), .B(n4316), .Z(n4310) );
  AND U4274 ( .A(n4317), .B(n4318), .Z(n4316) );
  XOR U4275 ( .A(n4220), .B(n4315), .Z(n4318) );
  XOR U4276 ( .A(n4315), .B(n4221), .Z(n4317) );
  XOR U4277 ( .A(n4319), .B(n4320), .Z(n4315) );
  AND U4278 ( .A(n4321), .B(n4322), .Z(n4320) );
  XOR U4279 ( .A(n4248), .B(n4319), .Z(n4322) );
  XOR U4280 ( .A(n4319), .B(n4249), .Z(n4321) );
  XOR U4281 ( .A(n4323), .B(n4324), .Z(n4319) );
  AND U4282 ( .A(n4325), .B(n4326), .Z(n4324) );
  XOR U4283 ( .A(n4323), .B(n4297), .Z(n4326) );
  XNOR U4284 ( .A(n4327), .B(n4328), .Z(n4151) );
  AND U4285 ( .A(n155), .B(n4329), .Z(n4328) );
  XNOR U4286 ( .A(n4330), .B(n4331), .Z(n155) );
  AND U4287 ( .A(n4332), .B(n4333), .Z(n4331) );
  XOR U4288 ( .A(n4330), .B(n4161), .Z(n4333) );
  XNOR U4289 ( .A(n4330), .B(n4121), .Z(n4332) );
  XOR U4290 ( .A(n4334), .B(n4335), .Z(n4330) );
  AND U4291 ( .A(n4336), .B(n4337), .Z(n4335) );
  XOR U4292 ( .A(n4334), .B(n4129), .Z(n4336) );
  XOR U4293 ( .A(n4338), .B(n4339), .Z(n4112) );
  AND U4294 ( .A(n159), .B(n4329), .Z(n4339) );
  XNOR U4295 ( .A(n4327), .B(n4338), .Z(n4329) );
  XNOR U4296 ( .A(n4340), .B(n4341), .Z(n159) );
  AND U4297 ( .A(n4342), .B(n4343), .Z(n4341) );
  XNOR U4298 ( .A(n4344), .B(n4340), .Z(n4343) );
  IV U4299 ( .A(n4161), .Z(n4344) );
  XOR U4300 ( .A(n4314), .B(n4345), .Z(n4161) );
  AND U4301 ( .A(n162), .B(n4346), .Z(n4345) );
  XOR U4302 ( .A(n4204), .B(n4201), .Z(n4346) );
  IV U4303 ( .A(n4314), .Z(n4204) );
  XNOR U4304 ( .A(n4121), .B(n4340), .Z(n4342) );
  XOR U4305 ( .A(n4347), .B(n4348), .Z(n4121) );
  AND U4306 ( .A(n178), .B(n4349), .Z(n4348) );
  XOR U4307 ( .A(n4334), .B(n4350), .Z(n4340) );
  AND U4308 ( .A(n4351), .B(n4337), .Z(n4350) );
  XNOR U4309 ( .A(n4171), .B(n4334), .Z(n4337) );
  XOR U4310 ( .A(n4221), .B(n4352), .Z(n4171) );
  AND U4311 ( .A(n162), .B(n4353), .Z(n4352) );
  XOR U4312 ( .A(n4217), .B(n4221), .Z(n4353) );
  XNOR U4313 ( .A(n4354), .B(n4334), .Z(n4351) );
  IV U4314 ( .A(n4129), .Z(n4354) );
  XOR U4315 ( .A(n4355), .B(n4356), .Z(n4129) );
  AND U4316 ( .A(n178), .B(n4357), .Z(n4356) );
  XOR U4317 ( .A(n4358), .B(n4359), .Z(n4334) );
  AND U4318 ( .A(n4360), .B(n4361), .Z(n4359) );
  XNOR U4319 ( .A(n4181), .B(n4358), .Z(n4361) );
  XOR U4320 ( .A(n4249), .B(n4362), .Z(n4181) );
  AND U4321 ( .A(n162), .B(n4363), .Z(n4362) );
  XOR U4322 ( .A(n4245), .B(n4249), .Z(n4363) );
  XOR U4323 ( .A(n4358), .B(n4138), .Z(n4360) );
  XOR U4324 ( .A(n4364), .B(n4365), .Z(n4138) );
  AND U4325 ( .A(n178), .B(n4366), .Z(n4365) );
  XOR U4326 ( .A(n4367), .B(n4368), .Z(n4358) );
  AND U4327 ( .A(n4369), .B(n4370), .Z(n4368) );
  XNOR U4328 ( .A(n4367), .B(n4189), .Z(n4370) );
  XOR U4329 ( .A(n4298), .B(n4371), .Z(n4189) );
  AND U4330 ( .A(n162), .B(n4372), .Z(n4371) );
  XOR U4331 ( .A(n4294), .B(n4298), .Z(n4372) );
  XNOR U4332 ( .A(n4373), .B(n4367), .Z(n4369) );
  IV U4333 ( .A(n4148), .Z(n4373) );
  XOR U4334 ( .A(n4374), .B(n4375), .Z(n4148) );
  AND U4335 ( .A(n178), .B(n4376), .Z(n4375) );
  AND U4336 ( .A(n4338), .B(n4327), .Z(n4367) );
  XNOR U4337 ( .A(n4377), .B(n4378), .Z(n4327) );
  AND U4338 ( .A(n162), .B(n4309), .Z(n4378) );
  XNOR U4339 ( .A(n4307), .B(n4377), .Z(n4309) );
  XNOR U4340 ( .A(n4379), .B(n4380), .Z(n162) );
  AND U4341 ( .A(n4381), .B(n4382), .Z(n4380) );
  XNOR U4342 ( .A(n4379), .B(n4201), .Z(n4382) );
  IV U4343 ( .A(n4205), .Z(n4201) );
  XOR U4344 ( .A(n4383), .B(n4384), .Z(n4205) );
  AND U4345 ( .A(n166), .B(n4385), .Z(n4384) );
  XOR U4346 ( .A(n4386), .B(n4383), .Z(n4385) );
  XNOR U4347 ( .A(n4379), .B(n4314), .Z(n4381) );
  XOR U4348 ( .A(n4387), .B(n4388), .Z(n4314) );
  AND U4349 ( .A(n174), .B(n4349), .Z(n4388) );
  XOR U4350 ( .A(n4347), .B(n4387), .Z(n4349) );
  XOR U4351 ( .A(n4389), .B(n4390), .Z(n4379) );
  AND U4352 ( .A(n4391), .B(n4392), .Z(n4390) );
  XNOR U4353 ( .A(n4389), .B(n4217), .Z(n4392) );
  IV U4354 ( .A(n4220), .Z(n4217) );
  XOR U4355 ( .A(n4393), .B(n4394), .Z(n4220) );
  AND U4356 ( .A(n166), .B(n4395), .Z(n4394) );
  XOR U4357 ( .A(n4396), .B(n4393), .Z(n4395) );
  XOR U4358 ( .A(n4221), .B(n4389), .Z(n4391) );
  XOR U4359 ( .A(n4397), .B(n4398), .Z(n4221) );
  AND U4360 ( .A(n174), .B(n4357), .Z(n4398) );
  XOR U4361 ( .A(n4397), .B(n4355), .Z(n4357) );
  XOR U4362 ( .A(n4399), .B(n4400), .Z(n4389) );
  AND U4363 ( .A(n4401), .B(n4402), .Z(n4400) );
  XNOR U4364 ( .A(n4399), .B(n4245), .Z(n4402) );
  IV U4365 ( .A(n4248), .Z(n4245) );
  XOR U4366 ( .A(n4403), .B(n4404), .Z(n4248) );
  AND U4367 ( .A(n166), .B(n4405), .Z(n4404) );
  XNOR U4368 ( .A(n4406), .B(n4403), .Z(n4405) );
  XOR U4369 ( .A(n4249), .B(n4399), .Z(n4401) );
  XOR U4370 ( .A(n4407), .B(n4408), .Z(n4249) );
  AND U4371 ( .A(n174), .B(n4366), .Z(n4408) );
  XOR U4372 ( .A(n4407), .B(n4364), .Z(n4366) );
  XOR U4373 ( .A(n4323), .B(n4409), .Z(n4399) );
  AND U4374 ( .A(n4325), .B(n4410), .Z(n4409) );
  XNOR U4375 ( .A(n4323), .B(n4294), .Z(n4410) );
  IV U4376 ( .A(n4297), .Z(n4294) );
  XOR U4377 ( .A(n4411), .B(n4412), .Z(n4297) );
  AND U4378 ( .A(n166), .B(n4413), .Z(n4412) );
  XOR U4379 ( .A(n4414), .B(n4411), .Z(n4413) );
  XOR U4380 ( .A(n4298), .B(n4323), .Z(n4325) );
  XOR U4381 ( .A(n4415), .B(n4416), .Z(n4298) );
  AND U4382 ( .A(n174), .B(n4376), .Z(n4416) );
  XOR U4383 ( .A(n4415), .B(n4374), .Z(n4376) );
  AND U4384 ( .A(n4377), .B(n4307), .Z(n4323) );
  XNOR U4385 ( .A(n4417), .B(n4418), .Z(n4307) );
  AND U4386 ( .A(n166), .B(n4419), .Z(n4418) );
  XNOR U4387 ( .A(n4420), .B(n4417), .Z(n4419) );
  XNOR U4388 ( .A(n4421), .B(n4422), .Z(n166) );
  AND U4389 ( .A(n4423), .B(n4424), .Z(n4422) );
  XOR U4390 ( .A(n4386), .B(n4421), .Z(n4424) );
  AND U4391 ( .A(n4425), .B(n4426), .Z(n4386) );
  XNOR U4392 ( .A(n4383), .B(n4421), .Z(n4423) );
  XNOR U4393 ( .A(n4427), .B(n4428), .Z(n4383) );
  AND U4394 ( .A(n170), .B(n4429), .Z(n4428) );
  XNOR U4395 ( .A(n4430), .B(n4431), .Z(n4429) );
  XOR U4396 ( .A(n4432), .B(n4433), .Z(n4421) );
  AND U4397 ( .A(n4434), .B(n4435), .Z(n4433) );
  XNOR U4398 ( .A(n4432), .B(n4425), .Z(n4435) );
  IV U4399 ( .A(n4396), .Z(n4425) );
  XOR U4400 ( .A(n4436), .B(n4437), .Z(n4396) );
  XOR U4401 ( .A(n4438), .B(n4426), .Z(n4437) );
  AND U4402 ( .A(n4406), .B(n4439), .Z(n4426) );
  AND U4403 ( .A(n4440), .B(n4441), .Z(n4438) );
  XOR U4404 ( .A(n4442), .B(n4436), .Z(n4440) );
  XNOR U4405 ( .A(n4393), .B(n4432), .Z(n4434) );
  XNOR U4406 ( .A(n4443), .B(n4444), .Z(n4393) );
  AND U4407 ( .A(n170), .B(n4445), .Z(n4444) );
  XNOR U4408 ( .A(n4446), .B(n4447), .Z(n4445) );
  XOR U4409 ( .A(n4448), .B(n4449), .Z(n4432) );
  AND U4410 ( .A(n4450), .B(n4451), .Z(n4449) );
  XNOR U4411 ( .A(n4448), .B(n4406), .Z(n4451) );
  XOR U4412 ( .A(n4452), .B(n4441), .Z(n4406) );
  XNOR U4413 ( .A(n4453), .B(n4436), .Z(n4441) );
  XOR U4414 ( .A(n4454), .B(n4455), .Z(n4436) );
  AND U4415 ( .A(n4456), .B(n4457), .Z(n4455) );
  XOR U4416 ( .A(n4458), .B(n4454), .Z(n4456) );
  XNOR U4417 ( .A(n4459), .B(n4460), .Z(n4453) );
  AND U4418 ( .A(n4461), .B(n4462), .Z(n4460) );
  XOR U4419 ( .A(n4459), .B(n4463), .Z(n4461) );
  XNOR U4420 ( .A(n4442), .B(n4439), .Z(n4452) );
  AND U4421 ( .A(n4464), .B(n4465), .Z(n4439) );
  XOR U4422 ( .A(n4466), .B(n4467), .Z(n4442) );
  AND U4423 ( .A(n4468), .B(n4469), .Z(n4467) );
  XOR U4424 ( .A(n4466), .B(n4470), .Z(n4468) );
  XNOR U4425 ( .A(n4403), .B(n4448), .Z(n4450) );
  XNOR U4426 ( .A(n4471), .B(n4472), .Z(n4403) );
  AND U4427 ( .A(n170), .B(n4473), .Z(n4472) );
  XNOR U4428 ( .A(n4474), .B(n4475), .Z(n4473) );
  XOR U4429 ( .A(n4476), .B(n4477), .Z(n4448) );
  AND U4430 ( .A(n4478), .B(n4479), .Z(n4477) );
  XNOR U4431 ( .A(n4476), .B(n4464), .Z(n4479) );
  IV U4432 ( .A(n4414), .Z(n4464) );
  XNOR U4433 ( .A(n4480), .B(n4457), .Z(n4414) );
  XNOR U4434 ( .A(n4481), .B(n4463), .Z(n4457) );
  XOR U4435 ( .A(n4482), .B(n4483), .Z(n4463) );
  NOR U4436 ( .A(n4484), .B(n4485), .Z(n4483) );
  XNOR U4437 ( .A(n4482), .B(n4486), .Z(n4484) );
  XNOR U4438 ( .A(n4462), .B(n4454), .Z(n4481) );
  XOR U4439 ( .A(n4487), .B(n4488), .Z(n4454) );
  AND U4440 ( .A(n4489), .B(n4490), .Z(n4488) );
  XNOR U4441 ( .A(n4487), .B(n4491), .Z(n4489) );
  XNOR U4442 ( .A(n4492), .B(n4459), .Z(n4462) );
  XOR U4443 ( .A(n4493), .B(n4494), .Z(n4459) );
  AND U4444 ( .A(n4495), .B(n4496), .Z(n4494) );
  XOR U4445 ( .A(n4493), .B(n4497), .Z(n4495) );
  XNOR U4446 ( .A(n4498), .B(n4499), .Z(n4492) );
  NOR U4447 ( .A(n4500), .B(n4501), .Z(n4499) );
  XOR U4448 ( .A(n4498), .B(n4502), .Z(n4500) );
  XNOR U4449 ( .A(n4458), .B(n4465), .Z(n4480) );
  NOR U4450 ( .A(n4420), .B(n4503), .Z(n4465) );
  XOR U4451 ( .A(n4470), .B(n4469), .Z(n4458) );
  XNOR U4452 ( .A(n4504), .B(n4466), .Z(n4469) );
  XOR U4453 ( .A(n4505), .B(n4506), .Z(n4466) );
  AND U4454 ( .A(n4507), .B(n4508), .Z(n4506) );
  XOR U4455 ( .A(n4505), .B(n4509), .Z(n4507) );
  XNOR U4456 ( .A(n4510), .B(n4511), .Z(n4504) );
  NOR U4457 ( .A(n4512), .B(n4513), .Z(n4511) );
  XNOR U4458 ( .A(n4510), .B(n4514), .Z(n4512) );
  XOR U4459 ( .A(n4515), .B(n4516), .Z(n4470) );
  NOR U4460 ( .A(n4517), .B(n4518), .Z(n4516) );
  XNOR U4461 ( .A(n4515), .B(n4519), .Z(n4517) );
  XNOR U4462 ( .A(n4411), .B(n4476), .Z(n4478) );
  XNOR U4463 ( .A(n4520), .B(n4521), .Z(n4411) );
  AND U4464 ( .A(n170), .B(n4522), .Z(n4521) );
  XNOR U4465 ( .A(n4523), .B(n4524), .Z(n4522) );
  AND U4466 ( .A(n4417), .B(n4420), .Z(n4476) );
  XOR U4467 ( .A(n4525), .B(n4503), .Z(n4420) );
  XNOR U4468 ( .A(p_input[256]), .B(p_input[80]), .Z(n4503) );
  XOR U4469 ( .A(n4491), .B(n4490), .Z(n4525) );
  XNOR U4470 ( .A(n4526), .B(n4497), .Z(n4490) );
  XNOR U4471 ( .A(n4486), .B(n4485), .Z(n4497) );
  XOR U4472 ( .A(n4527), .B(n4482), .Z(n4485) );
  XNOR U4473 ( .A(n3619), .B(p_input[90]), .Z(n4482) );
  XNOR U4474 ( .A(p_input[267]), .B(p_input[91]), .Z(n4527) );
  XOR U4475 ( .A(p_input[268]), .B(p_input[92]), .Z(n4486) );
  XNOR U4476 ( .A(n4496), .B(n4487), .Z(n4526) );
  XNOR U4477 ( .A(n3849), .B(p_input[81]), .Z(n4487) );
  XOR U4478 ( .A(n4528), .B(n4502), .Z(n4496) );
  XNOR U4479 ( .A(p_input[271]), .B(p_input[95]), .Z(n4502) );
  XOR U4480 ( .A(n4493), .B(n4501), .Z(n4528) );
  XOR U4481 ( .A(n4529), .B(n4498), .Z(n4501) );
  XOR U4482 ( .A(p_input[269]), .B(p_input[93]), .Z(n4498) );
  XNOR U4483 ( .A(p_input[270]), .B(p_input[94]), .Z(n4529) );
  XNOR U4484 ( .A(n3388), .B(p_input[89]), .Z(n4493) );
  XNOR U4485 ( .A(n4509), .B(n4508), .Z(n4491) );
  XNOR U4486 ( .A(n4530), .B(n4514), .Z(n4508) );
  XOR U4487 ( .A(p_input[264]), .B(p_input[88]), .Z(n4514) );
  XOR U4488 ( .A(n4505), .B(n4513), .Z(n4530) );
  XOR U4489 ( .A(n4531), .B(n4510), .Z(n4513) );
  XOR U4490 ( .A(p_input[262]), .B(p_input[86]), .Z(n4510) );
  XNOR U4491 ( .A(p_input[263]), .B(p_input[87]), .Z(n4531) );
  XNOR U4492 ( .A(n3391), .B(p_input[82]), .Z(n4505) );
  XNOR U4493 ( .A(n4519), .B(n4518), .Z(n4509) );
  XOR U4494 ( .A(n4532), .B(n4515), .Z(n4518) );
  XOR U4495 ( .A(p_input[259]), .B(p_input[83]), .Z(n4515) );
  XNOR U4496 ( .A(p_input[260]), .B(p_input[84]), .Z(n4532) );
  XOR U4497 ( .A(p_input[261]), .B(p_input[85]), .Z(n4519) );
  XNOR U4498 ( .A(n4533), .B(n4534), .Z(n4417) );
  AND U4499 ( .A(n170), .B(n4535), .Z(n4534) );
  XNOR U4500 ( .A(n4536), .B(n4537), .Z(n170) );
  AND U4501 ( .A(n4538), .B(n4539), .Z(n4537) );
  XOR U4502 ( .A(n4431), .B(n4536), .Z(n4539) );
  XNOR U4503 ( .A(n4540), .B(n4536), .Z(n4538) );
  XOR U4504 ( .A(n4541), .B(n4542), .Z(n4536) );
  AND U4505 ( .A(n4543), .B(n4544), .Z(n4542) );
  XOR U4506 ( .A(n4446), .B(n4541), .Z(n4544) );
  XOR U4507 ( .A(n4541), .B(n4447), .Z(n4543) );
  XOR U4508 ( .A(n4545), .B(n4546), .Z(n4541) );
  AND U4509 ( .A(n4547), .B(n4548), .Z(n4546) );
  XOR U4510 ( .A(n4474), .B(n4545), .Z(n4548) );
  XOR U4511 ( .A(n4545), .B(n4475), .Z(n4547) );
  XOR U4512 ( .A(n4549), .B(n4550), .Z(n4545) );
  AND U4513 ( .A(n4551), .B(n4552), .Z(n4550) );
  XOR U4514 ( .A(n4549), .B(n4523), .Z(n4552) );
  XNOR U4515 ( .A(n4553), .B(n4554), .Z(n4377) );
  AND U4516 ( .A(n174), .B(n4555), .Z(n4554) );
  XNOR U4517 ( .A(n4556), .B(n4557), .Z(n174) );
  AND U4518 ( .A(n4558), .B(n4559), .Z(n4557) );
  XOR U4519 ( .A(n4556), .B(n4387), .Z(n4559) );
  XNOR U4520 ( .A(n4556), .B(n4347), .Z(n4558) );
  XOR U4521 ( .A(n4560), .B(n4561), .Z(n4556) );
  AND U4522 ( .A(n4562), .B(n4563), .Z(n4561) );
  XOR U4523 ( .A(n4560), .B(n4355), .Z(n4562) );
  XOR U4524 ( .A(n4564), .B(n4565), .Z(n4338) );
  AND U4525 ( .A(n178), .B(n4555), .Z(n4565) );
  XNOR U4526 ( .A(n4553), .B(n4564), .Z(n4555) );
  XNOR U4527 ( .A(n4566), .B(n4567), .Z(n178) );
  AND U4528 ( .A(n4568), .B(n4569), .Z(n4567) );
  XNOR U4529 ( .A(n4570), .B(n4566), .Z(n4569) );
  IV U4530 ( .A(n4387), .Z(n4570) );
  XOR U4531 ( .A(n4540), .B(n4571), .Z(n4387) );
  AND U4532 ( .A(n181), .B(n4572), .Z(n4571) );
  XOR U4533 ( .A(n4430), .B(n4427), .Z(n4572) );
  IV U4534 ( .A(n4540), .Z(n4430) );
  XNOR U4535 ( .A(n4347), .B(n4566), .Z(n4568) );
  XOR U4536 ( .A(n4573), .B(n4574), .Z(n4347) );
  AND U4537 ( .A(n197), .B(n4575), .Z(n4574) );
  XOR U4538 ( .A(n4560), .B(n4576), .Z(n4566) );
  AND U4539 ( .A(n4577), .B(n4563), .Z(n4576) );
  XNOR U4540 ( .A(n4397), .B(n4560), .Z(n4563) );
  XOR U4541 ( .A(n4447), .B(n4578), .Z(n4397) );
  AND U4542 ( .A(n181), .B(n4579), .Z(n4578) );
  XOR U4543 ( .A(n4443), .B(n4447), .Z(n4579) );
  XNOR U4544 ( .A(n4580), .B(n4560), .Z(n4577) );
  IV U4545 ( .A(n4355), .Z(n4580) );
  XOR U4546 ( .A(n4581), .B(n4582), .Z(n4355) );
  AND U4547 ( .A(n197), .B(n4583), .Z(n4582) );
  XOR U4548 ( .A(n4584), .B(n4585), .Z(n4560) );
  AND U4549 ( .A(n4586), .B(n4587), .Z(n4585) );
  XNOR U4550 ( .A(n4407), .B(n4584), .Z(n4587) );
  XOR U4551 ( .A(n4475), .B(n4588), .Z(n4407) );
  AND U4552 ( .A(n181), .B(n4589), .Z(n4588) );
  XOR U4553 ( .A(n4471), .B(n4475), .Z(n4589) );
  XOR U4554 ( .A(n4584), .B(n4364), .Z(n4586) );
  XOR U4555 ( .A(n4590), .B(n4591), .Z(n4364) );
  AND U4556 ( .A(n197), .B(n4592), .Z(n4591) );
  XOR U4557 ( .A(n4593), .B(n4594), .Z(n4584) );
  AND U4558 ( .A(n4595), .B(n4596), .Z(n4594) );
  XNOR U4559 ( .A(n4593), .B(n4415), .Z(n4596) );
  XOR U4560 ( .A(n4524), .B(n4597), .Z(n4415) );
  AND U4561 ( .A(n181), .B(n4598), .Z(n4597) );
  XOR U4562 ( .A(n4520), .B(n4524), .Z(n4598) );
  XNOR U4563 ( .A(n4599), .B(n4593), .Z(n4595) );
  IV U4564 ( .A(n4374), .Z(n4599) );
  XOR U4565 ( .A(n4600), .B(n4601), .Z(n4374) );
  AND U4566 ( .A(n197), .B(n4602), .Z(n4601) );
  AND U4567 ( .A(n4564), .B(n4553), .Z(n4593) );
  XNOR U4568 ( .A(n4603), .B(n4604), .Z(n4553) );
  AND U4569 ( .A(n181), .B(n4535), .Z(n4604) );
  XNOR U4570 ( .A(n4533), .B(n4603), .Z(n4535) );
  XNOR U4571 ( .A(n4605), .B(n4606), .Z(n181) );
  AND U4572 ( .A(n4607), .B(n4608), .Z(n4606) );
  XNOR U4573 ( .A(n4605), .B(n4427), .Z(n4608) );
  IV U4574 ( .A(n4431), .Z(n4427) );
  XOR U4575 ( .A(n4609), .B(n4610), .Z(n4431) );
  AND U4576 ( .A(n185), .B(n4611), .Z(n4610) );
  XOR U4577 ( .A(n4612), .B(n4609), .Z(n4611) );
  XNOR U4578 ( .A(n4605), .B(n4540), .Z(n4607) );
  XOR U4579 ( .A(n4613), .B(n4614), .Z(n4540) );
  AND U4580 ( .A(n193), .B(n4575), .Z(n4614) );
  XOR U4581 ( .A(n4573), .B(n4613), .Z(n4575) );
  XOR U4582 ( .A(n4615), .B(n4616), .Z(n4605) );
  AND U4583 ( .A(n4617), .B(n4618), .Z(n4616) );
  XNOR U4584 ( .A(n4615), .B(n4443), .Z(n4618) );
  IV U4585 ( .A(n4446), .Z(n4443) );
  XOR U4586 ( .A(n4619), .B(n4620), .Z(n4446) );
  AND U4587 ( .A(n185), .B(n4621), .Z(n4620) );
  XOR U4588 ( .A(n4622), .B(n4619), .Z(n4621) );
  XOR U4589 ( .A(n4447), .B(n4615), .Z(n4617) );
  XOR U4590 ( .A(n4623), .B(n4624), .Z(n4447) );
  AND U4591 ( .A(n193), .B(n4583), .Z(n4624) );
  XOR U4592 ( .A(n4623), .B(n4581), .Z(n4583) );
  XOR U4593 ( .A(n4625), .B(n4626), .Z(n4615) );
  AND U4594 ( .A(n4627), .B(n4628), .Z(n4626) );
  XNOR U4595 ( .A(n4625), .B(n4471), .Z(n4628) );
  IV U4596 ( .A(n4474), .Z(n4471) );
  XOR U4597 ( .A(n4629), .B(n4630), .Z(n4474) );
  AND U4598 ( .A(n185), .B(n4631), .Z(n4630) );
  XNOR U4599 ( .A(n4632), .B(n4629), .Z(n4631) );
  XOR U4600 ( .A(n4475), .B(n4625), .Z(n4627) );
  XOR U4601 ( .A(n4633), .B(n4634), .Z(n4475) );
  AND U4602 ( .A(n193), .B(n4592), .Z(n4634) );
  XOR U4603 ( .A(n4633), .B(n4590), .Z(n4592) );
  XOR U4604 ( .A(n4549), .B(n4635), .Z(n4625) );
  AND U4605 ( .A(n4551), .B(n4636), .Z(n4635) );
  XNOR U4606 ( .A(n4549), .B(n4520), .Z(n4636) );
  IV U4607 ( .A(n4523), .Z(n4520) );
  XOR U4608 ( .A(n4637), .B(n4638), .Z(n4523) );
  AND U4609 ( .A(n185), .B(n4639), .Z(n4638) );
  XOR U4610 ( .A(n4640), .B(n4637), .Z(n4639) );
  XOR U4611 ( .A(n4524), .B(n4549), .Z(n4551) );
  XOR U4612 ( .A(n4641), .B(n4642), .Z(n4524) );
  AND U4613 ( .A(n193), .B(n4602), .Z(n4642) );
  XOR U4614 ( .A(n4641), .B(n4600), .Z(n4602) );
  AND U4615 ( .A(n4603), .B(n4533), .Z(n4549) );
  XNOR U4616 ( .A(n4643), .B(n4644), .Z(n4533) );
  AND U4617 ( .A(n185), .B(n4645), .Z(n4644) );
  XNOR U4618 ( .A(n4646), .B(n4643), .Z(n4645) );
  XNOR U4619 ( .A(n4647), .B(n4648), .Z(n185) );
  AND U4620 ( .A(n4649), .B(n4650), .Z(n4648) );
  XOR U4621 ( .A(n4612), .B(n4647), .Z(n4650) );
  AND U4622 ( .A(n4651), .B(n4652), .Z(n4612) );
  XNOR U4623 ( .A(n4609), .B(n4647), .Z(n4649) );
  XNOR U4624 ( .A(n4653), .B(n4654), .Z(n4609) );
  AND U4625 ( .A(n189), .B(n4655), .Z(n4654) );
  XNOR U4626 ( .A(n4656), .B(n4657), .Z(n4655) );
  XOR U4627 ( .A(n4658), .B(n4659), .Z(n4647) );
  AND U4628 ( .A(n4660), .B(n4661), .Z(n4659) );
  XNOR U4629 ( .A(n4658), .B(n4651), .Z(n4661) );
  IV U4630 ( .A(n4622), .Z(n4651) );
  XOR U4631 ( .A(n4662), .B(n4663), .Z(n4622) );
  XOR U4632 ( .A(n4664), .B(n4652), .Z(n4663) );
  AND U4633 ( .A(n4632), .B(n4665), .Z(n4652) );
  AND U4634 ( .A(n4666), .B(n4667), .Z(n4664) );
  XOR U4635 ( .A(n4668), .B(n4662), .Z(n4666) );
  XNOR U4636 ( .A(n4619), .B(n4658), .Z(n4660) );
  XNOR U4637 ( .A(n4669), .B(n4670), .Z(n4619) );
  AND U4638 ( .A(n189), .B(n4671), .Z(n4670) );
  XNOR U4639 ( .A(n4672), .B(n4673), .Z(n4671) );
  XOR U4640 ( .A(n4674), .B(n4675), .Z(n4658) );
  AND U4641 ( .A(n4676), .B(n4677), .Z(n4675) );
  XNOR U4642 ( .A(n4674), .B(n4632), .Z(n4677) );
  XOR U4643 ( .A(n4678), .B(n4667), .Z(n4632) );
  XNOR U4644 ( .A(n4679), .B(n4662), .Z(n4667) );
  XOR U4645 ( .A(n4680), .B(n4681), .Z(n4662) );
  AND U4646 ( .A(n4682), .B(n4683), .Z(n4681) );
  XOR U4647 ( .A(n4684), .B(n4680), .Z(n4682) );
  XNOR U4648 ( .A(n4685), .B(n4686), .Z(n4679) );
  AND U4649 ( .A(n4687), .B(n4688), .Z(n4686) );
  XOR U4650 ( .A(n4685), .B(n4689), .Z(n4687) );
  XNOR U4651 ( .A(n4668), .B(n4665), .Z(n4678) );
  AND U4652 ( .A(n4690), .B(n4691), .Z(n4665) );
  XOR U4653 ( .A(n4692), .B(n4693), .Z(n4668) );
  AND U4654 ( .A(n4694), .B(n4695), .Z(n4693) );
  XOR U4655 ( .A(n4692), .B(n4696), .Z(n4694) );
  XNOR U4656 ( .A(n4629), .B(n4674), .Z(n4676) );
  XNOR U4657 ( .A(n4697), .B(n4698), .Z(n4629) );
  AND U4658 ( .A(n189), .B(n4699), .Z(n4698) );
  XNOR U4659 ( .A(n4700), .B(n4701), .Z(n4699) );
  XOR U4660 ( .A(n4702), .B(n4703), .Z(n4674) );
  AND U4661 ( .A(n4704), .B(n4705), .Z(n4703) );
  XNOR U4662 ( .A(n4702), .B(n4690), .Z(n4705) );
  IV U4663 ( .A(n4640), .Z(n4690) );
  XNOR U4664 ( .A(n4706), .B(n4683), .Z(n4640) );
  XNOR U4665 ( .A(n4707), .B(n4689), .Z(n4683) );
  XNOR U4666 ( .A(n4708), .B(n4709), .Z(n4689) );
  NOR U4667 ( .A(n4710), .B(n4711), .Z(n4709) );
  XOR U4668 ( .A(n4708), .B(n4712), .Z(n4710) );
  XNOR U4669 ( .A(n4688), .B(n4680), .Z(n4707) );
  XOR U4670 ( .A(n4713), .B(n4714), .Z(n4680) );
  AND U4671 ( .A(n4715), .B(n4716), .Z(n4714) );
  XOR U4672 ( .A(n4713), .B(n4717), .Z(n4715) );
  XNOR U4673 ( .A(n4718), .B(n4685), .Z(n4688) );
  XOR U4674 ( .A(n4719), .B(n4720), .Z(n4685) );
  AND U4675 ( .A(n4721), .B(n4722), .Z(n4720) );
  XNOR U4676 ( .A(n4723), .B(n4724), .Z(n4721) );
  IV U4677 ( .A(n4719), .Z(n4723) );
  XNOR U4678 ( .A(n4725), .B(n4726), .Z(n4718) );
  NOR U4679 ( .A(n4727), .B(n4728), .Z(n4726) );
  XNOR U4680 ( .A(n4725), .B(n4729), .Z(n4727) );
  XNOR U4681 ( .A(n4684), .B(n4691), .Z(n4706) );
  NOR U4682 ( .A(n4646), .B(n4730), .Z(n4691) );
  XOR U4683 ( .A(n4696), .B(n4695), .Z(n4684) );
  XNOR U4684 ( .A(n4731), .B(n4692), .Z(n4695) );
  XOR U4685 ( .A(n4732), .B(n4733), .Z(n4692) );
  AND U4686 ( .A(n4734), .B(n4735), .Z(n4733) );
  XOR U4687 ( .A(n4732), .B(n4736), .Z(n4734) );
  XNOR U4688 ( .A(n4737), .B(n4738), .Z(n4731) );
  NOR U4689 ( .A(n4739), .B(n4740), .Z(n4738) );
  XNOR U4690 ( .A(n4737), .B(n4741), .Z(n4739) );
  XOR U4691 ( .A(n4742), .B(n4743), .Z(n4696) );
  NOR U4692 ( .A(n4744), .B(n4745), .Z(n4743) );
  XNOR U4693 ( .A(n4742), .B(n4746), .Z(n4744) );
  XNOR U4694 ( .A(n4637), .B(n4702), .Z(n4704) );
  XNOR U4695 ( .A(n4747), .B(n4748), .Z(n4637) );
  AND U4696 ( .A(n189), .B(n4749), .Z(n4748) );
  XNOR U4697 ( .A(n4750), .B(n4751), .Z(n4749) );
  AND U4698 ( .A(n4643), .B(n4646), .Z(n4702) );
  XOR U4699 ( .A(n4752), .B(n4730), .Z(n4646) );
  XNOR U4700 ( .A(p_input[256]), .B(p_input[96]), .Z(n4730) );
  XNOR U4701 ( .A(n4717), .B(n4716), .Z(n4752) );
  XNOR U4702 ( .A(n4753), .B(n4724), .Z(n4716) );
  XNOR U4703 ( .A(n4712), .B(n4711), .Z(n4724) );
  XNOR U4704 ( .A(n4754), .B(n4708), .Z(n4711) );
  XNOR U4705 ( .A(p_input[106]), .B(p_input[266]), .Z(n4708) );
  XOR U4706 ( .A(p_input[107]), .B(n3382), .Z(n4754) );
  XOR U4707 ( .A(p_input[108]), .B(p_input[268]), .Z(n4712) );
  XNOR U4708 ( .A(n4722), .B(n4713), .Z(n4753) );
  XNOR U4709 ( .A(n3849), .B(p_input[97]), .Z(n4713) );
  XNOR U4710 ( .A(n4755), .B(n4729), .Z(n4722) );
  XNOR U4711 ( .A(p_input[111]), .B(n3385), .Z(n4729) );
  XOR U4712 ( .A(n4719), .B(n4728), .Z(n4755) );
  XOR U4713 ( .A(n4756), .B(n4725), .Z(n4728) );
  XOR U4714 ( .A(p_input[109]), .B(p_input[269]), .Z(n4725) );
  XOR U4715 ( .A(p_input[110]), .B(n3387), .Z(n4756) );
  XOR U4716 ( .A(p_input[105]), .B(p_input[265]), .Z(n4719) );
  XOR U4717 ( .A(n4736), .B(n4735), .Z(n4717) );
  XNOR U4718 ( .A(n4757), .B(n4741), .Z(n4735) );
  XOR U4719 ( .A(p_input[104]), .B(p_input[264]), .Z(n4741) );
  XOR U4720 ( .A(n4732), .B(n4740), .Z(n4757) );
  XOR U4721 ( .A(n4758), .B(n4737), .Z(n4740) );
  XOR U4722 ( .A(p_input[102]), .B(p_input[262]), .Z(n4737) );
  XOR U4723 ( .A(p_input[103]), .B(n3625), .Z(n4758) );
  XNOR U4724 ( .A(n3391), .B(p_input[98]), .Z(n4732) );
  XNOR U4725 ( .A(n4746), .B(n4745), .Z(n4736) );
  XOR U4726 ( .A(n4759), .B(n4742), .Z(n4745) );
  XOR U4727 ( .A(p_input[259]), .B(p_input[99]), .Z(n4742) );
  XOR U4728 ( .A(p_input[100]), .B(n3627), .Z(n4759) );
  XOR U4729 ( .A(p_input[101]), .B(p_input[261]), .Z(n4746) );
  XNOR U4730 ( .A(n4760), .B(n4761), .Z(n4643) );
  AND U4731 ( .A(n189), .B(n4762), .Z(n4761) );
  XNOR U4732 ( .A(n4763), .B(n4764), .Z(n189) );
  AND U4733 ( .A(n4765), .B(n4766), .Z(n4764) );
  XOR U4734 ( .A(n4657), .B(n4763), .Z(n4766) );
  XNOR U4735 ( .A(n4767), .B(n4763), .Z(n4765) );
  XOR U4736 ( .A(n4768), .B(n4769), .Z(n4763) );
  AND U4737 ( .A(n4770), .B(n4771), .Z(n4769) );
  XOR U4738 ( .A(n4672), .B(n4768), .Z(n4771) );
  XOR U4739 ( .A(n4768), .B(n4673), .Z(n4770) );
  XOR U4740 ( .A(n4772), .B(n4773), .Z(n4768) );
  AND U4741 ( .A(n4774), .B(n4775), .Z(n4773) );
  XOR U4742 ( .A(n4700), .B(n4772), .Z(n4775) );
  XOR U4743 ( .A(n4772), .B(n4701), .Z(n4774) );
  XOR U4744 ( .A(n4776), .B(n4777), .Z(n4772) );
  AND U4745 ( .A(n4778), .B(n4779), .Z(n4777) );
  XOR U4746 ( .A(n4776), .B(n4750), .Z(n4779) );
  XNOR U4747 ( .A(n4780), .B(n4781), .Z(n4603) );
  AND U4748 ( .A(n193), .B(n4782), .Z(n4781) );
  XNOR U4749 ( .A(n4783), .B(n4784), .Z(n193) );
  AND U4750 ( .A(n4785), .B(n4786), .Z(n4784) );
  XOR U4751 ( .A(n4783), .B(n4613), .Z(n4786) );
  XNOR U4752 ( .A(n4783), .B(n4573), .Z(n4785) );
  XOR U4753 ( .A(n4787), .B(n4788), .Z(n4783) );
  AND U4754 ( .A(n4789), .B(n4790), .Z(n4788) );
  XOR U4755 ( .A(n4787), .B(n4581), .Z(n4789) );
  XOR U4756 ( .A(n4791), .B(n4792), .Z(n4564) );
  AND U4757 ( .A(n197), .B(n4782), .Z(n4792) );
  XNOR U4758 ( .A(n4780), .B(n4791), .Z(n4782) );
  XNOR U4759 ( .A(n4793), .B(n4794), .Z(n197) );
  AND U4760 ( .A(n4795), .B(n4796), .Z(n4794) );
  XNOR U4761 ( .A(n4797), .B(n4793), .Z(n4796) );
  IV U4762 ( .A(n4613), .Z(n4797) );
  XOR U4763 ( .A(n4767), .B(n4798), .Z(n4613) );
  AND U4764 ( .A(n200), .B(n4799), .Z(n4798) );
  XOR U4765 ( .A(n4656), .B(n4653), .Z(n4799) );
  IV U4766 ( .A(n4767), .Z(n4656) );
  XNOR U4767 ( .A(n4573), .B(n4793), .Z(n4795) );
  XOR U4768 ( .A(n4800), .B(n4801), .Z(n4573) );
  AND U4769 ( .A(n216), .B(n4802), .Z(n4801) );
  XOR U4770 ( .A(n4787), .B(n4803), .Z(n4793) );
  AND U4771 ( .A(n4804), .B(n4790), .Z(n4803) );
  XNOR U4772 ( .A(n4623), .B(n4787), .Z(n4790) );
  XOR U4773 ( .A(n4673), .B(n4805), .Z(n4623) );
  AND U4774 ( .A(n200), .B(n4806), .Z(n4805) );
  XOR U4775 ( .A(n4669), .B(n4673), .Z(n4806) );
  XNOR U4776 ( .A(n4807), .B(n4787), .Z(n4804) );
  IV U4777 ( .A(n4581), .Z(n4807) );
  XOR U4778 ( .A(n4808), .B(n4809), .Z(n4581) );
  AND U4779 ( .A(n216), .B(n4810), .Z(n4809) );
  XOR U4780 ( .A(n4811), .B(n4812), .Z(n4787) );
  AND U4781 ( .A(n4813), .B(n4814), .Z(n4812) );
  XNOR U4782 ( .A(n4633), .B(n4811), .Z(n4814) );
  XOR U4783 ( .A(n4701), .B(n4815), .Z(n4633) );
  AND U4784 ( .A(n200), .B(n4816), .Z(n4815) );
  XOR U4785 ( .A(n4697), .B(n4701), .Z(n4816) );
  XOR U4786 ( .A(n4811), .B(n4590), .Z(n4813) );
  XOR U4787 ( .A(n4817), .B(n4818), .Z(n4590) );
  AND U4788 ( .A(n216), .B(n4819), .Z(n4818) );
  XOR U4789 ( .A(n4820), .B(n4821), .Z(n4811) );
  AND U4790 ( .A(n4822), .B(n4823), .Z(n4821) );
  XNOR U4791 ( .A(n4820), .B(n4641), .Z(n4823) );
  XOR U4792 ( .A(n4751), .B(n4824), .Z(n4641) );
  AND U4793 ( .A(n200), .B(n4825), .Z(n4824) );
  XOR U4794 ( .A(n4747), .B(n4751), .Z(n4825) );
  XNOR U4795 ( .A(n4826), .B(n4820), .Z(n4822) );
  IV U4796 ( .A(n4600), .Z(n4826) );
  XOR U4797 ( .A(n4827), .B(n4828), .Z(n4600) );
  AND U4798 ( .A(n216), .B(n4829), .Z(n4828) );
  AND U4799 ( .A(n4791), .B(n4780), .Z(n4820) );
  XNOR U4800 ( .A(n4830), .B(n4831), .Z(n4780) );
  AND U4801 ( .A(n200), .B(n4762), .Z(n4831) );
  XNOR U4802 ( .A(n4760), .B(n4830), .Z(n4762) );
  XNOR U4803 ( .A(n4832), .B(n4833), .Z(n200) );
  AND U4804 ( .A(n4834), .B(n4835), .Z(n4833) );
  XNOR U4805 ( .A(n4832), .B(n4653), .Z(n4835) );
  IV U4806 ( .A(n4657), .Z(n4653) );
  XOR U4807 ( .A(n4836), .B(n4837), .Z(n4657) );
  AND U4808 ( .A(n204), .B(n4838), .Z(n4837) );
  XOR U4809 ( .A(n4839), .B(n4836), .Z(n4838) );
  XNOR U4810 ( .A(n4832), .B(n4767), .Z(n4834) );
  XOR U4811 ( .A(n4840), .B(n4841), .Z(n4767) );
  AND U4812 ( .A(n212), .B(n4802), .Z(n4841) );
  XOR U4813 ( .A(n4800), .B(n4840), .Z(n4802) );
  XOR U4814 ( .A(n4842), .B(n4843), .Z(n4832) );
  AND U4815 ( .A(n4844), .B(n4845), .Z(n4843) );
  XNOR U4816 ( .A(n4842), .B(n4669), .Z(n4845) );
  IV U4817 ( .A(n4672), .Z(n4669) );
  XOR U4818 ( .A(n4846), .B(n4847), .Z(n4672) );
  AND U4819 ( .A(n204), .B(n4848), .Z(n4847) );
  XOR U4820 ( .A(n4849), .B(n4846), .Z(n4848) );
  XOR U4821 ( .A(n4673), .B(n4842), .Z(n4844) );
  XOR U4822 ( .A(n4850), .B(n4851), .Z(n4673) );
  AND U4823 ( .A(n212), .B(n4810), .Z(n4851) );
  XOR U4824 ( .A(n4850), .B(n4808), .Z(n4810) );
  XOR U4825 ( .A(n4852), .B(n4853), .Z(n4842) );
  AND U4826 ( .A(n4854), .B(n4855), .Z(n4853) );
  XNOR U4827 ( .A(n4852), .B(n4697), .Z(n4855) );
  IV U4828 ( .A(n4700), .Z(n4697) );
  XOR U4829 ( .A(n4856), .B(n4857), .Z(n4700) );
  AND U4830 ( .A(n204), .B(n4858), .Z(n4857) );
  XNOR U4831 ( .A(n4859), .B(n4856), .Z(n4858) );
  XOR U4832 ( .A(n4701), .B(n4852), .Z(n4854) );
  XOR U4833 ( .A(n4860), .B(n4861), .Z(n4701) );
  AND U4834 ( .A(n212), .B(n4819), .Z(n4861) );
  XOR U4835 ( .A(n4860), .B(n4817), .Z(n4819) );
  XOR U4836 ( .A(n4776), .B(n4862), .Z(n4852) );
  AND U4837 ( .A(n4778), .B(n4863), .Z(n4862) );
  XNOR U4838 ( .A(n4776), .B(n4747), .Z(n4863) );
  IV U4839 ( .A(n4750), .Z(n4747) );
  XOR U4840 ( .A(n4864), .B(n4865), .Z(n4750) );
  AND U4841 ( .A(n204), .B(n4866), .Z(n4865) );
  XOR U4842 ( .A(n4867), .B(n4864), .Z(n4866) );
  XOR U4843 ( .A(n4751), .B(n4776), .Z(n4778) );
  XOR U4844 ( .A(n4868), .B(n4869), .Z(n4751) );
  AND U4845 ( .A(n212), .B(n4829), .Z(n4869) );
  XOR U4846 ( .A(n4868), .B(n4827), .Z(n4829) );
  AND U4847 ( .A(n4830), .B(n4760), .Z(n4776) );
  XNOR U4848 ( .A(n4870), .B(n4871), .Z(n4760) );
  AND U4849 ( .A(n204), .B(n4872), .Z(n4871) );
  XNOR U4850 ( .A(n4873), .B(n4870), .Z(n4872) );
  XNOR U4851 ( .A(n4874), .B(n4875), .Z(n204) );
  AND U4852 ( .A(n4876), .B(n4877), .Z(n4875) );
  XOR U4853 ( .A(n4839), .B(n4874), .Z(n4877) );
  AND U4854 ( .A(n4878), .B(n4879), .Z(n4839) );
  XNOR U4855 ( .A(n4836), .B(n4874), .Z(n4876) );
  XNOR U4856 ( .A(n4880), .B(n4881), .Z(n4836) );
  AND U4857 ( .A(n208), .B(n4882), .Z(n4881) );
  XNOR U4858 ( .A(n4883), .B(n4884), .Z(n4882) );
  XOR U4859 ( .A(n4885), .B(n4886), .Z(n4874) );
  AND U4860 ( .A(n4887), .B(n4888), .Z(n4886) );
  XNOR U4861 ( .A(n4885), .B(n4878), .Z(n4888) );
  IV U4862 ( .A(n4849), .Z(n4878) );
  XOR U4863 ( .A(n4889), .B(n4890), .Z(n4849) );
  XOR U4864 ( .A(n4891), .B(n4879), .Z(n4890) );
  AND U4865 ( .A(n4859), .B(n4892), .Z(n4879) );
  AND U4866 ( .A(n4893), .B(n4894), .Z(n4891) );
  XOR U4867 ( .A(n4895), .B(n4889), .Z(n4893) );
  XNOR U4868 ( .A(n4846), .B(n4885), .Z(n4887) );
  XNOR U4869 ( .A(n4896), .B(n4897), .Z(n4846) );
  AND U4870 ( .A(n208), .B(n4898), .Z(n4897) );
  XNOR U4871 ( .A(n4899), .B(n4900), .Z(n4898) );
  XOR U4872 ( .A(n4901), .B(n4902), .Z(n4885) );
  AND U4873 ( .A(n4903), .B(n4904), .Z(n4902) );
  XNOR U4874 ( .A(n4901), .B(n4859), .Z(n4904) );
  XOR U4875 ( .A(n4905), .B(n4894), .Z(n4859) );
  XNOR U4876 ( .A(n4906), .B(n4889), .Z(n4894) );
  XOR U4877 ( .A(n4907), .B(n4908), .Z(n4889) );
  AND U4878 ( .A(n4909), .B(n4910), .Z(n4908) );
  XOR U4879 ( .A(n4911), .B(n4907), .Z(n4909) );
  XNOR U4880 ( .A(n4912), .B(n4913), .Z(n4906) );
  AND U4881 ( .A(n4914), .B(n4915), .Z(n4913) );
  XOR U4882 ( .A(n4912), .B(n4916), .Z(n4914) );
  XNOR U4883 ( .A(n4895), .B(n4892), .Z(n4905) );
  AND U4884 ( .A(n4917), .B(n4918), .Z(n4892) );
  XOR U4885 ( .A(n4919), .B(n4920), .Z(n4895) );
  AND U4886 ( .A(n4921), .B(n4922), .Z(n4920) );
  XOR U4887 ( .A(n4919), .B(n4923), .Z(n4921) );
  XNOR U4888 ( .A(n4856), .B(n4901), .Z(n4903) );
  XNOR U4889 ( .A(n4924), .B(n4925), .Z(n4856) );
  AND U4890 ( .A(n208), .B(n4926), .Z(n4925) );
  XNOR U4891 ( .A(n4927), .B(n4928), .Z(n4926) );
  XOR U4892 ( .A(n4929), .B(n4930), .Z(n4901) );
  AND U4893 ( .A(n4931), .B(n4932), .Z(n4930) );
  XNOR U4894 ( .A(n4929), .B(n4917), .Z(n4932) );
  IV U4895 ( .A(n4867), .Z(n4917) );
  XNOR U4896 ( .A(n4933), .B(n4910), .Z(n4867) );
  XNOR U4897 ( .A(n4934), .B(n4916), .Z(n4910) );
  XNOR U4898 ( .A(n4935), .B(n4936), .Z(n4916) );
  NOR U4899 ( .A(n4937), .B(n4938), .Z(n4936) );
  XOR U4900 ( .A(n4935), .B(n4939), .Z(n4937) );
  XNOR U4901 ( .A(n4915), .B(n4907), .Z(n4934) );
  XOR U4902 ( .A(n4940), .B(n4941), .Z(n4907) );
  AND U4903 ( .A(n4942), .B(n4943), .Z(n4941) );
  XOR U4904 ( .A(n4940), .B(n4944), .Z(n4942) );
  XNOR U4905 ( .A(n4945), .B(n4912), .Z(n4915) );
  XOR U4906 ( .A(n4946), .B(n4947), .Z(n4912) );
  AND U4907 ( .A(n4948), .B(n4949), .Z(n4947) );
  XNOR U4908 ( .A(n4950), .B(n4951), .Z(n4948) );
  IV U4909 ( .A(n4946), .Z(n4950) );
  XNOR U4910 ( .A(n4952), .B(n4953), .Z(n4945) );
  NOR U4911 ( .A(n4954), .B(n4955), .Z(n4953) );
  XNOR U4912 ( .A(n4952), .B(n4956), .Z(n4954) );
  XNOR U4913 ( .A(n4911), .B(n4918), .Z(n4933) );
  NOR U4914 ( .A(n4873), .B(n4957), .Z(n4918) );
  XOR U4915 ( .A(n4923), .B(n4922), .Z(n4911) );
  XNOR U4916 ( .A(n4958), .B(n4919), .Z(n4922) );
  XOR U4917 ( .A(n4959), .B(n4960), .Z(n4919) );
  AND U4918 ( .A(n4961), .B(n4962), .Z(n4960) );
  XNOR U4919 ( .A(n4963), .B(n4964), .Z(n4961) );
  IV U4920 ( .A(n4959), .Z(n4963) );
  XNOR U4921 ( .A(n4965), .B(n4966), .Z(n4958) );
  NOR U4922 ( .A(n4967), .B(n4968), .Z(n4966) );
  XNOR U4923 ( .A(n4965), .B(n4969), .Z(n4967) );
  XOR U4924 ( .A(n4970), .B(n4971), .Z(n4923) );
  NOR U4925 ( .A(n4972), .B(n4973), .Z(n4971) );
  XNOR U4926 ( .A(n4970), .B(n4974), .Z(n4972) );
  XNOR U4927 ( .A(n4864), .B(n4929), .Z(n4931) );
  XNOR U4928 ( .A(n4975), .B(n4976), .Z(n4864) );
  AND U4929 ( .A(n208), .B(n4977), .Z(n4976) );
  XNOR U4930 ( .A(n4978), .B(n4979), .Z(n4977) );
  AND U4931 ( .A(n4870), .B(n4873), .Z(n4929) );
  XOR U4932 ( .A(n4980), .B(n4957), .Z(n4873) );
  XNOR U4933 ( .A(p_input[112]), .B(p_input[256]), .Z(n4957) );
  XNOR U4934 ( .A(n4944), .B(n4943), .Z(n4980) );
  XNOR U4935 ( .A(n4981), .B(n4951), .Z(n4943) );
  XNOR U4936 ( .A(n4939), .B(n4938), .Z(n4951) );
  XNOR U4937 ( .A(n4982), .B(n4935), .Z(n4938) );
  XNOR U4938 ( .A(p_input[122]), .B(p_input[266]), .Z(n4935) );
  XOR U4939 ( .A(p_input[123]), .B(n3382), .Z(n4982) );
  XOR U4940 ( .A(p_input[124]), .B(p_input[268]), .Z(n4939) );
  XOR U4941 ( .A(n4949), .B(n4983), .Z(n4981) );
  IV U4942 ( .A(n4940), .Z(n4983) );
  XOR U4943 ( .A(p_input[113]), .B(p_input[257]), .Z(n4940) );
  XNOR U4944 ( .A(n4984), .B(n4956), .Z(n4949) );
  XNOR U4945 ( .A(p_input[127]), .B(n3385), .Z(n4956) );
  XOR U4946 ( .A(n4946), .B(n4955), .Z(n4984) );
  XOR U4947 ( .A(n4985), .B(n4952), .Z(n4955) );
  XOR U4948 ( .A(p_input[125]), .B(p_input[269]), .Z(n4952) );
  XOR U4949 ( .A(p_input[126]), .B(n3387), .Z(n4985) );
  XOR U4950 ( .A(p_input[121]), .B(p_input[265]), .Z(n4946) );
  XOR U4951 ( .A(n4964), .B(n4962), .Z(n4944) );
  XNOR U4952 ( .A(n4986), .B(n4969), .Z(n4962) );
  XOR U4953 ( .A(p_input[120]), .B(p_input[264]), .Z(n4969) );
  XOR U4954 ( .A(n4959), .B(n4968), .Z(n4986) );
  XOR U4955 ( .A(n4987), .B(n4965), .Z(n4968) );
  XOR U4956 ( .A(p_input[118]), .B(p_input[262]), .Z(n4965) );
  XOR U4957 ( .A(p_input[119]), .B(n3625), .Z(n4987) );
  XOR U4958 ( .A(p_input[114]), .B(p_input[258]), .Z(n4959) );
  XNOR U4959 ( .A(n4974), .B(n4973), .Z(n4964) );
  XOR U4960 ( .A(n4988), .B(n4970), .Z(n4973) );
  XOR U4961 ( .A(p_input[115]), .B(p_input[259]), .Z(n4970) );
  XOR U4962 ( .A(p_input[116]), .B(n3627), .Z(n4988) );
  XOR U4963 ( .A(p_input[117]), .B(p_input[261]), .Z(n4974) );
  XNOR U4964 ( .A(n4989), .B(n4990), .Z(n4870) );
  AND U4965 ( .A(n208), .B(n4991), .Z(n4990) );
  XNOR U4966 ( .A(n4992), .B(n4993), .Z(n208) );
  AND U4967 ( .A(n4994), .B(n4995), .Z(n4993) );
  XOR U4968 ( .A(n4884), .B(n4992), .Z(n4995) );
  XNOR U4969 ( .A(n4996), .B(n4992), .Z(n4994) );
  XOR U4970 ( .A(n4997), .B(n4998), .Z(n4992) );
  AND U4971 ( .A(n4999), .B(n5000), .Z(n4998) );
  XOR U4972 ( .A(n4899), .B(n4997), .Z(n5000) );
  XOR U4973 ( .A(n4997), .B(n4900), .Z(n4999) );
  XOR U4974 ( .A(n5001), .B(n5002), .Z(n4997) );
  AND U4975 ( .A(n5003), .B(n5004), .Z(n5002) );
  XOR U4976 ( .A(n4927), .B(n5001), .Z(n5004) );
  XOR U4977 ( .A(n5001), .B(n4928), .Z(n5003) );
  XOR U4978 ( .A(n5005), .B(n5006), .Z(n5001) );
  AND U4979 ( .A(n5007), .B(n5008), .Z(n5006) );
  XOR U4980 ( .A(n5005), .B(n4978), .Z(n5008) );
  XNOR U4981 ( .A(n5009), .B(n5010), .Z(n4830) );
  AND U4982 ( .A(n212), .B(n5011), .Z(n5010) );
  XNOR U4983 ( .A(n5012), .B(n5013), .Z(n212) );
  AND U4984 ( .A(n5014), .B(n5015), .Z(n5013) );
  XOR U4985 ( .A(n5012), .B(n4840), .Z(n5015) );
  XNOR U4986 ( .A(n5012), .B(n4800), .Z(n5014) );
  XOR U4987 ( .A(n5016), .B(n5017), .Z(n5012) );
  AND U4988 ( .A(n5018), .B(n5019), .Z(n5017) );
  XOR U4989 ( .A(n5016), .B(n4808), .Z(n5018) );
  XOR U4990 ( .A(n5020), .B(n5021), .Z(n4791) );
  AND U4991 ( .A(n216), .B(n5011), .Z(n5021) );
  XNOR U4992 ( .A(n5009), .B(n5020), .Z(n5011) );
  XNOR U4993 ( .A(n5022), .B(n5023), .Z(n216) );
  AND U4994 ( .A(n5024), .B(n5025), .Z(n5023) );
  XNOR U4995 ( .A(n5026), .B(n5022), .Z(n5025) );
  IV U4996 ( .A(n4840), .Z(n5026) );
  XOR U4997 ( .A(n4996), .B(n5027), .Z(n4840) );
  AND U4998 ( .A(n219), .B(n5028), .Z(n5027) );
  XOR U4999 ( .A(n4883), .B(n4880), .Z(n5028) );
  XNOR U5000 ( .A(n4800), .B(n5022), .Z(n5024) );
  XNOR U5001 ( .A(n5029), .B(n5030), .Z(n4800) );
  AND U5002 ( .A(n235), .B(n5031), .Z(n5030) );
  XNOR U5003 ( .A(n5032), .B(n5033), .Z(n5031) );
  XOR U5004 ( .A(n5016), .B(n5034), .Z(n5022) );
  AND U5005 ( .A(n5035), .B(n5019), .Z(n5034) );
  XNOR U5006 ( .A(n4850), .B(n5016), .Z(n5019) );
  XOR U5007 ( .A(n4900), .B(n5036), .Z(n4850) );
  AND U5008 ( .A(n219), .B(n5037), .Z(n5036) );
  XOR U5009 ( .A(n4896), .B(n4900), .Z(n5037) );
  XNOR U5010 ( .A(n5038), .B(n5016), .Z(n5035) );
  IV U5011 ( .A(n4808), .Z(n5038) );
  XOR U5012 ( .A(n5039), .B(n5040), .Z(n4808) );
  AND U5013 ( .A(n235), .B(n5041), .Z(n5040) );
  XOR U5014 ( .A(n5042), .B(n5043), .Z(n5016) );
  AND U5015 ( .A(n5044), .B(n5045), .Z(n5043) );
  XNOR U5016 ( .A(n4860), .B(n5042), .Z(n5045) );
  XOR U5017 ( .A(n4928), .B(n5046), .Z(n4860) );
  AND U5018 ( .A(n219), .B(n5047), .Z(n5046) );
  XOR U5019 ( .A(n4924), .B(n4928), .Z(n5047) );
  XOR U5020 ( .A(n5042), .B(n4817), .Z(n5044) );
  XOR U5021 ( .A(n5048), .B(n5049), .Z(n4817) );
  AND U5022 ( .A(n235), .B(n5050), .Z(n5049) );
  XOR U5023 ( .A(n5051), .B(n5052), .Z(n5042) );
  AND U5024 ( .A(n5053), .B(n5054), .Z(n5052) );
  XNOR U5025 ( .A(n5051), .B(n4868), .Z(n5054) );
  XOR U5026 ( .A(n4979), .B(n5055), .Z(n4868) );
  AND U5027 ( .A(n219), .B(n5056), .Z(n5055) );
  XOR U5028 ( .A(n4975), .B(n4979), .Z(n5056) );
  XNOR U5029 ( .A(n5057), .B(n5051), .Z(n5053) );
  IV U5030 ( .A(n4827), .Z(n5057) );
  XOR U5031 ( .A(n5058), .B(n5059), .Z(n4827) );
  AND U5032 ( .A(n235), .B(n5060), .Z(n5059) );
  AND U5033 ( .A(n5020), .B(n5009), .Z(n5051) );
  XNOR U5034 ( .A(n5061), .B(n5062), .Z(n5009) );
  AND U5035 ( .A(n219), .B(n4991), .Z(n5062) );
  XNOR U5036 ( .A(n4989), .B(n5061), .Z(n4991) );
  XNOR U5037 ( .A(n5063), .B(n5064), .Z(n219) );
  AND U5038 ( .A(n5065), .B(n5066), .Z(n5064) );
  XNOR U5039 ( .A(n5063), .B(n4880), .Z(n5066) );
  IV U5040 ( .A(n4884), .Z(n4880) );
  XOR U5041 ( .A(n5067), .B(n5068), .Z(n4884) );
  AND U5042 ( .A(n223), .B(n5069), .Z(n5068) );
  XOR U5043 ( .A(n5070), .B(n5067), .Z(n5069) );
  XNOR U5044 ( .A(n5063), .B(n4996), .Z(n5065) );
  IV U5045 ( .A(n4883), .Z(n4996) );
  XOR U5046 ( .A(n5032), .B(n5071), .Z(n4883) );
  AND U5047 ( .A(n231), .B(n5072), .Z(n5071) );
  XOR U5048 ( .A(n5032), .B(n5029), .Z(n5072) );
  XOR U5049 ( .A(n5073), .B(n5074), .Z(n5063) );
  AND U5050 ( .A(n5075), .B(n5076), .Z(n5074) );
  XNOR U5051 ( .A(n5073), .B(n4896), .Z(n5076) );
  IV U5052 ( .A(n4899), .Z(n4896) );
  XOR U5053 ( .A(n5077), .B(n5078), .Z(n4899) );
  AND U5054 ( .A(n223), .B(n5079), .Z(n5078) );
  XOR U5055 ( .A(n5080), .B(n5077), .Z(n5079) );
  XOR U5056 ( .A(n4900), .B(n5073), .Z(n5075) );
  XOR U5057 ( .A(n5081), .B(n5082), .Z(n4900) );
  AND U5058 ( .A(n231), .B(n5041), .Z(n5082) );
  XOR U5059 ( .A(n5081), .B(n5039), .Z(n5041) );
  XOR U5060 ( .A(n5083), .B(n5084), .Z(n5073) );
  AND U5061 ( .A(n5085), .B(n5086), .Z(n5084) );
  XNOR U5062 ( .A(n5083), .B(n4924), .Z(n5086) );
  IV U5063 ( .A(n4927), .Z(n4924) );
  XOR U5064 ( .A(n5087), .B(n5088), .Z(n4927) );
  AND U5065 ( .A(n223), .B(n5089), .Z(n5088) );
  XNOR U5066 ( .A(n5090), .B(n5087), .Z(n5089) );
  XOR U5067 ( .A(n4928), .B(n5083), .Z(n5085) );
  XOR U5068 ( .A(n5091), .B(n5092), .Z(n4928) );
  AND U5069 ( .A(n231), .B(n5050), .Z(n5092) );
  XOR U5070 ( .A(n5091), .B(n5048), .Z(n5050) );
  XOR U5071 ( .A(n5005), .B(n5093), .Z(n5083) );
  AND U5072 ( .A(n5007), .B(n5094), .Z(n5093) );
  XNOR U5073 ( .A(n5005), .B(n4975), .Z(n5094) );
  IV U5074 ( .A(n4978), .Z(n4975) );
  XOR U5075 ( .A(n5095), .B(n5096), .Z(n4978) );
  AND U5076 ( .A(n223), .B(n5097), .Z(n5096) );
  XOR U5077 ( .A(n5098), .B(n5095), .Z(n5097) );
  XOR U5078 ( .A(n4979), .B(n5005), .Z(n5007) );
  XOR U5079 ( .A(n5099), .B(n5100), .Z(n4979) );
  AND U5080 ( .A(n231), .B(n5060), .Z(n5100) );
  XOR U5081 ( .A(n5099), .B(n5058), .Z(n5060) );
  AND U5082 ( .A(n5061), .B(n4989), .Z(n5005) );
  XNOR U5083 ( .A(n5101), .B(n5102), .Z(n4989) );
  AND U5084 ( .A(n223), .B(n5103), .Z(n5102) );
  XNOR U5085 ( .A(n5104), .B(n5101), .Z(n5103) );
  XNOR U5086 ( .A(n5105), .B(n5106), .Z(n223) );
  AND U5087 ( .A(n5107), .B(n5108), .Z(n5106) );
  XOR U5088 ( .A(n5070), .B(n5105), .Z(n5108) );
  AND U5089 ( .A(n5109), .B(n5110), .Z(n5070) );
  XNOR U5090 ( .A(n5067), .B(n5105), .Z(n5107) );
  XNOR U5091 ( .A(n5111), .B(n5112), .Z(n5067) );
  AND U5092 ( .A(n5113), .B(n227), .Z(n5112) );
  AND U5093 ( .A(n5111), .B(n5114), .Z(n5113) );
  XOR U5094 ( .A(n5115), .B(n5116), .Z(n5105) );
  AND U5095 ( .A(n5117), .B(n5118), .Z(n5116) );
  XNOR U5096 ( .A(n5115), .B(n5109), .Z(n5118) );
  IV U5097 ( .A(n5080), .Z(n5109) );
  XOR U5098 ( .A(n5119), .B(n5120), .Z(n5080) );
  XOR U5099 ( .A(n5121), .B(n5110), .Z(n5120) );
  AND U5100 ( .A(n5090), .B(n5122), .Z(n5110) );
  AND U5101 ( .A(n5123), .B(n5124), .Z(n5121) );
  XOR U5102 ( .A(n5125), .B(n5119), .Z(n5123) );
  XNOR U5103 ( .A(n5077), .B(n5115), .Z(n5117) );
  XNOR U5104 ( .A(n5126), .B(n5127), .Z(n5077) );
  AND U5105 ( .A(n227), .B(n5128), .Z(n5127) );
  XNOR U5106 ( .A(n5129), .B(n5130), .Z(n5128) );
  XOR U5107 ( .A(n5131), .B(n5132), .Z(n5115) );
  AND U5108 ( .A(n5133), .B(n5134), .Z(n5132) );
  XNOR U5109 ( .A(n5131), .B(n5090), .Z(n5134) );
  XOR U5110 ( .A(n5135), .B(n5124), .Z(n5090) );
  XNOR U5111 ( .A(n5136), .B(n5119), .Z(n5124) );
  XOR U5112 ( .A(n5137), .B(n5138), .Z(n5119) );
  AND U5113 ( .A(n5139), .B(n5140), .Z(n5138) );
  XOR U5114 ( .A(n5141), .B(n5137), .Z(n5139) );
  XNOR U5115 ( .A(n5142), .B(n5143), .Z(n5136) );
  AND U5116 ( .A(n5144), .B(n5145), .Z(n5143) );
  XOR U5117 ( .A(n5142), .B(n5146), .Z(n5144) );
  XNOR U5118 ( .A(n5125), .B(n5122), .Z(n5135) );
  AND U5119 ( .A(n5147), .B(n5148), .Z(n5122) );
  XOR U5120 ( .A(n5149), .B(n5150), .Z(n5125) );
  AND U5121 ( .A(n5151), .B(n5152), .Z(n5150) );
  XOR U5122 ( .A(n5149), .B(n5153), .Z(n5151) );
  XNOR U5123 ( .A(n5087), .B(n5131), .Z(n5133) );
  XNOR U5124 ( .A(n5154), .B(n5155), .Z(n5087) );
  AND U5125 ( .A(n227), .B(n5156), .Z(n5155) );
  XNOR U5126 ( .A(n5157), .B(n5158), .Z(n5156) );
  XOR U5127 ( .A(n5159), .B(n5160), .Z(n5131) );
  AND U5128 ( .A(n5161), .B(n5162), .Z(n5160) );
  XNOR U5129 ( .A(n5159), .B(n5147), .Z(n5162) );
  IV U5130 ( .A(n5098), .Z(n5147) );
  XNOR U5131 ( .A(n5163), .B(n5140), .Z(n5098) );
  XNOR U5132 ( .A(n5164), .B(n5146), .Z(n5140) );
  XNOR U5133 ( .A(n5165), .B(n5166), .Z(n5146) );
  NOR U5134 ( .A(n5167), .B(n5168), .Z(n5166) );
  XOR U5135 ( .A(n5165), .B(n5169), .Z(n5167) );
  XNOR U5136 ( .A(n5145), .B(n5137), .Z(n5164) );
  XOR U5137 ( .A(n5170), .B(n5171), .Z(n5137) );
  AND U5138 ( .A(n5172), .B(n5173), .Z(n5171) );
  XOR U5139 ( .A(n5170), .B(n5174), .Z(n5172) );
  XNOR U5140 ( .A(n5175), .B(n5142), .Z(n5145) );
  XOR U5141 ( .A(n5176), .B(n5177), .Z(n5142) );
  AND U5142 ( .A(n5178), .B(n5179), .Z(n5177) );
  XNOR U5143 ( .A(n5180), .B(n5181), .Z(n5178) );
  IV U5144 ( .A(n5176), .Z(n5180) );
  XNOR U5145 ( .A(n5182), .B(n5183), .Z(n5175) );
  NOR U5146 ( .A(n5184), .B(n5185), .Z(n5183) );
  XNOR U5147 ( .A(n5182), .B(n5186), .Z(n5184) );
  XNOR U5148 ( .A(n5141), .B(n5148), .Z(n5163) );
  NOR U5149 ( .A(n5104), .B(n5187), .Z(n5148) );
  XOR U5150 ( .A(n5153), .B(n5152), .Z(n5141) );
  XNOR U5151 ( .A(n5188), .B(n5149), .Z(n5152) );
  XOR U5152 ( .A(n5189), .B(n5190), .Z(n5149) );
  AND U5153 ( .A(n5191), .B(n5192), .Z(n5190) );
  XNOR U5154 ( .A(n5193), .B(n5194), .Z(n5191) );
  IV U5155 ( .A(n5189), .Z(n5193) );
  XNOR U5156 ( .A(n5195), .B(n5196), .Z(n5188) );
  NOR U5157 ( .A(n5197), .B(n5198), .Z(n5196) );
  XNOR U5158 ( .A(n5195), .B(n5199), .Z(n5197) );
  XOR U5159 ( .A(n5200), .B(n5201), .Z(n5153) );
  NOR U5160 ( .A(n5202), .B(n5203), .Z(n5201) );
  XNOR U5161 ( .A(n5200), .B(n5204), .Z(n5202) );
  XNOR U5162 ( .A(n5095), .B(n5159), .Z(n5161) );
  XNOR U5163 ( .A(n5205), .B(n5206), .Z(n5095) );
  AND U5164 ( .A(n227), .B(n5207), .Z(n5206) );
  XNOR U5165 ( .A(n5208), .B(n5209), .Z(n5207) );
  AND U5166 ( .A(n5101), .B(n5104), .Z(n5159) );
  XOR U5167 ( .A(n5210), .B(n5187), .Z(n5104) );
  XNOR U5168 ( .A(p_input[128]), .B(p_input[256]), .Z(n5187) );
  XNOR U5169 ( .A(n5174), .B(n5173), .Z(n5210) );
  XNOR U5170 ( .A(n5211), .B(n5181), .Z(n5173) );
  XNOR U5171 ( .A(n5169), .B(n5168), .Z(n5181) );
  XNOR U5172 ( .A(n5212), .B(n5165), .Z(n5168) );
  XNOR U5173 ( .A(p_input[138]), .B(p_input[266]), .Z(n5165) );
  XOR U5174 ( .A(p_input[139]), .B(n3382), .Z(n5212) );
  XOR U5175 ( .A(p_input[140]), .B(p_input[268]), .Z(n5169) );
  XOR U5176 ( .A(n5179), .B(n5213), .Z(n5211) );
  IV U5177 ( .A(n5170), .Z(n5213) );
  XOR U5178 ( .A(p_input[129]), .B(p_input[257]), .Z(n5170) );
  XNOR U5179 ( .A(n5214), .B(n5186), .Z(n5179) );
  XNOR U5180 ( .A(p_input[143]), .B(n3385), .Z(n5186) );
  XOR U5181 ( .A(n5176), .B(n5185), .Z(n5214) );
  XOR U5182 ( .A(n5215), .B(n5182), .Z(n5185) );
  XOR U5183 ( .A(p_input[141]), .B(p_input[269]), .Z(n5182) );
  XOR U5184 ( .A(p_input[142]), .B(n3387), .Z(n5215) );
  XOR U5185 ( .A(p_input[137]), .B(p_input[265]), .Z(n5176) );
  XOR U5186 ( .A(n5194), .B(n5192), .Z(n5174) );
  XNOR U5187 ( .A(n5216), .B(n5199), .Z(n5192) );
  XOR U5188 ( .A(p_input[136]), .B(p_input[264]), .Z(n5199) );
  XOR U5189 ( .A(n5189), .B(n5198), .Z(n5216) );
  XOR U5190 ( .A(n5217), .B(n5195), .Z(n5198) );
  XOR U5191 ( .A(p_input[134]), .B(p_input[262]), .Z(n5195) );
  XOR U5192 ( .A(p_input[135]), .B(n3625), .Z(n5217) );
  XOR U5193 ( .A(p_input[130]), .B(p_input[258]), .Z(n5189) );
  XNOR U5194 ( .A(n5204), .B(n5203), .Z(n5194) );
  XOR U5195 ( .A(n5218), .B(n5200), .Z(n5203) );
  XOR U5196 ( .A(p_input[131]), .B(p_input[259]), .Z(n5200) );
  XOR U5197 ( .A(p_input[132]), .B(n3627), .Z(n5218) );
  XOR U5198 ( .A(p_input[133]), .B(p_input[261]), .Z(n5204) );
  XNOR U5199 ( .A(n5219), .B(n5220), .Z(n5101) );
  AND U5200 ( .A(n227), .B(n5221), .Z(n5220) );
  XNOR U5201 ( .A(n5222), .B(n5223), .Z(n227) );
  AND U5202 ( .A(n5224), .B(n5225), .Z(n5223) );
  XNOR U5203 ( .A(n5111), .B(n5222), .Z(n5225) );
  XNOR U5204 ( .A(n5114), .B(n5222), .Z(n5224) );
  XOR U5205 ( .A(n5226), .B(n5227), .Z(n5222) );
  AND U5206 ( .A(n5228), .B(n5229), .Z(n5227) );
  XOR U5207 ( .A(n5129), .B(n5226), .Z(n5229) );
  XOR U5208 ( .A(n5226), .B(n5130), .Z(n5228) );
  XOR U5209 ( .A(n5230), .B(n5231), .Z(n5226) );
  AND U5210 ( .A(n5232), .B(n5233), .Z(n5231) );
  XOR U5211 ( .A(n5157), .B(n5230), .Z(n5233) );
  XOR U5212 ( .A(n5230), .B(n5158), .Z(n5232) );
  XOR U5213 ( .A(n5234), .B(n5235), .Z(n5230) );
  AND U5214 ( .A(n5236), .B(n5237), .Z(n5235) );
  XOR U5215 ( .A(n5234), .B(n5208), .Z(n5237) );
  XNOR U5216 ( .A(n5238), .B(n5239), .Z(n5061) );
  AND U5217 ( .A(n231), .B(n5240), .Z(n5239) );
  XNOR U5218 ( .A(n5241), .B(n5242), .Z(n231) );
  AND U5219 ( .A(n5243), .B(n5244), .Z(n5242) );
  XNOR U5220 ( .A(n5241), .B(n5032), .Z(n5244) );
  XOR U5221 ( .A(n5241), .B(n5029), .Z(n5243) );
  XOR U5222 ( .A(n5245), .B(n5246), .Z(n5241) );
  AND U5223 ( .A(n5247), .B(n5248), .Z(n5246) );
  XOR U5224 ( .A(n5245), .B(n5039), .Z(n5247) );
  XOR U5225 ( .A(n5249), .B(n5250), .Z(n5020) );
  AND U5226 ( .A(n235), .B(n5240), .Z(n5250) );
  XNOR U5227 ( .A(n5238), .B(n5249), .Z(n5240) );
  XNOR U5228 ( .A(n5251), .B(n5252), .Z(n235) );
  AND U5229 ( .A(n5253), .B(n5254), .Z(n5252) );
  XNOR U5230 ( .A(n5032), .B(n5251), .Z(n5254) );
  XNOR U5231 ( .A(n5114), .B(n5255), .Z(n5032) );
  AND U5232 ( .A(n5256), .B(n238), .Z(n5255) );
  NOR U5233 ( .A(n5257), .B(n5258), .Z(n5256) );
  XOR U5234 ( .A(n5251), .B(n5029), .Z(n5253) );
  IV U5235 ( .A(n5033), .Z(n5029) );
  AND U5236 ( .A(n5259), .B(n5260), .Z(n5033) );
  XOR U5237 ( .A(n5245), .B(n5261), .Z(n5251) );
  AND U5238 ( .A(n5262), .B(n5248), .Z(n5261) );
  XNOR U5239 ( .A(n5081), .B(n5245), .Z(n5248) );
  XOR U5240 ( .A(n5130), .B(n5263), .Z(n5081) );
  AND U5241 ( .A(n238), .B(n5264), .Z(n5263) );
  XOR U5242 ( .A(n5126), .B(n5130), .Z(n5264) );
  XNOR U5243 ( .A(n5265), .B(n5245), .Z(n5262) );
  IV U5244 ( .A(n5039), .Z(n5265) );
  XOR U5245 ( .A(n5266), .B(n5267), .Z(n5039) );
  AND U5246 ( .A(n254), .B(n5268), .Z(n5267) );
  XOR U5247 ( .A(n5269), .B(n5270), .Z(n5245) );
  AND U5248 ( .A(n5271), .B(n5272), .Z(n5270) );
  XNOR U5249 ( .A(n5091), .B(n5269), .Z(n5272) );
  XOR U5250 ( .A(n5158), .B(n5273), .Z(n5091) );
  AND U5251 ( .A(n238), .B(n5274), .Z(n5273) );
  XOR U5252 ( .A(n5154), .B(n5158), .Z(n5274) );
  XOR U5253 ( .A(n5269), .B(n5048), .Z(n5271) );
  XOR U5254 ( .A(n5275), .B(n5276), .Z(n5048) );
  AND U5255 ( .A(n254), .B(n5277), .Z(n5276) );
  XOR U5256 ( .A(n5278), .B(n5279), .Z(n5269) );
  AND U5257 ( .A(n5280), .B(n5281), .Z(n5279) );
  XNOR U5258 ( .A(n5278), .B(n5099), .Z(n5281) );
  XOR U5259 ( .A(n5209), .B(n5282), .Z(n5099) );
  AND U5260 ( .A(n238), .B(n5283), .Z(n5282) );
  XOR U5261 ( .A(n5205), .B(n5209), .Z(n5283) );
  XNOR U5262 ( .A(n5284), .B(n5278), .Z(n5280) );
  IV U5263 ( .A(n5058), .Z(n5284) );
  XOR U5264 ( .A(n5285), .B(n5286), .Z(n5058) );
  AND U5265 ( .A(n254), .B(n5287), .Z(n5286) );
  AND U5266 ( .A(n5249), .B(n5238), .Z(n5278) );
  XNOR U5267 ( .A(n5288), .B(n5289), .Z(n5238) );
  AND U5268 ( .A(n238), .B(n5221), .Z(n5289) );
  XNOR U5269 ( .A(n5219), .B(n5288), .Z(n5221) );
  XNOR U5270 ( .A(n5290), .B(n5291), .Z(n238) );
  AND U5271 ( .A(n5292), .B(n5293), .Z(n5291) );
  XNOR U5272 ( .A(n5111), .B(n5290), .Z(n5293) );
  IV U5273 ( .A(n5257), .Z(n5111) );
  AND U5274 ( .A(n5294), .B(n5295), .Z(n5257) );
  IV U5275 ( .A(n5296), .Z(n5294) );
  XNOR U5276 ( .A(n5114), .B(n5290), .Z(n5292) );
  IV U5277 ( .A(n5258), .Z(n5114) );
  NOR U5278 ( .A(n5259), .B(n5260), .Z(n5258) );
  XOR U5279 ( .A(n5297), .B(n5298), .Z(n5290) );
  AND U5280 ( .A(n5299), .B(n5300), .Z(n5298) );
  XNOR U5281 ( .A(n5297), .B(n5126), .Z(n5300) );
  IV U5282 ( .A(n5129), .Z(n5126) );
  XOR U5283 ( .A(n5301), .B(n5302), .Z(n5129) );
  AND U5284 ( .A(n242), .B(n5303), .Z(n5302) );
  XOR U5285 ( .A(n5304), .B(n5301), .Z(n5303) );
  XOR U5286 ( .A(n5130), .B(n5297), .Z(n5299) );
  XOR U5287 ( .A(n5305), .B(n5306), .Z(n5130) );
  AND U5288 ( .A(n250), .B(n5268), .Z(n5306) );
  XOR U5289 ( .A(n5305), .B(n5266), .Z(n5268) );
  XOR U5290 ( .A(n5307), .B(n5308), .Z(n5297) );
  AND U5291 ( .A(n5309), .B(n5310), .Z(n5308) );
  XNOR U5292 ( .A(n5307), .B(n5154), .Z(n5310) );
  IV U5293 ( .A(n5157), .Z(n5154) );
  XOR U5294 ( .A(n5311), .B(n5312), .Z(n5157) );
  AND U5295 ( .A(n242), .B(n5313), .Z(n5312) );
  XNOR U5296 ( .A(n5314), .B(n5311), .Z(n5313) );
  XOR U5297 ( .A(n5158), .B(n5307), .Z(n5309) );
  XOR U5298 ( .A(n5315), .B(n5316), .Z(n5158) );
  AND U5299 ( .A(n250), .B(n5277), .Z(n5316) );
  XOR U5300 ( .A(n5315), .B(n5275), .Z(n5277) );
  XOR U5301 ( .A(n5234), .B(n5317), .Z(n5307) );
  AND U5302 ( .A(n5236), .B(n5318), .Z(n5317) );
  XNOR U5303 ( .A(n5234), .B(n5205), .Z(n5318) );
  IV U5304 ( .A(n5208), .Z(n5205) );
  XOR U5305 ( .A(n5319), .B(n5320), .Z(n5208) );
  AND U5306 ( .A(n242), .B(n5321), .Z(n5320) );
  XOR U5307 ( .A(n5322), .B(n5319), .Z(n5321) );
  XOR U5308 ( .A(n5209), .B(n5234), .Z(n5236) );
  XOR U5309 ( .A(n5323), .B(n5324), .Z(n5209) );
  AND U5310 ( .A(n250), .B(n5287), .Z(n5324) );
  XOR U5311 ( .A(n5323), .B(n5285), .Z(n5287) );
  AND U5312 ( .A(n5288), .B(n5219), .Z(n5234) );
  XNOR U5313 ( .A(n5325), .B(n5326), .Z(n5219) );
  AND U5314 ( .A(n242), .B(n5327), .Z(n5326) );
  XNOR U5315 ( .A(n5328), .B(n5325), .Z(n5327) );
  XNOR U5316 ( .A(n5329), .B(n5330), .Z(n242) );
  NOR U5317 ( .A(n5331), .B(n5332), .Z(n5330) );
  XNOR U5318 ( .A(n5329), .B(n5296), .Z(n5332) );
  NOR U5319 ( .A(n5333), .B(n5334), .Z(n5296) );
  NOR U5320 ( .A(n5329), .B(n5295), .Z(n5331) );
  AND U5321 ( .A(n5335), .B(n5336), .Z(n5295) );
  XOR U5322 ( .A(n5337), .B(n5338), .Z(n5329) );
  AND U5323 ( .A(n5339), .B(n5340), .Z(n5338) );
  XNOR U5324 ( .A(n5337), .B(n5335), .Z(n5340) );
  IV U5325 ( .A(n5304), .Z(n5335) );
  XOR U5326 ( .A(n5341), .B(n5342), .Z(n5304) );
  XOR U5327 ( .A(n5343), .B(n5336), .Z(n5342) );
  AND U5328 ( .A(n5314), .B(n5344), .Z(n5336) );
  AND U5329 ( .A(n5345), .B(n5346), .Z(n5343) );
  XOR U5330 ( .A(n5347), .B(n5341), .Z(n5345) );
  XNOR U5331 ( .A(n5301), .B(n5337), .Z(n5339) );
  XNOR U5332 ( .A(n5348), .B(n5349), .Z(n5301) );
  AND U5333 ( .A(n246), .B(n5350), .Z(n5349) );
  XNOR U5334 ( .A(n5351), .B(n5352), .Z(n5350) );
  XOR U5335 ( .A(n5353), .B(n5354), .Z(n5337) );
  AND U5336 ( .A(n5355), .B(n5356), .Z(n5354) );
  XNOR U5337 ( .A(n5353), .B(n5314), .Z(n5356) );
  XOR U5338 ( .A(n5357), .B(n5346), .Z(n5314) );
  XNOR U5339 ( .A(n5358), .B(n5341), .Z(n5346) );
  XOR U5340 ( .A(n5359), .B(n5360), .Z(n5341) );
  AND U5341 ( .A(n5361), .B(n5362), .Z(n5360) );
  XOR U5342 ( .A(n5363), .B(n5359), .Z(n5361) );
  XNOR U5343 ( .A(n5364), .B(n5365), .Z(n5358) );
  AND U5344 ( .A(n5366), .B(n5367), .Z(n5365) );
  XOR U5345 ( .A(n5364), .B(n5368), .Z(n5366) );
  XNOR U5346 ( .A(n5347), .B(n5344), .Z(n5357) );
  AND U5347 ( .A(n5369), .B(n5370), .Z(n5344) );
  XOR U5348 ( .A(n5371), .B(n5372), .Z(n5347) );
  AND U5349 ( .A(n5373), .B(n5374), .Z(n5372) );
  XOR U5350 ( .A(n5371), .B(n5375), .Z(n5373) );
  XNOR U5351 ( .A(n5311), .B(n5353), .Z(n5355) );
  XNOR U5352 ( .A(n5376), .B(n5377), .Z(n5311) );
  AND U5353 ( .A(n246), .B(n5378), .Z(n5377) );
  XNOR U5354 ( .A(n5379), .B(n5380), .Z(n5378) );
  XOR U5355 ( .A(n5381), .B(n5382), .Z(n5353) );
  AND U5356 ( .A(n5383), .B(n5384), .Z(n5382) );
  XNOR U5357 ( .A(n5381), .B(n5369), .Z(n5384) );
  IV U5358 ( .A(n5322), .Z(n5369) );
  XNOR U5359 ( .A(n5385), .B(n5362), .Z(n5322) );
  XNOR U5360 ( .A(n5386), .B(n5368), .Z(n5362) );
  XNOR U5361 ( .A(n5387), .B(n5388), .Z(n5368) );
  NOR U5362 ( .A(n5389), .B(n5390), .Z(n5388) );
  XOR U5363 ( .A(n5387), .B(n5391), .Z(n5389) );
  XNOR U5364 ( .A(n5367), .B(n5359), .Z(n5386) );
  XOR U5365 ( .A(n5392), .B(n5393), .Z(n5359) );
  AND U5366 ( .A(n5394), .B(n5395), .Z(n5393) );
  XOR U5367 ( .A(n5392), .B(n5396), .Z(n5394) );
  XNOR U5368 ( .A(n5397), .B(n5364), .Z(n5367) );
  XOR U5369 ( .A(n5398), .B(n5399), .Z(n5364) );
  AND U5370 ( .A(n5400), .B(n5401), .Z(n5399) );
  XNOR U5371 ( .A(n5402), .B(n5403), .Z(n5400) );
  IV U5372 ( .A(n5398), .Z(n5402) );
  XNOR U5373 ( .A(n5404), .B(n5405), .Z(n5397) );
  NOR U5374 ( .A(n5406), .B(n5407), .Z(n5405) );
  XNOR U5375 ( .A(n5404), .B(n5408), .Z(n5406) );
  XNOR U5376 ( .A(n5363), .B(n5370), .Z(n5385) );
  NOR U5377 ( .A(n5328), .B(n5409), .Z(n5370) );
  XOR U5378 ( .A(n5375), .B(n5374), .Z(n5363) );
  XNOR U5379 ( .A(n5410), .B(n5371), .Z(n5374) );
  XOR U5380 ( .A(n5411), .B(n5412), .Z(n5371) );
  AND U5381 ( .A(n5413), .B(n5414), .Z(n5412) );
  XNOR U5382 ( .A(n5415), .B(n5416), .Z(n5413) );
  IV U5383 ( .A(n5411), .Z(n5415) );
  XNOR U5384 ( .A(n5417), .B(n5418), .Z(n5410) );
  NOR U5385 ( .A(n5419), .B(n5420), .Z(n5418) );
  XNOR U5386 ( .A(n5417), .B(n5421), .Z(n5419) );
  XOR U5387 ( .A(n5422), .B(n5423), .Z(n5375) );
  NOR U5388 ( .A(n5424), .B(n5425), .Z(n5423) );
  XNOR U5389 ( .A(n5422), .B(n5426), .Z(n5424) );
  XNOR U5390 ( .A(n5319), .B(n5381), .Z(n5383) );
  XNOR U5391 ( .A(n5427), .B(n5428), .Z(n5319) );
  AND U5392 ( .A(n246), .B(n5429), .Z(n5428) );
  XNOR U5393 ( .A(n5430), .B(n5431), .Z(n5429) );
  AND U5394 ( .A(n5325), .B(n5328), .Z(n5381) );
  XOR U5395 ( .A(n5432), .B(n5409), .Z(n5328) );
  XNOR U5396 ( .A(p_input[144]), .B(p_input[256]), .Z(n5409) );
  XNOR U5397 ( .A(n5396), .B(n5395), .Z(n5432) );
  XNOR U5398 ( .A(n5433), .B(n5403), .Z(n5395) );
  XNOR U5399 ( .A(n5391), .B(n5390), .Z(n5403) );
  XNOR U5400 ( .A(n5434), .B(n5387), .Z(n5390) );
  XNOR U5401 ( .A(p_input[154]), .B(p_input[266]), .Z(n5387) );
  XOR U5402 ( .A(p_input[155]), .B(n3382), .Z(n5434) );
  XOR U5403 ( .A(p_input[156]), .B(p_input[268]), .Z(n5391) );
  XOR U5404 ( .A(n5401), .B(n5435), .Z(n5433) );
  IV U5405 ( .A(n5392), .Z(n5435) );
  XOR U5406 ( .A(p_input[145]), .B(p_input[257]), .Z(n5392) );
  XNOR U5407 ( .A(n5436), .B(n5408), .Z(n5401) );
  XNOR U5408 ( .A(p_input[159]), .B(n3385), .Z(n5408) );
  XOR U5409 ( .A(n5398), .B(n5407), .Z(n5436) );
  XOR U5410 ( .A(n5437), .B(n5404), .Z(n5407) );
  XOR U5411 ( .A(p_input[157]), .B(p_input[269]), .Z(n5404) );
  XOR U5412 ( .A(p_input[158]), .B(n3387), .Z(n5437) );
  XOR U5413 ( .A(p_input[153]), .B(p_input[265]), .Z(n5398) );
  XOR U5414 ( .A(n5416), .B(n5414), .Z(n5396) );
  XNOR U5415 ( .A(n5438), .B(n5421), .Z(n5414) );
  XOR U5416 ( .A(p_input[152]), .B(p_input[264]), .Z(n5421) );
  XOR U5417 ( .A(n5411), .B(n5420), .Z(n5438) );
  XOR U5418 ( .A(n5439), .B(n5417), .Z(n5420) );
  XOR U5419 ( .A(p_input[150]), .B(p_input[262]), .Z(n5417) );
  XOR U5420 ( .A(p_input[151]), .B(n3625), .Z(n5439) );
  XOR U5421 ( .A(p_input[146]), .B(p_input[258]), .Z(n5411) );
  XNOR U5422 ( .A(n5426), .B(n5425), .Z(n5416) );
  XOR U5423 ( .A(n5440), .B(n5422), .Z(n5425) );
  XOR U5424 ( .A(p_input[147]), .B(p_input[259]), .Z(n5422) );
  XOR U5425 ( .A(p_input[148]), .B(n3627), .Z(n5440) );
  XOR U5426 ( .A(p_input[149]), .B(p_input[261]), .Z(n5426) );
  XNOR U5427 ( .A(n5441), .B(n5442), .Z(n5325) );
  AND U5428 ( .A(n246), .B(n5443), .Z(n5442) );
  XNOR U5429 ( .A(n5444), .B(n5445), .Z(n246) );
  NOR U5430 ( .A(n5446), .B(n5447), .Z(n5445) );
  XNOR U5431 ( .A(n5444), .B(n5448), .Z(n5447) );
  NOR U5432 ( .A(n5444), .B(n5334), .Z(n5446) );
  XOR U5433 ( .A(n5449), .B(n5450), .Z(n5444) );
  AND U5434 ( .A(n5451), .B(n5452), .Z(n5450) );
  XOR U5435 ( .A(n5351), .B(n5449), .Z(n5452) );
  XOR U5436 ( .A(n5449), .B(n5352), .Z(n5451) );
  XOR U5437 ( .A(n5453), .B(n5454), .Z(n5449) );
  AND U5438 ( .A(n5455), .B(n5456), .Z(n5454) );
  XOR U5439 ( .A(n5379), .B(n5453), .Z(n5456) );
  XOR U5440 ( .A(n5453), .B(n5380), .Z(n5455) );
  XOR U5441 ( .A(n5457), .B(n5458), .Z(n5453) );
  AND U5442 ( .A(n5459), .B(n5460), .Z(n5458) );
  XOR U5443 ( .A(n5457), .B(n5430), .Z(n5460) );
  XNOR U5444 ( .A(n5461), .B(n5462), .Z(n5288) );
  AND U5445 ( .A(n250), .B(n5463), .Z(n5462) );
  XNOR U5446 ( .A(n5464), .B(n5465), .Z(n250) );
  NOR U5447 ( .A(n5466), .B(n5467), .Z(n5465) );
  XOR U5448 ( .A(n5260), .B(n5464), .Z(n5467) );
  NOR U5449 ( .A(n5464), .B(n5259), .Z(n5466) );
  XOR U5450 ( .A(n5468), .B(n5469), .Z(n5464) );
  AND U5451 ( .A(n5470), .B(n5471), .Z(n5469) );
  XOR U5452 ( .A(n5468), .B(n5266), .Z(n5470) );
  XOR U5453 ( .A(n5472), .B(n5473), .Z(n5249) );
  AND U5454 ( .A(n254), .B(n5463), .Z(n5473) );
  XNOR U5455 ( .A(n5461), .B(n5472), .Z(n5463) );
  XNOR U5456 ( .A(n5474), .B(n5475), .Z(n254) );
  NOR U5457 ( .A(n5476), .B(n5477), .Z(n5475) );
  XNOR U5458 ( .A(n5260), .B(n5478), .Z(n5477) );
  IV U5459 ( .A(n5474), .Z(n5478) );
  AND U5460 ( .A(n5479), .B(n5480), .Z(n5260) );
  NOR U5461 ( .A(n5474), .B(n5259), .Z(n5476) );
  AND U5462 ( .A(n5334), .B(n5333), .Z(n5259) );
  IV U5463 ( .A(n5448), .Z(n5333) );
  XOR U5464 ( .A(n5468), .B(n5481), .Z(n5474) );
  AND U5465 ( .A(n5482), .B(n5471), .Z(n5481) );
  XNOR U5466 ( .A(n5305), .B(n5468), .Z(n5471) );
  XOR U5467 ( .A(n5352), .B(n5483), .Z(n5305) );
  AND U5468 ( .A(n257), .B(n5484), .Z(n5483) );
  XOR U5469 ( .A(n5348), .B(n5352), .Z(n5484) );
  XNOR U5470 ( .A(n5485), .B(n5468), .Z(n5482) );
  IV U5471 ( .A(n5266), .Z(n5485) );
  XOR U5472 ( .A(n5486), .B(n5487), .Z(n5266) );
  AND U5473 ( .A(n273), .B(n5488), .Z(n5487) );
  XOR U5474 ( .A(n5489), .B(n5490), .Z(n5468) );
  AND U5475 ( .A(n5491), .B(n5492), .Z(n5490) );
  XNOR U5476 ( .A(n5315), .B(n5489), .Z(n5492) );
  XOR U5477 ( .A(n5380), .B(n5493), .Z(n5315) );
  AND U5478 ( .A(n257), .B(n5494), .Z(n5493) );
  XOR U5479 ( .A(n5376), .B(n5380), .Z(n5494) );
  XOR U5480 ( .A(n5489), .B(n5275), .Z(n5491) );
  XOR U5481 ( .A(n5495), .B(n5496), .Z(n5275) );
  AND U5482 ( .A(n273), .B(n5497), .Z(n5496) );
  XOR U5483 ( .A(n5498), .B(n5499), .Z(n5489) );
  AND U5484 ( .A(n5500), .B(n5501), .Z(n5499) );
  XNOR U5485 ( .A(n5498), .B(n5323), .Z(n5501) );
  XOR U5486 ( .A(n5431), .B(n5502), .Z(n5323) );
  AND U5487 ( .A(n257), .B(n5503), .Z(n5502) );
  XOR U5488 ( .A(n5427), .B(n5431), .Z(n5503) );
  XNOR U5489 ( .A(n5504), .B(n5498), .Z(n5500) );
  IV U5490 ( .A(n5285), .Z(n5504) );
  XOR U5491 ( .A(n5505), .B(n5506), .Z(n5285) );
  AND U5492 ( .A(n273), .B(n5507), .Z(n5506) );
  AND U5493 ( .A(n5472), .B(n5461), .Z(n5498) );
  XNOR U5494 ( .A(n5508), .B(n5509), .Z(n5461) );
  AND U5495 ( .A(n257), .B(n5443), .Z(n5509) );
  XNOR U5496 ( .A(n5441), .B(n5508), .Z(n5443) );
  XNOR U5497 ( .A(n5510), .B(n5511), .Z(n257) );
  NOR U5498 ( .A(n5512), .B(n5513), .Z(n5511) );
  XNOR U5499 ( .A(n5510), .B(n5448), .Z(n5513) );
  NOR U5500 ( .A(n5479), .B(n5480), .Z(n5448) );
  NOR U5501 ( .A(n5510), .B(n5334), .Z(n5512) );
  AND U5502 ( .A(n5514), .B(n5515), .Z(n5334) );
  IV U5503 ( .A(n5516), .Z(n5514) );
  XOR U5504 ( .A(n5517), .B(n5518), .Z(n5510) );
  AND U5505 ( .A(n5519), .B(n5520), .Z(n5518) );
  XNOR U5506 ( .A(n5517), .B(n5348), .Z(n5520) );
  IV U5507 ( .A(n5351), .Z(n5348) );
  XOR U5508 ( .A(n5521), .B(n5522), .Z(n5351) );
  AND U5509 ( .A(n261), .B(n5523), .Z(n5522) );
  XOR U5510 ( .A(n5524), .B(n5521), .Z(n5523) );
  XOR U5511 ( .A(n5352), .B(n5517), .Z(n5519) );
  XOR U5512 ( .A(n5525), .B(n5526), .Z(n5352) );
  AND U5513 ( .A(n269), .B(n5488), .Z(n5526) );
  XOR U5514 ( .A(n5525), .B(n5486), .Z(n5488) );
  XOR U5515 ( .A(n5527), .B(n5528), .Z(n5517) );
  AND U5516 ( .A(n5529), .B(n5530), .Z(n5528) );
  XNOR U5517 ( .A(n5527), .B(n5376), .Z(n5530) );
  IV U5518 ( .A(n5379), .Z(n5376) );
  XOR U5519 ( .A(n5531), .B(n5532), .Z(n5379) );
  AND U5520 ( .A(n261), .B(n5533), .Z(n5532) );
  XNOR U5521 ( .A(n5534), .B(n5531), .Z(n5533) );
  XOR U5522 ( .A(n5380), .B(n5527), .Z(n5529) );
  XOR U5523 ( .A(n5535), .B(n5536), .Z(n5380) );
  AND U5524 ( .A(n269), .B(n5497), .Z(n5536) );
  XOR U5525 ( .A(n5535), .B(n5495), .Z(n5497) );
  XOR U5526 ( .A(n5457), .B(n5537), .Z(n5527) );
  AND U5527 ( .A(n5459), .B(n5538), .Z(n5537) );
  XNOR U5528 ( .A(n5457), .B(n5427), .Z(n5538) );
  IV U5529 ( .A(n5430), .Z(n5427) );
  XOR U5530 ( .A(n5539), .B(n5540), .Z(n5430) );
  AND U5531 ( .A(n261), .B(n5541), .Z(n5540) );
  XOR U5532 ( .A(n5542), .B(n5539), .Z(n5541) );
  XOR U5533 ( .A(n5431), .B(n5457), .Z(n5459) );
  XOR U5534 ( .A(n5543), .B(n5544), .Z(n5431) );
  AND U5535 ( .A(n269), .B(n5507), .Z(n5544) );
  XOR U5536 ( .A(n5543), .B(n5505), .Z(n5507) );
  AND U5537 ( .A(n5508), .B(n5441), .Z(n5457) );
  XNOR U5538 ( .A(n5545), .B(n5546), .Z(n5441) );
  AND U5539 ( .A(n261), .B(n5547), .Z(n5546) );
  XNOR U5540 ( .A(n5548), .B(n5545), .Z(n5547) );
  XNOR U5541 ( .A(n5549), .B(n5550), .Z(n261) );
  NOR U5542 ( .A(n5551), .B(n5552), .Z(n5550) );
  XNOR U5543 ( .A(n5549), .B(n5516), .Z(n5552) );
  NOR U5544 ( .A(n5553), .B(n5554), .Z(n5516) );
  NOR U5545 ( .A(n5549), .B(n5515), .Z(n5551) );
  AND U5546 ( .A(n5555), .B(n5556), .Z(n5515) );
  XOR U5547 ( .A(n5557), .B(n5558), .Z(n5549) );
  AND U5548 ( .A(n5559), .B(n5560), .Z(n5558) );
  XNOR U5549 ( .A(n5557), .B(n5555), .Z(n5560) );
  IV U5550 ( .A(n5524), .Z(n5555) );
  XOR U5551 ( .A(n5561), .B(n5562), .Z(n5524) );
  XOR U5552 ( .A(n5563), .B(n5556), .Z(n5562) );
  AND U5553 ( .A(n5534), .B(n5564), .Z(n5556) );
  AND U5554 ( .A(n5565), .B(n5566), .Z(n5563) );
  XOR U5555 ( .A(n5567), .B(n5561), .Z(n5565) );
  XNOR U5556 ( .A(n5521), .B(n5557), .Z(n5559) );
  XNOR U5557 ( .A(n5568), .B(n5569), .Z(n5521) );
  AND U5558 ( .A(n265), .B(n5570), .Z(n5569) );
  XNOR U5559 ( .A(n5571), .B(n5572), .Z(n5570) );
  XOR U5560 ( .A(n5573), .B(n5574), .Z(n5557) );
  AND U5561 ( .A(n5575), .B(n5576), .Z(n5574) );
  XNOR U5562 ( .A(n5573), .B(n5534), .Z(n5576) );
  XOR U5563 ( .A(n5577), .B(n5566), .Z(n5534) );
  XNOR U5564 ( .A(n5578), .B(n5561), .Z(n5566) );
  XOR U5565 ( .A(n5579), .B(n5580), .Z(n5561) );
  AND U5566 ( .A(n5581), .B(n5582), .Z(n5580) );
  XOR U5567 ( .A(n5583), .B(n5579), .Z(n5581) );
  XNOR U5568 ( .A(n5584), .B(n5585), .Z(n5578) );
  AND U5569 ( .A(n5586), .B(n5587), .Z(n5585) );
  XOR U5570 ( .A(n5584), .B(n5588), .Z(n5586) );
  XNOR U5571 ( .A(n5567), .B(n5564), .Z(n5577) );
  AND U5572 ( .A(n5589), .B(n5590), .Z(n5564) );
  XOR U5573 ( .A(n5591), .B(n5592), .Z(n5567) );
  AND U5574 ( .A(n5593), .B(n5594), .Z(n5592) );
  XOR U5575 ( .A(n5591), .B(n5595), .Z(n5593) );
  XNOR U5576 ( .A(n5531), .B(n5573), .Z(n5575) );
  XNOR U5577 ( .A(n5596), .B(n5597), .Z(n5531) );
  AND U5578 ( .A(n265), .B(n5598), .Z(n5597) );
  XNOR U5579 ( .A(n5599), .B(n5600), .Z(n5598) );
  XOR U5580 ( .A(n5601), .B(n5602), .Z(n5573) );
  AND U5581 ( .A(n5603), .B(n5604), .Z(n5602) );
  XNOR U5582 ( .A(n5601), .B(n5589), .Z(n5604) );
  IV U5583 ( .A(n5542), .Z(n5589) );
  XNOR U5584 ( .A(n5605), .B(n5582), .Z(n5542) );
  XNOR U5585 ( .A(n5606), .B(n5588), .Z(n5582) );
  XNOR U5586 ( .A(n5607), .B(n5608), .Z(n5588) );
  NOR U5587 ( .A(n5609), .B(n5610), .Z(n5608) );
  XOR U5588 ( .A(n5607), .B(n5611), .Z(n5609) );
  XNOR U5589 ( .A(n5587), .B(n5579), .Z(n5606) );
  XOR U5590 ( .A(n5612), .B(n5613), .Z(n5579) );
  AND U5591 ( .A(n5614), .B(n5615), .Z(n5613) );
  XOR U5592 ( .A(n5612), .B(n5616), .Z(n5614) );
  XNOR U5593 ( .A(n5617), .B(n5584), .Z(n5587) );
  XOR U5594 ( .A(n5618), .B(n5619), .Z(n5584) );
  AND U5595 ( .A(n5620), .B(n5621), .Z(n5619) );
  XNOR U5596 ( .A(n5622), .B(n5623), .Z(n5620) );
  IV U5597 ( .A(n5618), .Z(n5622) );
  XNOR U5598 ( .A(n5624), .B(n5625), .Z(n5617) );
  NOR U5599 ( .A(n5626), .B(n5627), .Z(n5625) );
  XNOR U5600 ( .A(n5624), .B(n5628), .Z(n5626) );
  XNOR U5601 ( .A(n5583), .B(n5590), .Z(n5605) );
  NOR U5602 ( .A(n5548), .B(n5629), .Z(n5590) );
  XOR U5603 ( .A(n5595), .B(n5594), .Z(n5583) );
  XNOR U5604 ( .A(n5630), .B(n5591), .Z(n5594) );
  XOR U5605 ( .A(n5631), .B(n5632), .Z(n5591) );
  AND U5606 ( .A(n5633), .B(n5634), .Z(n5632) );
  XNOR U5607 ( .A(n5635), .B(n5636), .Z(n5633) );
  IV U5608 ( .A(n5631), .Z(n5635) );
  XNOR U5609 ( .A(n5637), .B(n5638), .Z(n5630) );
  NOR U5610 ( .A(n5639), .B(n5640), .Z(n5638) );
  XNOR U5611 ( .A(n5637), .B(n5641), .Z(n5639) );
  XOR U5612 ( .A(n5642), .B(n5643), .Z(n5595) );
  NOR U5613 ( .A(n5644), .B(n5645), .Z(n5643) );
  XNOR U5614 ( .A(n5642), .B(n5646), .Z(n5644) );
  XNOR U5615 ( .A(n5539), .B(n5601), .Z(n5603) );
  XNOR U5616 ( .A(n5647), .B(n5648), .Z(n5539) );
  AND U5617 ( .A(n265), .B(n5649), .Z(n5648) );
  XNOR U5618 ( .A(n5650), .B(n5651), .Z(n5649) );
  AND U5619 ( .A(n5545), .B(n5548), .Z(n5601) );
  XOR U5620 ( .A(n5652), .B(n5629), .Z(n5548) );
  XNOR U5621 ( .A(p_input[160]), .B(p_input[256]), .Z(n5629) );
  XNOR U5622 ( .A(n5616), .B(n5615), .Z(n5652) );
  XNOR U5623 ( .A(n5653), .B(n5623), .Z(n5615) );
  XNOR U5624 ( .A(n5611), .B(n5610), .Z(n5623) );
  XNOR U5625 ( .A(n5654), .B(n5607), .Z(n5610) );
  XNOR U5626 ( .A(p_input[170]), .B(p_input[266]), .Z(n5607) );
  XOR U5627 ( .A(p_input[171]), .B(n3382), .Z(n5654) );
  XOR U5628 ( .A(p_input[172]), .B(p_input[268]), .Z(n5611) );
  XOR U5629 ( .A(n5621), .B(n5655), .Z(n5653) );
  IV U5630 ( .A(n5612), .Z(n5655) );
  XOR U5631 ( .A(p_input[161]), .B(p_input[257]), .Z(n5612) );
  XNOR U5632 ( .A(n5656), .B(n5628), .Z(n5621) );
  XNOR U5633 ( .A(p_input[175]), .B(n3385), .Z(n5628) );
  XOR U5634 ( .A(n5618), .B(n5627), .Z(n5656) );
  XOR U5635 ( .A(n5657), .B(n5624), .Z(n5627) );
  XOR U5636 ( .A(p_input[173]), .B(p_input[269]), .Z(n5624) );
  XOR U5637 ( .A(p_input[174]), .B(n3387), .Z(n5657) );
  XOR U5638 ( .A(p_input[169]), .B(p_input[265]), .Z(n5618) );
  XOR U5639 ( .A(n5636), .B(n5634), .Z(n5616) );
  XNOR U5640 ( .A(n5658), .B(n5641), .Z(n5634) );
  XOR U5641 ( .A(p_input[168]), .B(p_input[264]), .Z(n5641) );
  XOR U5642 ( .A(n5631), .B(n5640), .Z(n5658) );
  XOR U5643 ( .A(n5659), .B(n5637), .Z(n5640) );
  XOR U5644 ( .A(p_input[166]), .B(p_input[262]), .Z(n5637) );
  XOR U5645 ( .A(p_input[167]), .B(n3625), .Z(n5659) );
  XOR U5646 ( .A(p_input[162]), .B(p_input[258]), .Z(n5631) );
  XNOR U5647 ( .A(n5646), .B(n5645), .Z(n5636) );
  XOR U5648 ( .A(n5660), .B(n5642), .Z(n5645) );
  XOR U5649 ( .A(p_input[163]), .B(p_input[259]), .Z(n5642) );
  XOR U5650 ( .A(p_input[164]), .B(n3627), .Z(n5660) );
  XOR U5651 ( .A(p_input[165]), .B(p_input[261]), .Z(n5646) );
  XNOR U5652 ( .A(n5661), .B(n5662), .Z(n5545) );
  AND U5653 ( .A(n265), .B(n5663), .Z(n5662) );
  XNOR U5654 ( .A(n5664), .B(n5665), .Z(n265) );
  NOR U5655 ( .A(n5666), .B(n5667), .Z(n5665) );
  XNOR U5656 ( .A(n5664), .B(n5668), .Z(n5667) );
  NOR U5657 ( .A(n5664), .B(n5554), .Z(n5666) );
  XOR U5658 ( .A(n5669), .B(n5670), .Z(n5664) );
  AND U5659 ( .A(n5671), .B(n5672), .Z(n5670) );
  XOR U5660 ( .A(n5571), .B(n5669), .Z(n5672) );
  XOR U5661 ( .A(n5669), .B(n5572), .Z(n5671) );
  XOR U5662 ( .A(n5673), .B(n5674), .Z(n5669) );
  AND U5663 ( .A(n5675), .B(n5676), .Z(n5674) );
  XOR U5664 ( .A(n5599), .B(n5673), .Z(n5676) );
  XOR U5665 ( .A(n5673), .B(n5600), .Z(n5675) );
  XOR U5666 ( .A(n5677), .B(n5678), .Z(n5673) );
  AND U5667 ( .A(n5679), .B(n5680), .Z(n5678) );
  XOR U5668 ( .A(n5677), .B(n5650), .Z(n5680) );
  XNOR U5669 ( .A(n5681), .B(n5682), .Z(n5508) );
  AND U5670 ( .A(n269), .B(n5683), .Z(n5682) );
  XNOR U5671 ( .A(n5684), .B(n5685), .Z(n269) );
  NOR U5672 ( .A(n5686), .B(n5687), .Z(n5685) );
  XOR U5673 ( .A(n5480), .B(n5684), .Z(n5687) );
  NOR U5674 ( .A(n5684), .B(n5479), .Z(n5686) );
  XOR U5675 ( .A(n5688), .B(n5689), .Z(n5684) );
  AND U5676 ( .A(n5690), .B(n5691), .Z(n5689) );
  XOR U5677 ( .A(n5688), .B(n5486), .Z(n5690) );
  XOR U5678 ( .A(n5692), .B(n5693), .Z(n5472) );
  AND U5679 ( .A(n273), .B(n5683), .Z(n5693) );
  XNOR U5680 ( .A(n5681), .B(n5692), .Z(n5683) );
  XNOR U5681 ( .A(n5694), .B(n5695), .Z(n273) );
  NOR U5682 ( .A(n5696), .B(n5697), .Z(n5695) );
  XNOR U5683 ( .A(n5480), .B(n5698), .Z(n5697) );
  IV U5684 ( .A(n5694), .Z(n5698) );
  AND U5685 ( .A(n5699), .B(n5700), .Z(n5480) );
  NOR U5686 ( .A(n5694), .B(n5479), .Z(n5696) );
  AND U5687 ( .A(n5554), .B(n5553), .Z(n5479) );
  IV U5688 ( .A(n5668), .Z(n5553) );
  XOR U5689 ( .A(n5688), .B(n5701), .Z(n5694) );
  AND U5690 ( .A(n5702), .B(n5691), .Z(n5701) );
  XNOR U5691 ( .A(n5525), .B(n5688), .Z(n5691) );
  XOR U5692 ( .A(n5572), .B(n5703), .Z(n5525) );
  AND U5693 ( .A(n276), .B(n5704), .Z(n5703) );
  XOR U5694 ( .A(n5568), .B(n5572), .Z(n5704) );
  XNOR U5695 ( .A(n5705), .B(n5688), .Z(n5702) );
  IV U5696 ( .A(n5486), .Z(n5705) );
  XOR U5697 ( .A(n5706), .B(n5707), .Z(n5486) );
  AND U5698 ( .A(n292), .B(n5708), .Z(n5707) );
  XOR U5699 ( .A(n5709), .B(n5710), .Z(n5688) );
  AND U5700 ( .A(n5711), .B(n5712), .Z(n5710) );
  XNOR U5701 ( .A(n5535), .B(n5709), .Z(n5712) );
  XOR U5702 ( .A(n5600), .B(n5713), .Z(n5535) );
  AND U5703 ( .A(n276), .B(n5714), .Z(n5713) );
  XOR U5704 ( .A(n5596), .B(n5600), .Z(n5714) );
  XOR U5705 ( .A(n5709), .B(n5495), .Z(n5711) );
  XOR U5706 ( .A(n5715), .B(n5716), .Z(n5495) );
  AND U5707 ( .A(n292), .B(n5717), .Z(n5716) );
  XOR U5708 ( .A(n5718), .B(n5719), .Z(n5709) );
  AND U5709 ( .A(n5720), .B(n5721), .Z(n5719) );
  XNOR U5710 ( .A(n5718), .B(n5543), .Z(n5721) );
  XOR U5711 ( .A(n5651), .B(n5722), .Z(n5543) );
  AND U5712 ( .A(n276), .B(n5723), .Z(n5722) );
  XOR U5713 ( .A(n5647), .B(n5651), .Z(n5723) );
  XNOR U5714 ( .A(n5724), .B(n5718), .Z(n5720) );
  IV U5715 ( .A(n5505), .Z(n5724) );
  XOR U5716 ( .A(n5725), .B(n5726), .Z(n5505) );
  AND U5717 ( .A(n292), .B(n5727), .Z(n5726) );
  AND U5718 ( .A(n5692), .B(n5681), .Z(n5718) );
  XNOR U5719 ( .A(n5728), .B(n5729), .Z(n5681) );
  AND U5720 ( .A(n276), .B(n5663), .Z(n5729) );
  XNOR U5721 ( .A(n5661), .B(n5728), .Z(n5663) );
  XNOR U5722 ( .A(n5730), .B(n5731), .Z(n276) );
  NOR U5723 ( .A(n5732), .B(n5733), .Z(n5731) );
  XNOR U5724 ( .A(n5730), .B(n5668), .Z(n5733) );
  NOR U5725 ( .A(n5699), .B(n5700), .Z(n5668) );
  NOR U5726 ( .A(n5730), .B(n5554), .Z(n5732) );
  AND U5727 ( .A(n5734), .B(n5735), .Z(n5554) );
  IV U5728 ( .A(n5736), .Z(n5734) );
  XOR U5729 ( .A(n5737), .B(n5738), .Z(n5730) );
  AND U5730 ( .A(n5739), .B(n5740), .Z(n5738) );
  XNOR U5731 ( .A(n5737), .B(n5568), .Z(n5740) );
  IV U5732 ( .A(n5571), .Z(n5568) );
  XOR U5733 ( .A(n5741), .B(n5742), .Z(n5571) );
  AND U5734 ( .A(n280), .B(n5743), .Z(n5742) );
  XOR U5735 ( .A(n5744), .B(n5741), .Z(n5743) );
  XOR U5736 ( .A(n5572), .B(n5737), .Z(n5739) );
  XOR U5737 ( .A(n5745), .B(n5746), .Z(n5572) );
  AND U5738 ( .A(n288), .B(n5708), .Z(n5746) );
  XOR U5739 ( .A(n5745), .B(n5706), .Z(n5708) );
  XOR U5740 ( .A(n5747), .B(n5748), .Z(n5737) );
  AND U5741 ( .A(n5749), .B(n5750), .Z(n5748) );
  XNOR U5742 ( .A(n5747), .B(n5596), .Z(n5750) );
  IV U5743 ( .A(n5599), .Z(n5596) );
  XOR U5744 ( .A(n5751), .B(n5752), .Z(n5599) );
  AND U5745 ( .A(n280), .B(n5753), .Z(n5752) );
  XNOR U5746 ( .A(n5754), .B(n5751), .Z(n5753) );
  XOR U5747 ( .A(n5600), .B(n5747), .Z(n5749) );
  XOR U5748 ( .A(n5755), .B(n5756), .Z(n5600) );
  AND U5749 ( .A(n288), .B(n5717), .Z(n5756) );
  XOR U5750 ( .A(n5755), .B(n5715), .Z(n5717) );
  XOR U5751 ( .A(n5677), .B(n5757), .Z(n5747) );
  AND U5752 ( .A(n5679), .B(n5758), .Z(n5757) );
  XNOR U5753 ( .A(n5677), .B(n5647), .Z(n5758) );
  IV U5754 ( .A(n5650), .Z(n5647) );
  XOR U5755 ( .A(n5759), .B(n5760), .Z(n5650) );
  AND U5756 ( .A(n280), .B(n5761), .Z(n5760) );
  XOR U5757 ( .A(n5762), .B(n5759), .Z(n5761) );
  XOR U5758 ( .A(n5651), .B(n5677), .Z(n5679) );
  XOR U5759 ( .A(n5763), .B(n5764), .Z(n5651) );
  AND U5760 ( .A(n288), .B(n5727), .Z(n5764) );
  XOR U5761 ( .A(n5763), .B(n5725), .Z(n5727) );
  AND U5762 ( .A(n5728), .B(n5661), .Z(n5677) );
  XNOR U5763 ( .A(n5765), .B(n5766), .Z(n5661) );
  AND U5764 ( .A(n280), .B(n5767), .Z(n5766) );
  XNOR U5765 ( .A(n5768), .B(n5765), .Z(n5767) );
  XNOR U5766 ( .A(n5769), .B(n5770), .Z(n280) );
  NOR U5767 ( .A(n5771), .B(n5772), .Z(n5770) );
  XNOR U5768 ( .A(n5769), .B(n5736), .Z(n5772) );
  NOR U5769 ( .A(n5773), .B(n5774), .Z(n5736) );
  NOR U5770 ( .A(n5769), .B(n5735), .Z(n5771) );
  AND U5771 ( .A(n5775), .B(n5776), .Z(n5735) );
  XOR U5772 ( .A(n5777), .B(n5778), .Z(n5769) );
  AND U5773 ( .A(n5779), .B(n5780), .Z(n5778) );
  XNOR U5774 ( .A(n5777), .B(n5775), .Z(n5780) );
  IV U5775 ( .A(n5744), .Z(n5775) );
  XOR U5776 ( .A(n5781), .B(n5782), .Z(n5744) );
  XOR U5777 ( .A(n5783), .B(n5776), .Z(n5782) );
  AND U5778 ( .A(n5754), .B(n5784), .Z(n5776) );
  AND U5779 ( .A(n5785), .B(n5786), .Z(n5783) );
  XOR U5780 ( .A(n5787), .B(n5781), .Z(n5785) );
  XNOR U5781 ( .A(n5741), .B(n5777), .Z(n5779) );
  XNOR U5782 ( .A(n5788), .B(n5789), .Z(n5741) );
  AND U5783 ( .A(n284), .B(n5790), .Z(n5789) );
  XNOR U5784 ( .A(n5791), .B(n5792), .Z(n5790) );
  XOR U5785 ( .A(n5793), .B(n5794), .Z(n5777) );
  AND U5786 ( .A(n5795), .B(n5796), .Z(n5794) );
  XNOR U5787 ( .A(n5793), .B(n5754), .Z(n5796) );
  XOR U5788 ( .A(n5797), .B(n5786), .Z(n5754) );
  XNOR U5789 ( .A(n5798), .B(n5781), .Z(n5786) );
  XOR U5790 ( .A(n5799), .B(n5800), .Z(n5781) );
  AND U5791 ( .A(n5801), .B(n5802), .Z(n5800) );
  XOR U5792 ( .A(n5803), .B(n5799), .Z(n5801) );
  XNOR U5793 ( .A(n5804), .B(n5805), .Z(n5798) );
  AND U5794 ( .A(n5806), .B(n5807), .Z(n5805) );
  XOR U5795 ( .A(n5804), .B(n5808), .Z(n5806) );
  XNOR U5796 ( .A(n5787), .B(n5784), .Z(n5797) );
  AND U5797 ( .A(n5809), .B(n5810), .Z(n5784) );
  XOR U5798 ( .A(n5811), .B(n5812), .Z(n5787) );
  AND U5799 ( .A(n5813), .B(n5814), .Z(n5812) );
  XOR U5800 ( .A(n5811), .B(n5815), .Z(n5813) );
  XNOR U5801 ( .A(n5751), .B(n5793), .Z(n5795) );
  XNOR U5802 ( .A(n5816), .B(n5817), .Z(n5751) );
  AND U5803 ( .A(n284), .B(n5818), .Z(n5817) );
  XNOR U5804 ( .A(n5819), .B(n5820), .Z(n5818) );
  XOR U5805 ( .A(n5821), .B(n5822), .Z(n5793) );
  AND U5806 ( .A(n5823), .B(n5824), .Z(n5822) );
  XNOR U5807 ( .A(n5821), .B(n5809), .Z(n5824) );
  IV U5808 ( .A(n5762), .Z(n5809) );
  XNOR U5809 ( .A(n5825), .B(n5802), .Z(n5762) );
  XNOR U5810 ( .A(n5826), .B(n5808), .Z(n5802) );
  XNOR U5811 ( .A(n5827), .B(n5828), .Z(n5808) );
  NOR U5812 ( .A(n5829), .B(n5830), .Z(n5828) );
  XOR U5813 ( .A(n5827), .B(n5831), .Z(n5829) );
  XNOR U5814 ( .A(n5807), .B(n5799), .Z(n5826) );
  XOR U5815 ( .A(n5832), .B(n5833), .Z(n5799) );
  AND U5816 ( .A(n5834), .B(n5835), .Z(n5833) );
  XOR U5817 ( .A(n5832), .B(n5836), .Z(n5834) );
  XNOR U5818 ( .A(n5837), .B(n5804), .Z(n5807) );
  XOR U5819 ( .A(n5838), .B(n5839), .Z(n5804) );
  AND U5820 ( .A(n5840), .B(n5841), .Z(n5839) );
  XNOR U5821 ( .A(n5842), .B(n5843), .Z(n5840) );
  IV U5822 ( .A(n5838), .Z(n5842) );
  XNOR U5823 ( .A(n5844), .B(n5845), .Z(n5837) );
  NOR U5824 ( .A(n5846), .B(n5847), .Z(n5845) );
  XNOR U5825 ( .A(n5844), .B(n5848), .Z(n5846) );
  XNOR U5826 ( .A(n5803), .B(n5810), .Z(n5825) );
  NOR U5827 ( .A(n5768), .B(n5849), .Z(n5810) );
  XOR U5828 ( .A(n5815), .B(n5814), .Z(n5803) );
  XNOR U5829 ( .A(n5850), .B(n5811), .Z(n5814) );
  XOR U5830 ( .A(n5851), .B(n5852), .Z(n5811) );
  AND U5831 ( .A(n5853), .B(n5854), .Z(n5852) );
  XNOR U5832 ( .A(n5855), .B(n5856), .Z(n5853) );
  IV U5833 ( .A(n5851), .Z(n5855) );
  XNOR U5834 ( .A(n5857), .B(n5858), .Z(n5850) );
  NOR U5835 ( .A(n5859), .B(n5860), .Z(n5858) );
  XNOR U5836 ( .A(n5857), .B(n5861), .Z(n5859) );
  XOR U5837 ( .A(n5862), .B(n5863), .Z(n5815) );
  NOR U5838 ( .A(n5864), .B(n5865), .Z(n5863) );
  XNOR U5839 ( .A(n5862), .B(n5866), .Z(n5864) );
  XNOR U5840 ( .A(n5759), .B(n5821), .Z(n5823) );
  XNOR U5841 ( .A(n5867), .B(n5868), .Z(n5759) );
  AND U5842 ( .A(n284), .B(n5869), .Z(n5868) );
  XNOR U5843 ( .A(n5870), .B(n5871), .Z(n5869) );
  AND U5844 ( .A(n5765), .B(n5768), .Z(n5821) );
  XOR U5845 ( .A(n5872), .B(n5849), .Z(n5768) );
  XNOR U5846 ( .A(p_input[176]), .B(p_input[256]), .Z(n5849) );
  XNOR U5847 ( .A(n5836), .B(n5835), .Z(n5872) );
  XNOR U5848 ( .A(n5873), .B(n5843), .Z(n5835) );
  XNOR U5849 ( .A(n5831), .B(n5830), .Z(n5843) );
  XNOR U5850 ( .A(n5874), .B(n5827), .Z(n5830) );
  XNOR U5851 ( .A(p_input[186]), .B(p_input[266]), .Z(n5827) );
  XOR U5852 ( .A(p_input[187]), .B(n3382), .Z(n5874) );
  XOR U5853 ( .A(p_input[188]), .B(p_input[268]), .Z(n5831) );
  XOR U5854 ( .A(n5841), .B(n5875), .Z(n5873) );
  IV U5855 ( .A(n5832), .Z(n5875) );
  XOR U5856 ( .A(p_input[177]), .B(p_input[257]), .Z(n5832) );
  XNOR U5857 ( .A(n5876), .B(n5848), .Z(n5841) );
  XNOR U5858 ( .A(p_input[191]), .B(n3385), .Z(n5848) );
  XOR U5859 ( .A(n5838), .B(n5847), .Z(n5876) );
  XOR U5860 ( .A(n5877), .B(n5844), .Z(n5847) );
  XOR U5861 ( .A(p_input[189]), .B(p_input[269]), .Z(n5844) );
  XOR U5862 ( .A(p_input[190]), .B(n3387), .Z(n5877) );
  XOR U5863 ( .A(p_input[185]), .B(p_input[265]), .Z(n5838) );
  XOR U5864 ( .A(n5856), .B(n5854), .Z(n5836) );
  XNOR U5865 ( .A(n5878), .B(n5861), .Z(n5854) );
  XOR U5866 ( .A(p_input[184]), .B(p_input[264]), .Z(n5861) );
  XOR U5867 ( .A(n5851), .B(n5860), .Z(n5878) );
  XOR U5868 ( .A(n5879), .B(n5857), .Z(n5860) );
  XOR U5869 ( .A(p_input[182]), .B(p_input[262]), .Z(n5857) );
  XOR U5870 ( .A(p_input[183]), .B(n3625), .Z(n5879) );
  XOR U5871 ( .A(p_input[178]), .B(p_input[258]), .Z(n5851) );
  XNOR U5872 ( .A(n5866), .B(n5865), .Z(n5856) );
  XOR U5873 ( .A(n5880), .B(n5862), .Z(n5865) );
  XOR U5874 ( .A(p_input[179]), .B(p_input[259]), .Z(n5862) );
  XOR U5875 ( .A(p_input[180]), .B(n3627), .Z(n5880) );
  XOR U5876 ( .A(p_input[181]), .B(p_input[261]), .Z(n5866) );
  XNOR U5877 ( .A(n5881), .B(n5882), .Z(n5765) );
  AND U5878 ( .A(n284), .B(n5883), .Z(n5882) );
  XNOR U5879 ( .A(n5884), .B(n5885), .Z(n284) );
  NOR U5880 ( .A(n5886), .B(n5887), .Z(n5885) );
  XNOR U5881 ( .A(n5884), .B(n5888), .Z(n5887) );
  NOR U5882 ( .A(n5884), .B(n5774), .Z(n5886) );
  XOR U5883 ( .A(n5889), .B(n5890), .Z(n5884) );
  AND U5884 ( .A(n5891), .B(n5892), .Z(n5890) );
  XOR U5885 ( .A(n5791), .B(n5889), .Z(n5892) );
  XOR U5886 ( .A(n5889), .B(n5792), .Z(n5891) );
  XOR U5887 ( .A(n5893), .B(n5894), .Z(n5889) );
  AND U5888 ( .A(n5895), .B(n5896), .Z(n5894) );
  XOR U5889 ( .A(n5819), .B(n5893), .Z(n5896) );
  XOR U5890 ( .A(n5893), .B(n5820), .Z(n5895) );
  XOR U5891 ( .A(n5897), .B(n5898), .Z(n5893) );
  AND U5892 ( .A(n5899), .B(n5900), .Z(n5898) );
  XOR U5893 ( .A(n5897), .B(n5870), .Z(n5900) );
  XNOR U5894 ( .A(n5901), .B(n5902), .Z(n5728) );
  AND U5895 ( .A(n288), .B(n5903), .Z(n5902) );
  XNOR U5896 ( .A(n5904), .B(n5905), .Z(n288) );
  NOR U5897 ( .A(n5906), .B(n5907), .Z(n5905) );
  XOR U5898 ( .A(n5700), .B(n5904), .Z(n5907) );
  NOR U5899 ( .A(n5904), .B(n5699), .Z(n5906) );
  XOR U5900 ( .A(n5908), .B(n5909), .Z(n5904) );
  AND U5901 ( .A(n5910), .B(n5911), .Z(n5909) );
  XOR U5902 ( .A(n5908), .B(n5706), .Z(n5910) );
  XOR U5903 ( .A(n5912), .B(n5913), .Z(n5692) );
  AND U5904 ( .A(n292), .B(n5903), .Z(n5913) );
  XNOR U5905 ( .A(n5901), .B(n5912), .Z(n5903) );
  XNOR U5906 ( .A(n5914), .B(n5915), .Z(n292) );
  NOR U5907 ( .A(n5916), .B(n5917), .Z(n5915) );
  XNOR U5908 ( .A(n5700), .B(n5918), .Z(n5917) );
  IV U5909 ( .A(n5914), .Z(n5918) );
  AND U5910 ( .A(n5919), .B(n5920), .Z(n5700) );
  NOR U5911 ( .A(n5914), .B(n5699), .Z(n5916) );
  AND U5912 ( .A(n5774), .B(n5773), .Z(n5699) );
  IV U5913 ( .A(n5888), .Z(n5773) );
  XOR U5914 ( .A(n5908), .B(n5921), .Z(n5914) );
  AND U5915 ( .A(n5922), .B(n5911), .Z(n5921) );
  XNOR U5916 ( .A(n5745), .B(n5908), .Z(n5911) );
  XOR U5917 ( .A(n5792), .B(n5923), .Z(n5745) );
  AND U5918 ( .A(n295), .B(n5924), .Z(n5923) );
  XOR U5919 ( .A(n5788), .B(n5792), .Z(n5924) );
  XNOR U5920 ( .A(n5925), .B(n5908), .Z(n5922) );
  IV U5921 ( .A(n5706), .Z(n5925) );
  XOR U5922 ( .A(n5926), .B(n5927), .Z(n5706) );
  AND U5923 ( .A(n310), .B(n5928), .Z(n5927) );
  XOR U5924 ( .A(n5929), .B(n5930), .Z(n5908) );
  AND U5925 ( .A(n5931), .B(n5932), .Z(n5930) );
  XNOR U5926 ( .A(n5755), .B(n5929), .Z(n5932) );
  XOR U5927 ( .A(n5820), .B(n5933), .Z(n5755) );
  AND U5928 ( .A(n295), .B(n5934), .Z(n5933) );
  XOR U5929 ( .A(n5816), .B(n5820), .Z(n5934) );
  XOR U5930 ( .A(n5929), .B(n5715), .Z(n5931) );
  XOR U5931 ( .A(n5935), .B(n5936), .Z(n5715) );
  AND U5932 ( .A(n310), .B(n5937), .Z(n5936) );
  XOR U5933 ( .A(n5938), .B(n5939), .Z(n5929) );
  AND U5934 ( .A(n5940), .B(n5941), .Z(n5939) );
  XNOR U5935 ( .A(n5938), .B(n5763), .Z(n5941) );
  XOR U5936 ( .A(n5871), .B(n5942), .Z(n5763) );
  AND U5937 ( .A(n295), .B(n5943), .Z(n5942) );
  XOR U5938 ( .A(n5867), .B(n5871), .Z(n5943) );
  XNOR U5939 ( .A(n5944), .B(n5938), .Z(n5940) );
  IV U5940 ( .A(n5725), .Z(n5944) );
  XOR U5941 ( .A(n5945), .B(n5946), .Z(n5725) );
  AND U5942 ( .A(n310), .B(n5947), .Z(n5946) );
  AND U5943 ( .A(n5912), .B(n5901), .Z(n5938) );
  XNOR U5944 ( .A(n5948), .B(n5949), .Z(n5901) );
  AND U5945 ( .A(n295), .B(n5883), .Z(n5949) );
  XNOR U5946 ( .A(n5881), .B(n5948), .Z(n5883) );
  XNOR U5947 ( .A(n5950), .B(n5951), .Z(n295) );
  NOR U5948 ( .A(n5952), .B(n5953), .Z(n5951) );
  XNOR U5949 ( .A(n5950), .B(n5888), .Z(n5953) );
  NOR U5950 ( .A(n5919), .B(n5920), .Z(n5888) );
  NOR U5951 ( .A(n5950), .B(n5774), .Z(n5952) );
  AND U5952 ( .A(n5954), .B(n5955), .Z(n5774) );
  IV U5953 ( .A(n5956), .Z(n5954) );
  XOR U5954 ( .A(n5957), .B(n5958), .Z(n5950) );
  AND U5955 ( .A(n5959), .B(n5960), .Z(n5958) );
  XNOR U5956 ( .A(n5957), .B(n5788), .Z(n5960) );
  IV U5957 ( .A(n5791), .Z(n5788) );
  XOR U5958 ( .A(n5961), .B(n5962), .Z(n5791) );
  AND U5959 ( .A(n299), .B(n5963), .Z(n5962) );
  XOR U5960 ( .A(n5964), .B(n5961), .Z(n5963) );
  XOR U5961 ( .A(n5792), .B(n5957), .Z(n5959) );
  XOR U5962 ( .A(n5965), .B(n5966), .Z(n5792) );
  AND U5963 ( .A(n306), .B(n5928), .Z(n5966) );
  XOR U5964 ( .A(n5965), .B(n5926), .Z(n5928) );
  XOR U5965 ( .A(n5967), .B(n5968), .Z(n5957) );
  AND U5966 ( .A(n5969), .B(n5970), .Z(n5968) );
  XNOR U5967 ( .A(n5967), .B(n5816), .Z(n5970) );
  IV U5968 ( .A(n5819), .Z(n5816) );
  XOR U5969 ( .A(n5971), .B(n5972), .Z(n5819) );
  AND U5970 ( .A(n299), .B(n5973), .Z(n5972) );
  XNOR U5971 ( .A(n5974), .B(n5971), .Z(n5973) );
  XOR U5972 ( .A(n5820), .B(n5967), .Z(n5969) );
  XOR U5973 ( .A(n5975), .B(n5976), .Z(n5820) );
  AND U5974 ( .A(n306), .B(n5937), .Z(n5976) );
  XOR U5975 ( .A(n5975), .B(n5935), .Z(n5937) );
  XOR U5976 ( .A(n5897), .B(n5977), .Z(n5967) );
  AND U5977 ( .A(n5899), .B(n5978), .Z(n5977) );
  XNOR U5978 ( .A(n5897), .B(n5867), .Z(n5978) );
  IV U5979 ( .A(n5870), .Z(n5867) );
  XOR U5980 ( .A(n5979), .B(n5980), .Z(n5870) );
  AND U5981 ( .A(n299), .B(n5981), .Z(n5980) );
  XOR U5982 ( .A(n5982), .B(n5979), .Z(n5981) );
  XOR U5983 ( .A(n5871), .B(n5897), .Z(n5899) );
  XOR U5984 ( .A(n5983), .B(n5984), .Z(n5871) );
  AND U5985 ( .A(n306), .B(n5947), .Z(n5984) );
  XOR U5986 ( .A(n5983), .B(n5945), .Z(n5947) );
  AND U5987 ( .A(n5948), .B(n5881), .Z(n5897) );
  XNOR U5988 ( .A(n5985), .B(n5986), .Z(n5881) );
  AND U5989 ( .A(n299), .B(n5987), .Z(n5986) );
  XNOR U5990 ( .A(n5988), .B(n5985), .Z(n5987) );
  XNOR U5991 ( .A(n5989), .B(n5990), .Z(n299) );
  NOR U5992 ( .A(n5991), .B(n5992), .Z(n5990) );
  XNOR U5993 ( .A(n5989), .B(n5956), .Z(n5992) );
  NOR U5994 ( .A(n5993), .B(n5994), .Z(n5956) );
  NOR U5995 ( .A(n5989), .B(n5955), .Z(n5991) );
  AND U5996 ( .A(n5995), .B(n5996), .Z(n5955) );
  XOR U5997 ( .A(n5997), .B(n5998), .Z(n5989) );
  AND U5998 ( .A(n5999), .B(n6000), .Z(n5998) );
  XNOR U5999 ( .A(n5997), .B(n5995), .Z(n6000) );
  IV U6000 ( .A(n5964), .Z(n5995) );
  XOR U6001 ( .A(n6001), .B(n6002), .Z(n5964) );
  XOR U6002 ( .A(n6003), .B(n5996), .Z(n6002) );
  AND U6003 ( .A(n5974), .B(n6004), .Z(n5996) );
  AND U6004 ( .A(n6005), .B(n6006), .Z(n6003) );
  XOR U6005 ( .A(n6007), .B(n6001), .Z(n6005) );
  XNOR U6006 ( .A(n5961), .B(n5997), .Z(n5999) );
  XNOR U6007 ( .A(n6008), .B(n6009), .Z(n5961) );
  AND U6008 ( .A(n302), .B(n6010), .Z(n6009) );
  XOR U6009 ( .A(n6011), .B(n6012), .Z(n5997) );
  AND U6010 ( .A(n6013), .B(n6014), .Z(n6012) );
  XNOR U6011 ( .A(n6011), .B(n5974), .Z(n6014) );
  XOR U6012 ( .A(n6015), .B(n6006), .Z(n5974) );
  XNOR U6013 ( .A(n6016), .B(n6001), .Z(n6006) );
  XOR U6014 ( .A(n6017), .B(n6018), .Z(n6001) );
  AND U6015 ( .A(n6019), .B(n6020), .Z(n6018) );
  XOR U6016 ( .A(n6021), .B(n6017), .Z(n6019) );
  XNOR U6017 ( .A(n6022), .B(n6023), .Z(n6016) );
  AND U6018 ( .A(n6024), .B(n6025), .Z(n6023) );
  XOR U6019 ( .A(n6022), .B(n6026), .Z(n6024) );
  XNOR U6020 ( .A(n6007), .B(n6004), .Z(n6015) );
  AND U6021 ( .A(n6027), .B(n6028), .Z(n6004) );
  XOR U6022 ( .A(n6029), .B(n6030), .Z(n6007) );
  AND U6023 ( .A(n6031), .B(n6032), .Z(n6030) );
  XOR U6024 ( .A(n6029), .B(n6033), .Z(n6031) );
  XNOR U6025 ( .A(n5971), .B(n6011), .Z(n6013) );
  XNOR U6026 ( .A(n6034), .B(n6035), .Z(n5971) );
  AND U6027 ( .A(n302), .B(n6036), .Z(n6035) );
  XOR U6028 ( .A(n6037), .B(n6038), .Z(n6011) );
  AND U6029 ( .A(n6039), .B(n6040), .Z(n6038) );
  XNOR U6030 ( .A(n6037), .B(n6027), .Z(n6040) );
  IV U6031 ( .A(n5982), .Z(n6027) );
  XNOR U6032 ( .A(n6041), .B(n6020), .Z(n5982) );
  XNOR U6033 ( .A(n6042), .B(n6026), .Z(n6020) );
  XNOR U6034 ( .A(n6043), .B(n6044), .Z(n6026) );
  NOR U6035 ( .A(n6045), .B(n6046), .Z(n6044) );
  XOR U6036 ( .A(n6043), .B(n6047), .Z(n6045) );
  XNOR U6037 ( .A(n6025), .B(n6017), .Z(n6042) );
  XOR U6038 ( .A(n6048), .B(n6049), .Z(n6017) );
  AND U6039 ( .A(n6050), .B(n6051), .Z(n6049) );
  XOR U6040 ( .A(n6048), .B(n6052), .Z(n6050) );
  XNOR U6041 ( .A(n6053), .B(n6022), .Z(n6025) );
  XOR U6042 ( .A(n6054), .B(n6055), .Z(n6022) );
  AND U6043 ( .A(n6056), .B(n6057), .Z(n6055) );
  XNOR U6044 ( .A(n6058), .B(n6059), .Z(n6056) );
  IV U6045 ( .A(n6054), .Z(n6058) );
  XNOR U6046 ( .A(n6060), .B(n6061), .Z(n6053) );
  NOR U6047 ( .A(n6062), .B(n6063), .Z(n6061) );
  XNOR U6048 ( .A(n6060), .B(n6064), .Z(n6062) );
  XNOR U6049 ( .A(n6021), .B(n6028), .Z(n6041) );
  NOR U6050 ( .A(n5988), .B(n6065), .Z(n6028) );
  XOR U6051 ( .A(n6033), .B(n6032), .Z(n6021) );
  XNOR U6052 ( .A(n6066), .B(n6029), .Z(n6032) );
  XOR U6053 ( .A(n6067), .B(n6068), .Z(n6029) );
  AND U6054 ( .A(n6069), .B(n6070), .Z(n6068) );
  XNOR U6055 ( .A(n6071), .B(n6072), .Z(n6069) );
  IV U6056 ( .A(n6067), .Z(n6071) );
  XNOR U6057 ( .A(n6073), .B(n6074), .Z(n6066) );
  NOR U6058 ( .A(n6075), .B(n6076), .Z(n6074) );
  XNOR U6059 ( .A(n6073), .B(n6077), .Z(n6075) );
  XOR U6060 ( .A(n6078), .B(n6079), .Z(n6033) );
  NOR U6061 ( .A(n6080), .B(n6081), .Z(n6079) );
  XNOR U6062 ( .A(n6078), .B(n6082), .Z(n6080) );
  XNOR U6063 ( .A(n5979), .B(n6037), .Z(n6039) );
  XNOR U6064 ( .A(n6083), .B(n6084), .Z(n5979) );
  AND U6065 ( .A(n302), .B(n6085), .Z(n6084) );
  XNOR U6066 ( .A(n6086), .B(n6087), .Z(n6085) );
  AND U6067 ( .A(n5985), .B(n5988), .Z(n6037) );
  XOR U6068 ( .A(n6088), .B(n6065), .Z(n5988) );
  XNOR U6069 ( .A(p_input[192]), .B(p_input[256]), .Z(n6065) );
  XNOR U6070 ( .A(n6052), .B(n6051), .Z(n6088) );
  XNOR U6071 ( .A(n6089), .B(n6059), .Z(n6051) );
  XNOR U6072 ( .A(n6047), .B(n6046), .Z(n6059) );
  XNOR U6073 ( .A(n6090), .B(n6043), .Z(n6046) );
  XNOR U6074 ( .A(p_input[202]), .B(p_input[266]), .Z(n6043) );
  XOR U6075 ( .A(p_input[203]), .B(n3382), .Z(n6090) );
  XOR U6076 ( .A(p_input[204]), .B(p_input[268]), .Z(n6047) );
  XOR U6077 ( .A(n6057), .B(n6091), .Z(n6089) );
  IV U6078 ( .A(n6048), .Z(n6091) );
  XOR U6079 ( .A(p_input[193]), .B(p_input[257]), .Z(n6048) );
  XNOR U6080 ( .A(n6092), .B(n6064), .Z(n6057) );
  XNOR U6081 ( .A(p_input[207]), .B(n3385), .Z(n6064) );
  IV U6082 ( .A(p_input[271]), .Z(n3385) );
  XOR U6083 ( .A(n6054), .B(n6063), .Z(n6092) );
  XOR U6084 ( .A(n6093), .B(n6060), .Z(n6063) );
  XOR U6085 ( .A(p_input[205]), .B(p_input[269]), .Z(n6060) );
  XOR U6086 ( .A(p_input[206]), .B(n3387), .Z(n6093) );
  XOR U6087 ( .A(p_input[201]), .B(p_input[265]), .Z(n6054) );
  XOR U6088 ( .A(n6072), .B(n6070), .Z(n6052) );
  XNOR U6089 ( .A(n6094), .B(n6077), .Z(n6070) );
  XOR U6090 ( .A(p_input[200]), .B(p_input[264]), .Z(n6077) );
  XOR U6091 ( .A(n6067), .B(n6076), .Z(n6094) );
  XOR U6092 ( .A(n6095), .B(n6073), .Z(n6076) );
  XOR U6093 ( .A(p_input[198]), .B(p_input[262]), .Z(n6073) );
  XOR U6094 ( .A(p_input[199]), .B(n3625), .Z(n6095) );
  XOR U6095 ( .A(p_input[194]), .B(p_input[258]), .Z(n6067) );
  XNOR U6096 ( .A(n6082), .B(n6081), .Z(n6072) );
  XOR U6097 ( .A(n6096), .B(n6078), .Z(n6081) );
  XOR U6098 ( .A(p_input[195]), .B(p_input[259]), .Z(n6078) );
  XOR U6099 ( .A(p_input[196]), .B(n3627), .Z(n6096) );
  XOR U6100 ( .A(p_input[197]), .B(p_input[261]), .Z(n6082) );
  XNOR U6101 ( .A(n6097), .B(n6098), .Z(n5985) );
  AND U6102 ( .A(n302), .B(n6099), .Z(n6098) );
  XNOR U6103 ( .A(n6100), .B(n6101), .Z(n302) );
  NOR U6104 ( .A(n6102), .B(n6103), .Z(n6101) );
  XOR U6105 ( .A(n6100), .B(n5993), .Z(n6103) );
  XNOR U6106 ( .A(n6104), .B(n6105), .Z(n5948) );
  AND U6107 ( .A(n306), .B(n6106), .Z(n6105) );
  XNOR U6108 ( .A(n6107), .B(n6108), .Z(n306) );
  NOR U6109 ( .A(n6109), .B(n6110), .Z(n6108) );
  XOR U6110 ( .A(n5920), .B(n6107), .Z(n6110) );
  NOR U6111 ( .A(n6107), .B(n5919), .Z(n6109) );
  XOR U6112 ( .A(n6111), .B(n6112), .Z(n6107) );
  AND U6113 ( .A(n6113), .B(n6114), .Z(n6112) );
  XOR U6114 ( .A(n6111), .B(n5926), .Z(n6113) );
  XOR U6115 ( .A(n6115), .B(n6116), .Z(n5912) );
  AND U6116 ( .A(n310), .B(n6106), .Z(n6116) );
  XNOR U6117 ( .A(n6104), .B(n6115), .Z(n6106) );
  XNOR U6118 ( .A(n6117), .B(n6118), .Z(n310) );
  NOR U6119 ( .A(n6119), .B(n6120), .Z(n6118) );
  XNOR U6120 ( .A(n5920), .B(n6121), .Z(n6120) );
  IV U6121 ( .A(n6117), .Z(n6121) );
  AND U6122 ( .A(n6122), .B(n6123), .Z(n5920) );
  NOR U6123 ( .A(n6117), .B(n5919), .Z(n6119) );
  AND U6124 ( .A(n5993), .B(n5994), .Z(n5919) );
  IV U6125 ( .A(n6124), .Z(n5993) );
  XOR U6126 ( .A(n6111), .B(n6125), .Z(n6117) );
  AND U6127 ( .A(n6126), .B(n6114), .Z(n6125) );
  XNOR U6128 ( .A(n5965), .B(n6111), .Z(n6114) );
  XOR U6129 ( .A(n6127), .B(n6128), .Z(n5965) );
  AND U6130 ( .A(n313), .B(n6010), .Z(n6128) );
  XOR U6131 ( .A(n6008), .B(n6127), .Z(n6010) );
  XNOR U6132 ( .A(n6129), .B(n6111), .Z(n6126) );
  IV U6133 ( .A(n5926), .Z(n6129) );
  XOR U6134 ( .A(n6130), .B(n6131), .Z(n5926) );
  AND U6135 ( .A(n318), .B(n6132), .Z(n6131) );
  XOR U6136 ( .A(n6133), .B(n6134), .Z(n6111) );
  AND U6137 ( .A(n6135), .B(n6136), .Z(n6134) );
  XNOR U6138 ( .A(n5975), .B(n6133), .Z(n6136) );
  XOR U6139 ( .A(n6137), .B(n6138), .Z(n5975) );
  AND U6140 ( .A(n313), .B(n6036), .Z(n6138) );
  XOR U6141 ( .A(n6034), .B(n6137), .Z(n6036) );
  XOR U6142 ( .A(n6133), .B(n5935), .Z(n6135) );
  XOR U6143 ( .A(n6139), .B(n6140), .Z(n5935) );
  AND U6144 ( .A(n318), .B(n6141), .Z(n6140) );
  XOR U6145 ( .A(n6142), .B(n6143), .Z(n6133) );
  AND U6146 ( .A(n6144), .B(n6145), .Z(n6143) );
  XNOR U6147 ( .A(n6142), .B(n5983), .Z(n6145) );
  XOR U6148 ( .A(n6087), .B(n6146), .Z(n5983) );
  AND U6149 ( .A(n313), .B(n6147), .Z(n6146) );
  XOR U6150 ( .A(n6083), .B(n6087), .Z(n6147) );
  XNOR U6151 ( .A(n6148), .B(n6142), .Z(n6144) );
  IV U6152 ( .A(n5945), .Z(n6148) );
  XOR U6153 ( .A(n6149), .B(n6150), .Z(n5945) );
  AND U6154 ( .A(n318), .B(n6151), .Z(n6150) );
  AND U6155 ( .A(n6115), .B(n6104), .Z(n6142) );
  XNOR U6156 ( .A(n6152), .B(n6153), .Z(n6104) );
  AND U6157 ( .A(n313), .B(n6099), .Z(n6153) );
  XOR U6158 ( .A(n6154), .B(n6152), .Z(n6099) );
  XNOR U6159 ( .A(n6100), .B(n6155), .Z(n313) );
  NOR U6160 ( .A(n6102), .B(n6156), .Z(n6155) );
  XNOR U6161 ( .A(n6100), .B(n6124), .Z(n6156) );
  NOR U6162 ( .A(n6122), .B(n6123), .Z(n6124) );
  NOR U6163 ( .A(n6100), .B(n5994), .Z(n6102) );
  AND U6164 ( .A(n6008), .B(n6157), .Z(n5994) );
  XOR U6165 ( .A(n6158), .B(n6159), .Z(n6100) );
  AND U6166 ( .A(n6160), .B(n6161), .Z(n6159) );
  XNOR U6167 ( .A(n6008), .B(n6158), .Z(n6161) );
  XNOR U6168 ( .A(n6162), .B(n6163), .Z(n6008) );
  XOR U6169 ( .A(n6164), .B(n6157), .Z(n6163) );
  AND U6170 ( .A(n6034), .B(n6165), .Z(n6157) );
  AND U6171 ( .A(n6166), .B(n6167), .Z(n6164) );
  XOR U6172 ( .A(n6168), .B(n6162), .Z(n6166) );
  XOR U6173 ( .A(n6158), .B(n6127), .Z(n6160) );
  XOR U6174 ( .A(n6169), .B(n6170), .Z(n6127) );
  AND U6175 ( .A(n315), .B(n6132), .Z(n6170) );
  XOR U6176 ( .A(n6169), .B(n6130), .Z(n6132) );
  XOR U6177 ( .A(n6171), .B(n6172), .Z(n6158) );
  AND U6178 ( .A(n6173), .B(n6174), .Z(n6172) );
  XNOR U6179 ( .A(n6034), .B(n6171), .Z(n6174) );
  XOR U6180 ( .A(n6175), .B(n6167), .Z(n6034) );
  XNOR U6181 ( .A(n6176), .B(n6162), .Z(n6167) );
  XOR U6182 ( .A(n6177), .B(n6178), .Z(n6162) );
  AND U6183 ( .A(n6179), .B(n6180), .Z(n6178) );
  XOR U6184 ( .A(n6181), .B(n6177), .Z(n6179) );
  XNOR U6185 ( .A(n6182), .B(n6183), .Z(n6176) );
  AND U6186 ( .A(n6184), .B(n6185), .Z(n6183) );
  XOR U6187 ( .A(n6182), .B(n6186), .Z(n6184) );
  XNOR U6188 ( .A(n6168), .B(n6165), .Z(n6175) );
  AND U6189 ( .A(n6083), .B(n6187), .Z(n6165) );
  XOR U6190 ( .A(n6188), .B(n6189), .Z(n6168) );
  AND U6191 ( .A(n6190), .B(n6191), .Z(n6189) );
  XOR U6192 ( .A(n6188), .B(n6192), .Z(n6190) );
  XOR U6193 ( .A(n6171), .B(n6137), .Z(n6173) );
  XOR U6194 ( .A(n6193), .B(n6194), .Z(n6137) );
  AND U6195 ( .A(n315), .B(n6141), .Z(n6194) );
  XOR U6196 ( .A(n6193), .B(n6139), .Z(n6141) );
  XOR U6197 ( .A(n6195), .B(n6196), .Z(n6171) );
  AND U6198 ( .A(n6197), .B(n6198), .Z(n6196) );
  XNOR U6199 ( .A(n6195), .B(n6083), .Z(n6198) );
  IV U6200 ( .A(n6086), .Z(n6083) );
  XNOR U6201 ( .A(n6199), .B(n6180), .Z(n6086) );
  XNOR U6202 ( .A(n6200), .B(n6186), .Z(n6180) );
  XOR U6203 ( .A(n6201), .B(n6202), .Z(n6186) );
  NOR U6204 ( .A(n6203), .B(n6204), .Z(n6202) );
  XNOR U6205 ( .A(n6201), .B(n6205), .Z(n6203) );
  XNOR U6206 ( .A(n6185), .B(n6177), .Z(n6200) );
  XOR U6207 ( .A(n6206), .B(n6207), .Z(n6177) );
  AND U6208 ( .A(n6208), .B(n6209), .Z(n6207) );
  XNOR U6209 ( .A(n6206), .B(n6210), .Z(n6208) );
  XNOR U6210 ( .A(n6211), .B(n6182), .Z(n6185) );
  XOR U6211 ( .A(n6212), .B(n6213), .Z(n6182) );
  AND U6212 ( .A(n6214), .B(n6215), .Z(n6213) );
  XOR U6213 ( .A(n6212), .B(n6216), .Z(n6214) );
  XNOR U6214 ( .A(n6217), .B(n6218), .Z(n6211) );
  NOR U6215 ( .A(n6219), .B(n6220), .Z(n6218) );
  XOR U6216 ( .A(n6217), .B(n6221), .Z(n6219) );
  XNOR U6217 ( .A(n6181), .B(n6187), .Z(n6199) );
  AND U6218 ( .A(n6154), .B(n6222), .Z(n6187) );
  IV U6219 ( .A(n6097), .Z(n6154) );
  XOR U6220 ( .A(n6192), .B(n6191), .Z(n6181) );
  XNOR U6221 ( .A(n6223), .B(n6188), .Z(n6191) );
  XOR U6222 ( .A(n6224), .B(n6225), .Z(n6188) );
  AND U6223 ( .A(n6226), .B(n6227), .Z(n6225) );
  XOR U6224 ( .A(n6224), .B(n6228), .Z(n6226) );
  XNOR U6225 ( .A(n6229), .B(n6230), .Z(n6223) );
  NOR U6226 ( .A(n6231), .B(n6232), .Z(n6230) );
  XNOR U6227 ( .A(n6229), .B(n6233), .Z(n6231) );
  XOR U6228 ( .A(n6234), .B(n6235), .Z(n6192) );
  NOR U6229 ( .A(n6236), .B(n6237), .Z(n6235) );
  XNOR U6230 ( .A(n6234), .B(n6238), .Z(n6236) );
  XOR U6231 ( .A(n6087), .B(n6195), .Z(n6197) );
  XOR U6232 ( .A(n6239), .B(n6240), .Z(n6087) );
  AND U6233 ( .A(n315), .B(n6151), .Z(n6240) );
  XOR U6234 ( .A(n6239), .B(n6149), .Z(n6151) );
  AND U6235 ( .A(n6152), .B(n6097), .Z(n6195) );
  XNOR U6236 ( .A(n6241), .B(n6222), .Z(n6097) );
  XOR U6237 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(
        p_input[256]), .Z(n6222) );
  XOR U6238 ( .A(n6210), .B(n6209), .Z(n6241) );
  XNOR U6239 ( .A(n6242), .B(n6216), .Z(n6209) );
  XNOR U6240 ( .A(n6205), .B(n6204), .Z(n6216) );
  XOR U6241 ( .A(n6243), .B(n6201), .Z(n6204) );
  XNOR U6242 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n3619), 
        .Z(n6201) );
  XOR U6243 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n3382), 
        .Z(n6243) );
  XOR U6244 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(
        p_input[268]), .Z(n6205) );
  XNOR U6245 ( .A(n6215), .B(n6206), .Z(n6242) );
  XNOR U6246 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n3849), 
        .Z(n6206) );
  XOR U6247 ( .A(n6244), .B(n6221), .Z(n6215) );
  XNOR U6248 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(
        p_input[271]), .Z(n6221) );
  XOR U6249 ( .A(n6212), .B(n6220), .Z(n6244) );
  XOR U6250 ( .A(n6245), .B(n6217), .Z(n6220) );
  XOR U6251 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(
        p_input[269]), .Z(n6217) );
  XOR U6252 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n3387), 
        .Z(n6245) );
  XNOR U6253 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n3388), 
        .Z(n6212) );
  IV U6254 ( .A(p_input[265]), .Z(n3388) );
  XNOR U6255 ( .A(n6228), .B(n6227), .Z(n6210) );
  XNOR U6256 ( .A(n6246), .B(n6233), .Z(n6227) );
  XOR U6257 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(
        p_input[264]), .Z(n6233) );
  XOR U6258 ( .A(n6224), .B(n6232), .Z(n6246) );
  XOR U6259 ( .A(n6247), .B(n6229), .Z(n6232) );
  XOR U6260 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(
        p_input[262]), .Z(n6229) );
  XOR U6261 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n3625), 
        .Z(n6247) );
  XNOR U6262 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n3391), 
        .Z(n6224) );
  XNOR U6263 ( .A(n6238), .B(n6237), .Z(n6228) );
  XOR U6264 ( .A(n6248), .B(n6234), .Z(n6237) );
  XOR U6265 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(
        p_input[259]), .Z(n6234) );
  XOR U6266 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n3627), 
        .Z(n6248) );
  XOR U6267 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(
        p_input[261]), .Z(n6238) );
  XNOR U6268 ( .A(n6249), .B(n6250), .Z(n6152) );
  AND U6269 ( .A(n315), .B(n6251), .Z(n6250) );
  XNOR U6270 ( .A(n6252), .B(n6253), .Z(n315) );
  NOR U6271 ( .A(n6254), .B(n6255), .Z(n6253) );
  XOR U6272 ( .A(n6123), .B(n6252), .Z(n6255) );
  NOR U6273 ( .A(n6252), .B(n6122), .Z(n6254) );
  XOR U6274 ( .A(n6256), .B(n6257), .Z(n6252) );
  AND U6275 ( .A(n6258), .B(n6259), .Z(n6257) );
  XOR U6276 ( .A(n6256), .B(n6130), .Z(n6258) );
  XOR U6277 ( .A(n6260), .B(n6261), .Z(n6115) );
  AND U6278 ( .A(n318), .B(n6251), .Z(n6261) );
  XOR U6279 ( .A(n6262), .B(n6260), .Z(n6251) );
  XNOR U6280 ( .A(n6263), .B(n6264), .Z(n318) );
  NOR U6281 ( .A(n6265), .B(n6266), .Z(n6264) );
  XNOR U6282 ( .A(n6123), .B(n6267), .Z(n6266) );
  IV U6283 ( .A(n6263), .Z(n6267) );
  AND U6284 ( .A(n6130), .B(n6268), .Z(n6123) );
  NOR U6285 ( .A(n6263), .B(n6122), .Z(n6265) );
  AND U6286 ( .A(n6169), .B(n6269), .Z(n6122) );
  XOR U6287 ( .A(n6256), .B(n6270), .Z(n6263) );
  AND U6288 ( .A(n6271), .B(n6259), .Z(n6270) );
  XNOR U6289 ( .A(n6169), .B(n6256), .Z(n6259) );
  XNOR U6290 ( .A(n6272), .B(n6273), .Z(n6169) );
  XOR U6291 ( .A(n6274), .B(n6269), .Z(n6273) );
  AND U6292 ( .A(n6193), .B(n6275), .Z(n6269) );
  AND U6293 ( .A(n6276), .B(n6277), .Z(n6274) );
  XOR U6294 ( .A(n6278), .B(n6272), .Z(n6276) );
  XNOR U6295 ( .A(n6279), .B(n6256), .Z(n6271) );
  IV U6296 ( .A(n6130), .Z(n6279) );
  XNOR U6297 ( .A(n6280), .B(n6281), .Z(n6130) );
  XOR U6298 ( .A(n6282), .B(n6268), .Z(n6281) );
  AND U6299 ( .A(n6139), .B(n6283), .Z(n6268) );
  AND U6300 ( .A(n6284), .B(n6285), .Z(n6282) );
  XNOR U6301 ( .A(n6280), .B(n6286), .Z(n6284) );
  XOR U6302 ( .A(n6287), .B(n6288), .Z(n6256) );
  AND U6303 ( .A(n6289), .B(n6290), .Z(n6288) );
  XNOR U6304 ( .A(n6193), .B(n6287), .Z(n6290) );
  XOR U6305 ( .A(n6291), .B(n6277), .Z(n6193) );
  XNOR U6306 ( .A(n6292), .B(n6272), .Z(n6277) );
  XOR U6307 ( .A(n6293), .B(n6294), .Z(n6272) );
  AND U6308 ( .A(n6295), .B(n6296), .Z(n6294) );
  XOR U6309 ( .A(n6297), .B(n6293), .Z(n6295) );
  XNOR U6310 ( .A(n6298), .B(n6299), .Z(n6292) );
  AND U6311 ( .A(n6300), .B(n6301), .Z(n6299) );
  XOR U6312 ( .A(n6298), .B(n6302), .Z(n6300) );
  XNOR U6313 ( .A(n6278), .B(n6275), .Z(n6291) );
  AND U6314 ( .A(n6239), .B(n6303), .Z(n6275) );
  XOR U6315 ( .A(n6304), .B(n6305), .Z(n6278) );
  AND U6316 ( .A(n6306), .B(n6307), .Z(n6305) );
  XOR U6317 ( .A(n6304), .B(n6308), .Z(n6306) );
  XOR U6318 ( .A(n6287), .B(n6139), .Z(n6289) );
  XNOR U6319 ( .A(n6309), .B(n6286), .Z(n6139) );
  XNOR U6320 ( .A(n6310), .B(n6311), .Z(n6286) );
  AND U6321 ( .A(n6312), .B(n6313), .Z(n6311) );
  XOR U6322 ( .A(n6310), .B(n6314), .Z(n6312) );
  XNOR U6323 ( .A(n6285), .B(n6283), .Z(n6309) );
  AND U6324 ( .A(n6149), .B(n6315), .Z(n6283) );
  XNOR U6325 ( .A(n6316), .B(n6280), .Z(n6285) );
  XOR U6326 ( .A(n6317), .B(n6318), .Z(n6280) );
  AND U6327 ( .A(n6319), .B(n6320), .Z(n6318) );
  XOR U6328 ( .A(n6317), .B(n6321), .Z(n6319) );
  XNOR U6329 ( .A(n6322), .B(n6323), .Z(n6316) );
  AND U6330 ( .A(n6324), .B(n6325), .Z(n6323) );
  XNOR U6331 ( .A(n6322), .B(n6326), .Z(n6324) );
  XOR U6332 ( .A(n6327), .B(n6328), .Z(n6287) );
  AND U6333 ( .A(n6329), .B(n6330), .Z(n6328) );
  XNOR U6334 ( .A(n6327), .B(n6239), .Z(n6330) );
  XOR U6335 ( .A(n6331), .B(n6296), .Z(n6239) );
  XNOR U6336 ( .A(n6332), .B(n6302), .Z(n6296) );
  XOR U6337 ( .A(n6333), .B(n6334), .Z(n6302) );
  NOR U6338 ( .A(n6335), .B(n6336), .Z(n6334) );
  XNOR U6339 ( .A(n6333), .B(n6337), .Z(n6335) );
  XNOR U6340 ( .A(n6301), .B(n6293), .Z(n6332) );
  XOR U6341 ( .A(n6338), .B(n6339), .Z(n6293) );
  AND U6342 ( .A(n6340), .B(n6341), .Z(n6339) );
  XNOR U6343 ( .A(n6338), .B(n6342), .Z(n6340) );
  XNOR U6344 ( .A(n6343), .B(n6298), .Z(n6301) );
  XOR U6345 ( .A(n6344), .B(n6345), .Z(n6298) );
  AND U6346 ( .A(n6346), .B(n6347), .Z(n6345) );
  XOR U6347 ( .A(n6344), .B(n6348), .Z(n6346) );
  XNOR U6348 ( .A(n6349), .B(n6350), .Z(n6343) );
  NOR U6349 ( .A(n6351), .B(n6352), .Z(n6350) );
  XOR U6350 ( .A(n6349), .B(n6353), .Z(n6351) );
  XNOR U6351 ( .A(n6297), .B(n6303), .Z(n6331) );
  AND U6352 ( .A(n6262), .B(n6354), .Z(n6303) );
  IV U6353 ( .A(n6249), .Z(n6262) );
  XOR U6354 ( .A(n6308), .B(n6307), .Z(n6297) );
  XNOR U6355 ( .A(n6355), .B(n6304), .Z(n6307) );
  XOR U6356 ( .A(n6356), .B(n6357), .Z(n6304) );
  AND U6357 ( .A(n6358), .B(n6359), .Z(n6357) );
  XOR U6358 ( .A(n6356), .B(n6360), .Z(n6358) );
  XNOR U6359 ( .A(n6361), .B(n6362), .Z(n6355) );
  NOR U6360 ( .A(n6363), .B(n6364), .Z(n6362) );
  XNOR U6361 ( .A(n6361), .B(n6365), .Z(n6363) );
  XOR U6362 ( .A(n6366), .B(n6367), .Z(n6308) );
  NOR U6363 ( .A(n6368), .B(n6369), .Z(n6367) );
  XNOR U6364 ( .A(n6366), .B(n6370), .Z(n6368) );
  XNOR U6365 ( .A(n6371), .B(n6327), .Z(n6329) );
  IV U6366 ( .A(n6149), .Z(n6371) );
  XOR U6367 ( .A(n6372), .B(n6321), .Z(n6149) );
  XOR U6368 ( .A(n6314), .B(n6313), .Z(n6321) );
  XNOR U6369 ( .A(n6373), .B(n6310), .Z(n6313) );
  XOR U6370 ( .A(n6374), .B(n6375), .Z(n6310) );
  AND U6371 ( .A(n6376), .B(n6377), .Z(n6375) );
  XOR U6372 ( .A(n6374), .B(n6378), .Z(n6376) );
  XNOR U6373 ( .A(n6379), .B(n6380), .Z(n6373) );
  NOR U6374 ( .A(n6381), .B(n6382), .Z(n6380) );
  XNOR U6375 ( .A(n6379), .B(n6383), .Z(n6381) );
  XOR U6376 ( .A(n6384), .B(n6385), .Z(n6314) );
  NOR U6377 ( .A(n6386), .B(n6387), .Z(n6385) );
  XNOR U6378 ( .A(n6384), .B(n6388), .Z(n6386) );
  XNOR U6379 ( .A(n6320), .B(n6315), .Z(n6372) );
  AND U6380 ( .A(n6260), .B(n6389), .Z(n6315) );
  XOR U6381 ( .A(n6390), .B(n6326), .Z(n6320) );
  XNOR U6382 ( .A(n6391), .B(n6392), .Z(n6326) );
  NOR U6383 ( .A(n6393), .B(n6394), .Z(n6392) );
  XNOR U6384 ( .A(n6391), .B(n6395), .Z(n6393) );
  XNOR U6385 ( .A(n6325), .B(n6317), .Z(n6390) );
  XOR U6386 ( .A(n6396), .B(n6397), .Z(n6317) );
  AND U6387 ( .A(n6398), .B(n6399), .Z(n6397) );
  XOR U6388 ( .A(n6396), .B(n6400), .Z(n6398) );
  XNOR U6389 ( .A(n6401), .B(n6322), .Z(n6325) );
  XOR U6390 ( .A(n6402), .B(n6403), .Z(n6322) );
  AND U6391 ( .A(n6404), .B(n6405), .Z(n6403) );
  XOR U6392 ( .A(n6402), .B(n6406), .Z(n6404) );
  XNOR U6393 ( .A(n6407), .B(n6408), .Z(n6401) );
  NOR U6394 ( .A(n6409), .B(n6410), .Z(n6408) );
  XOR U6395 ( .A(n6407), .B(n6411), .Z(n6409) );
  AND U6396 ( .A(n6260), .B(n6249), .Z(n6327) );
  XNOR U6397 ( .A(n6412), .B(n6354), .Z(n6249) );
  XOR U6398 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(
        p_input[256]), .Z(n6354) );
  XOR U6399 ( .A(n6342), .B(n6341), .Z(n6412) );
  XNOR U6400 ( .A(n6413), .B(n6348), .Z(n6341) );
  XNOR U6401 ( .A(n6337), .B(n6336), .Z(n6348) );
  XOR U6402 ( .A(n6414), .B(n6333), .Z(n6336) );
  XNOR U6403 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(n3619), 
        .Z(n6333) );
  XOR U6404 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n3382), 
        .Z(n6414) );
  XOR U6405 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(
        p_input[268]), .Z(n6337) );
  XNOR U6406 ( .A(n6347), .B(n6338), .Z(n6413) );
  XNOR U6407 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(n3849), 
        .Z(n6338) );
  XOR U6408 ( .A(n6415), .B(n6353), .Z(n6347) );
  XNOR U6409 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(
        p_input[271]), .Z(n6353) );
  XOR U6410 ( .A(n6344), .B(n6352), .Z(n6415) );
  XOR U6411 ( .A(n6416), .B(n6349), .Z(n6352) );
  XOR U6412 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(
        p_input[269]), .Z(n6349) );
  XOR U6413 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(n3387), 
        .Z(n6416) );
  XNOR U6414 ( .A(n320), .B(p_input[265]), .Z(n6344) );
  IV U6415 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .Z(n320) );
  XNOR U6416 ( .A(n6360), .B(n6359), .Z(n6342) );
  XNOR U6417 ( .A(n6417), .B(n6365), .Z(n6359) );
  XNOR U6418 ( .A(n511), .B(p_input[264]), .Z(n6365) );
  IV U6419 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .Z(n511) );
  XOR U6420 ( .A(n6356), .B(n6364), .Z(n6417) );
  XOR U6421 ( .A(n6418), .B(n6361), .Z(n6364) );
  XNOR U6422 ( .A(n893), .B(p_input[262]), .Z(n6361) );
  IV U6423 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .Z(n893) );
  XOR U6424 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(n3625), 
        .Z(n6418) );
  XNOR U6425 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .B(n3391), 
        .Z(n6356) );
  XNOR U6426 ( .A(n6370), .B(n6369), .Z(n6360) );
  XOR U6427 ( .A(n6419), .B(n6366), .Z(n6369) );
  XNOR U6428 ( .A(n1468), .B(p_input[259]), .Z(n6366) );
  IV U6429 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .Z(n1468) );
  XOR U6430 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(n3627), 
        .Z(n6419) );
  XNOR U6431 ( .A(n1084), .B(p_input[261]), .Z(n6370) );
  IV U6432 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .Z(n1084) );
  XOR U6433 ( .A(n6420), .B(n6400), .Z(n6260) );
  XOR U6434 ( .A(n6378), .B(n6377), .Z(n6400) );
  XNOR U6435 ( .A(n6421), .B(n6383), .Z(n6377) );
  XNOR U6436 ( .A(n510), .B(p_input[264]), .Z(n6383) );
  IV U6437 ( .A(\knn_comb_/min_val_out[0][8] ), .Z(n510) );
  XOR U6438 ( .A(n6374), .B(n6382), .Z(n6421) );
  XOR U6439 ( .A(n6422), .B(n6379), .Z(n6382) );
  XNOR U6440 ( .A(n892), .B(p_input[262]), .Z(n6379) );
  IV U6441 ( .A(\knn_comb_/min_val_out[0][6] ), .Z(n892) );
  XOR U6442 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n3625), .Z(n6422) );
  IV U6443 ( .A(p_input[263]), .Z(n3625) );
  XNOR U6444 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n3391), .Z(n6374) );
  IV U6445 ( .A(p_input[258]), .Z(n3391) );
  XNOR U6446 ( .A(n6388), .B(n6387), .Z(n6378) );
  XOR U6447 ( .A(n6423), .B(n6384), .Z(n6387) );
  XNOR U6448 ( .A(n1467), .B(p_input[259]), .Z(n6384) );
  IV U6449 ( .A(\knn_comb_/min_val_out[0][3] ), .Z(n1467) );
  XOR U6450 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n3627), .Z(n6423) );
  IV U6451 ( .A(p_input[260]), .Z(n3627) );
  XNOR U6452 ( .A(n1083), .B(p_input[261]), .Z(n6388) );
  IV U6453 ( .A(\knn_comb_/min_val_out[0][5] ), .Z(n1083) );
  XNOR U6454 ( .A(n6399), .B(n6389), .Z(n6420) );
  XOR U6455 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[256]), .Z(n6389)
         );
  XNOR U6456 ( .A(n6424), .B(n6406), .Z(n6399) );
  XNOR U6457 ( .A(n6395), .B(n6394), .Z(n6406) );
  XOR U6458 ( .A(n6425), .B(n6391), .Z(n6394) );
  XNOR U6459 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n3619), .Z(n6391) );
  IV U6460 ( .A(p_input[266]), .Z(n3619) );
  XOR U6461 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n3382), .Z(n6425) );
  IV U6462 ( .A(p_input[267]), .Z(n3382) );
  XOR U6463 ( .A(\knn_comb_/min_val_out[0][12] ), .B(p_input[268]), .Z(n6395)
         );
  XNOR U6464 ( .A(n6405), .B(n6396), .Z(n6424) );
  XNOR U6465 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n3849), .Z(n6396) );
  IV U6466 ( .A(p_input[257]), .Z(n3849) );
  XOR U6467 ( .A(n6426), .B(n6411), .Z(n6405) );
  XNOR U6468 ( .A(\knn_comb_/min_val_out[0][15] ), .B(p_input[271]), .Z(n6411)
         );
  XOR U6469 ( .A(n6402), .B(n6410), .Z(n6426) );
  XOR U6470 ( .A(n6427), .B(n6407), .Z(n6410) );
  XOR U6471 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[269]), .Z(n6407)
         );
  XOR U6472 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n3387), .Z(n6427) );
  IV U6473 ( .A(p_input[270]), .Z(n3387) );
  XNOR U6474 ( .A(n319), .B(p_input[265]), .Z(n6402) );
  IV U6475 ( .A(\knn_comb_/min_val_out[0][9] ), .Z(n319) );
endmodule

