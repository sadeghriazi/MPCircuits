
module knn_comb_BMR_W32_K2_N16 ( p_input, o );
  input [543:0] p_input;
  output [63:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/min_val_out[0][16] , \knn_comb_/min_val_out[0][17] ,
         \knn_comb_/min_val_out[0][18] , \knn_comb_/min_val_out[0][19] ,
         \knn_comb_/min_val_out[0][20] , \knn_comb_/min_val_out[0][21] ,
         \knn_comb_/min_val_out[0][22] , \knn_comb_/min_val_out[0][23] ,
         \knn_comb_/min_val_out[0][24] , \knn_comb_/min_val_out[0][25] ,
         \knn_comb_/min_val_out[0][26] , \knn_comb_/min_val_out[0][27] ,
         \knn_comb_/min_val_out[0][28] , \knn_comb_/min_val_out[0][29] ,
         \knn_comb_/min_val_out[0][30] , \knn_comb_/min_val_out[0][31] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][31] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123;
  assign \knn_comb_/min_val_out[0][0]  = p_input[480];
  assign \knn_comb_/min_val_out[0][1]  = p_input[481];
  assign \knn_comb_/min_val_out[0][2]  = p_input[482];
  assign \knn_comb_/min_val_out[0][3]  = p_input[483];
  assign \knn_comb_/min_val_out[0][4]  = p_input[484];
  assign \knn_comb_/min_val_out[0][5]  = p_input[485];
  assign \knn_comb_/min_val_out[0][6]  = p_input[486];
  assign \knn_comb_/min_val_out[0][7]  = p_input[487];
  assign \knn_comb_/min_val_out[0][8]  = p_input[488];
  assign \knn_comb_/min_val_out[0][9]  = p_input[489];
  assign \knn_comb_/min_val_out[0][10]  = p_input[490];
  assign \knn_comb_/min_val_out[0][11]  = p_input[491];
  assign \knn_comb_/min_val_out[0][12]  = p_input[492];
  assign \knn_comb_/min_val_out[0][13]  = p_input[493];
  assign \knn_comb_/min_val_out[0][14]  = p_input[494];
  assign \knn_comb_/min_val_out[0][15]  = p_input[495];
  assign \knn_comb_/min_val_out[0][16]  = p_input[496];
  assign \knn_comb_/min_val_out[0][17]  = p_input[497];
  assign \knn_comb_/min_val_out[0][18]  = p_input[498];
  assign \knn_comb_/min_val_out[0][19]  = p_input[499];
  assign \knn_comb_/min_val_out[0][20]  = p_input[500];
  assign \knn_comb_/min_val_out[0][21]  = p_input[501];
  assign \knn_comb_/min_val_out[0][22]  = p_input[502];
  assign \knn_comb_/min_val_out[0][23]  = p_input[503];
  assign \knn_comb_/min_val_out[0][24]  = p_input[504];
  assign \knn_comb_/min_val_out[0][25]  = p_input[505];
  assign \knn_comb_/min_val_out[0][26]  = p_input[506];
  assign \knn_comb_/min_val_out[0][27]  = p_input[507];
  assign \knn_comb_/min_val_out[0][28]  = p_input[508];
  assign \knn_comb_/min_val_out[0][29]  = p_input[509];
  assign \knn_comb_/min_val_out[0][30]  = p_input[510];
  assign \knn_comb_/min_val_out[0][31]  = p_input[511];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][0]  = p_input[448];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][1]  = p_input[449];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][2]  = p_input[450];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][3]  = p_input[451];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][4]  = p_input[452];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][5]  = p_input[453];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][6]  = p_input[454];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][7]  = p_input[455];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][8]  = p_input[456];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][9]  = p_input[457];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][10]  = p_input[458];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][11]  = p_input[459];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][12]  = p_input[460];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][13]  = p_input[461];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][14]  = p_input[462];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][15]  = p_input[463];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][16]  = p_input[464];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][17]  = p_input[465];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][18]  = p_input[466];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][19]  = p_input[467];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][20]  = p_input[468];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][21]  = p_input[469];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][22]  = p_input[470];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][23]  = p_input[471];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][24]  = p_input[472];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][25]  = p_input[473];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][26]  = p_input[474];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][27]  = p_input[475];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][28]  = p_input[476];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][29]  = p_input[477];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][30]  = p_input[478];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][31]  = p_input[479];

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  XOR U2 ( .A(n3), .B(n4), .Z(o[8]) );
  XOR U3 ( .A(n5), .B(n6), .Z(o[7]) );
  XOR U4 ( .A(n7), .B(n8), .Z(o[6]) );
  XOR U5 ( .A(n9), .B(n10), .Z(o[63]) );
  XOR U6 ( .A(n11), .B(n12), .Z(o[62]) );
  XOR U7 ( .A(n13), .B(n14), .Z(o[61]) );
  XOR U8 ( .A(n15), .B(n16), .Z(o[60]) );
  XOR U9 ( .A(n17), .B(n18), .Z(o[5]) );
  XOR U10 ( .A(n19), .B(n20), .Z(o[59]) );
  XOR U11 ( .A(n21), .B(n22), .Z(o[58]) );
  XOR U12 ( .A(n23), .B(n24), .Z(o[57]) );
  XOR U13 ( .A(n25), .B(n26), .Z(o[56]) );
  XOR U14 ( .A(n27), .B(n28), .Z(o[55]) );
  XOR U15 ( .A(n29), .B(n30), .Z(o[54]) );
  XOR U16 ( .A(n31), .B(n32), .Z(o[53]) );
  XOR U17 ( .A(n33), .B(n34), .Z(o[52]) );
  XOR U18 ( .A(n35), .B(n36), .Z(o[51]) );
  XOR U19 ( .A(n37), .B(n38), .Z(o[50]) );
  XOR U20 ( .A(n39), .B(n40), .Z(o[4]) );
  XOR U21 ( .A(n41), .B(n42), .Z(o[49]) );
  XOR U22 ( .A(n43), .B(n44), .Z(o[48]) );
  XOR U23 ( .A(n45), .B(n46), .Z(o[47]) );
  XOR U24 ( .A(n47), .B(n48), .Z(o[46]) );
  XOR U25 ( .A(n49), .B(n50), .Z(o[45]) );
  XOR U26 ( .A(n51), .B(n52), .Z(o[44]) );
  XOR U27 ( .A(n53), .B(n54), .Z(o[43]) );
  XOR U28 ( .A(n55), .B(n56), .Z(o[42]) );
  XOR U29 ( .A(n1), .B(n57), .Z(o[41]) );
  AND U30 ( .A(n58), .B(n59), .Z(n1) );
  XOR U31 ( .A(n2), .B(n57), .Z(n59) );
  XOR U32 ( .A(n60), .B(n61), .Z(n57) );
  AND U33 ( .A(n62), .B(n63), .Z(n61) );
  XOR U34 ( .A(p_input[9]), .B(n60), .Z(n63) );
  XOR U35 ( .A(n64), .B(n65), .Z(n60) );
  AND U36 ( .A(n66), .B(n67), .Z(n65) );
  XOR U37 ( .A(n68), .B(n69), .Z(n2) );
  AND U38 ( .A(n70), .B(n67), .Z(n69) );
  XNOR U39 ( .A(n71), .B(n64), .Z(n67) );
  XOR U40 ( .A(n72), .B(n73), .Z(n64) );
  AND U41 ( .A(n74), .B(n75), .Z(n73) );
  XOR U42 ( .A(p_input[41]), .B(n72), .Z(n75) );
  XOR U43 ( .A(n76), .B(n77), .Z(n72) );
  AND U44 ( .A(n78), .B(n79), .Z(n77) );
  IV U45 ( .A(n68), .Z(n71) );
  XNOR U46 ( .A(n80), .B(n81), .Z(n68) );
  AND U47 ( .A(n82), .B(n79), .Z(n81) );
  XNOR U48 ( .A(n80), .B(n76), .Z(n79) );
  XOR U49 ( .A(n83), .B(n84), .Z(n76) );
  AND U50 ( .A(n85), .B(n86), .Z(n84) );
  XOR U51 ( .A(p_input[73]), .B(n83), .Z(n86) );
  XOR U52 ( .A(n87), .B(n88), .Z(n83) );
  AND U53 ( .A(n89), .B(n90), .Z(n88) );
  XOR U54 ( .A(n91), .B(n92), .Z(n80) );
  AND U55 ( .A(n93), .B(n90), .Z(n92) );
  XNOR U56 ( .A(n91), .B(n87), .Z(n90) );
  XOR U57 ( .A(n94), .B(n95), .Z(n87) );
  AND U58 ( .A(n96), .B(n97), .Z(n95) );
  XOR U59 ( .A(p_input[105]), .B(n94), .Z(n97) );
  XOR U60 ( .A(n98), .B(n99), .Z(n94) );
  AND U61 ( .A(n100), .B(n101), .Z(n99) );
  XOR U62 ( .A(n102), .B(n103), .Z(n91) );
  AND U63 ( .A(n104), .B(n101), .Z(n103) );
  XNOR U64 ( .A(n102), .B(n98), .Z(n101) );
  XOR U65 ( .A(n105), .B(n106), .Z(n98) );
  AND U66 ( .A(n107), .B(n108), .Z(n106) );
  XOR U67 ( .A(p_input[137]), .B(n105), .Z(n108) );
  XOR U68 ( .A(n109), .B(n110), .Z(n105) );
  AND U69 ( .A(n111), .B(n112), .Z(n110) );
  XOR U70 ( .A(n113), .B(n114), .Z(n102) );
  AND U71 ( .A(n115), .B(n112), .Z(n114) );
  XNOR U72 ( .A(n113), .B(n109), .Z(n112) );
  XOR U73 ( .A(n116), .B(n117), .Z(n109) );
  AND U74 ( .A(n118), .B(n119), .Z(n117) );
  XOR U75 ( .A(p_input[169]), .B(n116), .Z(n119) );
  XOR U76 ( .A(n120), .B(n121), .Z(n116) );
  AND U77 ( .A(n122), .B(n123), .Z(n121) );
  XOR U78 ( .A(n124), .B(n125), .Z(n113) );
  AND U79 ( .A(n126), .B(n123), .Z(n125) );
  XNOR U80 ( .A(n124), .B(n120), .Z(n123) );
  XOR U81 ( .A(n127), .B(n128), .Z(n120) );
  AND U82 ( .A(n129), .B(n130), .Z(n128) );
  XOR U83 ( .A(p_input[201]), .B(n127), .Z(n130) );
  XOR U84 ( .A(n131), .B(n132), .Z(n127) );
  AND U85 ( .A(n133), .B(n134), .Z(n132) );
  XOR U86 ( .A(n135), .B(n136), .Z(n124) );
  AND U87 ( .A(n137), .B(n134), .Z(n136) );
  XNOR U88 ( .A(n135), .B(n131), .Z(n134) );
  XOR U89 ( .A(n138), .B(n139), .Z(n131) );
  AND U90 ( .A(n140), .B(n141), .Z(n139) );
  XOR U91 ( .A(p_input[233]), .B(n138), .Z(n141) );
  XOR U92 ( .A(n142), .B(n143), .Z(n138) );
  AND U93 ( .A(n144), .B(n145), .Z(n143) );
  XOR U94 ( .A(n146), .B(n147), .Z(n135) );
  AND U95 ( .A(n148), .B(n145), .Z(n147) );
  XNOR U96 ( .A(n146), .B(n142), .Z(n145) );
  XOR U97 ( .A(n149), .B(n150), .Z(n142) );
  AND U98 ( .A(n151), .B(n152), .Z(n150) );
  XOR U99 ( .A(p_input[265]), .B(n149), .Z(n152) );
  XOR U100 ( .A(n153), .B(n154), .Z(n149) );
  AND U101 ( .A(n155), .B(n156), .Z(n154) );
  XOR U102 ( .A(n157), .B(n158), .Z(n146) );
  AND U103 ( .A(n159), .B(n156), .Z(n158) );
  XNOR U104 ( .A(n157), .B(n153), .Z(n156) );
  XOR U105 ( .A(n160), .B(n161), .Z(n153) );
  AND U106 ( .A(n162), .B(n163), .Z(n161) );
  XOR U107 ( .A(p_input[297]), .B(n160), .Z(n163) );
  XOR U108 ( .A(n164), .B(n165), .Z(n160) );
  AND U109 ( .A(n166), .B(n167), .Z(n165) );
  XOR U110 ( .A(n168), .B(n169), .Z(n157) );
  AND U111 ( .A(n170), .B(n167), .Z(n169) );
  XNOR U112 ( .A(n168), .B(n164), .Z(n167) );
  XOR U113 ( .A(n171), .B(n172), .Z(n164) );
  AND U114 ( .A(n173), .B(n174), .Z(n172) );
  XOR U115 ( .A(p_input[329]), .B(n171), .Z(n174) );
  XOR U116 ( .A(n175), .B(n176), .Z(n171) );
  AND U117 ( .A(n177), .B(n178), .Z(n176) );
  XOR U118 ( .A(n179), .B(n180), .Z(n168) );
  AND U119 ( .A(n181), .B(n178), .Z(n180) );
  XNOR U120 ( .A(n179), .B(n175), .Z(n178) );
  XOR U121 ( .A(n182), .B(n183), .Z(n175) );
  AND U122 ( .A(n184), .B(n185), .Z(n183) );
  XOR U123 ( .A(p_input[361]), .B(n182), .Z(n185) );
  XOR U124 ( .A(n186), .B(n187), .Z(n182) );
  AND U125 ( .A(n188), .B(n189), .Z(n187) );
  XOR U126 ( .A(n190), .B(n191), .Z(n179) );
  AND U127 ( .A(n192), .B(n189), .Z(n191) );
  XNOR U128 ( .A(n190), .B(n186), .Z(n189) );
  XOR U129 ( .A(n193), .B(n194), .Z(n186) );
  AND U130 ( .A(n195), .B(n196), .Z(n194) );
  XOR U131 ( .A(p_input[393]), .B(n193), .Z(n196) );
  XOR U132 ( .A(n197), .B(n198), .Z(n193) );
  AND U133 ( .A(n199), .B(n200), .Z(n198) );
  XOR U134 ( .A(n201), .B(n202), .Z(n190) );
  AND U135 ( .A(n203), .B(n200), .Z(n202) );
  XNOR U136 ( .A(n201), .B(n197), .Z(n200) );
  XOR U137 ( .A(n204), .B(n205), .Z(n197) );
  AND U138 ( .A(n206), .B(n207), .Z(n205) );
  XOR U139 ( .A(p_input[425]), .B(n204), .Z(n207) );
  XNOR U140 ( .A(n208), .B(n209), .Z(n204) );
  AND U141 ( .A(n210), .B(n211), .Z(n209) );
  XNOR U142 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n212), .Z(n201) );
  AND U143 ( .A(n213), .B(n211), .Z(n212) );
  XOR U144 ( .A(n214), .B(n208), .Z(n211) );
  XOR U145 ( .A(n3), .B(n215), .Z(o[40]) );
  AND U146 ( .A(n58), .B(n216), .Z(n3) );
  XOR U147 ( .A(n4), .B(n215), .Z(n216) );
  XOR U148 ( .A(n217), .B(n218), .Z(n215) );
  AND U149 ( .A(n62), .B(n219), .Z(n218) );
  XOR U150 ( .A(p_input[8]), .B(n217), .Z(n219) );
  XOR U151 ( .A(n220), .B(n221), .Z(n217) );
  AND U152 ( .A(n66), .B(n222), .Z(n221) );
  XOR U153 ( .A(n223), .B(n224), .Z(n4) );
  AND U154 ( .A(n70), .B(n222), .Z(n224) );
  XNOR U155 ( .A(n225), .B(n220), .Z(n222) );
  XOR U156 ( .A(n226), .B(n227), .Z(n220) );
  AND U157 ( .A(n74), .B(n228), .Z(n227) );
  XOR U158 ( .A(p_input[40]), .B(n226), .Z(n228) );
  XOR U159 ( .A(n229), .B(n230), .Z(n226) );
  AND U160 ( .A(n78), .B(n231), .Z(n230) );
  IV U161 ( .A(n223), .Z(n225) );
  XNOR U162 ( .A(n232), .B(n233), .Z(n223) );
  AND U163 ( .A(n82), .B(n231), .Z(n233) );
  XNOR U164 ( .A(n232), .B(n229), .Z(n231) );
  XOR U165 ( .A(n234), .B(n235), .Z(n229) );
  AND U166 ( .A(n85), .B(n236), .Z(n235) );
  XOR U167 ( .A(p_input[72]), .B(n234), .Z(n236) );
  XOR U168 ( .A(n237), .B(n238), .Z(n234) );
  AND U169 ( .A(n89), .B(n239), .Z(n238) );
  XOR U170 ( .A(n240), .B(n241), .Z(n232) );
  AND U171 ( .A(n93), .B(n239), .Z(n241) );
  XNOR U172 ( .A(n240), .B(n237), .Z(n239) );
  XOR U173 ( .A(n242), .B(n243), .Z(n237) );
  AND U174 ( .A(n96), .B(n244), .Z(n243) );
  XOR U175 ( .A(p_input[104]), .B(n242), .Z(n244) );
  XOR U176 ( .A(n245), .B(n246), .Z(n242) );
  AND U177 ( .A(n100), .B(n247), .Z(n246) );
  XOR U178 ( .A(n248), .B(n249), .Z(n240) );
  AND U179 ( .A(n104), .B(n247), .Z(n249) );
  XNOR U180 ( .A(n248), .B(n245), .Z(n247) );
  XOR U181 ( .A(n250), .B(n251), .Z(n245) );
  AND U182 ( .A(n107), .B(n252), .Z(n251) );
  XOR U183 ( .A(p_input[136]), .B(n250), .Z(n252) );
  XOR U184 ( .A(n253), .B(n254), .Z(n250) );
  AND U185 ( .A(n111), .B(n255), .Z(n254) );
  XOR U186 ( .A(n256), .B(n257), .Z(n248) );
  AND U187 ( .A(n115), .B(n255), .Z(n257) );
  XNOR U188 ( .A(n256), .B(n253), .Z(n255) );
  XOR U189 ( .A(n258), .B(n259), .Z(n253) );
  AND U190 ( .A(n118), .B(n260), .Z(n259) );
  XOR U191 ( .A(p_input[168]), .B(n258), .Z(n260) );
  XOR U192 ( .A(n261), .B(n262), .Z(n258) );
  AND U193 ( .A(n122), .B(n263), .Z(n262) );
  XOR U194 ( .A(n264), .B(n265), .Z(n256) );
  AND U195 ( .A(n126), .B(n263), .Z(n265) );
  XNOR U196 ( .A(n264), .B(n261), .Z(n263) );
  XOR U197 ( .A(n266), .B(n267), .Z(n261) );
  AND U198 ( .A(n129), .B(n268), .Z(n267) );
  XOR U199 ( .A(p_input[200]), .B(n266), .Z(n268) );
  XOR U200 ( .A(n269), .B(n270), .Z(n266) );
  AND U201 ( .A(n133), .B(n271), .Z(n270) );
  XOR U202 ( .A(n272), .B(n273), .Z(n264) );
  AND U203 ( .A(n137), .B(n271), .Z(n273) );
  XNOR U204 ( .A(n272), .B(n269), .Z(n271) );
  XOR U205 ( .A(n274), .B(n275), .Z(n269) );
  AND U206 ( .A(n140), .B(n276), .Z(n275) );
  XOR U207 ( .A(p_input[232]), .B(n274), .Z(n276) );
  XOR U208 ( .A(n277), .B(n278), .Z(n274) );
  AND U209 ( .A(n144), .B(n279), .Z(n278) );
  XOR U210 ( .A(n280), .B(n281), .Z(n272) );
  AND U211 ( .A(n148), .B(n279), .Z(n281) );
  XNOR U212 ( .A(n280), .B(n277), .Z(n279) );
  XOR U213 ( .A(n282), .B(n283), .Z(n277) );
  AND U214 ( .A(n151), .B(n284), .Z(n283) );
  XOR U215 ( .A(p_input[264]), .B(n282), .Z(n284) );
  XOR U216 ( .A(n285), .B(n286), .Z(n282) );
  AND U217 ( .A(n155), .B(n287), .Z(n286) );
  XOR U218 ( .A(n288), .B(n289), .Z(n280) );
  AND U219 ( .A(n159), .B(n287), .Z(n289) );
  XNOR U220 ( .A(n288), .B(n285), .Z(n287) );
  XOR U221 ( .A(n290), .B(n291), .Z(n285) );
  AND U222 ( .A(n162), .B(n292), .Z(n291) );
  XOR U223 ( .A(p_input[296]), .B(n290), .Z(n292) );
  XOR U224 ( .A(n293), .B(n294), .Z(n290) );
  AND U225 ( .A(n166), .B(n295), .Z(n294) );
  XOR U226 ( .A(n296), .B(n297), .Z(n288) );
  AND U227 ( .A(n170), .B(n295), .Z(n297) );
  XNOR U228 ( .A(n296), .B(n293), .Z(n295) );
  XOR U229 ( .A(n298), .B(n299), .Z(n293) );
  AND U230 ( .A(n173), .B(n300), .Z(n299) );
  XOR U231 ( .A(p_input[328]), .B(n298), .Z(n300) );
  XOR U232 ( .A(n301), .B(n302), .Z(n298) );
  AND U233 ( .A(n177), .B(n303), .Z(n302) );
  XOR U234 ( .A(n304), .B(n305), .Z(n296) );
  AND U235 ( .A(n181), .B(n303), .Z(n305) );
  XNOR U236 ( .A(n304), .B(n301), .Z(n303) );
  XOR U237 ( .A(n306), .B(n307), .Z(n301) );
  AND U238 ( .A(n184), .B(n308), .Z(n307) );
  XOR U239 ( .A(p_input[360]), .B(n306), .Z(n308) );
  XOR U240 ( .A(n309), .B(n310), .Z(n306) );
  AND U241 ( .A(n188), .B(n311), .Z(n310) );
  XOR U242 ( .A(n312), .B(n313), .Z(n304) );
  AND U243 ( .A(n192), .B(n311), .Z(n313) );
  XNOR U244 ( .A(n312), .B(n309), .Z(n311) );
  XOR U245 ( .A(n314), .B(n315), .Z(n309) );
  AND U246 ( .A(n195), .B(n316), .Z(n315) );
  XOR U247 ( .A(p_input[392]), .B(n314), .Z(n316) );
  XOR U248 ( .A(n317), .B(n318), .Z(n314) );
  AND U249 ( .A(n199), .B(n319), .Z(n318) );
  XOR U250 ( .A(n320), .B(n321), .Z(n312) );
  AND U251 ( .A(n203), .B(n319), .Z(n321) );
  XNOR U252 ( .A(n320), .B(n317), .Z(n319) );
  XOR U253 ( .A(n322), .B(n323), .Z(n317) );
  AND U254 ( .A(n206), .B(n324), .Z(n323) );
  XOR U255 ( .A(p_input[424]), .B(n322), .Z(n324) );
  XNOR U256 ( .A(n325), .B(n326), .Z(n322) );
  AND U257 ( .A(n210), .B(n327), .Z(n326) );
  XNOR U258 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n328), .Z(n320) );
  AND U259 ( .A(n213), .B(n327), .Z(n328) );
  XOR U260 ( .A(n329), .B(n325), .Z(n327) );
  IV U261 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .Z(n325) );
  IV U262 ( .A(\knn_comb_/min_val_out[0][8] ), .Z(n329) );
  XOR U263 ( .A(n330), .B(n331), .Z(o[3]) );
  XOR U264 ( .A(n5), .B(n332), .Z(o[39]) );
  AND U265 ( .A(n58), .B(n333), .Z(n5) );
  XOR U266 ( .A(n6), .B(n332), .Z(n333) );
  XOR U267 ( .A(n334), .B(n335), .Z(n332) );
  AND U268 ( .A(n62), .B(n336), .Z(n335) );
  XOR U269 ( .A(p_input[7]), .B(n334), .Z(n336) );
  XOR U270 ( .A(n337), .B(n338), .Z(n334) );
  AND U271 ( .A(n66), .B(n339), .Z(n338) );
  XOR U272 ( .A(n340), .B(n341), .Z(n6) );
  AND U273 ( .A(n70), .B(n339), .Z(n341) );
  XNOR U274 ( .A(n342), .B(n337), .Z(n339) );
  XOR U275 ( .A(n343), .B(n344), .Z(n337) );
  AND U276 ( .A(n74), .B(n345), .Z(n344) );
  XOR U277 ( .A(p_input[39]), .B(n343), .Z(n345) );
  XOR U278 ( .A(n346), .B(n347), .Z(n343) );
  AND U279 ( .A(n78), .B(n348), .Z(n347) );
  IV U280 ( .A(n340), .Z(n342) );
  XNOR U281 ( .A(n349), .B(n350), .Z(n340) );
  AND U282 ( .A(n82), .B(n348), .Z(n350) );
  XNOR U283 ( .A(n349), .B(n346), .Z(n348) );
  XOR U284 ( .A(n351), .B(n352), .Z(n346) );
  AND U285 ( .A(n85), .B(n353), .Z(n352) );
  XOR U286 ( .A(p_input[71]), .B(n351), .Z(n353) );
  XOR U287 ( .A(n354), .B(n355), .Z(n351) );
  AND U288 ( .A(n89), .B(n356), .Z(n355) );
  XOR U289 ( .A(n357), .B(n358), .Z(n349) );
  AND U290 ( .A(n93), .B(n356), .Z(n358) );
  XNOR U291 ( .A(n357), .B(n354), .Z(n356) );
  XOR U292 ( .A(n359), .B(n360), .Z(n354) );
  AND U293 ( .A(n96), .B(n361), .Z(n360) );
  XOR U294 ( .A(p_input[103]), .B(n359), .Z(n361) );
  XOR U295 ( .A(n362), .B(n363), .Z(n359) );
  AND U296 ( .A(n100), .B(n364), .Z(n363) );
  XOR U297 ( .A(n365), .B(n366), .Z(n357) );
  AND U298 ( .A(n104), .B(n364), .Z(n366) );
  XNOR U299 ( .A(n365), .B(n362), .Z(n364) );
  XOR U300 ( .A(n367), .B(n368), .Z(n362) );
  AND U301 ( .A(n107), .B(n369), .Z(n368) );
  XOR U302 ( .A(p_input[135]), .B(n367), .Z(n369) );
  XOR U303 ( .A(n370), .B(n371), .Z(n367) );
  AND U304 ( .A(n111), .B(n372), .Z(n371) );
  XOR U305 ( .A(n373), .B(n374), .Z(n365) );
  AND U306 ( .A(n115), .B(n372), .Z(n374) );
  XNOR U307 ( .A(n373), .B(n370), .Z(n372) );
  XOR U308 ( .A(n375), .B(n376), .Z(n370) );
  AND U309 ( .A(n118), .B(n377), .Z(n376) );
  XOR U310 ( .A(p_input[167]), .B(n375), .Z(n377) );
  XOR U311 ( .A(n378), .B(n379), .Z(n375) );
  AND U312 ( .A(n122), .B(n380), .Z(n379) );
  XOR U313 ( .A(n381), .B(n382), .Z(n373) );
  AND U314 ( .A(n126), .B(n380), .Z(n382) );
  XNOR U315 ( .A(n381), .B(n378), .Z(n380) );
  XOR U316 ( .A(n383), .B(n384), .Z(n378) );
  AND U317 ( .A(n129), .B(n385), .Z(n384) );
  XOR U318 ( .A(p_input[199]), .B(n383), .Z(n385) );
  XOR U319 ( .A(n386), .B(n387), .Z(n383) );
  AND U320 ( .A(n133), .B(n388), .Z(n387) );
  XOR U321 ( .A(n389), .B(n390), .Z(n381) );
  AND U322 ( .A(n137), .B(n388), .Z(n390) );
  XNOR U323 ( .A(n389), .B(n386), .Z(n388) );
  XOR U324 ( .A(n391), .B(n392), .Z(n386) );
  AND U325 ( .A(n140), .B(n393), .Z(n392) );
  XOR U326 ( .A(p_input[231]), .B(n391), .Z(n393) );
  XOR U327 ( .A(n394), .B(n395), .Z(n391) );
  AND U328 ( .A(n144), .B(n396), .Z(n395) );
  XOR U329 ( .A(n397), .B(n398), .Z(n389) );
  AND U330 ( .A(n148), .B(n396), .Z(n398) );
  XNOR U331 ( .A(n397), .B(n394), .Z(n396) );
  XOR U332 ( .A(n399), .B(n400), .Z(n394) );
  AND U333 ( .A(n151), .B(n401), .Z(n400) );
  XOR U334 ( .A(p_input[263]), .B(n399), .Z(n401) );
  XOR U335 ( .A(n402), .B(n403), .Z(n399) );
  AND U336 ( .A(n155), .B(n404), .Z(n403) );
  XOR U337 ( .A(n405), .B(n406), .Z(n397) );
  AND U338 ( .A(n159), .B(n404), .Z(n406) );
  XNOR U339 ( .A(n405), .B(n402), .Z(n404) );
  XOR U340 ( .A(n407), .B(n408), .Z(n402) );
  AND U341 ( .A(n162), .B(n409), .Z(n408) );
  XOR U342 ( .A(p_input[295]), .B(n407), .Z(n409) );
  XOR U343 ( .A(n410), .B(n411), .Z(n407) );
  AND U344 ( .A(n166), .B(n412), .Z(n411) );
  XOR U345 ( .A(n413), .B(n414), .Z(n405) );
  AND U346 ( .A(n170), .B(n412), .Z(n414) );
  XNOR U347 ( .A(n413), .B(n410), .Z(n412) );
  XOR U348 ( .A(n415), .B(n416), .Z(n410) );
  AND U349 ( .A(n173), .B(n417), .Z(n416) );
  XOR U350 ( .A(p_input[327]), .B(n415), .Z(n417) );
  XOR U351 ( .A(n418), .B(n419), .Z(n415) );
  AND U352 ( .A(n177), .B(n420), .Z(n419) );
  XOR U353 ( .A(n421), .B(n422), .Z(n413) );
  AND U354 ( .A(n181), .B(n420), .Z(n422) );
  XNOR U355 ( .A(n421), .B(n418), .Z(n420) );
  XOR U356 ( .A(n423), .B(n424), .Z(n418) );
  AND U357 ( .A(n184), .B(n425), .Z(n424) );
  XOR U358 ( .A(p_input[359]), .B(n423), .Z(n425) );
  XOR U359 ( .A(n426), .B(n427), .Z(n423) );
  AND U360 ( .A(n188), .B(n428), .Z(n427) );
  XOR U361 ( .A(n429), .B(n430), .Z(n421) );
  AND U362 ( .A(n192), .B(n428), .Z(n430) );
  XNOR U363 ( .A(n429), .B(n426), .Z(n428) );
  XOR U364 ( .A(n431), .B(n432), .Z(n426) );
  AND U365 ( .A(n195), .B(n433), .Z(n432) );
  XOR U366 ( .A(p_input[391]), .B(n431), .Z(n433) );
  XOR U367 ( .A(n434), .B(n435), .Z(n431) );
  AND U368 ( .A(n199), .B(n436), .Z(n435) );
  XOR U369 ( .A(n437), .B(n438), .Z(n429) );
  AND U370 ( .A(n203), .B(n436), .Z(n438) );
  XNOR U371 ( .A(n437), .B(n434), .Z(n436) );
  XOR U372 ( .A(n439), .B(n440), .Z(n434) );
  AND U373 ( .A(n206), .B(n441), .Z(n440) );
  XOR U374 ( .A(p_input[423]), .B(n439), .Z(n441) );
  XNOR U375 ( .A(n442), .B(n443), .Z(n439) );
  AND U376 ( .A(n210), .B(n444), .Z(n443) );
  XNOR U377 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n445), .Z(n437) );
  AND U378 ( .A(n213), .B(n444), .Z(n445) );
  XOR U379 ( .A(n446), .B(n442), .Z(n444) );
  XOR U380 ( .A(n7), .B(n447), .Z(o[38]) );
  AND U381 ( .A(n58), .B(n448), .Z(n7) );
  XOR U382 ( .A(n8), .B(n447), .Z(n448) );
  XOR U383 ( .A(n449), .B(n450), .Z(n447) );
  AND U384 ( .A(n62), .B(n451), .Z(n450) );
  XOR U385 ( .A(p_input[6]), .B(n449), .Z(n451) );
  XOR U386 ( .A(n452), .B(n453), .Z(n449) );
  AND U387 ( .A(n66), .B(n454), .Z(n453) );
  XOR U388 ( .A(n455), .B(n456), .Z(n8) );
  AND U389 ( .A(n70), .B(n454), .Z(n456) );
  XNOR U390 ( .A(n457), .B(n452), .Z(n454) );
  XOR U391 ( .A(n458), .B(n459), .Z(n452) );
  AND U392 ( .A(n74), .B(n460), .Z(n459) );
  XOR U393 ( .A(p_input[38]), .B(n458), .Z(n460) );
  XOR U394 ( .A(n461), .B(n462), .Z(n458) );
  AND U395 ( .A(n78), .B(n463), .Z(n462) );
  IV U396 ( .A(n455), .Z(n457) );
  XNOR U397 ( .A(n464), .B(n465), .Z(n455) );
  AND U398 ( .A(n82), .B(n463), .Z(n465) );
  XNOR U399 ( .A(n464), .B(n461), .Z(n463) );
  XOR U400 ( .A(n466), .B(n467), .Z(n461) );
  AND U401 ( .A(n85), .B(n468), .Z(n467) );
  XOR U402 ( .A(p_input[70]), .B(n466), .Z(n468) );
  XOR U403 ( .A(n469), .B(n470), .Z(n466) );
  AND U404 ( .A(n89), .B(n471), .Z(n470) );
  XOR U405 ( .A(n472), .B(n473), .Z(n464) );
  AND U406 ( .A(n93), .B(n471), .Z(n473) );
  XNOR U407 ( .A(n472), .B(n469), .Z(n471) );
  XOR U408 ( .A(n474), .B(n475), .Z(n469) );
  AND U409 ( .A(n96), .B(n476), .Z(n475) );
  XOR U410 ( .A(p_input[102]), .B(n474), .Z(n476) );
  XOR U411 ( .A(n477), .B(n478), .Z(n474) );
  AND U412 ( .A(n100), .B(n479), .Z(n478) );
  XOR U413 ( .A(n480), .B(n481), .Z(n472) );
  AND U414 ( .A(n104), .B(n479), .Z(n481) );
  XNOR U415 ( .A(n480), .B(n477), .Z(n479) );
  XOR U416 ( .A(n482), .B(n483), .Z(n477) );
  AND U417 ( .A(n107), .B(n484), .Z(n483) );
  XOR U418 ( .A(p_input[134]), .B(n482), .Z(n484) );
  XOR U419 ( .A(n485), .B(n486), .Z(n482) );
  AND U420 ( .A(n111), .B(n487), .Z(n486) );
  XOR U421 ( .A(n488), .B(n489), .Z(n480) );
  AND U422 ( .A(n115), .B(n487), .Z(n489) );
  XNOR U423 ( .A(n488), .B(n485), .Z(n487) );
  XOR U424 ( .A(n490), .B(n491), .Z(n485) );
  AND U425 ( .A(n118), .B(n492), .Z(n491) );
  XOR U426 ( .A(p_input[166]), .B(n490), .Z(n492) );
  XOR U427 ( .A(n493), .B(n494), .Z(n490) );
  AND U428 ( .A(n122), .B(n495), .Z(n494) );
  XOR U429 ( .A(n496), .B(n497), .Z(n488) );
  AND U430 ( .A(n126), .B(n495), .Z(n497) );
  XNOR U431 ( .A(n496), .B(n493), .Z(n495) );
  XOR U432 ( .A(n498), .B(n499), .Z(n493) );
  AND U433 ( .A(n129), .B(n500), .Z(n499) );
  XOR U434 ( .A(p_input[198]), .B(n498), .Z(n500) );
  XOR U435 ( .A(n501), .B(n502), .Z(n498) );
  AND U436 ( .A(n133), .B(n503), .Z(n502) );
  XOR U437 ( .A(n504), .B(n505), .Z(n496) );
  AND U438 ( .A(n137), .B(n503), .Z(n505) );
  XNOR U439 ( .A(n504), .B(n501), .Z(n503) );
  XOR U440 ( .A(n506), .B(n507), .Z(n501) );
  AND U441 ( .A(n140), .B(n508), .Z(n507) );
  XOR U442 ( .A(p_input[230]), .B(n506), .Z(n508) );
  XOR U443 ( .A(n509), .B(n510), .Z(n506) );
  AND U444 ( .A(n144), .B(n511), .Z(n510) );
  XOR U445 ( .A(n512), .B(n513), .Z(n504) );
  AND U446 ( .A(n148), .B(n511), .Z(n513) );
  XNOR U447 ( .A(n512), .B(n509), .Z(n511) );
  XOR U448 ( .A(n514), .B(n515), .Z(n509) );
  AND U449 ( .A(n151), .B(n516), .Z(n515) );
  XOR U450 ( .A(p_input[262]), .B(n514), .Z(n516) );
  XOR U451 ( .A(n517), .B(n518), .Z(n514) );
  AND U452 ( .A(n155), .B(n519), .Z(n518) );
  XOR U453 ( .A(n520), .B(n521), .Z(n512) );
  AND U454 ( .A(n159), .B(n519), .Z(n521) );
  XNOR U455 ( .A(n520), .B(n517), .Z(n519) );
  XOR U456 ( .A(n522), .B(n523), .Z(n517) );
  AND U457 ( .A(n162), .B(n524), .Z(n523) );
  XOR U458 ( .A(p_input[294]), .B(n522), .Z(n524) );
  XOR U459 ( .A(n525), .B(n526), .Z(n522) );
  AND U460 ( .A(n166), .B(n527), .Z(n526) );
  XOR U461 ( .A(n528), .B(n529), .Z(n520) );
  AND U462 ( .A(n170), .B(n527), .Z(n529) );
  XNOR U463 ( .A(n528), .B(n525), .Z(n527) );
  XOR U464 ( .A(n530), .B(n531), .Z(n525) );
  AND U465 ( .A(n173), .B(n532), .Z(n531) );
  XOR U466 ( .A(p_input[326]), .B(n530), .Z(n532) );
  XOR U467 ( .A(n533), .B(n534), .Z(n530) );
  AND U468 ( .A(n177), .B(n535), .Z(n534) );
  XOR U469 ( .A(n536), .B(n537), .Z(n528) );
  AND U470 ( .A(n181), .B(n535), .Z(n537) );
  XNOR U471 ( .A(n536), .B(n533), .Z(n535) );
  XOR U472 ( .A(n538), .B(n539), .Z(n533) );
  AND U473 ( .A(n184), .B(n540), .Z(n539) );
  XOR U474 ( .A(p_input[358]), .B(n538), .Z(n540) );
  XOR U475 ( .A(n541), .B(n542), .Z(n538) );
  AND U476 ( .A(n188), .B(n543), .Z(n542) );
  XOR U477 ( .A(n544), .B(n545), .Z(n536) );
  AND U478 ( .A(n192), .B(n543), .Z(n545) );
  XNOR U479 ( .A(n544), .B(n541), .Z(n543) );
  XOR U480 ( .A(n546), .B(n547), .Z(n541) );
  AND U481 ( .A(n195), .B(n548), .Z(n547) );
  XOR U482 ( .A(p_input[390]), .B(n546), .Z(n548) );
  XOR U483 ( .A(n549), .B(n550), .Z(n546) );
  AND U484 ( .A(n199), .B(n551), .Z(n550) );
  XOR U485 ( .A(n552), .B(n553), .Z(n544) );
  AND U486 ( .A(n203), .B(n551), .Z(n553) );
  XNOR U487 ( .A(n552), .B(n549), .Z(n551) );
  XOR U488 ( .A(n554), .B(n555), .Z(n549) );
  AND U489 ( .A(n206), .B(n556), .Z(n555) );
  XOR U490 ( .A(p_input[422]), .B(n554), .Z(n556) );
  XNOR U491 ( .A(n557), .B(n558), .Z(n554) );
  AND U492 ( .A(n210), .B(n559), .Z(n558) );
  XNOR U493 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n560), .Z(n552) );
  AND U494 ( .A(n213), .B(n559), .Z(n560) );
  XOR U495 ( .A(n561), .B(n557), .Z(n559) );
  XOR U496 ( .A(n17), .B(n562), .Z(o[37]) );
  AND U497 ( .A(n58), .B(n563), .Z(n17) );
  XOR U498 ( .A(n18), .B(n562), .Z(n563) );
  XOR U499 ( .A(n564), .B(n565), .Z(n562) );
  AND U500 ( .A(n62), .B(n566), .Z(n565) );
  XOR U501 ( .A(p_input[5]), .B(n564), .Z(n566) );
  XOR U502 ( .A(n567), .B(n568), .Z(n564) );
  AND U503 ( .A(n66), .B(n569), .Z(n568) );
  XOR U504 ( .A(n570), .B(n571), .Z(n18) );
  AND U505 ( .A(n70), .B(n569), .Z(n571) );
  XNOR U506 ( .A(n572), .B(n567), .Z(n569) );
  XOR U507 ( .A(n573), .B(n574), .Z(n567) );
  AND U508 ( .A(n74), .B(n575), .Z(n574) );
  XOR U509 ( .A(p_input[37]), .B(n573), .Z(n575) );
  XOR U510 ( .A(n576), .B(n577), .Z(n573) );
  AND U511 ( .A(n78), .B(n578), .Z(n577) );
  IV U512 ( .A(n570), .Z(n572) );
  XNOR U513 ( .A(n579), .B(n580), .Z(n570) );
  AND U514 ( .A(n82), .B(n578), .Z(n580) );
  XNOR U515 ( .A(n579), .B(n576), .Z(n578) );
  XOR U516 ( .A(n581), .B(n582), .Z(n576) );
  AND U517 ( .A(n85), .B(n583), .Z(n582) );
  XOR U518 ( .A(p_input[69]), .B(n581), .Z(n583) );
  XOR U519 ( .A(n584), .B(n585), .Z(n581) );
  AND U520 ( .A(n89), .B(n586), .Z(n585) );
  XOR U521 ( .A(n587), .B(n588), .Z(n579) );
  AND U522 ( .A(n93), .B(n586), .Z(n588) );
  XNOR U523 ( .A(n587), .B(n584), .Z(n586) );
  XOR U524 ( .A(n589), .B(n590), .Z(n584) );
  AND U525 ( .A(n96), .B(n591), .Z(n590) );
  XOR U526 ( .A(p_input[101]), .B(n589), .Z(n591) );
  XOR U527 ( .A(n592), .B(n593), .Z(n589) );
  AND U528 ( .A(n100), .B(n594), .Z(n593) );
  XOR U529 ( .A(n595), .B(n596), .Z(n587) );
  AND U530 ( .A(n104), .B(n594), .Z(n596) );
  XNOR U531 ( .A(n595), .B(n592), .Z(n594) );
  XOR U532 ( .A(n597), .B(n598), .Z(n592) );
  AND U533 ( .A(n107), .B(n599), .Z(n598) );
  XOR U534 ( .A(p_input[133]), .B(n597), .Z(n599) );
  XOR U535 ( .A(n600), .B(n601), .Z(n597) );
  AND U536 ( .A(n111), .B(n602), .Z(n601) );
  XOR U537 ( .A(n603), .B(n604), .Z(n595) );
  AND U538 ( .A(n115), .B(n602), .Z(n604) );
  XNOR U539 ( .A(n603), .B(n600), .Z(n602) );
  XOR U540 ( .A(n605), .B(n606), .Z(n600) );
  AND U541 ( .A(n118), .B(n607), .Z(n606) );
  XOR U542 ( .A(p_input[165]), .B(n605), .Z(n607) );
  XOR U543 ( .A(n608), .B(n609), .Z(n605) );
  AND U544 ( .A(n122), .B(n610), .Z(n609) );
  XOR U545 ( .A(n611), .B(n612), .Z(n603) );
  AND U546 ( .A(n126), .B(n610), .Z(n612) );
  XNOR U547 ( .A(n611), .B(n608), .Z(n610) );
  XOR U548 ( .A(n613), .B(n614), .Z(n608) );
  AND U549 ( .A(n129), .B(n615), .Z(n614) );
  XOR U550 ( .A(p_input[197]), .B(n613), .Z(n615) );
  XOR U551 ( .A(n616), .B(n617), .Z(n613) );
  AND U552 ( .A(n133), .B(n618), .Z(n617) );
  XOR U553 ( .A(n619), .B(n620), .Z(n611) );
  AND U554 ( .A(n137), .B(n618), .Z(n620) );
  XNOR U555 ( .A(n619), .B(n616), .Z(n618) );
  XOR U556 ( .A(n621), .B(n622), .Z(n616) );
  AND U557 ( .A(n140), .B(n623), .Z(n622) );
  XOR U558 ( .A(p_input[229]), .B(n621), .Z(n623) );
  XOR U559 ( .A(n624), .B(n625), .Z(n621) );
  AND U560 ( .A(n144), .B(n626), .Z(n625) );
  XOR U561 ( .A(n627), .B(n628), .Z(n619) );
  AND U562 ( .A(n148), .B(n626), .Z(n628) );
  XNOR U563 ( .A(n627), .B(n624), .Z(n626) );
  XOR U564 ( .A(n629), .B(n630), .Z(n624) );
  AND U565 ( .A(n151), .B(n631), .Z(n630) );
  XOR U566 ( .A(p_input[261]), .B(n629), .Z(n631) );
  XOR U567 ( .A(n632), .B(n633), .Z(n629) );
  AND U568 ( .A(n155), .B(n634), .Z(n633) );
  XOR U569 ( .A(n635), .B(n636), .Z(n627) );
  AND U570 ( .A(n159), .B(n634), .Z(n636) );
  XNOR U571 ( .A(n635), .B(n632), .Z(n634) );
  XOR U572 ( .A(n637), .B(n638), .Z(n632) );
  AND U573 ( .A(n162), .B(n639), .Z(n638) );
  XOR U574 ( .A(p_input[293]), .B(n637), .Z(n639) );
  XOR U575 ( .A(n640), .B(n641), .Z(n637) );
  AND U576 ( .A(n166), .B(n642), .Z(n641) );
  XOR U577 ( .A(n643), .B(n644), .Z(n635) );
  AND U578 ( .A(n170), .B(n642), .Z(n644) );
  XNOR U579 ( .A(n643), .B(n640), .Z(n642) );
  XOR U580 ( .A(n645), .B(n646), .Z(n640) );
  AND U581 ( .A(n173), .B(n647), .Z(n646) );
  XOR U582 ( .A(p_input[325]), .B(n645), .Z(n647) );
  XOR U583 ( .A(n648), .B(n649), .Z(n645) );
  AND U584 ( .A(n177), .B(n650), .Z(n649) );
  XOR U585 ( .A(n651), .B(n652), .Z(n643) );
  AND U586 ( .A(n181), .B(n650), .Z(n652) );
  XNOR U587 ( .A(n651), .B(n648), .Z(n650) );
  XOR U588 ( .A(n653), .B(n654), .Z(n648) );
  AND U589 ( .A(n184), .B(n655), .Z(n654) );
  XOR U590 ( .A(p_input[357]), .B(n653), .Z(n655) );
  XOR U591 ( .A(n656), .B(n657), .Z(n653) );
  AND U592 ( .A(n188), .B(n658), .Z(n657) );
  XOR U593 ( .A(n659), .B(n660), .Z(n651) );
  AND U594 ( .A(n192), .B(n658), .Z(n660) );
  XNOR U595 ( .A(n659), .B(n656), .Z(n658) );
  XOR U596 ( .A(n661), .B(n662), .Z(n656) );
  AND U597 ( .A(n195), .B(n663), .Z(n662) );
  XOR U598 ( .A(p_input[389]), .B(n661), .Z(n663) );
  XOR U599 ( .A(n664), .B(n665), .Z(n661) );
  AND U600 ( .A(n199), .B(n666), .Z(n665) );
  XOR U601 ( .A(n667), .B(n668), .Z(n659) );
  AND U602 ( .A(n203), .B(n666), .Z(n668) );
  XNOR U603 ( .A(n667), .B(n664), .Z(n666) );
  XOR U604 ( .A(n669), .B(n670), .Z(n664) );
  AND U605 ( .A(n206), .B(n671), .Z(n670) );
  XOR U606 ( .A(p_input[421]), .B(n669), .Z(n671) );
  XNOR U607 ( .A(n672), .B(n673), .Z(n669) );
  AND U608 ( .A(n210), .B(n674), .Z(n673) );
  XNOR U609 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n675), .Z(n667) );
  AND U610 ( .A(n213), .B(n674), .Z(n675) );
  XOR U611 ( .A(n676), .B(n672), .Z(n674) );
  IV U612 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .Z(n672) );
  IV U613 ( .A(\knn_comb_/min_val_out[0][5] ), .Z(n676) );
  XOR U614 ( .A(n39), .B(n677), .Z(o[36]) );
  AND U615 ( .A(n58), .B(n678), .Z(n39) );
  XOR U616 ( .A(n40), .B(n677), .Z(n678) );
  XOR U617 ( .A(n679), .B(n680), .Z(n677) );
  AND U618 ( .A(n62), .B(n681), .Z(n680) );
  XOR U619 ( .A(p_input[4]), .B(n679), .Z(n681) );
  XOR U620 ( .A(n682), .B(n683), .Z(n679) );
  AND U621 ( .A(n66), .B(n684), .Z(n683) );
  XOR U622 ( .A(n685), .B(n686), .Z(n40) );
  AND U623 ( .A(n70), .B(n684), .Z(n686) );
  XNOR U624 ( .A(n687), .B(n682), .Z(n684) );
  XOR U625 ( .A(n688), .B(n689), .Z(n682) );
  AND U626 ( .A(n74), .B(n690), .Z(n689) );
  XOR U627 ( .A(p_input[36]), .B(n688), .Z(n690) );
  XOR U628 ( .A(n691), .B(n692), .Z(n688) );
  AND U629 ( .A(n78), .B(n693), .Z(n692) );
  IV U630 ( .A(n685), .Z(n687) );
  XNOR U631 ( .A(n694), .B(n695), .Z(n685) );
  AND U632 ( .A(n82), .B(n693), .Z(n695) );
  XNOR U633 ( .A(n694), .B(n691), .Z(n693) );
  XOR U634 ( .A(n696), .B(n697), .Z(n691) );
  AND U635 ( .A(n85), .B(n698), .Z(n697) );
  XOR U636 ( .A(p_input[68]), .B(n696), .Z(n698) );
  XOR U637 ( .A(n699), .B(n700), .Z(n696) );
  AND U638 ( .A(n89), .B(n701), .Z(n700) );
  XOR U639 ( .A(n702), .B(n703), .Z(n694) );
  AND U640 ( .A(n93), .B(n701), .Z(n703) );
  XNOR U641 ( .A(n702), .B(n699), .Z(n701) );
  XOR U642 ( .A(n704), .B(n705), .Z(n699) );
  AND U643 ( .A(n96), .B(n706), .Z(n705) );
  XOR U644 ( .A(p_input[100]), .B(n704), .Z(n706) );
  XOR U645 ( .A(n707), .B(n708), .Z(n704) );
  AND U646 ( .A(n100), .B(n709), .Z(n708) );
  XOR U647 ( .A(n710), .B(n711), .Z(n702) );
  AND U648 ( .A(n104), .B(n709), .Z(n711) );
  XNOR U649 ( .A(n710), .B(n707), .Z(n709) );
  XOR U650 ( .A(n712), .B(n713), .Z(n707) );
  AND U651 ( .A(n107), .B(n714), .Z(n713) );
  XOR U652 ( .A(p_input[132]), .B(n712), .Z(n714) );
  XOR U653 ( .A(n715), .B(n716), .Z(n712) );
  AND U654 ( .A(n111), .B(n717), .Z(n716) );
  XOR U655 ( .A(n718), .B(n719), .Z(n710) );
  AND U656 ( .A(n115), .B(n717), .Z(n719) );
  XNOR U657 ( .A(n718), .B(n715), .Z(n717) );
  XOR U658 ( .A(n720), .B(n721), .Z(n715) );
  AND U659 ( .A(n118), .B(n722), .Z(n721) );
  XOR U660 ( .A(p_input[164]), .B(n720), .Z(n722) );
  XOR U661 ( .A(n723), .B(n724), .Z(n720) );
  AND U662 ( .A(n122), .B(n725), .Z(n724) );
  XOR U663 ( .A(n726), .B(n727), .Z(n718) );
  AND U664 ( .A(n126), .B(n725), .Z(n727) );
  XNOR U665 ( .A(n726), .B(n723), .Z(n725) );
  XOR U666 ( .A(n728), .B(n729), .Z(n723) );
  AND U667 ( .A(n129), .B(n730), .Z(n729) );
  XOR U668 ( .A(p_input[196]), .B(n728), .Z(n730) );
  XOR U669 ( .A(n731), .B(n732), .Z(n728) );
  AND U670 ( .A(n133), .B(n733), .Z(n732) );
  XOR U671 ( .A(n734), .B(n735), .Z(n726) );
  AND U672 ( .A(n137), .B(n733), .Z(n735) );
  XNOR U673 ( .A(n734), .B(n731), .Z(n733) );
  XOR U674 ( .A(n736), .B(n737), .Z(n731) );
  AND U675 ( .A(n140), .B(n738), .Z(n737) );
  XOR U676 ( .A(p_input[228]), .B(n736), .Z(n738) );
  XOR U677 ( .A(n739), .B(n740), .Z(n736) );
  AND U678 ( .A(n144), .B(n741), .Z(n740) );
  XOR U679 ( .A(n742), .B(n743), .Z(n734) );
  AND U680 ( .A(n148), .B(n741), .Z(n743) );
  XNOR U681 ( .A(n742), .B(n739), .Z(n741) );
  XOR U682 ( .A(n744), .B(n745), .Z(n739) );
  AND U683 ( .A(n151), .B(n746), .Z(n745) );
  XOR U684 ( .A(p_input[260]), .B(n744), .Z(n746) );
  XOR U685 ( .A(n747), .B(n748), .Z(n744) );
  AND U686 ( .A(n155), .B(n749), .Z(n748) );
  XOR U687 ( .A(n750), .B(n751), .Z(n742) );
  AND U688 ( .A(n159), .B(n749), .Z(n751) );
  XNOR U689 ( .A(n750), .B(n747), .Z(n749) );
  XOR U690 ( .A(n752), .B(n753), .Z(n747) );
  AND U691 ( .A(n162), .B(n754), .Z(n753) );
  XOR U692 ( .A(p_input[292]), .B(n752), .Z(n754) );
  XOR U693 ( .A(n755), .B(n756), .Z(n752) );
  AND U694 ( .A(n166), .B(n757), .Z(n756) );
  XOR U695 ( .A(n758), .B(n759), .Z(n750) );
  AND U696 ( .A(n170), .B(n757), .Z(n759) );
  XNOR U697 ( .A(n758), .B(n755), .Z(n757) );
  XOR U698 ( .A(n760), .B(n761), .Z(n755) );
  AND U699 ( .A(n173), .B(n762), .Z(n761) );
  XOR U700 ( .A(p_input[324]), .B(n760), .Z(n762) );
  XOR U701 ( .A(n763), .B(n764), .Z(n760) );
  AND U702 ( .A(n177), .B(n765), .Z(n764) );
  XOR U703 ( .A(n766), .B(n767), .Z(n758) );
  AND U704 ( .A(n181), .B(n765), .Z(n767) );
  XNOR U705 ( .A(n766), .B(n763), .Z(n765) );
  XOR U706 ( .A(n768), .B(n769), .Z(n763) );
  AND U707 ( .A(n184), .B(n770), .Z(n769) );
  XOR U708 ( .A(p_input[356]), .B(n768), .Z(n770) );
  XOR U709 ( .A(n771), .B(n772), .Z(n768) );
  AND U710 ( .A(n188), .B(n773), .Z(n772) );
  XOR U711 ( .A(n774), .B(n775), .Z(n766) );
  AND U712 ( .A(n192), .B(n773), .Z(n775) );
  XNOR U713 ( .A(n774), .B(n771), .Z(n773) );
  XOR U714 ( .A(n776), .B(n777), .Z(n771) );
  AND U715 ( .A(n195), .B(n778), .Z(n777) );
  XOR U716 ( .A(p_input[388]), .B(n776), .Z(n778) );
  XOR U717 ( .A(n779), .B(n780), .Z(n776) );
  AND U718 ( .A(n199), .B(n781), .Z(n780) );
  XOR U719 ( .A(n782), .B(n783), .Z(n774) );
  AND U720 ( .A(n203), .B(n781), .Z(n783) );
  XNOR U721 ( .A(n782), .B(n779), .Z(n781) );
  XOR U722 ( .A(n784), .B(n785), .Z(n779) );
  AND U723 ( .A(n206), .B(n786), .Z(n785) );
  XOR U724 ( .A(p_input[420]), .B(n784), .Z(n786) );
  XNOR U725 ( .A(n787), .B(n788), .Z(n784) );
  AND U726 ( .A(n210), .B(n789), .Z(n788) );
  XNOR U727 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n790), .Z(n782) );
  AND U728 ( .A(n213), .B(n789), .Z(n790) );
  XOR U729 ( .A(n791), .B(n787), .Z(n789) );
  XOR U730 ( .A(n330), .B(n792), .Z(o[35]) );
  AND U731 ( .A(n58), .B(n793), .Z(n330) );
  XOR U732 ( .A(n331), .B(n792), .Z(n793) );
  XOR U733 ( .A(n794), .B(n795), .Z(n792) );
  AND U734 ( .A(n62), .B(n796), .Z(n795) );
  XOR U735 ( .A(p_input[3]), .B(n794), .Z(n796) );
  XOR U736 ( .A(n797), .B(n798), .Z(n794) );
  AND U737 ( .A(n66), .B(n799), .Z(n798) );
  XOR U738 ( .A(n800), .B(n801), .Z(n331) );
  AND U739 ( .A(n70), .B(n799), .Z(n801) );
  XNOR U740 ( .A(n802), .B(n797), .Z(n799) );
  XOR U741 ( .A(n803), .B(n804), .Z(n797) );
  AND U742 ( .A(n74), .B(n805), .Z(n804) );
  XOR U743 ( .A(p_input[35]), .B(n803), .Z(n805) );
  XOR U744 ( .A(n806), .B(n807), .Z(n803) );
  AND U745 ( .A(n78), .B(n808), .Z(n807) );
  IV U746 ( .A(n800), .Z(n802) );
  XNOR U747 ( .A(n809), .B(n810), .Z(n800) );
  AND U748 ( .A(n82), .B(n808), .Z(n810) );
  XNOR U749 ( .A(n809), .B(n806), .Z(n808) );
  XOR U750 ( .A(n811), .B(n812), .Z(n806) );
  AND U751 ( .A(n85), .B(n813), .Z(n812) );
  XOR U752 ( .A(p_input[67]), .B(n811), .Z(n813) );
  XOR U753 ( .A(n814), .B(n815), .Z(n811) );
  AND U754 ( .A(n89), .B(n816), .Z(n815) );
  XOR U755 ( .A(n817), .B(n818), .Z(n809) );
  AND U756 ( .A(n93), .B(n816), .Z(n818) );
  XNOR U757 ( .A(n817), .B(n814), .Z(n816) );
  XOR U758 ( .A(n819), .B(n820), .Z(n814) );
  AND U759 ( .A(n96), .B(n821), .Z(n820) );
  XOR U760 ( .A(p_input[99]), .B(n819), .Z(n821) );
  XOR U761 ( .A(n822), .B(n823), .Z(n819) );
  AND U762 ( .A(n100), .B(n824), .Z(n823) );
  XOR U763 ( .A(n825), .B(n826), .Z(n817) );
  AND U764 ( .A(n104), .B(n824), .Z(n826) );
  XNOR U765 ( .A(n825), .B(n822), .Z(n824) );
  XOR U766 ( .A(n827), .B(n828), .Z(n822) );
  AND U767 ( .A(n107), .B(n829), .Z(n828) );
  XOR U768 ( .A(p_input[131]), .B(n827), .Z(n829) );
  XOR U769 ( .A(n830), .B(n831), .Z(n827) );
  AND U770 ( .A(n111), .B(n832), .Z(n831) );
  XOR U771 ( .A(n833), .B(n834), .Z(n825) );
  AND U772 ( .A(n115), .B(n832), .Z(n834) );
  XNOR U773 ( .A(n833), .B(n830), .Z(n832) );
  XOR U774 ( .A(n835), .B(n836), .Z(n830) );
  AND U775 ( .A(n118), .B(n837), .Z(n836) );
  XOR U776 ( .A(p_input[163]), .B(n835), .Z(n837) );
  XOR U777 ( .A(n838), .B(n839), .Z(n835) );
  AND U778 ( .A(n122), .B(n840), .Z(n839) );
  XOR U779 ( .A(n841), .B(n842), .Z(n833) );
  AND U780 ( .A(n126), .B(n840), .Z(n842) );
  XNOR U781 ( .A(n841), .B(n838), .Z(n840) );
  XOR U782 ( .A(n843), .B(n844), .Z(n838) );
  AND U783 ( .A(n129), .B(n845), .Z(n844) );
  XOR U784 ( .A(p_input[195]), .B(n843), .Z(n845) );
  XOR U785 ( .A(n846), .B(n847), .Z(n843) );
  AND U786 ( .A(n133), .B(n848), .Z(n847) );
  XOR U787 ( .A(n849), .B(n850), .Z(n841) );
  AND U788 ( .A(n137), .B(n848), .Z(n850) );
  XNOR U789 ( .A(n849), .B(n846), .Z(n848) );
  XOR U790 ( .A(n851), .B(n852), .Z(n846) );
  AND U791 ( .A(n140), .B(n853), .Z(n852) );
  XOR U792 ( .A(p_input[227]), .B(n851), .Z(n853) );
  XOR U793 ( .A(n854), .B(n855), .Z(n851) );
  AND U794 ( .A(n144), .B(n856), .Z(n855) );
  XOR U795 ( .A(n857), .B(n858), .Z(n849) );
  AND U796 ( .A(n148), .B(n856), .Z(n858) );
  XNOR U797 ( .A(n857), .B(n854), .Z(n856) );
  XOR U798 ( .A(n859), .B(n860), .Z(n854) );
  AND U799 ( .A(n151), .B(n861), .Z(n860) );
  XOR U800 ( .A(p_input[259]), .B(n859), .Z(n861) );
  XOR U801 ( .A(n862), .B(n863), .Z(n859) );
  AND U802 ( .A(n155), .B(n864), .Z(n863) );
  XOR U803 ( .A(n865), .B(n866), .Z(n857) );
  AND U804 ( .A(n159), .B(n864), .Z(n866) );
  XNOR U805 ( .A(n865), .B(n862), .Z(n864) );
  XOR U806 ( .A(n867), .B(n868), .Z(n862) );
  AND U807 ( .A(n162), .B(n869), .Z(n868) );
  XOR U808 ( .A(p_input[291]), .B(n867), .Z(n869) );
  XOR U809 ( .A(n870), .B(n871), .Z(n867) );
  AND U810 ( .A(n166), .B(n872), .Z(n871) );
  XOR U811 ( .A(n873), .B(n874), .Z(n865) );
  AND U812 ( .A(n170), .B(n872), .Z(n874) );
  XNOR U813 ( .A(n873), .B(n870), .Z(n872) );
  XOR U814 ( .A(n875), .B(n876), .Z(n870) );
  AND U815 ( .A(n173), .B(n877), .Z(n876) );
  XOR U816 ( .A(p_input[323]), .B(n875), .Z(n877) );
  XOR U817 ( .A(n878), .B(n879), .Z(n875) );
  AND U818 ( .A(n177), .B(n880), .Z(n879) );
  XOR U819 ( .A(n881), .B(n882), .Z(n873) );
  AND U820 ( .A(n181), .B(n880), .Z(n882) );
  XNOR U821 ( .A(n881), .B(n878), .Z(n880) );
  XOR U822 ( .A(n883), .B(n884), .Z(n878) );
  AND U823 ( .A(n184), .B(n885), .Z(n884) );
  XOR U824 ( .A(p_input[355]), .B(n883), .Z(n885) );
  XOR U825 ( .A(n886), .B(n887), .Z(n883) );
  AND U826 ( .A(n188), .B(n888), .Z(n887) );
  XOR U827 ( .A(n889), .B(n890), .Z(n881) );
  AND U828 ( .A(n192), .B(n888), .Z(n890) );
  XNOR U829 ( .A(n889), .B(n886), .Z(n888) );
  XOR U830 ( .A(n891), .B(n892), .Z(n886) );
  AND U831 ( .A(n195), .B(n893), .Z(n892) );
  XOR U832 ( .A(p_input[387]), .B(n891), .Z(n893) );
  XOR U833 ( .A(n894), .B(n895), .Z(n891) );
  AND U834 ( .A(n199), .B(n896), .Z(n895) );
  XOR U835 ( .A(n897), .B(n898), .Z(n889) );
  AND U836 ( .A(n203), .B(n896), .Z(n898) );
  XNOR U837 ( .A(n897), .B(n894), .Z(n896) );
  XOR U838 ( .A(n899), .B(n900), .Z(n894) );
  AND U839 ( .A(n206), .B(n901), .Z(n900) );
  XOR U840 ( .A(p_input[419]), .B(n899), .Z(n901) );
  XNOR U841 ( .A(n902), .B(n903), .Z(n899) );
  AND U842 ( .A(n210), .B(n904), .Z(n903) );
  XNOR U843 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n905), .Z(n897) );
  AND U844 ( .A(n213), .B(n904), .Z(n905) );
  XOR U845 ( .A(n906), .B(n902), .Z(n904) );
  XOR U846 ( .A(n907), .B(n908), .Z(o[34]) );
  XOR U847 ( .A(n909), .B(n910), .Z(o[33]) );
  XOR U848 ( .A(n911), .B(n912), .Z(o[32]) );
  XOR U849 ( .A(n9), .B(n913), .Z(o[31]) );
  AND U850 ( .A(n58), .B(n914), .Z(n9) );
  XOR U851 ( .A(n10), .B(n913), .Z(n914) );
  XOR U852 ( .A(n915), .B(n916), .Z(n913) );
  AND U853 ( .A(n70), .B(n917), .Z(n916) );
  XOR U854 ( .A(n918), .B(n919), .Z(n10) );
  AND U855 ( .A(n62), .B(n920), .Z(n919) );
  XOR U856 ( .A(p_input[31]), .B(n918), .Z(n920) );
  XNOR U857 ( .A(n921), .B(n922), .Z(n918) );
  AND U858 ( .A(n66), .B(n917), .Z(n922) );
  XNOR U859 ( .A(n921), .B(n915), .Z(n917) );
  XOR U860 ( .A(n923), .B(n924), .Z(n915) );
  AND U861 ( .A(n82), .B(n925), .Z(n924) );
  XNOR U862 ( .A(n926), .B(n927), .Z(n921) );
  AND U863 ( .A(n74), .B(n928), .Z(n927) );
  XOR U864 ( .A(p_input[63]), .B(n926), .Z(n928) );
  XNOR U865 ( .A(n929), .B(n930), .Z(n926) );
  AND U866 ( .A(n78), .B(n925), .Z(n930) );
  XNOR U867 ( .A(n929), .B(n923), .Z(n925) );
  XOR U868 ( .A(n931), .B(n932), .Z(n923) );
  AND U869 ( .A(n93), .B(n933), .Z(n932) );
  XNOR U870 ( .A(n934), .B(n935), .Z(n929) );
  AND U871 ( .A(n85), .B(n936), .Z(n935) );
  XOR U872 ( .A(p_input[95]), .B(n934), .Z(n936) );
  XNOR U873 ( .A(n937), .B(n938), .Z(n934) );
  AND U874 ( .A(n89), .B(n933), .Z(n938) );
  XNOR U875 ( .A(n937), .B(n931), .Z(n933) );
  XOR U876 ( .A(n939), .B(n940), .Z(n931) );
  AND U877 ( .A(n104), .B(n941), .Z(n940) );
  XNOR U878 ( .A(n942), .B(n943), .Z(n937) );
  AND U879 ( .A(n96), .B(n944), .Z(n943) );
  XOR U880 ( .A(p_input[127]), .B(n942), .Z(n944) );
  XNOR U881 ( .A(n945), .B(n946), .Z(n942) );
  AND U882 ( .A(n100), .B(n941), .Z(n946) );
  XNOR U883 ( .A(n945), .B(n939), .Z(n941) );
  XOR U884 ( .A(n947), .B(n948), .Z(n939) );
  AND U885 ( .A(n115), .B(n949), .Z(n948) );
  XNOR U886 ( .A(n950), .B(n951), .Z(n945) );
  AND U887 ( .A(n107), .B(n952), .Z(n951) );
  XOR U888 ( .A(p_input[159]), .B(n950), .Z(n952) );
  XNOR U889 ( .A(n953), .B(n954), .Z(n950) );
  AND U890 ( .A(n111), .B(n949), .Z(n954) );
  XNOR U891 ( .A(n953), .B(n947), .Z(n949) );
  XOR U892 ( .A(n955), .B(n956), .Z(n947) );
  AND U893 ( .A(n126), .B(n957), .Z(n956) );
  XNOR U894 ( .A(n958), .B(n959), .Z(n953) );
  AND U895 ( .A(n118), .B(n960), .Z(n959) );
  XOR U896 ( .A(p_input[191]), .B(n958), .Z(n960) );
  XNOR U897 ( .A(n961), .B(n962), .Z(n958) );
  AND U898 ( .A(n122), .B(n957), .Z(n962) );
  XNOR U899 ( .A(n961), .B(n955), .Z(n957) );
  XOR U900 ( .A(n963), .B(n964), .Z(n955) );
  AND U901 ( .A(n137), .B(n965), .Z(n964) );
  XNOR U902 ( .A(n966), .B(n967), .Z(n961) );
  AND U903 ( .A(n129), .B(n968), .Z(n967) );
  XOR U904 ( .A(p_input[223]), .B(n966), .Z(n968) );
  XNOR U905 ( .A(n969), .B(n970), .Z(n966) );
  AND U906 ( .A(n133), .B(n965), .Z(n970) );
  XNOR U907 ( .A(n969), .B(n963), .Z(n965) );
  XOR U908 ( .A(n971), .B(n972), .Z(n963) );
  AND U909 ( .A(n148), .B(n973), .Z(n972) );
  XNOR U910 ( .A(n974), .B(n975), .Z(n969) );
  AND U911 ( .A(n140), .B(n976), .Z(n975) );
  XOR U912 ( .A(p_input[255]), .B(n974), .Z(n976) );
  XNOR U913 ( .A(n977), .B(n978), .Z(n974) );
  AND U914 ( .A(n144), .B(n973), .Z(n978) );
  XNOR U915 ( .A(n977), .B(n971), .Z(n973) );
  XOR U916 ( .A(n979), .B(n980), .Z(n971) );
  AND U917 ( .A(n159), .B(n981), .Z(n980) );
  XNOR U918 ( .A(n982), .B(n983), .Z(n977) );
  AND U919 ( .A(n151), .B(n984), .Z(n983) );
  XOR U920 ( .A(p_input[287]), .B(n982), .Z(n984) );
  XNOR U921 ( .A(n985), .B(n986), .Z(n982) );
  AND U922 ( .A(n155), .B(n981), .Z(n986) );
  XNOR U923 ( .A(n985), .B(n979), .Z(n981) );
  XOR U924 ( .A(n987), .B(n988), .Z(n979) );
  AND U925 ( .A(n170), .B(n989), .Z(n988) );
  XNOR U926 ( .A(n990), .B(n991), .Z(n985) );
  AND U927 ( .A(n162), .B(n992), .Z(n991) );
  XOR U928 ( .A(p_input[319]), .B(n990), .Z(n992) );
  XNOR U929 ( .A(n993), .B(n994), .Z(n990) );
  AND U930 ( .A(n166), .B(n989), .Z(n994) );
  XNOR U931 ( .A(n993), .B(n987), .Z(n989) );
  XOR U932 ( .A(n995), .B(n996), .Z(n987) );
  AND U933 ( .A(n181), .B(n997), .Z(n996) );
  XNOR U934 ( .A(n998), .B(n999), .Z(n993) );
  AND U935 ( .A(n173), .B(n1000), .Z(n999) );
  XOR U936 ( .A(p_input[351]), .B(n998), .Z(n1000) );
  XNOR U937 ( .A(n1001), .B(n1002), .Z(n998) );
  AND U938 ( .A(n177), .B(n997), .Z(n1002) );
  XNOR U939 ( .A(n1001), .B(n995), .Z(n997) );
  XOR U940 ( .A(n1003), .B(n1004), .Z(n995) );
  AND U941 ( .A(n192), .B(n1005), .Z(n1004) );
  XNOR U942 ( .A(n1006), .B(n1007), .Z(n1001) );
  AND U943 ( .A(n184), .B(n1008), .Z(n1007) );
  XOR U944 ( .A(p_input[383]), .B(n1006), .Z(n1008) );
  XNOR U945 ( .A(n1009), .B(n1010), .Z(n1006) );
  AND U946 ( .A(n188), .B(n1005), .Z(n1010) );
  XNOR U947 ( .A(n1009), .B(n1003), .Z(n1005) );
  XOR U948 ( .A(n1011), .B(n1012), .Z(n1003) );
  AND U949 ( .A(n203), .B(n1013), .Z(n1012) );
  XNOR U950 ( .A(n1014), .B(n1015), .Z(n1009) );
  AND U951 ( .A(n195), .B(n1016), .Z(n1015) );
  XOR U952 ( .A(p_input[415]), .B(n1014), .Z(n1016) );
  XNOR U953 ( .A(n1017), .B(n1018), .Z(n1014) );
  AND U954 ( .A(n199), .B(n1013), .Z(n1018) );
  XNOR U955 ( .A(n1017), .B(n1011), .Z(n1013) );
  XOR U956 ( .A(\knn_comb_/min_val_out[0][31] ), .B(n1019), .Z(n1011) );
  AND U957 ( .A(n213), .B(n1020), .Z(n1019) );
  XNOR U958 ( .A(n1021), .B(n1022), .Z(n1017) );
  AND U959 ( .A(n206), .B(n1023), .Z(n1022) );
  XOR U960 ( .A(p_input[447]), .B(n1021), .Z(n1023) );
  XNOR U961 ( .A(n1024), .B(n1025), .Z(n1021) );
  AND U962 ( .A(n210), .B(n1020), .Z(n1025) );
  XOR U963 ( .A(n1026), .B(n1024), .Z(n1020) );
  IV U964 ( .A(\knn_comb_/min_val_out[0][31] ), .Z(n1026) );
  IV U965 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .Z(n1024) );
  XOR U966 ( .A(n11), .B(n1027), .Z(o[30]) );
  AND U967 ( .A(n58), .B(n1028), .Z(n11) );
  XOR U968 ( .A(n12), .B(n1027), .Z(n1028) );
  XOR U969 ( .A(n1029), .B(n1030), .Z(n1027) );
  AND U970 ( .A(n70), .B(n1031), .Z(n1030) );
  XOR U971 ( .A(n1032), .B(n1033), .Z(n12) );
  AND U972 ( .A(n62), .B(n1034), .Z(n1033) );
  XOR U973 ( .A(p_input[30]), .B(n1032), .Z(n1034) );
  XNOR U974 ( .A(n1035), .B(n1036), .Z(n1032) );
  AND U975 ( .A(n66), .B(n1031), .Z(n1036) );
  XNOR U976 ( .A(n1035), .B(n1029), .Z(n1031) );
  XOR U977 ( .A(n1037), .B(n1038), .Z(n1029) );
  AND U978 ( .A(n82), .B(n1039), .Z(n1038) );
  XNOR U979 ( .A(n1040), .B(n1041), .Z(n1035) );
  AND U980 ( .A(n74), .B(n1042), .Z(n1041) );
  XOR U981 ( .A(p_input[62]), .B(n1040), .Z(n1042) );
  XNOR U982 ( .A(n1043), .B(n1044), .Z(n1040) );
  AND U983 ( .A(n78), .B(n1039), .Z(n1044) );
  XNOR U984 ( .A(n1043), .B(n1037), .Z(n1039) );
  XOR U985 ( .A(n1045), .B(n1046), .Z(n1037) );
  AND U986 ( .A(n93), .B(n1047), .Z(n1046) );
  XNOR U987 ( .A(n1048), .B(n1049), .Z(n1043) );
  AND U988 ( .A(n85), .B(n1050), .Z(n1049) );
  XOR U989 ( .A(p_input[94]), .B(n1048), .Z(n1050) );
  XNOR U990 ( .A(n1051), .B(n1052), .Z(n1048) );
  AND U991 ( .A(n89), .B(n1047), .Z(n1052) );
  XNOR U992 ( .A(n1051), .B(n1045), .Z(n1047) );
  XOR U993 ( .A(n1053), .B(n1054), .Z(n1045) );
  AND U994 ( .A(n104), .B(n1055), .Z(n1054) );
  XNOR U995 ( .A(n1056), .B(n1057), .Z(n1051) );
  AND U996 ( .A(n96), .B(n1058), .Z(n1057) );
  XOR U997 ( .A(p_input[126]), .B(n1056), .Z(n1058) );
  XNOR U998 ( .A(n1059), .B(n1060), .Z(n1056) );
  AND U999 ( .A(n100), .B(n1055), .Z(n1060) );
  XNOR U1000 ( .A(n1059), .B(n1053), .Z(n1055) );
  XOR U1001 ( .A(n1061), .B(n1062), .Z(n1053) );
  AND U1002 ( .A(n115), .B(n1063), .Z(n1062) );
  XNOR U1003 ( .A(n1064), .B(n1065), .Z(n1059) );
  AND U1004 ( .A(n107), .B(n1066), .Z(n1065) );
  XOR U1005 ( .A(p_input[158]), .B(n1064), .Z(n1066) );
  XNOR U1006 ( .A(n1067), .B(n1068), .Z(n1064) );
  AND U1007 ( .A(n111), .B(n1063), .Z(n1068) );
  XNOR U1008 ( .A(n1067), .B(n1061), .Z(n1063) );
  XOR U1009 ( .A(n1069), .B(n1070), .Z(n1061) );
  AND U1010 ( .A(n126), .B(n1071), .Z(n1070) );
  XNOR U1011 ( .A(n1072), .B(n1073), .Z(n1067) );
  AND U1012 ( .A(n118), .B(n1074), .Z(n1073) );
  XOR U1013 ( .A(p_input[190]), .B(n1072), .Z(n1074) );
  XNOR U1014 ( .A(n1075), .B(n1076), .Z(n1072) );
  AND U1015 ( .A(n122), .B(n1071), .Z(n1076) );
  XNOR U1016 ( .A(n1075), .B(n1069), .Z(n1071) );
  XOR U1017 ( .A(n1077), .B(n1078), .Z(n1069) );
  AND U1018 ( .A(n137), .B(n1079), .Z(n1078) );
  XNOR U1019 ( .A(n1080), .B(n1081), .Z(n1075) );
  AND U1020 ( .A(n129), .B(n1082), .Z(n1081) );
  XOR U1021 ( .A(p_input[222]), .B(n1080), .Z(n1082) );
  XNOR U1022 ( .A(n1083), .B(n1084), .Z(n1080) );
  AND U1023 ( .A(n133), .B(n1079), .Z(n1084) );
  XNOR U1024 ( .A(n1083), .B(n1077), .Z(n1079) );
  XOR U1025 ( .A(n1085), .B(n1086), .Z(n1077) );
  AND U1026 ( .A(n148), .B(n1087), .Z(n1086) );
  XNOR U1027 ( .A(n1088), .B(n1089), .Z(n1083) );
  AND U1028 ( .A(n140), .B(n1090), .Z(n1089) );
  XOR U1029 ( .A(p_input[254]), .B(n1088), .Z(n1090) );
  XNOR U1030 ( .A(n1091), .B(n1092), .Z(n1088) );
  AND U1031 ( .A(n144), .B(n1087), .Z(n1092) );
  XNOR U1032 ( .A(n1091), .B(n1085), .Z(n1087) );
  XOR U1033 ( .A(n1093), .B(n1094), .Z(n1085) );
  AND U1034 ( .A(n159), .B(n1095), .Z(n1094) );
  XNOR U1035 ( .A(n1096), .B(n1097), .Z(n1091) );
  AND U1036 ( .A(n151), .B(n1098), .Z(n1097) );
  XOR U1037 ( .A(p_input[286]), .B(n1096), .Z(n1098) );
  XNOR U1038 ( .A(n1099), .B(n1100), .Z(n1096) );
  AND U1039 ( .A(n155), .B(n1095), .Z(n1100) );
  XNOR U1040 ( .A(n1099), .B(n1093), .Z(n1095) );
  XOR U1041 ( .A(n1101), .B(n1102), .Z(n1093) );
  AND U1042 ( .A(n170), .B(n1103), .Z(n1102) );
  XNOR U1043 ( .A(n1104), .B(n1105), .Z(n1099) );
  AND U1044 ( .A(n162), .B(n1106), .Z(n1105) );
  XOR U1045 ( .A(p_input[318]), .B(n1104), .Z(n1106) );
  XNOR U1046 ( .A(n1107), .B(n1108), .Z(n1104) );
  AND U1047 ( .A(n166), .B(n1103), .Z(n1108) );
  XNOR U1048 ( .A(n1107), .B(n1101), .Z(n1103) );
  XOR U1049 ( .A(n1109), .B(n1110), .Z(n1101) );
  AND U1050 ( .A(n181), .B(n1111), .Z(n1110) );
  XNOR U1051 ( .A(n1112), .B(n1113), .Z(n1107) );
  AND U1052 ( .A(n173), .B(n1114), .Z(n1113) );
  XOR U1053 ( .A(p_input[350]), .B(n1112), .Z(n1114) );
  XNOR U1054 ( .A(n1115), .B(n1116), .Z(n1112) );
  AND U1055 ( .A(n177), .B(n1111), .Z(n1116) );
  XNOR U1056 ( .A(n1115), .B(n1109), .Z(n1111) );
  XOR U1057 ( .A(n1117), .B(n1118), .Z(n1109) );
  AND U1058 ( .A(n192), .B(n1119), .Z(n1118) );
  XNOR U1059 ( .A(n1120), .B(n1121), .Z(n1115) );
  AND U1060 ( .A(n184), .B(n1122), .Z(n1121) );
  XOR U1061 ( .A(p_input[382]), .B(n1120), .Z(n1122) );
  XNOR U1062 ( .A(n1123), .B(n1124), .Z(n1120) );
  AND U1063 ( .A(n188), .B(n1119), .Z(n1124) );
  XNOR U1064 ( .A(n1123), .B(n1117), .Z(n1119) );
  XOR U1065 ( .A(n1125), .B(n1126), .Z(n1117) );
  AND U1066 ( .A(n203), .B(n1127), .Z(n1126) );
  XNOR U1067 ( .A(n1128), .B(n1129), .Z(n1123) );
  AND U1068 ( .A(n195), .B(n1130), .Z(n1129) );
  XOR U1069 ( .A(p_input[414]), .B(n1128), .Z(n1130) );
  XNOR U1070 ( .A(n1131), .B(n1132), .Z(n1128) );
  AND U1071 ( .A(n199), .B(n1127), .Z(n1132) );
  XNOR U1072 ( .A(n1131), .B(n1125), .Z(n1127) );
  XOR U1073 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n1133), .Z(n1125) );
  AND U1074 ( .A(n213), .B(n1134), .Z(n1133) );
  XNOR U1075 ( .A(n1135), .B(n1136), .Z(n1131) );
  AND U1076 ( .A(n206), .B(n1137), .Z(n1136) );
  XOR U1077 ( .A(p_input[446]), .B(n1135), .Z(n1137) );
  XNOR U1078 ( .A(n1138), .B(n1139), .Z(n1135) );
  AND U1079 ( .A(n210), .B(n1134), .Z(n1139) );
  XOR U1080 ( .A(n1140), .B(n1138), .Z(n1134) );
  IV U1081 ( .A(\knn_comb_/min_val_out[0][30] ), .Z(n1140) );
  IV U1082 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .Z(n1138) );
  XOR U1083 ( .A(n907), .B(n1141), .Z(o[2]) );
  AND U1084 ( .A(n58), .B(n1142), .Z(n907) );
  XOR U1085 ( .A(n908), .B(n1141), .Z(n1142) );
  XOR U1086 ( .A(n1143), .B(n1144), .Z(n1141) );
  AND U1087 ( .A(n70), .B(n1145), .Z(n1144) );
  XOR U1088 ( .A(n1146), .B(n1147), .Z(n908) );
  AND U1089 ( .A(n62), .B(n1148), .Z(n1147) );
  XOR U1090 ( .A(p_input[2]), .B(n1146), .Z(n1148) );
  XNOR U1091 ( .A(n1149), .B(n1150), .Z(n1146) );
  AND U1092 ( .A(n66), .B(n1145), .Z(n1150) );
  XNOR U1093 ( .A(n1149), .B(n1143), .Z(n1145) );
  XOR U1094 ( .A(n1151), .B(n1152), .Z(n1143) );
  AND U1095 ( .A(n82), .B(n1153), .Z(n1152) );
  XNOR U1096 ( .A(n1154), .B(n1155), .Z(n1149) );
  AND U1097 ( .A(n74), .B(n1156), .Z(n1155) );
  XOR U1098 ( .A(p_input[34]), .B(n1154), .Z(n1156) );
  XNOR U1099 ( .A(n1157), .B(n1158), .Z(n1154) );
  AND U1100 ( .A(n78), .B(n1153), .Z(n1158) );
  XNOR U1101 ( .A(n1157), .B(n1151), .Z(n1153) );
  XOR U1102 ( .A(n1159), .B(n1160), .Z(n1151) );
  AND U1103 ( .A(n93), .B(n1161), .Z(n1160) );
  XNOR U1104 ( .A(n1162), .B(n1163), .Z(n1157) );
  AND U1105 ( .A(n85), .B(n1164), .Z(n1163) );
  XOR U1106 ( .A(p_input[66]), .B(n1162), .Z(n1164) );
  XNOR U1107 ( .A(n1165), .B(n1166), .Z(n1162) );
  AND U1108 ( .A(n89), .B(n1161), .Z(n1166) );
  XNOR U1109 ( .A(n1165), .B(n1159), .Z(n1161) );
  XOR U1110 ( .A(n1167), .B(n1168), .Z(n1159) );
  AND U1111 ( .A(n104), .B(n1169), .Z(n1168) );
  XNOR U1112 ( .A(n1170), .B(n1171), .Z(n1165) );
  AND U1113 ( .A(n96), .B(n1172), .Z(n1171) );
  XOR U1114 ( .A(p_input[98]), .B(n1170), .Z(n1172) );
  XNOR U1115 ( .A(n1173), .B(n1174), .Z(n1170) );
  AND U1116 ( .A(n100), .B(n1169), .Z(n1174) );
  XNOR U1117 ( .A(n1173), .B(n1167), .Z(n1169) );
  XOR U1118 ( .A(n1175), .B(n1176), .Z(n1167) );
  AND U1119 ( .A(n115), .B(n1177), .Z(n1176) );
  XNOR U1120 ( .A(n1178), .B(n1179), .Z(n1173) );
  AND U1121 ( .A(n107), .B(n1180), .Z(n1179) );
  XOR U1122 ( .A(p_input[130]), .B(n1178), .Z(n1180) );
  XNOR U1123 ( .A(n1181), .B(n1182), .Z(n1178) );
  AND U1124 ( .A(n111), .B(n1177), .Z(n1182) );
  XNOR U1125 ( .A(n1181), .B(n1175), .Z(n1177) );
  XOR U1126 ( .A(n1183), .B(n1184), .Z(n1175) );
  AND U1127 ( .A(n126), .B(n1185), .Z(n1184) );
  XNOR U1128 ( .A(n1186), .B(n1187), .Z(n1181) );
  AND U1129 ( .A(n118), .B(n1188), .Z(n1187) );
  XOR U1130 ( .A(p_input[162]), .B(n1186), .Z(n1188) );
  XNOR U1131 ( .A(n1189), .B(n1190), .Z(n1186) );
  AND U1132 ( .A(n122), .B(n1185), .Z(n1190) );
  XNOR U1133 ( .A(n1189), .B(n1183), .Z(n1185) );
  XOR U1134 ( .A(n1191), .B(n1192), .Z(n1183) );
  AND U1135 ( .A(n137), .B(n1193), .Z(n1192) );
  XNOR U1136 ( .A(n1194), .B(n1195), .Z(n1189) );
  AND U1137 ( .A(n129), .B(n1196), .Z(n1195) );
  XOR U1138 ( .A(p_input[194]), .B(n1194), .Z(n1196) );
  XNOR U1139 ( .A(n1197), .B(n1198), .Z(n1194) );
  AND U1140 ( .A(n133), .B(n1193), .Z(n1198) );
  XNOR U1141 ( .A(n1197), .B(n1191), .Z(n1193) );
  XOR U1142 ( .A(n1199), .B(n1200), .Z(n1191) );
  AND U1143 ( .A(n148), .B(n1201), .Z(n1200) );
  XNOR U1144 ( .A(n1202), .B(n1203), .Z(n1197) );
  AND U1145 ( .A(n140), .B(n1204), .Z(n1203) );
  XOR U1146 ( .A(p_input[226]), .B(n1202), .Z(n1204) );
  XNOR U1147 ( .A(n1205), .B(n1206), .Z(n1202) );
  AND U1148 ( .A(n144), .B(n1201), .Z(n1206) );
  XNOR U1149 ( .A(n1205), .B(n1199), .Z(n1201) );
  XOR U1150 ( .A(n1207), .B(n1208), .Z(n1199) );
  AND U1151 ( .A(n159), .B(n1209), .Z(n1208) );
  XNOR U1152 ( .A(n1210), .B(n1211), .Z(n1205) );
  AND U1153 ( .A(n151), .B(n1212), .Z(n1211) );
  XOR U1154 ( .A(p_input[258]), .B(n1210), .Z(n1212) );
  XNOR U1155 ( .A(n1213), .B(n1214), .Z(n1210) );
  AND U1156 ( .A(n155), .B(n1209), .Z(n1214) );
  XNOR U1157 ( .A(n1213), .B(n1207), .Z(n1209) );
  XOR U1158 ( .A(n1215), .B(n1216), .Z(n1207) );
  AND U1159 ( .A(n170), .B(n1217), .Z(n1216) );
  XNOR U1160 ( .A(n1218), .B(n1219), .Z(n1213) );
  AND U1161 ( .A(n162), .B(n1220), .Z(n1219) );
  XOR U1162 ( .A(p_input[290]), .B(n1218), .Z(n1220) );
  XNOR U1163 ( .A(n1221), .B(n1222), .Z(n1218) );
  AND U1164 ( .A(n166), .B(n1217), .Z(n1222) );
  XNOR U1165 ( .A(n1221), .B(n1215), .Z(n1217) );
  XOR U1166 ( .A(n1223), .B(n1224), .Z(n1215) );
  AND U1167 ( .A(n181), .B(n1225), .Z(n1224) );
  XNOR U1168 ( .A(n1226), .B(n1227), .Z(n1221) );
  AND U1169 ( .A(n173), .B(n1228), .Z(n1227) );
  XOR U1170 ( .A(p_input[322]), .B(n1226), .Z(n1228) );
  XNOR U1171 ( .A(n1229), .B(n1230), .Z(n1226) );
  AND U1172 ( .A(n177), .B(n1225), .Z(n1230) );
  XNOR U1173 ( .A(n1229), .B(n1223), .Z(n1225) );
  XOR U1174 ( .A(n1231), .B(n1232), .Z(n1223) );
  AND U1175 ( .A(n192), .B(n1233), .Z(n1232) );
  XNOR U1176 ( .A(n1234), .B(n1235), .Z(n1229) );
  AND U1177 ( .A(n184), .B(n1236), .Z(n1235) );
  XOR U1178 ( .A(p_input[354]), .B(n1234), .Z(n1236) );
  XNOR U1179 ( .A(n1237), .B(n1238), .Z(n1234) );
  AND U1180 ( .A(n188), .B(n1233), .Z(n1238) );
  XNOR U1181 ( .A(n1237), .B(n1231), .Z(n1233) );
  XOR U1182 ( .A(n1239), .B(n1240), .Z(n1231) );
  AND U1183 ( .A(n203), .B(n1241), .Z(n1240) );
  XNOR U1184 ( .A(n1242), .B(n1243), .Z(n1237) );
  AND U1185 ( .A(n195), .B(n1244), .Z(n1243) );
  XOR U1186 ( .A(p_input[386]), .B(n1242), .Z(n1244) );
  XNOR U1187 ( .A(n1245), .B(n1246), .Z(n1242) );
  AND U1188 ( .A(n199), .B(n1241), .Z(n1246) );
  XNOR U1189 ( .A(n1245), .B(n1239), .Z(n1241) );
  XOR U1190 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n1247), .Z(n1239) );
  AND U1191 ( .A(n213), .B(n1248), .Z(n1247) );
  XNOR U1192 ( .A(n1249), .B(n1250), .Z(n1245) );
  AND U1193 ( .A(n206), .B(n1251), .Z(n1250) );
  XOR U1194 ( .A(p_input[418]), .B(n1249), .Z(n1251) );
  XNOR U1195 ( .A(n1252), .B(n1253), .Z(n1249) );
  AND U1196 ( .A(n210), .B(n1248), .Z(n1253) );
  XOR U1197 ( .A(\knn_comb_/min_val_out[0][2] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n1248) );
  XOR U1198 ( .A(n13), .B(n1254), .Z(o[29]) );
  AND U1199 ( .A(n58), .B(n1255), .Z(n13) );
  XOR U1200 ( .A(n14), .B(n1254), .Z(n1255) );
  XOR U1201 ( .A(n1256), .B(n1257), .Z(n1254) );
  AND U1202 ( .A(n70), .B(n1258), .Z(n1257) );
  XOR U1203 ( .A(n1259), .B(n1260), .Z(n14) );
  AND U1204 ( .A(n62), .B(n1261), .Z(n1260) );
  XOR U1205 ( .A(p_input[29]), .B(n1259), .Z(n1261) );
  XNOR U1206 ( .A(n1262), .B(n1263), .Z(n1259) );
  AND U1207 ( .A(n66), .B(n1258), .Z(n1263) );
  XNOR U1208 ( .A(n1262), .B(n1256), .Z(n1258) );
  XOR U1209 ( .A(n1264), .B(n1265), .Z(n1256) );
  AND U1210 ( .A(n82), .B(n1266), .Z(n1265) );
  XNOR U1211 ( .A(n1267), .B(n1268), .Z(n1262) );
  AND U1212 ( .A(n74), .B(n1269), .Z(n1268) );
  XOR U1213 ( .A(p_input[61]), .B(n1267), .Z(n1269) );
  XNOR U1214 ( .A(n1270), .B(n1271), .Z(n1267) );
  AND U1215 ( .A(n78), .B(n1266), .Z(n1271) );
  XNOR U1216 ( .A(n1270), .B(n1264), .Z(n1266) );
  XOR U1217 ( .A(n1272), .B(n1273), .Z(n1264) );
  AND U1218 ( .A(n93), .B(n1274), .Z(n1273) );
  XNOR U1219 ( .A(n1275), .B(n1276), .Z(n1270) );
  AND U1220 ( .A(n85), .B(n1277), .Z(n1276) );
  XOR U1221 ( .A(p_input[93]), .B(n1275), .Z(n1277) );
  XNOR U1222 ( .A(n1278), .B(n1279), .Z(n1275) );
  AND U1223 ( .A(n89), .B(n1274), .Z(n1279) );
  XNOR U1224 ( .A(n1278), .B(n1272), .Z(n1274) );
  XOR U1225 ( .A(n1280), .B(n1281), .Z(n1272) );
  AND U1226 ( .A(n104), .B(n1282), .Z(n1281) );
  XNOR U1227 ( .A(n1283), .B(n1284), .Z(n1278) );
  AND U1228 ( .A(n96), .B(n1285), .Z(n1284) );
  XOR U1229 ( .A(p_input[125]), .B(n1283), .Z(n1285) );
  XNOR U1230 ( .A(n1286), .B(n1287), .Z(n1283) );
  AND U1231 ( .A(n100), .B(n1282), .Z(n1287) );
  XNOR U1232 ( .A(n1286), .B(n1280), .Z(n1282) );
  XOR U1233 ( .A(n1288), .B(n1289), .Z(n1280) );
  AND U1234 ( .A(n115), .B(n1290), .Z(n1289) );
  XNOR U1235 ( .A(n1291), .B(n1292), .Z(n1286) );
  AND U1236 ( .A(n107), .B(n1293), .Z(n1292) );
  XOR U1237 ( .A(p_input[157]), .B(n1291), .Z(n1293) );
  XNOR U1238 ( .A(n1294), .B(n1295), .Z(n1291) );
  AND U1239 ( .A(n111), .B(n1290), .Z(n1295) );
  XNOR U1240 ( .A(n1294), .B(n1288), .Z(n1290) );
  XOR U1241 ( .A(n1296), .B(n1297), .Z(n1288) );
  AND U1242 ( .A(n126), .B(n1298), .Z(n1297) );
  XNOR U1243 ( .A(n1299), .B(n1300), .Z(n1294) );
  AND U1244 ( .A(n118), .B(n1301), .Z(n1300) );
  XOR U1245 ( .A(p_input[189]), .B(n1299), .Z(n1301) );
  XNOR U1246 ( .A(n1302), .B(n1303), .Z(n1299) );
  AND U1247 ( .A(n122), .B(n1298), .Z(n1303) );
  XNOR U1248 ( .A(n1302), .B(n1296), .Z(n1298) );
  XOR U1249 ( .A(n1304), .B(n1305), .Z(n1296) );
  AND U1250 ( .A(n137), .B(n1306), .Z(n1305) );
  XNOR U1251 ( .A(n1307), .B(n1308), .Z(n1302) );
  AND U1252 ( .A(n129), .B(n1309), .Z(n1308) );
  XOR U1253 ( .A(p_input[221]), .B(n1307), .Z(n1309) );
  XNOR U1254 ( .A(n1310), .B(n1311), .Z(n1307) );
  AND U1255 ( .A(n133), .B(n1306), .Z(n1311) );
  XNOR U1256 ( .A(n1310), .B(n1304), .Z(n1306) );
  XOR U1257 ( .A(n1312), .B(n1313), .Z(n1304) );
  AND U1258 ( .A(n148), .B(n1314), .Z(n1313) );
  XNOR U1259 ( .A(n1315), .B(n1316), .Z(n1310) );
  AND U1260 ( .A(n140), .B(n1317), .Z(n1316) );
  XOR U1261 ( .A(p_input[253]), .B(n1315), .Z(n1317) );
  XNOR U1262 ( .A(n1318), .B(n1319), .Z(n1315) );
  AND U1263 ( .A(n144), .B(n1314), .Z(n1319) );
  XNOR U1264 ( .A(n1318), .B(n1312), .Z(n1314) );
  XOR U1265 ( .A(n1320), .B(n1321), .Z(n1312) );
  AND U1266 ( .A(n159), .B(n1322), .Z(n1321) );
  XNOR U1267 ( .A(n1323), .B(n1324), .Z(n1318) );
  AND U1268 ( .A(n151), .B(n1325), .Z(n1324) );
  XOR U1269 ( .A(p_input[285]), .B(n1323), .Z(n1325) );
  XNOR U1270 ( .A(n1326), .B(n1327), .Z(n1323) );
  AND U1271 ( .A(n155), .B(n1322), .Z(n1327) );
  XNOR U1272 ( .A(n1326), .B(n1320), .Z(n1322) );
  XOR U1273 ( .A(n1328), .B(n1329), .Z(n1320) );
  AND U1274 ( .A(n170), .B(n1330), .Z(n1329) );
  XNOR U1275 ( .A(n1331), .B(n1332), .Z(n1326) );
  AND U1276 ( .A(n162), .B(n1333), .Z(n1332) );
  XOR U1277 ( .A(p_input[317]), .B(n1331), .Z(n1333) );
  XNOR U1278 ( .A(n1334), .B(n1335), .Z(n1331) );
  AND U1279 ( .A(n166), .B(n1330), .Z(n1335) );
  XNOR U1280 ( .A(n1334), .B(n1328), .Z(n1330) );
  XOR U1281 ( .A(n1336), .B(n1337), .Z(n1328) );
  AND U1282 ( .A(n181), .B(n1338), .Z(n1337) );
  XNOR U1283 ( .A(n1339), .B(n1340), .Z(n1334) );
  AND U1284 ( .A(n173), .B(n1341), .Z(n1340) );
  XOR U1285 ( .A(p_input[349]), .B(n1339), .Z(n1341) );
  XNOR U1286 ( .A(n1342), .B(n1343), .Z(n1339) );
  AND U1287 ( .A(n177), .B(n1338), .Z(n1343) );
  XNOR U1288 ( .A(n1342), .B(n1336), .Z(n1338) );
  XOR U1289 ( .A(n1344), .B(n1345), .Z(n1336) );
  AND U1290 ( .A(n192), .B(n1346), .Z(n1345) );
  XNOR U1291 ( .A(n1347), .B(n1348), .Z(n1342) );
  AND U1292 ( .A(n184), .B(n1349), .Z(n1348) );
  XOR U1293 ( .A(p_input[381]), .B(n1347), .Z(n1349) );
  XNOR U1294 ( .A(n1350), .B(n1351), .Z(n1347) );
  AND U1295 ( .A(n188), .B(n1346), .Z(n1351) );
  XNOR U1296 ( .A(n1350), .B(n1344), .Z(n1346) );
  XOR U1297 ( .A(n1352), .B(n1353), .Z(n1344) );
  AND U1298 ( .A(n203), .B(n1354), .Z(n1353) );
  XNOR U1299 ( .A(n1355), .B(n1356), .Z(n1350) );
  AND U1300 ( .A(n195), .B(n1357), .Z(n1356) );
  XOR U1301 ( .A(p_input[413]), .B(n1355), .Z(n1357) );
  XNOR U1302 ( .A(n1358), .B(n1359), .Z(n1355) );
  AND U1303 ( .A(n199), .B(n1354), .Z(n1359) );
  XNOR U1304 ( .A(n1358), .B(n1352), .Z(n1354) );
  XOR U1305 ( .A(\knn_comb_/min_val_out[0][29] ), .B(n1360), .Z(n1352) );
  AND U1306 ( .A(n213), .B(n1361), .Z(n1360) );
  XNOR U1307 ( .A(n1362), .B(n1363), .Z(n1358) );
  AND U1308 ( .A(n206), .B(n1364), .Z(n1363) );
  XOR U1309 ( .A(p_input[445]), .B(n1362), .Z(n1364) );
  XNOR U1310 ( .A(n1365), .B(n1366), .Z(n1362) );
  AND U1311 ( .A(n210), .B(n1361), .Z(n1366) );
  XOR U1312 ( .A(\knn_comb_/min_val_out[0][29] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .Z(n1361) );
  XOR U1313 ( .A(n15), .B(n1367), .Z(o[28]) );
  AND U1314 ( .A(n58), .B(n1368), .Z(n15) );
  XOR U1315 ( .A(n16), .B(n1367), .Z(n1368) );
  XOR U1316 ( .A(n1369), .B(n1370), .Z(n1367) );
  AND U1317 ( .A(n70), .B(n1371), .Z(n1370) );
  XOR U1318 ( .A(n1372), .B(n1373), .Z(n16) );
  AND U1319 ( .A(n62), .B(n1374), .Z(n1373) );
  XOR U1320 ( .A(p_input[28]), .B(n1372), .Z(n1374) );
  XNOR U1321 ( .A(n1375), .B(n1376), .Z(n1372) );
  AND U1322 ( .A(n66), .B(n1371), .Z(n1376) );
  XNOR U1323 ( .A(n1375), .B(n1369), .Z(n1371) );
  XOR U1324 ( .A(n1377), .B(n1378), .Z(n1369) );
  AND U1325 ( .A(n82), .B(n1379), .Z(n1378) );
  XNOR U1326 ( .A(n1380), .B(n1381), .Z(n1375) );
  AND U1327 ( .A(n74), .B(n1382), .Z(n1381) );
  XOR U1328 ( .A(p_input[60]), .B(n1380), .Z(n1382) );
  XNOR U1329 ( .A(n1383), .B(n1384), .Z(n1380) );
  AND U1330 ( .A(n78), .B(n1379), .Z(n1384) );
  XNOR U1331 ( .A(n1383), .B(n1377), .Z(n1379) );
  XOR U1332 ( .A(n1385), .B(n1386), .Z(n1377) );
  AND U1333 ( .A(n93), .B(n1387), .Z(n1386) );
  XNOR U1334 ( .A(n1388), .B(n1389), .Z(n1383) );
  AND U1335 ( .A(n85), .B(n1390), .Z(n1389) );
  XOR U1336 ( .A(p_input[92]), .B(n1388), .Z(n1390) );
  XNOR U1337 ( .A(n1391), .B(n1392), .Z(n1388) );
  AND U1338 ( .A(n89), .B(n1387), .Z(n1392) );
  XNOR U1339 ( .A(n1391), .B(n1385), .Z(n1387) );
  XOR U1340 ( .A(n1393), .B(n1394), .Z(n1385) );
  AND U1341 ( .A(n104), .B(n1395), .Z(n1394) );
  XNOR U1342 ( .A(n1396), .B(n1397), .Z(n1391) );
  AND U1343 ( .A(n96), .B(n1398), .Z(n1397) );
  XOR U1344 ( .A(p_input[124]), .B(n1396), .Z(n1398) );
  XNOR U1345 ( .A(n1399), .B(n1400), .Z(n1396) );
  AND U1346 ( .A(n100), .B(n1395), .Z(n1400) );
  XNOR U1347 ( .A(n1399), .B(n1393), .Z(n1395) );
  XOR U1348 ( .A(n1401), .B(n1402), .Z(n1393) );
  AND U1349 ( .A(n115), .B(n1403), .Z(n1402) );
  XNOR U1350 ( .A(n1404), .B(n1405), .Z(n1399) );
  AND U1351 ( .A(n107), .B(n1406), .Z(n1405) );
  XOR U1352 ( .A(p_input[156]), .B(n1404), .Z(n1406) );
  XNOR U1353 ( .A(n1407), .B(n1408), .Z(n1404) );
  AND U1354 ( .A(n111), .B(n1403), .Z(n1408) );
  XNOR U1355 ( .A(n1407), .B(n1401), .Z(n1403) );
  XOR U1356 ( .A(n1409), .B(n1410), .Z(n1401) );
  AND U1357 ( .A(n126), .B(n1411), .Z(n1410) );
  XNOR U1358 ( .A(n1412), .B(n1413), .Z(n1407) );
  AND U1359 ( .A(n118), .B(n1414), .Z(n1413) );
  XOR U1360 ( .A(p_input[188]), .B(n1412), .Z(n1414) );
  XNOR U1361 ( .A(n1415), .B(n1416), .Z(n1412) );
  AND U1362 ( .A(n122), .B(n1411), .Z(n1416) );
  XNOR U1363 ( .A(n1415), .B(n1409), .Z(n1411) );
  XOR U1364 ( .A(n1417), .B(n1418), .Z(n1409) );
  AND U1365 ( .A(n137), .B(n1419), .Z(n1418) );
  XNOR U1366 ( .A(n1420), .B(n1421), .Z(n1415) );
  AND U1367 ( .A(n129), .B(n1422), .Z(n1421) );
  XOR U1368 ( .A(p_input[220]), .B(n1420), .Z(n1422) );
  XNOR U1369 ( .A(n1423), .B(n1424), .Z(n1420) );
  AND U1370 ( .A(n133), .B(n1419), .Z(n1424) );
  XNOR U1371 ( .A(n1423), .B(n1417), .Z(n1419) );
  XOR U1372 ( .A(n1425), .B(n1426), .Z(n1417) );
  AND U1373 ( .A(n148), .B(n1427), .Z(n1426) );
  XNOR U1374 ( .A(n1428), .B(n1429), .Z(n1423) );
  AND U1375 ( .A(n140), .B(n1430), .Z(n1429) );
  XOR U1376 ( .A(p_input[252]), .B(n1428), .Z(n1430) );
  XNOR U1377 ( .A(n1431), .B(n1432), .Z(n1428) );
  AND U1378 ( .A(n144), .B(n1427), .Z(n1432) );
  XNOR U1379 ( .A(n1431), .B(n1425), .Z(n1427) );
  XOR U1380 ( .A(n1433), .B(n1434), .Z(n1425) );
  AND U1381 ( .A(n159), .B(n1435), .Z(n1434) );
  XNOR U1382 ( .A(n1436), .B(n1437), .Z(n1431) );
  AND U1383 ( .A(n151), .B(n1438), .Z(n1437) );
  XOR U1384 ( .A(p_input[284]), .B(n1436), .Z(n1438) );
  XNOR U1385 ( .A(n1439), .B(n1440), .Z(n1436) );
  AND U1386 ( .A(n155), .B(n1435), .Z(n1440) );
  XNOR U1387 ( .A(n1439), .B(n1433), .Z(n1435) );
  XOR U1388 ( .A(n1441), .B(n1442), .Z(n1433) );
  AND U1389 ( .A(n170), .B(n1443), .Z(n1442) );
  XNOR U1390 ( .A(n1444), .B(n1445), .Z(n1439) );
  AND U1391 ( .A(n162), .B(n1446), .Z(n1445) );
  XOR U1392 ( .A(p_input[316]), .B(n1444), .Z(n1446) );
  XNOR U1393 ( .A(n1447), .B(n1448), .Z(n1444) );
  AND U1394 ( .A(n166), .B(n1443), .Z(n1448) );
  XNOR U1395 ( .A(n1447), .B(n1441), .Z(n1443) );
  XOR U1396 ( .A(n1449), .B(n1450), .Z(n1441) );
  AND U1397 ( .A(n181), .B(n1451), .Z(n1450) );
  XNOR U1398 ( .A(n1452), .B(n1453), .Z(n1447) );
  AND U1399 ( .A(n173), .B(n1454), .Z(n1453) );
  XOR U1400 ( .A(p_input[348]), .B(n1452), .Z(n1454) );
  XNOR U1401 ( .A(n1455), .B(n1456), .Z(n1452) );
  AND U1402 ( .A(n177), .B(n1451), .Z(n1456) );
  XNOR U1403 ( .A(n1455), .B(n1449), .Z(n1451) );
  XOR U1404 ( .A(n1457), .B(n1458), .Z(n1449) );
  AND U1405 ( .A(n192), .B(n1459), .Z(n1458) );
  XNOR U1406 ( .A(n1460), .B(n1461), .Z(n1455) );
  AND U1407 ( .A(n184), .B(n1462), .Z(n1461) );
  XOR U1408 ( .A(p_input[380]), .B(n1460), .Z(n1462) );
  XNOR U1409 ( .A(n1463), .B(n1464), .Z(n1460) );
  AND U1410 ( .A(n188), .B(n1459), .Z(n1464) );
  XNOR U1411 ( .A(n1463), .B(n1457), .Z(n1459) );
  XOR U1412 ( .A(n1465), .B(n1466), .Z(n1457) );
  AND U1413 ( .A(n203), .B(n1467), .Z(n1466) );
  XNOR U1414 ( .A(n1468), .B(n1469), .Z(n1463) );
  AND U1415 ( .A(n195), .B(n1470), .Z(n1469) );
  XOR U1416 ( .A(p_input[412]), .B(n1468), .Z(n1470) );
  XNOR U1417 ( .A(n1471), .B(n1472), .Z(n1468) );
  AND U1418 ( .A(n199), .B(n1467), .Z(n1472) );
  XNOR U1419 ( .A(n1471), .B(n1465), .Z(n1467) );
  XOR U1420 ( .A(\knn_comb_/min_val_out[0][28] ), .B(n1473), .Z(n1465) );
  AND U1421 ( .A(n213), .B(n1474), .Z(n1473) );
  XNOR U1422 ( .A(n1475), .B(n1476), .Z(n1471) );
  AND U1423 ( .A(n206), .B(n1477), .Z(n1476) );
  XOR U1424 ( .A(p_input[444]), .B(n1475), .Z(n1477) );
  XNOR U1425 ( .A(n1478), .B(n1479), .Z(n1475) );
  AND U1426 ( .A(n210), .B(n1474), .Z(n1479) );
  XOR U1427 ( .A(\knn_comb_/min_val_out[0][28] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .Z(n1474) );
  XOR U1428 ( .A(n19), .B(n1480), .Z(o[27]) );
  AND U1429 ( .A(n58), .B(n1481), .Z(n19) );
  XOR U1430 ( .A(n20), .B(n1480), .Z(n1481) );
  XOR U1431 ( .A(n1482), .B(n1483), .Z(n1480) );
  AND U1432 ( .A(n70), .B(n1484), .Z(n1483) );
  XOR U1433 ( .A(n1485), .B(n1486), .Z(n20) );
  AND U1434 ( .A(n62), .B(n1487), .Z(n1486) );
  XOR U1435 ( .A(p_input[27]), .B(n1485), .Z(n1487) );
  XNOR U1436 ( .A(n1488), .B(n1489), .Z(n1485) );
  AND U1437 ( .A(n66), .B(n1484), .Z(n1489) );
  XNOR U1438 ( .A(n1488), .B(n1482), .Z(n1484) );
  XOR U1439 ( .A(n1490), .B(n1491), .Z(n1482) );
  AND U1440 ( .A(n82), .B(n1492), .Z(n1491) );
  XNOR U1441 ( .A(n1493), .B(n1494), .Z(n1488) );
  AND U1442 ( .A(n74), .B(n1495), .Z(n1494) );
  XOR U1443 ( .A(p_input[59]), .B(n1493), .Z(n1495) );
  XNOR U1444 ( .A(n1496), .B(n1497), .Z(n1493) );
  AND U1445 ( .A(n78), .B(n1492), .Z(n1497) );
  XNOR U1446 ( .A(n1496), .B(n1490), .Z(n1492) );
  XOR U1447 ( .A(n1498), .B(n1499), .Z(n1490) );
  AND U1448 ( .A(n93), .B(n1500), .Z(n1499) );
  XNOR U1449 ( .A(n1501), .B(n1502), .Z(n1496) );
  AND U1450 ( .A(n85), .B(n1503), .Z(n1502) );
  XOR U1451 ( .A(p_input[91]), .B(n1501), .Z(n1503) );
  XNOR U1452 ( .A(n1504), .B(n1505), .Z(n1501) );
  AND U1453 ( .A(n89), .B(n1500), .Z(n1505) );
  XNOR U1454 ( .A(n1504), .B(n1498), .Z(n1500) );
  XOR U1455 ( .A(n1506), .B(n1507), .Z(n1498) );
  AND U1456 ( .A(n104), .B(n1508), .Z(n1507) );
  XNOR U1457 ( .A(n1509), .B(n1510), .Z(n1504) );
  AND U1458 ( .A(n96), .B(n1511), .Z(n1510) );
  XOR U1459 ( .A(p_input[123]), .B(n1509), .Z(n1511) );
  XNOR U1460 ( .A(n1512), .B(n1513), .Z(n1509) );
  AND U1461 ( .A(n100), .B(n1508), .Z(n1513) );
  XNOR U1462 ( .A(n1512), .B(n1506), .Z(n1508) );
  XOR U1463 ( .A(n1514), .B(n1515), .Z(n1506) );
  AND U1464 ( .A(n115), .B(n1516), .Z(n1515) );
  XNOR U1465 ( .A(n1517), .B(n1518), .Z(n1512) );
  AND U1466 ( .A(n107), .B(n1519), .Z(n1518) );
  XOR U1467 ( .A(p_input[155]), .B(n1517), .Z(n1519) );
  XNOR U1468 ( .A(n1520), .B(n1521), .Z(n1517) );
  AND U1469 ( .A(n111), .B(n1516), .Z(n1521) );
  XNOR U1470 ( .A(n1520), .B(n1514), .Z(n1516) );
  XOR U1471 ( .A(n1522), .B(n1523), .Z(n1514) );
  AND U1472 ( .A(n126), .B(n1524), .Z(n1523) );
  XNOR U1473 ( .A(n1525), .B(n1526), .Z(n1520) );
  AND U1474 ( .A(n118), .B(n1527), .Z(n1526) );
  XOR U1475 ( .A(p_input[187]), .B(n1525), .Z(n1527) );
  XNOR U1476 ( .A(n1528), .B(n1529), .Z(n1525) );
  AND U1477 ( .A(n122), .B(n1524), .Z(n1529) );
  XNOR U1478 ( .A(n1528), .B(n1522), .Z(n1524) );
  XOR U1479 ( .A(n1530), .B(n1531), .Z(n1522) );
  AND U1480 ( .A(n137), .B(n1532), .Z(n1531) );
  XNOR U1481 ( .A(n1533), .B(n1534), .Z(n1528) );
  AND U1482 ( .A(n129), .B(n1535), .Z(n1534) );
  XOR U1483 ( .A(p_input[219]), .B(n1533), .Z(n1535) );
  XNOR U1484 ( .A(n1536), .B(n1537), .Z(n1533) );
  AND U1485 ( .A(n133), .B(n1532), .Z(n1537) );
  XNOR U1486 ( .A(n1536), .B(n1530), .Z(n1532) );
  XOR U1487 ( .A(n1538), .B(n1539), .Z(n1530) );
  AND U1488 ( .A(n148), .B(n1540), .Z(n1539) );
  XNOR U1489 ( .A(n1541), .B(n1542), .Z(n1536) );
  AND U1490 ( .A(n140), .B(n1543), .Z(n1542) );
  XOR U1491 ( .A(p_input[251]), .B(n1541), .Z(n1543) );
  XNOR U1492 ( .A(n1544), .B(n1545), .Z(n1541) );
  AND U1493 ( .A(n144), .B(n1540), .Z(n1545) );
  XNOR U1494 ( .A(n1544), .B(n1538), .Z(n1540) );
  XOR U1495 ( .A(n1546), .B(n1547), .Z(n1538) );
  AND U1496 ( .A(n159), .B(n1548), .Z(n1547) );
  XNOR U1497 ( .A(n1549), .B(n1550), .Z(n1544) );
  AND U1498 ( .A(n151), .B(n1551), .Z(n1550) );
  XOR U1499 ( .A(p_input[283]), .B(n1549), .Z(n1551) );
  XNOR U1500 ( .A(n1552), .B(n1553), .Z(n1549) );
  AND U1501 ( .A(n155), .B(n1548), .Z(n1553) );
  XNOR U1502 ( .A(n1552), .B(n1546), .Z(n1548) );
  XOR U1503 ( .A(n1554), .B(n1555), .Z(n1546) );
  AND U1504 ( .A(n170), .B(n1556), .Z(n1555) );
  XNOR U1505 ( .A(n1557), .B(n1558), .Z(n1552) );
  AND U1506 ( .A(n162), .B(n1559), .Z(n1558) );
  XOR U1507 ( .A(p_input[315]), .B(n1557), .Z(n1559) );
  XNOR U1508 ( .A(n1560), .B(n1561), .Z(n1557) );
  AND U1509 ( .A(n166), .B(n1556), .Z(n1561) );
  XNOR U1510 ( .A(n1560), .B(n1554), .Z(n1556) );
  XOR U1511 ( .A(n1562), .B(n1563), .Z(n1554) );
  AND U1512 ( .A(n181), .B(n1564), .Z(n1563) );
  XNOR U1513 ( .A(n1565), .B(n1566), .Z(n1560) );
  AND U1514 ( .A(n173), .B(n1567), .Z(n1566) );
  XOR U1515 ( .A(p_input[347]), .B(n1565), .Z(n1567) );
  XNOR U1516 ( .A(n1568), .B(n1569), .Z(n1565) );
  AND U1517 ( .A(n177), .B(n1564), .Z(n1569) );
  XNOR U1518 ( .A(n1568), .B(n1562), .Z(n1564) );
  XOR U1519 ( .A(n1570), .B(n1571), .Z(n1562) );
  AND U1520 ( .A(n192), .B(n1572), .Z(n1571) );
  XNOR U1521 ( .A(n1573), .B(n1574), .Z(n1568) );
  AND U1522 ( .A(n184), .B(n1575), .Z(n1574) );
  XOR U1523 ( .A(p_input[379]), .B(n1573), .Z(n1575) );
  XNOR U1524 ( .A(n1576), .B(n1577), .Z(n1573) );
  AND U1525 ( .A(n188), .B(n1572), .Z(n1577) );
  XNOR U1526 ( .A(n1576), .B(n1570), .Z(n1572) );
  XOR U1527 ( .A(n1578), .B(n1579), .Z(n1570) );
  AND U1528 ( .A(n203), .B(n1580), .Z(n1579) );
  XNOR U1529 ( .A(n1581), .B(n1582), .Z(n1576) );
  AND U1530 ( .A(n195), .B(n1583), .Z(n1582) );
  XOR U1531 ( .A(p_input[411]), .B(n1581), .Z(n1583) );
  XNOR U1532 ( .A(n1584), .B(n1585), .Z(n1581) );
  AND U1533 ( .A(n199), .B(n1580), .Z(n1585) );
  XNOR U1534 ( .A(n1584), .B(n1578), .Z(n1580) );
  XOR U1535 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n1586), .Z(n1578) );
  AND U1536 ( .A(n213), .B(n1587), .Z(n1586) );
  XNOR U1537 ( .A(n1588), .B(n1589), .Z(n1584) );
  AND U1538 ( .A(n206), .B(n1590), .Z(n1589) );
  XOR U1539 ( .A(p_input[443]), .B(n1588), .Z(n1590) );
  XNOR U1540 ( .A(n1591), .B(n1592), .Z(n1588) );
  AND U1541 ( .A(n210), .B(n1587), .Z(n1592) );
  XOR U1542 ( .A(n1593), .B(n1591), .Z(n1587) );
  IV U1543 ( .A(\knn_comb_/min_val_out[0][27] ), .Z(n1593) );
  IV U1544 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .Z(n1591) );
  XOR U1545 ( .A(n21), .B(n1594), .Z(o[26]) );
  AND U1546 ( .A(n58), .B(n1595), .Z(n21) );
  XOR U1547 ( .A(n22), .B(n1594), .Z(n1595) );
  XOR U1548 ( .A(n1596), .B(n1597), .Z(n1594) );
  AND U1549 ( .A(n70), .B(n1598), .Z(n1597) );
  XOR U1550 ( .A(n1599), .B(n1600), .Z(n22) );
  AND U1551 ( .A(n62), .B(n1601), .Z(n1600) );
  XOR U1552 ( .A(p_input[26]), .B(n1599), .Z(n1601) );
  XNOR U1553 ( .A(n1602), .B(n1603), .Z(n1599) );
  AND U1554 ( .A(n66), .B(n1598), .Z(n1603) );
  XNOR U1555 ( .A(n1602), .B(n1596), .Z(n1598) );
  XOR U1556 ( .A(n1604), .B(n1605), .Z(n1596) );
  AND U1557 ( .A(n82), .B(n1606), .Z(n1605) );
  XNOR U1558 ( .A(n1607), .B(n1608), .Z(n1602) );
  AND U1559 ( .A(n74), .B(n1609), .Z(n1608) );
  XOR U1560 ( .A(p_input[58]), .B(n1607), .Z(n1609) );
  XNOR U1561 ( .A(n1610), .B(n1611), .Z(n1607) );
  AND U1562 ( .A(n78), .B(n1606), .Z(n1611) );
  XNOR U1563 ( .A(n1610), .B(n1604), .Z(n1606) );
  XOR U1564 ( .A(n1612), .B(n1613), .Z(n1604) );
  AND U1565 ( .A(n93), .B(n1614), .Z(n1613) );
  XNOR U1566 ( .A(n1615), .B(n1616), .Z(n1610) );
  AND U1567 ( .A(n85), .B(n1617), .Z(n1616) );
  XOR U1568 ( .A(p_input[90]), .B(n1615), .Z(n1617) );
  XNOR U1569 ( .A(n1618), .B(n1619), .Z(n1615) );
  AND U1570 ( .A(n89), .B(n1614), .Z(n1619) );
  XNOR U1571 ( .A(n1618), .B(n1612), .Z(n1614) );
  XOR U1572 ( .A(n1620), .B(n1621), .Z(n1612) );
  AND U1573 ( .A(n104), .B(n1622), .Z(n1621) );
  XNOR U1574 ( .A(n1623), .B(n1624), .Z(n1618) );
  AND U1575 ( .A(n96), .B(n1625), .Z(n1624) );
  XOR U1576 ( .A(p_input[122]), .B(n1623), .Z(n1625) );
  XNOR U1577 ( .A(n1626), .B(n1627), .Z(n1623) );
  AND U1578 ( .A(n100), .B(n1622), .Z(n1627) );
  XNOR U1579 ( .A(n1626), .B(n1620), .Z(n1622) );
  XOR U1580 ( .A(n1628), .B(n1629), .Z(n1620) );
  AND U1581 ( .A(n115), .B(n1630), .Z(n1629) );
  XNOR U1582 ( .A(n1631), .B(n1632), .Z(n1626) );
  AND U1583 ( .A(n107), .B(n1633), .Z(n1632) );
  XOR U1584 ( .A(p_input[154]), .B(n1631), .Z(n1633) );
  XNOR U1585 ( .A(n1634), .B(n1635), .Z(n1631) );
  AND U1586 ( .A(n111), .B(n1630), .Z(n1635) );
  XNOR U1587 ( .A(n1634), .B(n1628), .Z(n1630) );
  XOR U1588 ( .A(n1636), .B(n1637), .Z(n1628) );
  AND U1589 ( .A(n126), .B(n1638), .Z(n1637) );
  XNOR U1590 ( .A(n1639), .B(n1640), .Z(n1634) );
  AND U1591 ( .A(n118), .B(n1641), .Z(n1640) );
  XOR U1592 ( .A(p_input[186]), .B(n1639), .Z(n1641) );
  XNOR U1593 ( .A(n1642), .B(n1643), .Z(n1639) );
  AND U1594 ( .A(n122), .B(n1638), .Z(n1643) );
  XNOR U1595 ( .A(n1642), .B(n1636), .Z(n1638) );
  XOR U1596 ( .A(n1644), .B(n1645), .Z(n1636) );
  AND U1597 ( .A(n137), .B(n1646), .Z(n1645) );
  XNOR U1598 ( .A(n1647), .B(n1648), .Z(n1642) );
  AND U1599 ( .A(n129), .B(n1649), .Z(n1648) );
  XOR U1600 ( .A(p_input[218]), .B(n1647), .Z(n1649) );
  XNOR U1601 ( .A(n1650), .B(n1651), .Z(n1647) );
  AND U1602 ( .A(n133), .B(n1646), .Z(n1651) );
  XNOR U1603 ( .A(n1650), .B(n1644), .Z(n1646) );
  XOR U1604 ( .A(n1652), .B(n1653), .Z(n1644) );
  AND U1605 ( .A(n148), .B(n1654), .Z(n1653) );
  XNOR U1606 ( .A(n1655), .B(n1656), .Z(n1650) );
  AND U1607 ( .A(n140), .B(n1657), .Z(n1656) );
  XOR U1608 ( .A(p_input[250]), .B(n1655), .Z(n1657) );
  XNOR U1609 ( .A(n1658), .B(n1659), .Z(n1655) );
  AND U1610 ( .A(n144), .B(n1654), .Z(n1659) );
  XNOR U1611 ( .A(n1658), .B(n1652), .Z(n1654) );
  XOR U1612 ( .A(n1660), .B(n1661), .Z(n1652) );
  AND U1613 ( .A(n159), .B(n1662), .Z(n1661) );
  XNOR U1614 ( .A(n1663), .B(n1664), .Z(n1658) );
  AND U1615 ( .A(n151), .B(n1665), .Z(n1664) );
  XOR U1616 ( .A(p_input[282]), .B(n1663), .Z(n1665) );
  XNOR U1617 ( .A(n1666), .B(n1667), .Z(n1663) );
  AND U1618 ( .A(n155), .B(n1662), .Z(n1667) );
  XNOR U1619 ( .A(n1666), .B(n1660), .Z(n1662) );
  XOR U1620 ( .A(n1668), .B(n1669), .Z(n1660) );
  AND U1621 ( .A(n170), .B(n1670), .Z(n1669) );
  XNOR U1622 ( .A(n1671), .B(n1672), .Z(n1666) );
  AND U1623 ( .A(n162), .B(n1673), .Z(n1672) );
  XOR U1624 ( .A(p_input[314]), .B(n1671), .Z(n1673) );
  XNOR U1625 ( .A(n1674), .B(n1675), .Z(n1671) );
  AND U1626 ( .A(n166), .B(n1670), .Z(n1675) );
  XNOR U1627 ( .A(n1674), .B(n1668), .Z(n1670) );
  XOR U1628 ( .A(n1676), .B(n1677), .Z(n1668) );
  AND U1629 ( .A(n181), .B(n1678), .Z(n1677) );
  XNOR U1630 ( .A(n1679), .B(n1680), .Z(n1674) );
  AND U1631 ( .A(n173), .B(n1681), .Z(n1680) );
  XOR U1632 ( .A(p_input[346]), .B(n1679), .Z(n1681) );
  XNOR U1633 ( .A(n1682), .B(n1683), .Z(n1679) );
  AND U1634 ( .A(n177), .B(n1678), .Z(n1683) );
  XNOR U1635 ( .A(n1682), .B(n1676), .Z(n1678) );
  XOR U1636 ( .A(n1684), .B(n1685), .Z(n1676) );
  AND U1637 ( .A(n192), .B(n1686), .Z(n1685) );
  XNOR U1638 ( .A(n1687), .B(n1688), .Z(n1682) );
  AND U1639 ( .A(n184), .B(n1689), .Z(n1688) );
  XOR U1640 ( .A(p_input[378]), .B(n1687), .Z(n1689) );
  XNOR U1641 ( .A(n1690), .B(n1691), .Z(n1687) );
  AND U1642 ( .A(n188), .B(n1686), .Z(n1691) );
  XNOR U1643 ( .A(n1690), .B(n1684), .Z(n1686) );
  XOR U1644 ( .A(n1692), .B(n1693), .Z(n1684) );
  AND U1645 ( .A(n203), .B(n1694), .Z(n1693) );
  XNOR U1646 ( .A(n1695), .B(n1696), .Z(n1690) );
  AND U1647 ( .A(n195), .B(n1697), .Z(n1696) );
  XOR U1648 ( .A(p_input[410]), .B(n1695), .Z(n1697) );
  XNOR U1649 ( .A(n1698), .B(n1699), .Z(n1695) );
  AND U1650 ( .A(n199), .B(n1694), .Z(n1699) );
  XNOR U1651 ( .A(n1698), .B(n1692), .Z(n1694) );
  XOR U1652 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n1700), .Z(n1692) );
  AND U1653 ( .A(n213), .B(n1701), .Z(n1700) );
  XNOR U1654 ( .A(n1702), .B(n1703), .Z(n1698) );
  AND U1655 ( .A(n206), .B(n1704), .Z(n1703) );
  XOR U1656 ( .A(p_input[442]), .B(n1702), .Z(n1704) );
  XNOR U1657 ( .A(n1705), .B(n1706), .Z(n1702) );
  AND U1658 ( .A(n210), .B(n1701), .Z(n1706) );
  XOR U1659 ( .A(\knn_comb_/min_val_out[0][26] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .Z(n1701) );
  XOR U1660 ( .A(n23), .B(n1707), .Z(o[25]) );
  AND U1661 ( .A(n58), .B(n1708), .Z(n23) );
  XOR U1662 ( .A(n24), .B(n1707), .Z(n1708) );
  XOR U1663 ( .A(n1709), .B(n1710), .Z(n1707) );
  AND U1664 ( .A(n70), .B(n1711), .Z(n1710) );
  XOR U1665 ( .A(n1712), .B(n1713), .Z(n24) );
  AND U1666 ( .A(n62), .B(n1714), .Z(n1713) );
  XOR U1667 ( .A(p_input[25]), .B(n1712), .Z(n1714) );
  XNOR U1668 ( .A(n1715), .B(n1716), .Z(n1712) );
  AND U1669 ( .A(n66), .B(n1711), .Z(n1716) );
  XNOR U1670 ( .A(n1715), .B(n1709), .Z(n1711) );
  XOR U1671 ( .A(n1717), .B(n1718), .Z(n1709) );
  AND U1672 ( .A(n82), .B(n1719), .Z(n1718) );
  XNOR U1673 ( .A(n1720), .B(n1721), .Z(n1715) );
  AND U1674 ( .A(n74), .B(n1722), .Z(n1721) );
  XOR U1675 ( .A(p_input[57]), .B(n1720), .Z(n1722) );
  XNOR U1676 ( .A(n1723), .B(n1724), .Z(n1720) );
  AND U1677 ( .A(n78), .B(n1719), .Z(n1724) );
  XNOR U1678 ( .A(n1723), .B(n1717), .Z(n1719) );
  XOR U1679 ( .A(n1725), .B(n1726), .Z(n1717) );
  AND U1680 ( .A(n93), .B(n1727), .Z(n1726) );
  XNOR U1681 ( .A(n1728), .B(n1729), .Z(n1723) );
  AND U1682 ( .A(n85), .B(n1730), .Z(n1729) );
  XOR U1683 ( .A(p_input[89]), .B(n1728), .Z(n1730) );
  XNOR U1684 ( .A(n1731), .B(n1732), .Z(n1728) );
  AND U1685 ( .A(n89), .B(n1727), .Z(n1732) );
  XNOR U1686 ( .A(n1731), .B(n1725), .Z(n1727) );
  XOR U1687 ( .A(n1733), .B(n1734), .Z(n1725) );
  AND U1688 ( .A(n104), .B(n1735), .Z(n1734) );
  XNOR U1689 ( .A(n1736), .B(n1737), .Z(n1731) );
  AND U1690 ( .A(n96), .B(n1738), .Z(n1737) );
  XOR U1691 ( .A(p_input[121]), .B(n1736), .Z(n1738) );
  XNOR U1692 ( .A(n1739), .B(n1740), .Z(n1736) );
  AND U1693 ( .A(n100), .B(n1735), .Z(n1740) );
  XNOR U1694 ( .A(n1739), .B(n1733), .Z(n1735) );
  XOR U1695 ( .A(n1741), .B(n1742), .Z(n1733) );
  AND U1696 ( .A(n115), .B(n1743), .Z(n1742) );
  XNOR U1697 ( .A(n1744), .B(n1745), .Z(n1739) );
  AND U1698 ( .A(n107), .B(n1746), .Z(n1745) );
  XOR U1699 ( .A(p_input[153]), .B(n1744), .Z(n1746) );
  XNOR U1700 ( .A(n1747), .B(n1748), .Z(n1744) );
  AND U1701 ( .A(n111), .B(n1743), .Z(n1748) );
  XNOR U1702 ( .A(n1747), .B(n1741), .Z(n1743) );
  XOR U1703 ( .A(n1749), .B(n1750), .Z(n1741) );
  AND U1704 ( .A(n126), .B(n1751), .Z(n1750) );
  XNOR U1705 ( .A(n1752), .B(n1753), .Z(n1747) );
  AND U1706 ( .A(n118), .B(n1754), .Z(n1753) );
  XOR U1707 ( .A(p_input[185]), .B(n1752), .Z(n1754) );
  XNOR U1708 ( .A(n1755), .B(n1756), .Z(n1752) );
  AND U1709 ( .A(n122), .B(n1751), .Z(n1756) );
  XNOR U1710 ( .A(n1755), .B(n1749), .Z(n1751) );
  XOR U1711 ( .A(n1757), .B(n1758), .Z(n1749) );
  AND U1712 ( .A(n137), .B(n1759), .Z(n1758) );
  XNOR U1713 ( .A(n1760), .B(n1761), .Z(n1755) );
  AND U1714 ( .A(n129), .B(n1762), .Z(n1761) );
  XOR U1715 ( .A(p_input[217]), .B(n1760), .Z(n1762) );
  XNOR U1716 ( .A(n1763), .B(n1764), .Z(n1760) );
  AND U1717 ( .A(n133), .B(n1759), .Z(n1764) );
  XNOR U1718 ( .A(n1763), .B(n1757), .Z(n1759) );
  XOR U1719 ( .A(n1765), .B(n1766), .Z(n1757) );
  AND U1720 ( .A(n148), .B(n1767), .Z(n1766) );
  XNOR U1721 ( .A(n1768), .B(n1769), .Z(n1763) );
  AND U1722 ( .A(n140), .B(n1770), .Z(n1769) );
  XOR U1723 ( .A(p_input[249]), .B(n1768), .Z(n1770) );
  XNOR U1724 ( .A(n1771), .B(n1772), .Z(n1768) );
  AND U1725 ( .A(n144), .B(n1767), .Z(n1772) );
  XNOR U1726 ( .A(n1771), .B(n1765), .Z(n1767) );
  XOR U1727 ( .A(n1773), .B(n1774), .Z(n1765) );
  AND U1728 ( .A(n159), .B(n1775), .Z(n1774) );
  XNOR U1729 ( .A(n1776), .B(n1777), .Z(n1771) );
  AND U1730 ( .A(n151), .B(n1778), .Z(n1777) );
  XOR U1731 ( .A(p_input[281]), .B(n1776), .Z(n1778) );
  XNOR U1732 ( .A(n1779), .B(n1780), .Z(n1776) );
  AND U1733 ( .A(n155), .B(n1775), .Z(n1780) );
  XNOR U1734 ( .A(n1779), .B(n1773), .Z(n1775) );
  XOR U1735 ( .A(n1781), .B(n1782), .Z(n1773) );
  AND U1736 ( .A(n170), .B(n1783), .Z(n1782) );
  XNOR U1737 ( .A(n1784), .B(n1785), .Z(n1779) );
  AND U1738 ( .A(n162), .B(n1786), .Z(n1785) );
  XOR U1739 ( .A(p_input[313]), .B(n1784), .Z(n1786) );
  XNOR U1740 ( .A(n1787), .B(n1788), .Z(n1784) );
  AND U1741 ( .A(n166), .B(n1783), .Z(n1788) );
  XNOR U1742 ( .A(n1787), .B(n1781), .Z(n1783) );
  XOR U1743 ( .A(n1789), .B(n1790), .Z(n1781) );
  AND U1744 ( .A(n181), .B(n1791), .Z(n1790) );
  XNOR U1745 ( .A(n1792), .B(n1793), .Z(n1787) );
  AND U1746 ( .A(n173), .B(n1794), .Z(n1793) );
  XOR U1747 ( .A(p_input[345]), .B(n1792), .Z(n1794) );
  XNOR U1748 ( .A(n1795), .B(n1796), .Z(n1792) );
  AND U1749 ( .A(n177), .B(n1791), .Z(n1796) );
  XNOR U1750 ( .A(n1795), .B(n1789), .Z(n1791) );
  XOR U1751 ( .A(n1797), .B(n1798), .Z(n1789) );
  AND U1752 ( .A(n192), .B(n1799), .Z(n1798) );
  XNOR U1753 ( .A(n1800), .B(n1801), .Z(n1795) );
  AND U1754 ( .A(n184), .B(n1802), .Z(n1801) );
  XOR U1755 ( .A(p_input[377]), .B(n1800), .Z(n1802) );
  XNOR U1756 ( .A(n1803), .B(n1804), .Z(n1800) );
  AND U1757 ( .A(n188), .B(n1799), .Z(n1804) );
  XNOR U1758 ( .A(n1803), .B(n1797), .Z(n1799) );
  XOR U1759 ( .A(n1805), .B(n1806), .Z(n1797) );
  AND U1760 ( .A(n203), .B(n1807), .Z(n1806) );
  XNOR U1761 ( .A(n1808), .B(n1809), .Z(n1803) );
  AND U1762 ( .A(n195), .B(n1810), .Z(n1809) );
  XOR U1763 ( .A(p_input[409]), .B(n1808), .Z(n1810) );
  XNOR U1764 ( .A(n1811), .B(n1812), .Z(n1808) );
  AND U1765 ( .A(n199), .B(n1807), .Z(n1812) );
  XNOR U1766 ( .A(n1811), .B(n1805), .Z(n1807) );
  XOR U1767 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n1813), .Z(n1805) );
  AND U1768 ( .A(n213), .B(n1814), .Z(n1813) );
  XNOR U1769 ( .A(n1815), .B(n1816), .Z(n1811) );
  AND U1770 ( .A(n206), .B(n1817), .Z(n1816) );
  XOR U1771 ( .A(p_input[441]), .B(n1815), .Z(n1817) );
  XNOR U1772 ( .A(n1818), .B(n1819), .Z(n1815) );
  AND U1773 ( .A(n210), .B(n1814), .Z(n1819) );
  XOR U1774 ( .A(\knn_comb_/min_val_out[0][25] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .Z(n1814) );
  XOR U1775 ( .A(n25), .B(n1820), .Z(o[24]) );
  AND U1776 ( .A(n58), .B(n1821), .Z(n25) );
  XOR U1777 ( .A(n26), .B(n1820), .Z(n1821) );
  XOR U1778 ( .A(n1822), .B(n1823), .Z(n1820) );
  AND U1779 ( .A(n70), .B(n1824), .Z(n1823) );
  XOR U1780 ( .A(n1825), .B(n1826), .Z(n26) );
  AND U1781 ( .A(n62), .B(n1827), .Z(n1826) );
  XOR U1782 ( .A(p_input[24]), .B(n1825), .Z(n1827) );
  XNOR U1783 ( .A(n1828), .B(n1829), .Z(n1825) );
  AND U1784 ( .A(n66), .B(n1824), .Z(n1829) );
  XNOR U1785 ( .A(n1828), .B(n1822), .Z(n1824) );
  XOR U1786 ( .A(n1830), .B(n1831), .Z(n1822) );
  AND U1787 ( .A(n82), .B(n1832), .Z(n1831) );
  XNOR U1788 ( .A(n1833), .B(n1834), .Z(n1828) );
  AND U1789 ( .A(n74), .B(n1835), .Z(n1834) );
  XOR U1790 ( .A(p_input[56]), .B(n1833), .Z(n1835) );
  XNOR U1791 ( .A(n1836), .B(n1837), .Z(n1833) );
  AND U1792 ( .A(n78), .B(n1832), .Z(n1837) );
  XNOR U1793 ( .A(n1836), .B(n1830), .Z(n1832) );
  XOR U1794 ( .A(n1838), .B(n1839), .Z(n1830) );
  AND U1795 ( .A(n93), .B(n1840), .Z(n1839) );
  XNOR U1796 ( .A(n1841), .B(n1842), .Z(n1836) );
  AND U1797 ( .A(n85), .B(n1843), .Z(n1842) );
  XOR U1798 ( .A(p_input[88]), .B(n1841), .Z(n1843) );
  XNOR U1799 ( .A(n1844), .B(n1845), .Z(n1841) );
  AND U1800 ( .A(n89), .B(n1840), .Z(n1845) );
  XNOR U1801 ( .A(n1844), .B(n1838), .Z(n1840) );
  XOR U1802 ( .A(n1846), .B(n1847), .Z(n1838) );
  AND U1803 ( .A(n104), .B(n1848), .Z(n1847) );
  XNOR U1804 ( .A(n1849), .B(n1850), .Z(n1844) );
  AND U1805 ( .A(n96), .B(n1851), .Z(n1850) );
  XOR U1806 ( .A(p_input[120]), .B(n1849), .Z(n1851) );
  XNOR U1807 ( .A(n1852), .B(n1853), .Z(n1849) );
  AND U1808 ( .A(n100), .B(n1848), .Z(n1853) );
  XNOR U1809 ( .A(n1852), .B(n1846), .Z(n1848) );
  XOR U1810 ( .A(n1854), .B(n1855), .Z(n1846) );
  AND U1811 ( .A(n115), .B(n1856), .Z(n1855) );
  XNOR U1812 ( .A(n1857), .B(n1858), .Z(n1852) );
  AND U1813 ( .A(n107), .B(n1859), .Z(n1858) );
  XOR U1814 ( .A(p_input[152]), .B(n1857), .Z(n1859) );
  XNOR U1815 ( .A(n1860), .B(n1861), .Z(n1857) );
  AND U1816 ( .A(n111), .B(n1856), .Z(n1861) );
  XNOR U1817 ( .A(n1860), .B(n1854), .Z(n1856) );
  XOR U1818 ( .A(n1862), .B(n1863), .Z(n1854) );
  AND U1819 ( .A(n126), .B(n1864), .Z(n1863) );
  XNOR U1820 ( .A(n1865), .B(n1866), .Z(n1860) );
  AND U1821 ( .A(n118), .B(n1867), .Z(n1866) );
  XOR U1822 ( .A(p_input[184]), .B(n1865), .Z(n1867) );
  XNOR U1823 ( .A(n1868), .B(n1869), .Z(n1865) );
  AND U1824 ( .A(n122), .B(n1864), .Z(n1869) );
  XNOR U1825 ( .A(n1868), .B(n1862), .Z(n1864) );
  XOR U1826 ( .A(n1870), .B(n1871), .Z(n1862) );
  AND U1827 ( .A(n137), .B(n1872), .Z(n1871) );
  XNOR U1828 ( .A(n1873), .B(n1874), .Z(n1868) );
  AND U1829 ( .A(n129), .B(n1875), .Z(n1874) );
  XOR U1830 ( .A(p_input[216]), .B(n1873), .Z(n1875) );
  XNOR U1831 ( .A(n1876), .B(n1877), .Z(n1873) );
  AND U1832 ( .A(n133), .B(n1872), .Z(n1877) );
  XNOR U1833 ( .A(n1876), .B(n1870), .Z(n1872) );
  XOR U1834 ( .A(n1878), .B(n1879), .Z(n1870) );
  AND U1835 ( .A(n148), .B(n1880), .Z(n1879) );
  XNOR U1836 ( .A(n1881), .B(n1882), .Z(n1876) );
  AND U1837 ( .A(n140), .B(n1883), .Z(n1882) );
  XOR U1838 ( .A(p_input[248]), .B(n1881), .Z(n1883) );
  XNOR U1839 ( .A(n1884), .B(n1885), .Z(n1881) );
  AND U1840 ( .A(n144), .B(n1880), .Z(n1885) );
  XNOR U1841 ( .A(n1884), .B(n1878), .Z(n1880) );
  XOR U1842 ( .A(n1886), .B(n1887), .Z(n1878) );
  AND U1843 ( .A(n159), .B(n1888), .Z(n1887) );
  XNOR U1844 ( .A(n1889), .B(n1890), .Z(n1884) );
  AND U1845 ( .A(n151), .B(n1891), .Z(n1890) );
  XOR U1846 ( .A(p_input[280]), .B(n1889), .Z(n1891) );
  XNOR U1847 ( .A(n1892), .B(n1893), .Z(n1889) );
  AND U1848 ( .A(n155), .B(n1888), .Z(n1893) );
  XNOR U1849 ( .A(n1892), .B(n1886), .Z(n1888) );
  XOR U1850 ( .A(n1894), .B(n1895), .Z(n1886) );
  AND U1851 ( .A(n170), .B(n1896), .Z(n1895) );
  XNOR U1852 ( .A(n1897), .B(n1898), .Z(n1892) );
  AND U1853 ( .A(n162), .B(n1899), .Z(n1898) );
  XOR U1854 ( .A(p_input[312]), .B(n1897), .Z(n1899) );
  XNOR U1855 ( .A(n1900), .B(n1901), .Z(n1897) );
  AND U1856 ( .A(n166), .B(n1896), .Z(n1901) );
  XNOR U1857 ( .A(n1900), .B(n1894), .Z(n1896) );
  XOR U1858 ( .A(n1902), .B(n1903), .Z(n1894) );
  AND U1859 ( .A(n181), .B(n1904), .Z(n1903) );
  XNOR U1860 ( .A(n1905), .B(n1906), .Z(n1900) );
  AND U1861 ( .A(n173), .B(n1907), .Z(n1906) );
  XOR U1862 ( .A(p_input[344]), .B(n1905), .Z(n1907) );
  XNOR U1863 ( .A(n1908), .B(n1909), .Z(n1905) );
  AND U1864 ( .A(n177), .B(n1904), .Z(n1909) );
  XNOR U1865 ( .A(n1908), .B(n1902), .Z(n1904) );
  XOR U1866 ( .A(n1910), .B(n1911), .Z(n1902) );
  AND U1867 ( .A(n192), .B(n1912), .Z(n1911) );
  XNOR U1868 ( .A(n1913), .B(n1914), .Z(n1908) );
  AND U1869 ( .A(n184), .B(n1915), .Z(n1914) );
  XOR U1870 ( .A(p_input[376]), .B(n1913), .Z(n1915) );
  XNOR U1871 ( .A(n1916), .B(n1917), .Z(n1913) );
  AND U1872 ( .A(n188), .B(n1912), .Z(n1917) );
  XNOR U1873 ( .A(n1916), .B(n1910), .Z(n1912) );
  XOR U1874 ( .A(n1918), .B(n1919), .Z(n1910) );
  AND U1875 ( .A(n203), .B(n1920), .Z(n1919) );
  XNOR U1876 ( .A(n1921), .B(n1922), .Z(n1916) );
  AND U1877 ( .A(n195), .B(n1923), .Z(n1922) );
  XOR U1878 ( .A(p_input[408]), .B(n1921), .Z(n1923) );
  XNOR U1879 ( .A(n1924), .B(n1925), .Z(n1921) );
  AND U1880 ( .A(n199), .B(n1920), .Z(n1925) );
  XNOR U1881 ( .A(n1924), .B(n1918), .Z(n1920) );
  XOR U1882 ( .A(\knn_comb_/min_val_out[0][24] ), .B(n1926), .Z(n1918) );
  AND U1883 ( .A(n213), .B(n1927), .Z(n1926) );
  XNOR U1884 ( .A(n1928), .B(n1929), .Z(n1924) );
  AND U1885 ( .A(n206), .B(n1930), .Z(n1929) );
  XOR U1886 ( .A(p_input[440]), .B(n1928), .Z(n1930) );
  XNOR U1887 ( .A(n1931), .B(n1932), .Z(n1928) );
  AND U1888 ( .A(n210), .B(n1927), .Z(n1932) );
  XOR U1889 ( .A(\knn_comb_/min_val_out[0][24] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .Z(n1927) );
  XOR U1890 ( .A(n27), .B(n1933), .Z(o[23]) );
  AND U1891 ( .A(n58), .B(n1934), .Z(n27) );
  XOR U1892 ( .A(n28), .B(n1933), .Z(n1934) );
  XOR U1893 ( .A(n1935), .B(n1936), .Z(n1933) );
  AND U1894 ( .A(n70), .B(n1937), .Z(n1936) );
  XOR U1895 ( .A(n1938), .B(n1939), .Z(n28) );
  AND U1896 ( .A(n62), .B(n1940), .Z(n1939) );
  XOR U1897 ( .A(p_input[23]), .B(n1938), .Z(n1940) );
  XNOR U1898 ( .A(n1941), .B(n1942), .Z(n1938) );
  AND U1899 ( .A(n66), .B(n1937), .Z(n1942) );
  XNOR U1900 ( .A(n1941), .B(n1935), .Z(n1937) );
  XOR U1901 ( .A(n1943), .B(n1944), .Z(n1935) );
  AND U1902 ( .A(n82), .B(n1945), .Z(n1944) );
  XNOR U1903 ( .A(n1946), .B(n1947), .Z(n1941) );
  AND U1904 ( .A(n74), .B(n1948), .Z(n1947) );
  XOR U1905 ( .A(p_input[55]), .B(n1946), .Z(n1948) );
  XNOR U1906 ( .A(n1949), .B(n1950), .Z(n1946) );
  AND U1907 ( .A(n78), .B(n1945), .Z(n1950) );
  XNOR U1908 ( .A(n1949), .B(n1943), .Z(n1945) );
  XOR U1909 ( .A(n1951), .B(n1952), .Z(n1943) );
  AND U1910 ( .A(n93), .B(n1953), .Z(n1952) );
  XNOR U1911 ( .A(n1954), .B(n1955), .Z(n1949) );
  AND U1912 ( .A(n85), .B(n1956), .Z(n1955) );
  XOR U1913 ( .A(p_input[87]), .B(n1954), .Z(n1956) );
  XNOR U1914 ( .A(n1957), .B(n1958), .Z(n1954) );
  AND U1915 ( .A(n89), .B(n1953), .Z(n1958) );
  XNOR U1916 ( .A(n1957), .B(n1951), .Z(n1953) );
  XOR U1917 ( .A(n1959), .B(n1960), .Z(n1951) );
  AND U1918 ( .A(n104), .B(n1961), .Z(n1960) );
  XNOR U1919 ( .A(n1962), .B(n1963), .Z(n1957) );
  AND U1920 ( .A(n96), .B(n1964), .Z(n1963) );
  XOR U1921 ( .A(p_input[119]), .B(n1962), .Z(n1964) );
  XNOR U1922 ( .A(n1965), .B(n1966), .Z(n1962) );
  AND U1923 ( .A(n100), .B(n1961), .Z(n1966) );
  XNOR U1924 ( .A(n1965), .B(n1959), .Z(n1961) );
  XOR U1925 ( .A(n1967), .B(n1968), .Z(n1959) );
  AND U1926 ( .A(n115), .B(n1969), .Z(n1968) );
  XNOR U1927 ( .A(n1970), .B(n1971), .Z(n1965) );
  AND U1928 ( .A(n107), .B(n1972), .Z(n1971) );
  XOR U1929 ( .A(p_input[151]), .B(n1970), .Z(n1972) );
  XNOR U1930 ( .A(n1973), .B(n1974), .Z(n1970) );
  AND U1931 ( .A(n111), .B(n1969), .Z(n1974) );
  XNOR U1932 ( .A(n1973), .B(n1967), .Z(n1969) );
  XOR U1933 ( .A(n1975), .B(n1976), .Z(n1967) );
  AND U1934 ( .A(n126), .B(n1977), .Z(n1976) );
  XNOR U1935 ( .A(n1978), .B(n1979), .Z(n1973) );
  AND U1936 ( .A(n118), .B(n1980), .Z(n1979) );
  XOR U1937 ( .A(p_input[183]), .B(n1978), .Z(n1980) );
  XNOR U1938 ( .A(n1981), .B(n1982), .Z(n1978) );
  AND U1939 ( .A(n122), .B(n1977), .Z(n1982) );
  XNOR U1940 ( .A(n1981), .B(n1975), .Z(n1977) );
  XOR U1941 ( .A(n1983), .B(n1984), .Z(n1975) );
  AND U1942 ( .A(n137), .B(n1985), .Z(n1984) );
  XNOR U1943 ( .A(n1986), .B(n1987), .Z(n1981) );
  AND U1944 ( .A(n129), .B(n1988), .Z(n1987) );
  XOR U1945 ( .A(p_input[215]), .B(n1986), .Z(n1988) );
  XNOR U1946 ( .A(n1989), .B(n1990), .Z(n1986) );
  AND U1947 ( .A(n133), .B(n1985), .Z(n1990) );
  XNOR U1948 ( .A(n1989), .B(n1983), .Z(n1985) );
  XOR U1949 ( .A(n1991), .B(n1992), .Z(n1983) );
  AND U1950 ( .A(n148), .B(n1993), .Z(n1992) );
  XNOR U1951 ( .A(n1994), .B(n1995), .Z(n1989) );
  AND U1952 ( .A(n140), .B(n1996), .Z(n1995) );
  XOR U1953 ( .A(p_input[247]), .B(n1994), .Z(n1996) );
  XNOR U1954 ( .A(n1997), .B(n1998), .Z(n1994) );
  AND U1955 ( .A(n144), .B(n1993), .Z(n1998) );
  XNOR U1956 ( .A(n1997), .B(n1991), .Z(n1993) );
  XOR U1957 ( .A(n1999), .B(n2000), .Z(n1991) );
  AND U1958 ( .A(n159), .B(n2001), .Z(n2000) );
  XNOR U1959 ( .A(n2002), .B(n2003), .Z(n1997) );
  AND U1960 ( .A(n151), .B(n2004), .Z(n2003) );
  XOR U1961 ( .A(p_input[279]), .B(n2002), .Z(n2004) );
  XNOR U1962 ( .A(n2005), .B(n2006), .Z(n2002) );
  AND U1963 ( .A(n155), .B(n2001), .Z(n2006) );
  XNOR U1964 ( .A(n2005), .B(n1999), .Z(n2001) );
  XOR U1965 ( .A(n2007), .B(n2008), .Z(n1999) );
  AND U1966 ( .A(n170), .B(n2009), .Z(n2008) );
  XNOR U1967 ( .A(n2010), .B(n2011), .Z(n2005) );
  AND U1968 ( .A(n162), .B(n2012), .Z(n2011) );
  XOR U1969 ( .A(p_input[311]), .B(n2010), .Z(n2012) );
  XNOR U1970 ( .A(n2013), .B(n2014), .Z(n2010) );
  AND U1971 ( .A(n166), .B(n2009), .Z(n2014) );
  XNOR U1972 ( .A(n2013), .B(n2007), .Z(n2009) );
  XOR U1973 ( .A(n2015), .B(n2016), .Z(n2007) );
  AND U1974 ( .A(n181), .B(n2017), .Z(n2016) );
  XNOR U1975 ( .A(n2018), .B(n2019), .Z(n2013) );
  AND U1976 ( .A(n173), .B(n2020), .Z(n2019) );
  XOR U1977 ( .A(p_input[343]), .B(n2018), .Z(n2020) );
  XNOR U1978 ( .A(n2021), .B(n2022), .Z(n2018) );
  AND U1979 ( .A(n177), .B(n2017), .Z(n2022) );
  XNOR U1980 ( .A(n2021), .B(n2015), .Z(n2017) );
  XOR U1981 ( .A(n2023), .B(n2024), .Z(n2015) );
  AND U1982 ( .A(n192), .B(n2025), .Z(n2024) );
  XNOR U1983 ( .A(n2026), .B(n2027), .Z(n2021) );
  AND U1984 ( .A(n184), .B(n2028), .Z(n2027) );
  XOR U1985 ( .A(p_input[375]), .B(n2026), .Z(n2028) );
  XNOR U1986 ( .A(n2029), .B(n2030), .Z(n2026) );
  AND U1987 ( .A(n188), .B(n2025), .Z(n2030) );
  XNOR U1988 ( .A(n2029), .B(n2023), .Z(n2025) );
  XOR U1989 ( .A(n2031), .B(n2032), .Z(n2023) );
  AND U1990 ( .A(n203), .B(n2033), .Z(n2032) );
  XNOR U1991 ( .A(n2034), .B(n2035), .Z(n2029) );
  AND U1992 ( .A(n195), .B(n2036), .Z(n2035) );
  XOR U1993 ( .A(p_input[407]), .B(n2034), .Z(n2036) );
  XNOR U1994 ( .A(n2037), .B(n2038), .Z(n2034) );
  AND U1995 ( .A(n199), .B(n2033), .Z(n2038) );
  XNOR U1996 ( .A(n2037), .B(n2031), .Z(n2033) );
  XOR U1997 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n2039), .Z(n2031) );
  AND U1998 ( .A(n213), .B(n2040), .Z(n2039) );
  XNOR U1999 ( .A(n2041), .B(n2042), .Z(n2037) );
  AND U2000 ( .A(n206), .B(n2043), .Z(n2042) );
  XOR U2001 ( .A(p_input[439]), .B(n2041), .Z(n2043) );
  XNOR U2002 ( .A(n2044), .B(n2045), .Z(n2041) );
  AND U2003 ( .A(n210), .B(n2040), .Z(n2045) );
  XOR U2004 ( .A(n2046), .B(n2044), .Z(n2040) );
  IV U2005 ( .A(\knn_comb_/min_val_out[0][23] ), .Z(n2046) );
  IV U2006 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .Z(n2044) );
  XOR U2007 ( .A(n29), .B(n2047), .Z(o[22]) );
  AND U2008 ( .A(n58), .B(n2048), .Z(n29) );
  XOR U2009 ( .A(n30), .B(n2047), .Z(n2048) );
  XOR U2010 ( .A(n2049), .B(n2050), .Z(n2047) );
  AND U2011 ( .A(n70), .B(n2051), .Z(n2050) );
  XOR U2012 ( .A(n2052), .B(n2053), .Z(n30) );
  AND U2013 ( .A(n62), .B(n2054), .Z(n2053) );
  XOR U2014 ( .A(p_input[22]), .B(n2052), .Z(n2054) );
  XNOR U2015 ( .A(n2055), .B(n2056), .Z(n2052) );
  AND U2016 ( .A(n66), .B(n2051), .Z(n2056) );
  XNOR U2017 ( .A(n2055), .B(n2049), .Z(n2051) );
  XOR U2018 ( .A(n2057), .B(n2058), .Z(n2049) );
  AND U2019 ( .A(n82), .B(n2059), .Z(n2058) );
  XNOR U2020 ( .A(n2060), .B(n2061), .Z(n2055) );
  AND U2021 ( .A(n74), .B(n2062), .Z(n2061) );
  XOR U2022 ( .A(p_input[54]), .B(n2060), .Z(n2062) );
  XNOR U2023 ( .A(n2063), .B(n2064), .Z(n2060) );
  AND U2024 ( .A(n78), .B(n2059), .Z(n2064) );
  XNOR U2025 ( .A(n2063), .B(n2057), .Z(n2059) );
  XOR U2026 ( .A(n2065), .B(n2066), .Z(n2057) );
  AND U2027 ( .A(n93), .B(n2067), .Z(n2066) );
  XNOR U2028 ( .A(n2068), .B(n2069), .Z(n2063) );
  AND U2029 ( .A(n85), .B(n2070), .Z(n2069) );
  XOR U2030 ( .A(p_input[86]), .B(n2068), .Z(n2070) );
  XNOR U2031 ( .A(n2071), .B(n2072), .Z(n2068) );
  AND U2032 ( .A(n89), .B(n2067), .Z(n2072) );
  XNOR U2033 ( .A(n2071), .B(n2065), .Z(n2067) );
  XOR U2034 ( .A(n2073), .B(n2074), .Z(n2065) );
  AND U2035 ( .A(n104), .B(n2075), .Z(n2074) );
  XNOR U2036 ( .A(n2076), .B(n2077), .Z(n2071) );
  AND U2037 ( .A(n96), .B(n2078), .Z(n2077) );
  XOR U2038 ( .A(p_input[118]), .B(n2076), .Z(n2078) );
  XNOR U2039 ( .A(n2079), .B(n2080), .Z(n2076) );
  AND U2040 ( .A(n100), .B(n2075), .Z(n2080) );
  XNOR U2041 ( .A(n2079), .B(n2073), .Z(n2075) );
  XOR U2042 ( .A(n2081), .B(n2082), .Z(n2073) );
  AND U2043 ( .A(n115), .B(n2083), .Z(n2082) );
  XNOR U2044 ( .A(n2084), .B(n2085), .Z(n2079) );
  AND U2045 ( .A(n107), .B(n2086), .Z(n2085) );
  XOR U2046 ( .A(p_input[150]), .B(n2084), .Z(n2086) );
  XNOR U2047 ( .A(n2087), .B(n2088), .Z(n2084) );
  AND U2048 ( .A(n111), .B(n2083), .Z(n2088) );
  XNOR U2049 ( .A(n2087), .B(n2081), .Z(n2083) );
  XOR U2050 ( .A(n2089), .B(n2090), .Z(n2081) );
  AND U2051 ( .A(n126), .B(n2091), .Z(n2090) );
  XNOR U2052 ( .A(n2092), .B(n2093), .Z(n2087) );
  AND U2053 ( .A(n118), .B(n2094), .Z(n2093) );
  XOR U2054 ( .A(p_input[182]), .B(n2092), .Z(n2094) );
  XNOR U2055 ( .A(n2095), .B(n2096), .Z(n2092) );
  AND U2056 ( .A(n122), .B(n2091), .Z(n2096) );
  XNOR U2057 ( .A(n2095), .B(n2089), .Z(n2091) );
  XOR U2058 ( .A(n2097), .B(n2098), .Z(n2089) );
  AND U2059 ( .A(n137), .B(n2099), .Z(n2098) );
  XNOR U2060 ( .A(n2100), .B(n2101), .Z(n2095) );
  AND U2061 ( .A(n129), .B(n2102), .Z(n2101) );
  XOR U2062 ( .A(p_input[214]), .B(n2100), .Z(n2102) );
  XNOR U2063 ( .A(n2103), .B(n2104), .Z(n2100) );
  AND U2064 ( .A(n133), .B(n2099), .Z(n2104) );
  XNOR U2065 ( .A(n2103), .B(n2097), .Z(n2099) );
  XOR U2066 ( .A(n2105), .B(n2106), .Z(n2097) );
  AND U2067 ( .A(n148), .B(n2107), .Z(n2106) );
  XNOR U2068 ( .A(n2108), .B(n2109), .Z(n2103) );
  AND U2069 ( .A(n140), .B(n2110), .Z(n2109) );
  XOR U2070 ( .A(p_input[246]), .B(n2108), .Z(n2110) );
  XNOR U2071 ( .A(n2111), .B(n2112), .Z(n2108) );
  AND U2072 ( .A(n144), .B(n2107), .Z(n2112) );
  XNOR U2073 ( .A(n2111), .B(n2105), .Z(n2107) );
  XOR U2074 ( .A(n2113), .B(n2114), .Z(n2105) );
  AND U2075 ( .A(n159), .B(n2115), .Z(n2114) );
  XNOR U2076 ( .A(n2116), .B(n2117), .Z(n2111) );
  AND U2077 ( .A(n151), .B(n2118), .Z(n2117) );
  XOR U2078 ( .A(p_input[278]), .B(n2116), .Z(n2118) );
  XNOR U2079 ( .A(n2119), .B(n2120), .Z(n2116) );
  AND U2080 ( .A(n155), .B(n2115), .Z(n2120) );
  XNOR U2081 ( .A(n2119), .B(n2113), .Z(n2115) );
  XOR U2082 ( .A(n2121), .B(n2122), .Z(n2113) );
  AND U2083 ( .A(n170), .B(n2123), .Z(n2122) );
  XNOR U2084 ( .A(n2124), .B(n2125), .Z(n2119) );
  AND U2085 ( .A(n162), .B(n2126), .Z(n2125) );
  XOR U2086 ( .A(p_input[310]), .B(n2124), .Z(n2126) );
  XNOR U2087 ( .A(n2127), .B(n2128), .Z(n2124) );
  AND U2088 ( .A(n166), .B(n2123), .Z(n2128) );
  XNOR U2089 ( .A(n2127), .B(n2121), .Z(n2123) );
  XOR U2090 ( .A(n2129), .B(n2130), .Z(n2121) );
  AND U2091 ( .A(n181), .B(n2131), .Z(n2130) );
  XNOR U2092 ( .A(n2132), .B(n2133), .Z(n2127) );
  AND U2093 ( .A(n173), .B(n2134), .Z(n2133) );
  XOR U2094 ( .A(p_input[342]), .B(n2132), .Z(n2134) );
  XNOR U2095 ( .A(n2135), .B(n2136), .Z(n2132) );
  AND U2096 ( .A(n177), .B(n2131), .Z(n2136) );
  XNOR U2097 ( .A(n2135), .B(n2129), .Z(n2131) );
  XOR U2098 ( .A(n2137), .B(n2138), .Z(n2129) );
  AND U2099 ( .A(n192), .B(n2139), .Z(n2138) );
  XNOR U2100 ( .A(n2140), .B(n2141), .Z(n2135) );
  AND U2101 ( .A(n184), .B(n2142), .Z(n2141) );
  XOR U2102 ( .A(p_input[374]), .B(n2140), .Z(n2142) );
  XNOR U2103 ( .A(n2143), .B(n2144), .Z(n2140) );
  AND U2104 ( .A(n188), .B(n2139), .Z(n2144) );
  XNOR U2105 ( .A(n2143), .B(n2137), .Z(n2139) );
  XOR U2106 ( .A(n2145), .B(n2146), .Z(n2137) );
  AND U2107 ( .A(n203), .B(n2147), .Z(n2146) );
  XNOR U2108 ( .A(n2148), .B(n2149), .Z(n2143) );
  AND U2109 ( .A(n195), .B(n2150), .Z(n2149) );
  XOR U2110 ( .A(p_input[406]), .B(n2148), .Z(n2150) );
  XNOR U2111 ( .A(n2151), .B(n2152), .Z(n2148) );
  AND U2112 ( .A(n199), .B(n2147), .Z(n2152) );
  XNOR U2113 ( .A(n2151), .B(n2145), .Z(n2147) );
  XOR U2114 ( .A(\knn_comb_/min_val_out[0][22] ), .B(n2153), .Z(n2145) );
  AND U2115 ( .A(n213), .B(n2154), .Z(n2153) );
  XNOR U2116 ( .A(n2155), .B(n2156), .Z(n2151) );
  AND U2117 ( .A(n206), .B(n2157), .Z(n2156) );
  XOR U2118 ( .A(p_input[438]), .B(n2155), .Z(n2157) );
  XNOR U2119 ( .A(n2158), .B(n2159), .Z(n2155) );
  AND U2120 ( .A(n210), .B(n2154), .Z(n2159) );
  XOR U2121 ( .A(\knn_comb_/min_val_out[0][22] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .Z(n2154) );
  XOR U2122 ( .A(n31), .B(n2160), .Z(o[21]) );
  AND U2123 ( .A(n58), .B(n2161), .Z(n31) );
  XOR U2124 ( .A(n32), .B(n2160), .Z(n2161) );
  XOR U2125 ( .A(n2162), .B(n2163), .Z(n2160) );
  AND U2126 ( .A(n70), .B(n2164), .Z(n2163) );
  XOR U2127 ( .A(n2165), .B(n2166), .Z(n32) );
  AND U2128 ( .A(n62), .B(n2167), .Z(n2166) );
  XOR U2129 ( .A(p_input[21]), .B(n2165), .Z(n2167) );
  XNOR U2130 ( .A(n2168), .B(n2169), .Z(n2165) );
  AND U2131 ( .A(n66), .B(n2164), .Z(n2169) );
  XNOR U2132 ( .A(n2168), .B(n2162), .Z(n2164) );
  XOR U2133 ( .A(n2170), .B(n2171), .Z(n2162) );
  AND U2134 ( .A(n82), .B(n2172), .Z(n2171) );
  XNOR U2135 ( .A(n2173), .B(n2174), .Z(n2168) );
  AND U2136 ( .A(n74), .B(n2175), .Z(n2174) );
  XOR U2137 ( .A(p_input[53]), .B(n2173), .Z(n2175) );
  XNOR U2138 ( .A(n2176), .B(n2177), .Z(n2173) );
  AND U2139 ( .A(n78), .B(n2172), .Z(n2177) );
  XNOR U2140 ( .A(n2176), .B(n2170), .Z(n2172) );
  XOR U2141 ( .A(n2178), .B(n2179), .Z(n2170) );
  AND U2142 ( .A(n93), .B(n2180), .Z(n2179) );
  XNOR U2143 ( .A(n2181), .B(n2182), .Z(n2176) );
  AND U2144 ( .A(n85), .B(n2183), .Z(n2182) );
  XOR U2145 ( .A(p_input[85]), .B(n2181), .Z(n2183) );
  XNOR U2146 ( .A(n2184), .B(n2185), .Z(n2181) );
  AND U2147 ( .A(n89), .B(n2180), .Z(n2185) );
  XNOR U2148 ( .A(n2184), .B(n2178), .Z(n2180) );
  XOR U2149 ( .A(n2186), .B(n2187), .Z(n2178) );
  AND U2150 ( .A(n104), .B(n2188), .Z(n2187) );
  XNOR U2151 ( .A(n2189), .B(n2190), .Z(n2184) );
  AND U2152 ( .A(n96), .B(n2191), .Z(n2190) );
  XOR U2153 ( .A(p_input[117]), .B(n2189), .Z(n2191) );
  XNOR U2154 ( .A(n2192), .B(n2193), .Z(n2189) );
  AND U2155 ( .A(n100), .B(n2188), .Z(n2193) );
  XNOR U2156 ( .A(n2192), .B(n2186), .Z(n2188) );
  XOR U2157 ( .A(n2194), .B(n2195), .Z(n2186) );
  AND U2158 ( .A(n115), .B(n2196), .Z(n2195) );
  XNOR U2159 ( .A(n2197), .B(n2198), .Z(n2192) );
  AND U2160 ( .A(n107), .B(n2199), .Z(n2198) );
  XOR U2161 ( .A(p_input[149]), .B(n2197), .Z(n2199) );
  XNOR U2162 ( .A(n2200), .B(n2201), .Z(n2197) );
  AND U2163 ( .A(n111), .B(n2196), .Z(n2201) );
  XNOR U2164 ( .A(n2200), .B(n2194), .Z(n2196) );
  XOR U2165 ( .A(n2202), .B(n2203), .Z(n2194) );
  AND U2166 ( .A(n126), .B(n2204), .Z(n2203) );
  XNOR U2167 ( .A(n2205), .B(n2206), .Z(n2200) );
  AND U2168 ( .A(n118), .B(n2207), .Z(n2206) );
  XOR U2169 ( .A(p_input[181]), .B(n2205), .Z(n2207) );
  XNOR U2170 ( .A(n2208), .B(n2209), .Z(n2205) );
  AND U2171 ( .A(n122), .B(n2204), .Z(n2209) );
  XNOR U2172 ( .A(n2208), .B(n2202), .Z(n2204) );
  XOR U2173 ( .A(n2210), .B(n2211), .Z(n2202) );
  AND U2174 ( .A(n137), .B(n2212), .Z(n2211) );
  XNOR U2175 ( .A(n2213), .B(n2214), .Z(n2208) );
  AND U2176 ( .A(n129), .B(n2215), .Z(n2214) );
  XOR U2177 ( .A(p_input[213]), .B(n2213), .Z(n2215) );
  XNOR U2178 ( .A(n2216), .B(n2217), .Z(n2213) );
  AND U2179 ( .A(n133), .B(n2212), .Z(n2217) );
  XNOR U2180 ( .A(n2216), .B(n2210), .Z(n2212) );
  XOR U2181 ( .A(n2218), .B(n2219), .Z(n2210) );
  AND U2182 ( .A(n148), .B(n2220), .Z(n2219) );
  XNOR U2183 ( .A(n2221), .B(n2222), .Z(n2216) );
  AND U2184 ( .A(n140), .B(n2223), .Z(n2222) );
  XOR U2185 ( .A(p_input[245]), .B(n2221), .Z(n2223) );
  XNOR U2186 ( .A(n2224), .B(n2225), .Z(n2221) );
  AND U2187 ( .A(n144), .B(n2220), .Z(n2225) );
  XNOR U2188 ( .A(n2224), .B(n2218), .Z(n2220) );
  XOR U2189 ( .A(n2226), .B(n2227), .Z(n2218) );
  AND U2190 ( .A(n159), .B(n2228), .Z(n2227) );
  XNOR U2191 ( .A(n2229), .B(n2230), .Z(n2224) );
  AND U2192 ( .A(n151), .B(n2231), .Z(n2230) );
  XOR U2193 ( .A(p_input[277]), .B(n2229), .Z(n2231) );
  XNOR U2194 ( .A(n2232), .B(n2233), .Z(n2229) );
  AND U2195 ( .A(n155), .B(n2228), .Z(n2233) );
  XNOR U2196 ( .A(n2232), .B(n2226), .Z(n2228) );
  XOR U2197 ( .A(n2234), .B(n2235), .Z(n2226) );
  AND U2198 ( .A(n170), .B(n2236), .Z(n2235) );
  XNOR U2199 ( .A(n2237), .B(n2238), .Z(n2232) );
  AND U2200 ( .A(n162), .B(n2239), .Z(n2238) );
  XOR U2201 ( .A(p_input[309]), .B(n2237), .Z(n2239) );
  XNOR U2202 ( .A(n2240), .B(n2241), .Z(n2237) );
  AND U2203 ( .A(n166), .B(n2236), .Z(n2241) );
  XNOR U2204 ( .A(n2240), .B(n2234), .Z(n2236) );
  XOR U2205 ( .A(n2242), .B(n2243), .Z(n2234) );
  AND U2206 ( .A(n181), .B(n2244), .Z(n2243) );
  XNOR U2207 ( .A(n2245), .B(n2246), .Z(n2240) );
  AND U2208 ( .A(n173), .B(n2247), .Z(n2246) );
  XOR U2209 ( .A(p_input[341]), .B(n2245), .Z(n2247) );
  XNOR U2210 ( .A(n2248), .B(n2249), .Z(n2245) );
  AND U2211 ( .A(n177), .B(n2244), .Z(n2249) );
  XNOR U2212 ( .A(n2248), .B(n2242), .Z(n2244) );
  XOR U2213 ( .A(n2250), .B(n2251), .Z(n2242) );
  AND U2214 ( .A(n192), .B(n2252), .Z(n2251) );
  XNOR U2215 ( .A(n2253), .B(n2254), .Z(n2248) );
  AND U2216 ( .A(n184), .B(n2255), .Z(n2254) );
  XOR U2217 ( .A(p_input[373]), .B(n2253), .Z(n2255) );
  XNOR U2218 ( .A(n2256), .B(n2257), .Z(n2253) );
  AND U2219 ( .A(n188), .B(n2252), .Z(n2257) );
  XNOR U2220 ( .A(n2256), .B(n2250), .Z(n2252) );
  XOR U2221 ( .A(n2258), .B(n2259), .Z(n2250) );
  AND U2222 ( .A(n203), .B(n2260), .Z(n2259) );
  XNOR U2223 ( .A(n2261), .B(n2262), .Z(n2256) );
  AND U2224 ( .A(n195), .B(n2263), .Z(n2262) );
  XOR U2225 ( .A(p_input[405]), .B(n2261), .Z(n2263) );
  XNOR U2226 ( .A(n2264), .B(n2265), .Z(n2261) );
  AND U2227 ( .A(n199), .B(n2260), .Z(n2265) );
  XNOR U2228 ( .A(n2264), .B(n2258), .Z(n2260) );
  XOR U2229 ( .A(\knn_comb_/min_val_out[0][21] ), .B(n2266), .Z(n2258) );
  AND U2230 ( .A(n213), .B(n2267), .Z(n2266) );
  XNOR U2231 ( .A(n2268), .B(n2269), .Z(n2264) );
  AND U2232 ( .A(n206), .B(n2270), .Z(n2269) );
  XOR U2233 ( .A(p_input[437]), .B(n2268), .Z(n2270) );
  XNOR U2234 ( .A(n2271), .B(n2272), .Z(n2268) );
  AND U2235 ( .A(n210), .B(n2267), .Z(n2272) );
  XOR U2236 ( .A(\knn_comb_/min_val_out[0][21] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .Z(n2267) );
  XOR U2237 ( .A(n33), .B(n2273), .Z(o[20]) );
  AND U2238 ( .A(n58), .B(n2274), .Z(n33) );
  XOR U2239 ( .A(n34), .B(n2273), .Z(n2274) );
  XOR U2240 ( .A(n2275), .B(n2276), .Z(n2273) );
  AND U2241 ( .A(n70), .B(n2277), .Z(n2276) );
  XOR U2242 ( .A(n2278), .B(n2279), .Z(n34) );
  AND U2243 ( .A(n62), .B(n2280), .Z(n2279) );
  XOR U2244 ( .A(p_input[20]), .B(n2278), .Z(n2280) );
  XNOR U2245 ( .A(n2281), .B(n2282), .Z(n2278) );
  AND U2246 ( .A(n66), .B(n2277), .Z(n2282) );
  XNOR U2247 ( .A(n2281), .B(n2275), .Z(n2277) );
  XOR U2248 ( .A(n2283), .B(n2284), .Z(n2275) );
  AND U2249 ( .A(n82), .B(n2285), .Z(n2284) );
  XNOR U2250 ( .A(n2286), .B(n2287), .Z(n2281) );
  AND U2251 ( .A(n74), .B(n2288), .Z(n2287) );
  XOR U2252 ( .A(p_input[52]), .B(n2286), .Z(n2288) );
  XNOR U2253 ( .A(n2289), .B(n2290), .Z(n2286) );
  AND U2254 ( .A(n78), .B(n2285), .Z(n2290) );
  XNOR U2255 ( .A(n2289), .B(n2283), .Z(n2285) );
  XOR U2256 ( .A(n2291), .B(n2292), .Z(n2283) );
  AND U2257 ( .A(n93), .B(n2293), .Z(n2292) );
  XNOR U2258 ( .A(n2294), .B(n2295), .Z(n2289) );
  AND U2259 ( .A(n85), .B(n2296), .Z(n2295) );
  XOR U2260 ( .A(p_input[84]), .B(n2294), .Z(n2296) );
  XNOR U2261 ( .A(n2297), .B(n2298), .Z(n2294) );
  AND U2262 ( .A(n89), .B(n2293), .Z(n2298) );
  XNOR U2263 ( .A(n2297), .B(n2291), .Z(n2293) );
  XOR U2264 ( .A(n2299), .B(n2300), .Z(n2291) );
  AND U2265 ( .A(n104), .B(n2301), .Z(n2300) );
  XNOR U2266 ( .A(n2302), .B(n2303), .Z(n2297) );
  AND U2267 ( .A(n96), .B(n2304), .Z(n2303) );
  XOR U2268 ( .A(p_input[116]), .B(n2302), .Z(n2304) );
  XNOR U2269 ( .A(n2305), .B(n2306), .Z(n2302) );
  AND U2270 ( .A(n100), .B(n2301), .Z(n2306) );
  XNOR U2271 ( .A(n2305), .B(n2299), .Z(n2301) );
  XOR U2272 ( .A(n2307), .B(n2308), .Z(n2299) );
  AND U2273 ( .A(n115), .B(n2309), .Z(n2308) );
  XNOR U2274 ( .A(n2310), .B(n2311), .Z(n2305) );
  AND U2275 ( .A(n107), .B(n2312), .Z(n2311) );
  XOR U2276 ( .A(p_input[148]), .B(n2310), .Z(n2312) );
  XNOR U2277 ( .A(n2313), .B(n2314), .Z(n2310) );
  AND U2278 ( .A(n111), .B(n2309), .Z(n2314) );
  XNOR U2279 ( .A(n2313), .B(n2307), .Z(n2309) );
  XOR U2280 ( .A(n2315), .B(n2316), .Z(n2307) );
  AND U2281 ( .A(n126), .B(n2317), .Z(n2316) );
  XNOR U2282 ( .A(n2318), .B(n2319), .Z(n2313) );
  AND U2283 ( .A(n118), .B(n2320), .Z(n2319) );
  XOR U2284 ( .A(p_input[180]), .B(n2318), .Z(n2320) );
  XNOR U2285 ( .A(n2321), .B(n2322), .Z(n2318) );
  AND U2286 ( .A(n122), .B(n2317), .Z(n2322) );
  XNOR U2287 ( .A(n2321), .B(n2315), .Z(n2317) );
  XOR U2288 ( .A(n2323), .B(n2324), .Z(n2315) );
  AND U2289 ( .A(n137), .B(n2325), .Z(n2324) );
  XNOR U2290 ( .A(n2326), .B(n2327), .Z(n2321) );
  AND U2291 ( .A(n129), .B(n2328), .Z(n2327) );
  XOR U2292 ( .A(p_input[212]), .B(n2326), .Z(n2328) );
  XNOR U2293 ( .A(n2329), .B(n2330), .Z(n2326) );
  AND U2294 ( .A(n133), .B(n2325), .Z(n2330) );
  XNOR U2295 ( .A(n2329), .B(n2323), .Z(n2325) );
  XOR U2296 ( .A(n2331), .B(n2332), .Z(n2323) );
  AND U2297 ( .A(n148), .B(n2333), .Z(n2332) );
  XNOR U2298 ( .A(n2334), .B(n2335), .Z(n2329) );
  AND U2299 ( .A(n140), .B(n2336), .Z(n2335) );
  XOR U2300 ( .A(p_input[244]), .B(n2334), .Z(n2336) );
  XNOR U2301 ( .A(n2337), .B(n2338), .Z(n2334) );
  AND U2302 ( .A(n144), .B(n2333), .Z(n2338) );
  XNOR U2303 ( .A(n2337), .B(n2331), .Z(n2333) );
  XOR U2304 ( .A(n2339), .B(n2340), .Z(n2331) );
  AND U2305 ( .A(n159), .B(n2341), .Z(n2340) );
  XNOR U2306 ( .A(n2342), .B(n2343), .Z(n2337) );
  AND U2307 ( .A(n151), .B(n2344), .Z(n2343) );
  XOR U2308 ( .A(p_input[276]), .B(n2342), .Z(n2344) );
  XNOR U2309 ( .A(n2345), .B(n2346), .Z(n2342) );
  AND U2310 ( .A(n155), .B(n2341), .Z(n2346) );
  XNOR U2311 ( .A(n2345), .B(n2339), .Z(n2341) );
  XOR U2312 ( .A(n2347), .B(n2348), .Z(n2339) );
  AND U2313 ( .A(n170), .B(n2349), .Z(n2348) );
  XNOR U2314 ( .A(n2350), .B(n2351), .Z(n2345) );
  AND U2315 ( .A(n162), .B(n2352), .Z(n2351) );
  XOR U2316 ( .A(p_input[308]), .B(n2350), .Z(n2352) );
  XNOR U2317 ( .A(n2353), .B(n2354), .Z(n2350) );
  AND U2318 ( .A(n166), .B(n2349), .Z(n2354) );
  XNOR U2319 ( .A(n2353), .B(n2347), .Z(n2349) );
  XOR U2320 ( .A(n2355), .B(n2356), .Z(n2347) );
  AND U2321 ( .A(n181), .B(n2357), .Z(n2356) );
  XNOR U2322 ( .A(n2358), .B(n2359), .Z(n2353) );
  AND U2323 ( .A(n173), .B(n2360), .Z(n2359) );
  XOR U2324 ( .A(p_input[340]), .B(n2358), .Z(n2360) );
  XNOR U2325 ( .A(n2361), .B(n2362), .Z(n2358) );
  AND U2326 ( .A(n177), .B(n2357), .Z(n2362) );
  XNOR U2327 ( .A(n2361), .B(n2355), .Z(n2357) );
  XOR U2328 ( .A(n2363), .B(n2364), .Z(n2355) );
  AND U2329 ( .A(n192), .B(n2365), .Z(n2364) );
  XNOR U2330 ( .A(n2366), .B(n2367), .Z(n2361) );
  AND U2331 ( .A(n184), .B(n2368), .Z(n2367) );
  XOR U2332 ( .A(p_input[372]), .B(n2366), .Z(n2368) );
  XNOR U2333 ( .A(n2369), .B(n2370), .Z(n2366) );
  AND U2334 ( .A(n188), .B(n2365), .Z(n2370) );
  XNOR U2335 ( .A(n2369), .B(n2363), .Z(n2365) );
  XOR U2336 ( .A(n2371), .B(n2372), .Z(n2363) );
  AND U2337 ( .A(n203), .B(n2373), .Z(n2372) );
  XNOR U2338 ( .A(n2374), .B(n2375), .Z(n2369) );
  AND U2339 ( .A(n195), .B(n2376), .Z(n2375) );
  XOR U2340 ( .A(p_input[404]), .B(n2374), .Z(n2376) );
  XNOR U2341 ( .A(n2377), .B(n2378), .Z(n2374) );
  AND U2342 ( .A(n199), .B(n2373), .Z(n2378) );
  XNOR U2343 ( .A(n2377), .B(n2371), .Z(n2373) );
  XOR U2344 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n2379), .Z(n2371) );
  AND U2345 ( .A(n213), .B(n2380), .Z(n2379) );
  XNOR U2346 ( .A(n2381), .B(n2382), .Z(n2377) );
  AND U2347 ( .A(n206), .B(n2383), .Z(n2382) );
  XOR U2348 ( .A(p_input[436]), .B(n2381), .Z(n2383) );
  XNOR U2349 ( .A(n2384), .B(n2385), .Z(n2381) );
  AND U2350 ( .A(n210), .B(n2380), .Z(n2385) );
  XOR U2351 ( .A(n2386), .B(n2384), .Z(n2380) );
  IV U2352 ( .A(\knn_comb_/min_val_out[0][20] ), .Z(n2386) );
  IV U2353 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .Z(n2384) );
  XOR U2354 ( .A(n909), .B(n2387), .Z(o[1]) );
  AND U2355 ( .A(n58), .B(n2388), .Z(n909) );
  XOR U2356 ( .A(n910), .B(n2387), .Z(n2388) );
  XOR U2357 ( .A(n2389), .B(n2390), .Z(n2387) );
  AND U2358 ( .A(n70), .B(n2391), .Z(n2390) );
  XOR U2359 ( .A(n2392), .B(n2393), .Z(n910) );
  AND U2360 ( .A(n62), .B(n2394), .Z(n2393) );
  XOR U2361 ( .A(p_input[1]), .B(n2392), .Z(n2394) );
  XNOR U2362 ( .A(n2395), .B(n2396), .Z(n2392) );
  AND U2363 ( .A(n66), .B(n2391), .Z(n2396) );
  XNOR U2364 ( .A(n2395), .B(n2389), .Z(n2391) );
  XOR U2365 ( .A(n2397), .B(n2398), .Z(n2389) );
  AND U2366 ( .A(n82), .B(n2399), .Z(n2398) );
  XNOR U2367 ( .A(n2400), .B(n2401), .Z(n2395) );
  AND U2368 ( .A(n74), .B(n2402), .Z(n2401) );
  XOR U2369 ( .A(p_input[33]), .B(n2400), .Z(n2402) );
  XNOR U2370 ( .A(n2403), .B(n2404), .Z(n2400) );
  AND U2371 ( .A(n78), .B(n2399), .Z(n2404) );
  XNOR U2372 ( .A(n2403), .B(n2397), .Z(n2399) );
  XOR U2373 ( .A(n2405), .B(n2406), .Z(n2397) );
  AND U2374 ( .A(n93), .B(n2407), .Z(n2406) );
  XNOR U2375 ( .A(n2408), .B(n2409), .Z(n2403) );
  AND U2376 ( .A(n85), .B(n2410), .Z(n2409) );
  XOR U2377 ( .A(p_input[65]), .B(n2408), .Z(n2410) );
  XNOR U2378 ( .A(n2411), .B(n2412), .Z(n2408) );
  AND U2379 ( .A(n89), .B(n2407), .Z(n2412) );
  XNOR U2380 ( .A(n2411), .B(n2405), .Z(n2407) );
  XOR U2381 ( .A(n2413), .B(n2414), .Z(n2405) );
  AND U2382 ( .A(n104), .B(n2415), .Z(n2414) );
  XNOR U2383 ( .A(n2416), .B(n2417), .Z(n2411) );
  AND U2384 ( .A(n96), .B(n2418), .Z(n2417) );
  XOR U2385 ( .A(p_input[97]), .B(n2416), .Z(n2418) );
  XNOR U2386 ( .A(n2419), .B(n2420), .Z(n2416) );
  AND U2387 ( .A(n100), .B(n2415), .Z(n2420) );
  XNOR U2388 ( .A(n2419), .B(n2413), .Z(n2415) );
  XOR U2389 ( .A(n2421), .B(n2422), .Z(n2413) );
  AND U2390 ( .A(n115), .B(n2423), .Z(n2422) );
  XNOR U2391 ( .A(n2424), .B(n2425), .Z(n2419) );
  AND U2392 ( .A(n107), .B(n2426), .Z(n2425) );
  XOR U2393 ( .A(p_input[129]), .B(n2424), .Z(n2426) );
  XNOR U2394 ( .A(n2427), .B(n2428), .Z(n2424) );
  AND U2395 ( .A(n111), .B(n2423), .Z(n2428) );
  XNOR U2396 ( .A(n2427), .B(n2421), .Z(n2423) );
  XOR U2397 ( .A(n2429), .B(n2430), .Z(n2421) );
  AND U2398 ( .A(n126), .B(n2431), .Z(n2430) );
  XNOR U2399 ( .A(n2432), .B(n2433), .Z(n2427) );
  AND U2400 ( .A(n118), .B(n2434), .Z(n2433) );
  XOR U2401 ( .A(p_input[161]), .B(n2432), .Z(n2434) );
  XNOR U2402 ( .A(n2435), .B(n2436), .Z(n2432) );
  AND U2403 ( .A(n122), .B(n2431), .Z(n2436) );
  XNOR U2404 ( .A(n2435), .B(n2429), .Z(n2431) );
  XOR U2405 ( .A(n2437), .B(n2438), .Z(n2429) );
  AND U2406 ( .A(n137), .B(n2439), .Z(n2438) );
  XNOR U2407 ( .A(n2440), .B(n2441), .Z(n2435) );
  AND U2408 ( .A(n129), .B(n2442), .Z(n2441) );
  XOR U2409 ( .A(p_input[193]), .B(n2440), .Z(n2442) );
  XNOR U2410 ( .A(n2443), .B(n2444), .Z(n2440) );
  AND U2411 ( .A(n133), .B(n2439), .Z(n2444) );
  XNOR U2412 ( .A(n2443), .B(n2437), .Z(n2439) );
  XOR U2413 ( .A(n2445), .B(n2446), .Z(n2437) );
  AND U2414 ( .A(n148), .B(n2447), .Z(n2446) );
  XNOR U2415 ( .A(n2448), .B(n2449), .Z(n2443) );
  AND U2416 ( .A(n140), .B(n2450), .Z(n2449) );
  XOR U2417 ( .A(p_input[225]), .B(n2448), .Z(n2450) );
  XNOR U2418 ( .A(n2451), .B(n2452), .Z(n2448) );
  AND U2419 ( .A(n144), .B(n2447), .Z(n2452) );
  XNOR U2420 ( .A(n2451), .B(n2445), .Z(n2447) );
  XOR U2421 ( .A(n2453), .B(n2454), .Z(n2445) );
  AND U2422 ( .A(n159), .B(n2455), .Z(n2454) );
  XNOR U2423 ( .A(n2456), .B(n2457), .Z(n2451) );
  AND U2424 ( .A(n151), .B(n2458), .Z(n2457) );
  XOR U2425 ( .A(p_input[257]), .B(n2456), .Z(n2458) );
  XNOR U2426 ( .A(n2459), .B(n2460), .Z(n2456) );
  AND U2427 ( .A(n155), .B(n2455), .Z(n2460) );
  XNOR U2428 ( .A(n2459), .B(n2453), .Z(n2455) );
  XOR U2429 ( .A(n2461), .B(n2462), .Z(n2453) );
  AND U2430 ( .A(n170), .B(n2463), .Z(n2462) );
  XNOR U2431 ( .A(n2464), .B(n2465), .Z(n2459) );
  AND U2432 ( .A(n162), .B(n2466), .Z(n2465) );
  XOR U2433 ( .A(p_input[289]), .B(n2464), .Z(n2466) );
  XNOR U2434 ( .A(n2467), .B(n2468), .Z(n2464) );
  AND U2435 ( .A(n166), .B(n2463), .Z(n2468) );
  XNOR U2436 ( .A(n2467), .B(n2461), .Z(n2463) );
  XOR U2437 ( .A(n2469), .B(n2470), .Z(n2461) );
  AND U2438 ( .A(n181), .B(n2471), .Z(n2470) );
  XNOR U2439 ( .A(n2472), .B(n2473), .Z(n2467) );
  AND U2440 ( .A(n173), .B(n2474), .Z(n2473) );
  XOR U2441 ( .A(p_input[321]), .B(n2472), .Z(n2474) );
  XNOR U2442 ( .A(n2475), .B(n2476), .Z(n2472) );
  AND U2443 ( .A(n177), .B(n2471), .Z(n2476) );
  XNOR U2444 ( .A(n2475), .B(n2469), .Z(n2471) );
  XOR U2445 ( .A(n2477), .B(n2478), .Z(n2469) );
  AND U2446 ( .A(n192), .B(n2479), .Z(n2478) );
  XNOR U2447 ( .A(n2480), .B(n2481), .Z(n2475) );
  AND U2448 ( .A(n184), .B(n2482), .Z(n2481) );
  XOR U2449 ( .A(p_input[353]), .B(n2480), .Z(n2482) );
  XNOR U2450 ( .A(n2483), .B(n2484), .Z(n2480) );
  AND U2451 ( .A(n188), .B(n2479), .Z(n2484) );
  XNOR U2452 ( .A(n2483), .B(n2477), .Z(n2479) );
  XOR U2453 ( .A(n2485), .B(n2486), .Z(n2477) );
  AND U2454 ( .A(n203), .B(n2487), .Z(n2486) );
  XNOR U2455 ( .A(n2488), .B(n2489), .Z(n2483) );
  AND U2456 ( .A(n195), .B(n2490), .Z(n2489) );
  XOR U2457 ( .A(p_input[385]), .B(n2488), .Z(n2490) );
  XNOR U2458 ( .A(n2491), .B(n2492), .Z(n2488) );
  AND U2459 ( .A(n199), .B(n2487), .Z(n2492) );
  XNOR U2460 ( .A(n2491), .B(n2485), .Z(n2487) );
  XOR U2461 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n2493), .Z(n2485) );
  AND U2462 ( .A(n213), .B(n2494), .Z(n2493) );
  XNOR U2463 ( .A(n2495), .B(n2496), .Z(n2491) );
  AND U2464 ( .A(n206), .B(n2497), .Z(n2496) );
  XOR U2465 ( .A(p_input[417]), .B(n2495), .Z(n2497) );
  XNOR U2466 ( .A(n2498), .B(n2499), .Z(n2495) );
  AND U2467 ( .A(n210), .B(n2494), .Z(n2499) );
  XOR U2468 ( .A(\knn_comb_/min_val_out[0][1] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n2494) );
  XOR U2469 ( .A(n35), .B(n2500), .Z(o[19]) );
  AND U2470 ( .A(n58), .B(n2501), .Z(n35) );
  XOR U2471 ( .A(n36), .B(n2500), .Z(n2501) );
  XOR U2472 ( .A(n2502), .B(n2503), .Z(n2500) );
  AND U2473 ( .A(n70), .B(n2504), .Z(n2503) );
  XOR U2474 ( .A(n2505), .B(n2506), .Z(n36) );
  AND U2475 ( .A(n62), .B(n2507), .Z(n2506) );
  XOR U2476 ( .A(p_input[19]), .B(n2505), .Z(n2507) );
  XNOR U2477 ( .A(n2508), .B(n2509), .Z(n2505) );
  AND U2478 ( .A(n66), .B(n2504), .Z(n2509) );
  XNOR U2479 ( .A(n2508), .B(n2502), .Z(n2504) );
  XOR U2480 ( .A(n2510), .B(n2511), .Z(n2502) );
  AND U2481 ( .A(n82), .B(n2512), .Z(n2511) );
  XNOR U2482 ( .A(n2513), .B(n2514), .Z(n2508) );
  AND U2483 ( .A(n74), .B(n2515), .Z(n2514) );
  XOR U2484 ( .A(p_input[51]), .B(n2513), .Z(n2515) );
  XNOR U2485 ( .A(n2516), .B(n2517), .Z(n2513) );
  AND U2486 ( .A(n78), .B(n2512), .Z(n2517) );
  XNOR U2487 ( .A(n2516), .B(n2510), .Z(n2512) );
  XOR U2488 ( .A(n2518), .B(n2519), .Z(n2510) );
  AND U2489 ( .A(n93), .B(n2520), .Z(n2519) );
  XNOR U2490 ( .A(n2521), .B(n2522), .Z(n2516) );
  AND U2491 ( .A(n85), .B(n2523), .Z(n2522) );
  XOR U2492 ( .A(p_input[83]), .B(n2521), .Z(n2523) );
  XNOR U2493 ( .A(n2524), .B(n2525), .Z(n2521) );
  AND U2494 ( .A(n89), .B(n2520), .Z(n2525) );
  XNOR U2495 ( .A(n2524), .B(n2518), .Z(n2520) );
  XOR U2496 ( .A(n2526), .B(n2527), .Z(n2518) );
  AND U2497 ( .A(n104), .B(n2528), .Z(n2527) );
  XNOR U2498 ( .A(n2529), .B(n2530), .Z(n2524) );
  AND U2499 ( .A(n96), .B(n2531), .Z(n2530) );
  XOR U2500 ( .A(p_input[115]), .B(n2529), .Z(n2531) );
  XNOR U2501 ( .A(n2532), .B(n2533), .Z(n2529) );
  AND U2502 ( .A(n100), .B(n2528), .Z(n2533) );
  XNOR U2503 ( .A(n2532), .B(n2526), .Z(n2528) );
  XOR U2504 ( .A(n2534), .B(n2535), .Z(n2526) );
  AND U2505 ( .A(n115), .B(n2536), .Z(n2535) );
  XNOR U2506 ( .A(n2537), .B(n2538), .Z(n2532) );
  AND U2507 ( .A(n107), .B(n2539), .Z(n2538) );
  XOR U2508 ( .A(p_input[147]), .B(n2537), .Z(n2539) );
  XNOR U2509 ( .A(n2540), .B(n2541), .Z(n2537) );
  AND U2510 ( .A(n111), .B(n2536), .Z(n2541) );
  XNOR U2511 ( .A(n2540), .B(n2534), .Z(n2536) );
  XOR U2512 ( .A(n2542), .B(n2543), .Z(n2534) );
  AND U2513 ( .A(n126), .B(n2544), .Z(n2543) );
  XNOR U2514 ( .A(n2545), .B(n2546), .Z(n2540) );
  AND U2515 ( .A(n118), .B(n2547), .Z(n2546) );
  XOR U2516 ( .A(p_input[179]), .B(n2545), .Z(n2547) );
  XNOR U2517 ( .A(n2548), .B(n2549), .Z(n2545) );
  AND U2518 ( .A(n122), .B(n2544), .Z(n2549) );
  XNOR U2519 ( .A(n2548), .B(n2542), .Z(n2544) );
  XOR U2520 ( .A(n2550), .B(n2551), .Z(n2542) );
  AND U2521 ( .A(n137), .B(n2552), .Z(n2551) );
  XNOR U2522 ( .A(n2553), .B(n2554), .Z(n2548) );
  AND U2523 ( .A(n129), .B(n2555), .Z(n2554) );
  XOR U2524 ( .A(p_input[211]), .B(n2553), .Z(n2555) );
  XNOR U2525 ( .A(n2556), .B(n2557), .Z(n2553) );
  AND U2526 ( .A(n133), .B(n2552), .Z(n2557) );
  XNOR U2527 ( .A(n2556), .B(n2550), .Z(n2552) );
  XOR U2528 ( .A(n2558), .B(n2559), .Z(n2550) );
  AND U2529 ( .A(n148), .B(n2560), .Z(n2559) );
  XNOR U2530 ( .A(n2561), .B(n2562), .Z(n2556) );
  AND U2531 ( .A(n140), .B(n2563), .Z(n2562) );
  XOR U2532 ( .A(p_input[243]), .B(n2561), .Z(n2563) );
  XNOR U2533 ( .A(n2564), .B(n2565), .Z(n2561) );
  AND U2534 ( .A(n144), .B(n2560), .Z(n2565) );
  XNOR U2535 ( .A(n2564), .B(n2558), .Z(n2560) );
  XOR U2536 ( .A(n2566), .B(n2567), .Z(n2558) );
  AND U2537 ( .A(n159), .B(n2568), .Z(n2567) );
  XNOR U2538 ( .A(n2569), .B(n2570), .Z(n2564) );
  AND U2539 ( .A(n151), .B(n2571), .Z(n2570) );
  XOR U2540 ( .A(p_input[275]), .B(n2569), .Z(n2571) );
  XNOR U2541 ( .A(n2572), .B(n2573), .Z(n2569) );
  AND U2542 ( .A(n155), .B(n2568), .Z(n2573) );
  XNOR U2543 ( .A(n2572), .B(n2566), .Z(n2568) );
  XOR U2544 ( .A(n2574), .B(n2575), .Z(n2566) );
  AND U2545 ( .A(n170), .B(n2576), .Z(n2575) );
  XNOR U2546 ( .A(n2577), .B(n2578), .Z(n2572) );
  AND U2547 ( .A(n162), .B(n2579), .Z(n2578) );
  XOR U2548 ( .A(p_input[307]), .B(n2577), .Z(n2579) );
  XNOR U2549 ( .A(n2580), .B(n2581), .Z(n2577) );
  AND U2550 ( .A(n166), .B(n2576), .Z(n2581) );
  XNOR U2551 ( .A(n2580), .B(n2574), .Z(n2576) );
  XOR U2552 ( .A(n2582), .B(n2583), .Z(n2574) );
  AND U2553 ( .A(n181), .B(n2584), .Z(n2583) );
  XNOR U2554 ( .A(n2585), .B(n2586), .Z(n2580) );
  AND U2555 ( .A(n173), .B(n2587), .Z(n2586) );
  XOR U2556 ( .A(p_input[339]), .B(n2585), .Z(n2587) );
  XNOR U2557 ( .A(n2588), .B(n2589), .Z(n2585) );
  AND U2558 ( .A(n177), .B(n2584), .Z(n2589) );
  XNOR U2559 ( .A(n2588), .B(n2582), .Z(n2584) );
  XOR U2560 ( .A(n2590), .B(n2591), .Z(n2582) );
  AND U2561 ( .A(n192), .B(n2592), .Z(n2591) );
  XNOR U2562 ( .A(n2593), .B(n2594), .Z(n2588) );
  AND U2563 ( .A(n184), .B(n2595), .Z(n2594) );
  XOR U2564 ( .A(p_input[371]), .B(n2593), .Z(n2595) );
  XNOR U2565 ( .A(n2596), .B(n2597), .Z(n2593) );
  AND U2566 ( .A(n188), .B(n2592), .Z(n2597) );
  XNOR U2567 ( .A(n2596), .B(n2590), .Z(n2592) );
  XOR U2568 ( .A(n2598), .B(n2599), .Z(n2590) );
  AND U2569 ( .A(n203), .B(n2600), .Z(n2599) );
  XNOR U2570 ( .A(n2601), .B(n2602), .Z(n2596) );
  AND U2571 ( .A(n195), .B(n2603), .Z(n2602) );
  XOR U2572 ( .A(p_input[403]), .B(n2601), .Z(n2603) );
  XNOR U2573 ( .A(n2604), .B(n2605), .Z(n2601) );
  AND U2574 ( .A(n199), .B(n2600), .Z(n2605) );
  XNOR U2575 ( .A(n2604), .B(n2598), .Z(n2600) );
  XOR U2576 ( .A(\knn_comb_/min_val_out[0][19] ), .B(n2606), .Z(n2598) );
  AND U2577 ( .A(n213), .B(n2607), .Z(n2606) );
  XNOR U2578 ( .A(n2608), .B(n2609), .Z(n2604) );
  AND U2579 ( .A(n206), .B(n2610), .Z(n2609) );
  XOR U2580 ( .A(p_input[435]), .B(n2608), .Z(n2610) );
  XNOR U2581 ( .A(n2611), .B(n2612), .Z(n2608) );
  AND U2582 ( .A(n210), .B(n2607), .Z(n2612) );
  XOR U2583 ( .A(\knn_comb_/min_val_out[0][19] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .Z(n2607) );
  XOR U2584 ( .A(n37), .B(n2613), .Z(o[18]) );
  AND U2585 ( .A(n58), .B(n2614), .Z(n37) );
  XOR U2586 ( .A(n38), .B(n2613), .Z(n2614) );
  XOR U2587 ( .A(n2615), .B(n2616), .Z(n2613) );
  AND U2588 ( .A(n70), .B(n2617), .Z(n2616) );
  XOR U2589 ( .A(n2618), .B(n2619), .Z(n38) );
  AND U2590 ( .A(n62), .B(n2620), .Z(n2619) );
  XOR U2591 ( .A(p_input[18]), .B(n2618), .Z(n2620) );
  XNOR U2592 ( .A(n2621), .B(n2622), .Z(n2618) );
  AND U2593 ( .A(n66), .B(n2617), .Z(n2622) );
  XNOR U2594 ( .A(n2621), .B(n2615), .Z(n2617) );
  XOR U2595 ( .A(n2623), .B(n2624), .Z(n2615) );
  AND U2596 ( .A(n82), .B(n2625), .Z(n2624) );
  XNOR U2597 ( .A(n2626), .B(n2627), .Z(n2621) );
  AND U2598 ( .A(n74), .B(n2628), .Z(n2627) );
  XOR U2599 ( .A(p_input[50]), .B(n2626), .Z(n2628) );
  XNOR U2600 ( .A(n2629), .B(n2630), .Z(n2626) );
  AND U2601 ( .A(n78), .B(n2625), .Z(n2630) );
  XNOR U2602 ( .A(n2629), .B(n2623), .Z(n2625) );
  XOR U2603 ( .A(n2631), .B(n2632), .Z(n2623) );
  AND U2604 ( .A(n93), .B(n2633), .Z(n2632) );
  XNOR U2605 ( .A(n2634), .B(n2635), .Z(n2629) );
  AND U2606 ( .A(n85), .B(n2636), .Z(n2635) );
  XOR U2607 ( .A(p_input[82]), .B(n2634), .Z(n2636) );
  XNOR U2608 ( .A(n2637), .B(n2638), .Z(n2634) );
  AND U2609 ( .A(n89), .B(n2633), .Z(n2638) );
  XNOR U2610 ( .A(n2637), .B(n2631), .Z(n2633) );
  XOR U2611 ( .A(n2639), .B(n2640), .Z(n2631) );
  AND U2612 ( .A(n104), .B(n2641), .Z(n2640) );
  XNOR U2613 ( .A(n2642), .B(n2643), .Z(n2637) );
  AND U2614 ( .A(n96), .B(n2644), .Z(n2643) );
  XOR U2615 ( .A(p_input[114]), .B(n2642), .Z(n2644) );
  XNOR U2616 ( .A(n2645), .B(n2646), .Z(n2642) );
  AND U2617 ( .A(n100), .B(n2641), .Z(n2646) );
  XNOR U2618 ( .A(n2645), .B(n2639), .Z(n2641) );
  XOR U2619 ( .A(n2647), .B(n2648), .Z(n2639) );
  AND U2620 ( .A(n115), .B(n2649), .Z(n2648) );
  XNOR U2621 ( .A(n2650), .B(n2651), .Z(n2645) );
  AND U2622 ( .A(n107), .B(n2652), .Z(n2651) );
  XOR U2623 ( .A(p_input[146]), .B(n2650), .Z(n2652) );
  XNOR U2624 ( .A(n2653), .B(n2654), .Z(n2650) );
  AND U2625 ( .A(n111), .B(n2649), .Z(n2654) );
  XNOR U2626 ( .A(n2653), .B(n2647), .Z(n2649) );
  XOR U2627 ( .A(n2655), .B(n2656), .Z(n2647) );
  AND U2628 ( .A(n126), .B(n2657), .Z(n2656) );
  XNOR U2629 ( .A(n2658), .B(n2659), .Z(n2653) );
  AND U2630 ( .A(n118), .B(n2660), .Z(n2659) );
  XOR U2631 ( .A(p_input[178]), .B(n2658), .Z(n2660) );
  XNOR U2632 ( .A(n2661), .B(n2662), .Z(n2658) );
  AND U2633 ( .A(n122), .B(n2657), .Z(n2662) );
  XNOR U2634 ( .A(n2661), .B(n2655), .Z(n2657) );
  XOR U2635 ( .A(n2663), .B(n2664), .Z(n2655) );
  AND U2636 ( .A(n137), .B(n2665), .Z(n2664) );
  XNOR U2637 ( .A(n2666), .B(n2667), .Z(n2661) );
  AND U2638 ( .A(n129), .B(n2668), .Z(n2667) );
  XOR U2639 ( .A(p_input[210]), .B(n2666), .Z(n2668) );
  XNOR U2640 ( .A(n2669), .B(n2670), .Z(n2666) );
  AND U2641 ( .A(n133), .B(n2665), .Z(n2670) );
  XNOR U2642 ( .A(n2669), .B(n2663), .Z(n2665) );
  XOR U2643 ( .A(n2671), .B(n2672), .Z(n2663) );
  AND U2644 ( .A(n148), .B(n2673), .Z(n2672) );
  XNOR U2645 ( .A(n2674), .B(n2675), .Z(n2669) );
  AND U2646 ( .A(n140), .B(n2676), .Z(n2675) );
  XOR U2647 ( .A(p_input[242]), .B(n2674), .Z(n2676) );
  XNOR U2648 ( .A(n2677), .B(n2678), .Z(n2674) );
  AND U2649 ( .A(n144), .B(n2673), .Z(n2678) );
  XNOR U2650 ( .A(n2677), .B(n2671), .Z(n2673) );
  XOR U2651 ( .A(n2679), .B(n2680), .Z(n2671) );
  AND U2652 ( .A(n159), .B(n2681), .Z(n2680) );
  XNOR U2653 ( .A(n2682), .B(n2683), .Z(n2677) );
  AND U2654 ( .A(n151), .B(n2684), .Z(n2683) );
  XOR U2655 ( .A(p_input[274]), .B(n2682), .Z(n2684) );
  XNOR U2656 ( .A(n2685), .B(n2686), .Z(n2682) );
  AND U2657 ( .A(n155), .B(n2681), .Z(n2686) );
  XNOR U2658 ( .A(n2685), .B(n2679), .Z(n2681) );
  XOR U2659 ( .A(n2687), .B(n2688), .Z(n2679) );
  AND U2660 ( .A(n170), .B(n2689), .Z(n2688) );
  XNOR U2661 ( .A(n2690), .B(n2691), .Z(n2685) );
  AND U2662 ( .A(n162), .B(n2692), .Z(n2691) );
  XOR U2663 ( .A(p_input[306]), .B(n2690), .Z(n2692) );
  XNOR U2664 ( .A(n2693), .B(n2694), .Z(n2690) );
  AND U2665 ( .A(n166), .B(n2689), .Z(n2694) );
  XNOR U2666 ( .A(n2693), .B(n2687), .Z(n2689) );
  XOR U2667 ( .A(n2695), .B(n2696), .Z(n2687) );
  AND U2668 ( .A(n181), .B(n2697), .Z(n2696) );
  XNOR U2669 ( .A(n2698), .B(n2699), .Z(n2693) );
  AND U2670 ( .A(n173), .B(n2700), .Z(n2699) );
  XOR U2671 ( .A(p_input[338]), .B(n2698), .Z(n2700) );
  XNOR U2672 ( .A(n2701), .B(n2702), .Z(n2698) );
  AND U2673 ( .A(n177), .B(n2697), .Z(n2702) );
  XNOR U2674 ( .A(n2701), .B(n2695), .Z(n2697) );
  XOR U2675 ( .A(n2703), .B(n2704), .Z(n2695) );
  AND U2676 ( .A(n192), .B(n2705), .Z(n2704) );
  XNOR U2677 ( .A(n2706), .B(n2707), .Z(n2701) );
  AND U2678 ( .A(n184), .B(n2708), .Z(n2707) );
  XOR U2679 ( .A(p_input[370]), .B(n2706), .Z(n2708) );
  XNOR U2680 ( .A(n2709), .B(n2710), .Z(n2706) );
  AND U2681 ( .A(n188), .B(n2705), .Z(n2710) );
  XNOR U2682 ( .A(n2709), .B(n2703), .Z(n2705) );
  XOR U2683 ( .A(n2711), .B(n2712), .Z(n2703) );
  AND U2684 ( .A(n203), .B(n2713), .Z(n2712) );
  XNOR U2685 ( .A(n2714), .B(n2715), .Z(n2709) );
  AND U2686 ( .A(n195), .B(n2716), .Z(n2715) );
  XOR U2687 ( .A(p_input[402]), .B(n2714), .Z(n2716) );
  XNOR U2688 ( .A(n2717), .B(n2718), .Z(n2714) );
  AND U2689 ( .A(n199), .B(n2713), .Z(n2718) );
  XNOR U2690 ( .A(n2717), .B(n2711), .Z(n2713) );
  XOR U2691 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n2719), .Z(n2711) );
  AND U2692 ( .A(n213), .B(n2720), .Z(n2719) );
  XNOR U2693 ( .A(n2721), .B(n2722), .Z(n2717) );
  AND U2694 ( .A(n206), .B(n2723), .Z(n2722) );
  XOR U2695 ( .A(p_input[434]), .B(n2721), .Z(n2723) );
  XNOR U2696 ( .A(n2724), .B(n2725), .Z(n2721) );
  AND U2697 ( .A(n210), .B(n2720), .Z(n2725) );
  XOR U2698 ( .A(\knn_comb_/min_val_out[0][18] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .Z(n2720) );
  XOR U2699 ( .A(n41), .B(n2726), .Z(o[17]) );
  AND U2700 ( .A(n58), .B(n2727), .Z(n41) );
  XOR U2701 ( .A(n42), .B(n2726), .Z(n2727) );
  XOR U2702 ( .A(n2728), .B(n2729), .Z(n2726) );
  AND U2703 ( .A(n70), .B(n2730), .Z(n2729) );
  XOR U2704 ( .A(n2731), .B(n2732), .Z(n42) );
  AND U2705 ( .A(n62), .B(n2733), .Z(n2732) );
  XOR U2706 ( .A(p_input[17]), .B(n2731), .Z(n2733) );
  XNOR U2707 ( .A(n2734), .B(n2735), .Z(n2731) );
  AND U2708 ( .A(n66), .B(n2730), .Z(n2735) );
  XNOR U2709 ( .A(n2734), .B(n2728), .Z(n2730) );
  XOR U2710 ( .A(n2736), .B(n2737), .Z(n2728) );
  AND U2711 ( .A(n82), .B(n2738), .Z(n2737) );
  XNOR U2712 ( .A(n2739), .B(n2740), .Z(n2734) );
  AND U2713 ( .A(n74), .B(n2741), .Z(n2740) );
  XOR U2714 ( .A(p_input[49]), .B(n2739), .Z(n2741) );
  XNOR U2715 ( .A(n2742), .B(n2743), .Z(n2739) );
  AND U2716 ( .A(n78), .B(n2738), .Z(n2743) );
  XNOR U2717 ( .A(n2742), .B(n2736), .Z(n2738) );
  XOR U2718 ( .A(n2744), .B(n2745), .Z(n2736) );
  AND U2719 ( .A(n93), .B(n2746), .Z(n2745) );
  XNOR U2720 ( .A(n2747), .B(n2748), .Z(n2742) );
  AND U2721 ( .A(n85), .B(n2749), .Z(n2748) );
  XOR U2722 ( .A(p_input[81]), .B(n2747), .Z(n2749) );
  XNOR U2723 ( .A(n2750), .B(n2751), .Z(n2747) );
  AND U2724 ( .A(n89), .B(n2746), .Z(n2751) );
  XNOR U2725 ( .A(n2750), .B(n2744), .Z(n2746) );
  XOR U2726 ( .A(n2752), .B(n2753), .Z(n2744) );
  AND U2727 ( .A(n104), .B(n2754), .Z(n2753) );
  XNOR U2728 ( .A(n2755), .B(n2756), .Z(n2750) );
  AND U2729 ( .A(n96), .B(n2757), .Z(n2756) );
  XOR U2730 ( .A(p_input[113]), .B(n2755), .Z(n2757) );
  XNOR U2731 ( .A(n2758), .B(n2759), .Z(n2755) );
  AND U2732 ( .A(n100), .B(n2754), .Z(n2759) );
  XNOR U2733 ( .A(n2758), .B(n2752), .Z(n2754) );
  XOR U2734 ( .A(n2760), .B(n2761), .Z(n2752) );
  AND U2735 ( .A(n115), .B(n2762), .Z(n2761) );
  XNOR U2736 ( .A(n2763), .B(n2764), .Z(n2758) );
  AND U2737 ( .A(n107), .B(n2765), .Z(n2764) );
  XOR U2738 ( .A(p_input[145]), .B(n2763), .Z(n2765) );
  XNOR U2739 ( .A(n2766), .B(n2767), .Z(n2763) );
  AND U2740 ( .A(n111), .B(n2762), .Z(n2767) );
  XNOR U2741 ( .A(n2766), .B(n2760), .Z(n2762) );
  XOR U2742 ( .A(n2768), .B(n2769), .Z(n2760) );
  AND U2743 ( .A(n126), .B(n2770), .Z(n2769) );
  XNOR U2744 ( .A(n2771), .B(n2772), .Z(n2766) );
  AND U2745 ( .A(n118), .B(n2773), .Z(n2772) );
  XOR U2746 ( .A(p_input[177]), .B(n2771), .Z(n2773) );
  XNOR U2747 ( .A(n2774), .B(n2775), .Z(n2771) );
  AND U2748 ( .A(n122), .B(n2770), .Z(n2775) );
  XNOR U2749 ( .A(n2774), .B(n2768), .Z(n2770) );
  XOR U2750 ( .A(n2776), .B(n2777), .Z(n2768) );
  AND U2751 ( .A(n137), .B(n2778), .Z(n2777) );
  XNOR U2752 ( .A(n2779), .B(n2780), .Z(n2774) );
  AND U2753 ( .A(n129), .B(n2781), .Z(n2780) );
  XOR U2754 ( .A(p_input[209]), .B(n2779), .Z(n2781) );
  XNOR U2755 ( .A(n2782), .B(n2783), .Z(n2779) );
  AND U2756 ( .A(n133), .B(n2778), .Z(n2783) );
  XNOR U2757 ( .A(n2782), .B(n2776), .Z(n2778) );
  XOR U2758 ( .A(n2784), .B(n2785), .Z(n2776) );
  AND U2759 ( .A(n148), .B(n2786), .Z(n2785) );
  XNOR U2760 ( .A(n2787), .B(n2788), .Z(n2782) );
  AND U2761 ( .A(n140), .B(n2789), .Z(n2788) );
  XOR U2762 ( .A(p_input[241]), .B(n2787), .Z(n2789) );
  XNOR U2763 ( .A(n2790), .B(n2791), .Z(n2787) );
  AND U2764 ( .A(n144), .B(n2786), .Z(n2791) );
  XNOR U2765 ( .A(n2790), .B(n2784), .Z(n2786) );
  XOR U2766 ( .A(n2792), .B(n2793), .Z(n2784) );
  AND U2767 ( .A(n159), .B(n2794), .Z(n2793) );
  XNOR U2768 ( .A(n2795), .B(n2796), .Z(n2790) );
  AND U2769 ( .A(n151), .B(n2797), .Z(n2796) );
  XOR U2770 ( .A(p_input[273]), .B(n2795), .Z(n2797) );
  XNOR U2771 ( .A(n2798), .B(n2799), .Z(n2795) );
  AND U2772 ( .A(n155), .B(n2794), .Z(n2799) );
  XNOR U2773 ( .A(n2798), .B(n2792), .Z(n2794) );
  XOR U2774 ( .A(n2800), .B(n2801), .Z(n2792) );
  AND U2775 ( .A(n170), .B(n2802), .Z(n2801) );
  XNOR U2776 ( .A(n2803), .B(n2804), .Z(n2798) );
  AND U2777 ( .A(n162), .B(n2805), .Z(n2804) );
  XOR U2778 ( .A(p_input[305]), .B(n2803), .Z(n2805) );
  XNOR U2779 ( .A(n2806), .B(n2807), .Z(n2803) );
  AND U2780 ( .A(n166), .B(n2802), .Z(n2807) );
  XNOR U2781 ( .A(n2806), .B(n2800), .Z(n2802) );
  XOR U2782 ( .A(n2808), .B(n2809), .Z(n2800) );
  AND U2783 ( .A(n181), .B(n2810), .Z(n2809) );
  XNOR U2784 ( .A(n2811), .B(n2812), .Z(n2806) );
  AND U2785 ( .A(n173), .B(n2813), .Z(n2812) );
  XOR U2786 ( .A(p_input[337]), .B(n2811), .Z(n2813) );
  XNOR U2787 ( .A(n2814), .B(n2815), .Z(n2811) );
  AND U2788 ( .A(n177), .B(n2810), .Z(n2815) );
  XNOR U2789 ( .A(n2814), .B(n2808), .Z(n2810) );
  XOR U2790 ( .A(n2816), .B(n2817), .Z(n2808) );
  AND U2791 ( .A(n192), .B(n2818), .Z(n2817) );
  XNOR U2792 ( .A(n2819), .B(n2820), .Z(n2814) );
  AND U2793 ( .A(n184), .B(n2821), .Z(n2820) );
  XOR U2794 ( .A(p_input[369]), .B(n2819), .Z(n2821) );
  XNOR U2795 ( .A(n2822), .B(n2823), .Z(n2819) );
  AND U2796 ( .A(n188), .B(n2818), .Z(n2823) );
  XNOR U2797 ( .A(n2822), .B(n2816), .Z(n2818) );
  XOR U2798 ( .A(n2824), .B(n2825), .Z(n2816) );
  AND U2799 ( .A(n203), .B(n2826), .Z(n2825) );
  XNOR U2800 ( .A(n2827), .B(n2828), .Z(n2822) );
  AND U2801 ( .A(n195), .B(n2829), .Z(n2828) );
  XOR U2802 ( .A(p_input[401]), .B(n2827), .Z(n2829) );
  XNOR U2803 ( .A(n2830), .B(n2831), .Z(n2827) );
  AND U2804 ( .A(n199), .B(n2826), .Z(n2831) );
  XNOR U2805 ( .A(n2830), .B(n2824), .Z(n2826) );
  XOR U2806 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n2832), .Z(n2824) );
  AND U2807 ( .A(n213), .B(n2833), .Z(n2832) );
  XNOR U2808 ( .A(n2834), .B(n2835), .Z(n2830) );
  AND U2809 ( .A(n206), .B(n2836), .Z(n2835) );
  XOR U2810 ( .A(p_input[433]), .B(n2834), .Z(n2836) );
  XNOR U2811 ( .A(n2837), .B(n2838), .Z(n2834) );
  AND U2812 ( .A(n210), .B(n2833), .Z(n2838) );
  XOR U2813 ( .A(\knn_comb_/min_val_out[0][17] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .Z(n2833) );
  XOR U2814 ( .A(n43), .B(n2839), .Z(o[16]) );
  AND U2815 ( .A(n58), .B(n2840), .Z(n43) );
  XOR U2816 ( .A(n44), .B(n2839), .Z(n2840) );
  XOR U2817 ( .A(n2841), .B(n2842), .Z(n2839) );
  AND U2818 ( .A(n70), .B(n2843), .Z(n2842) );
  XOR U2819 ( .A(n2844), .B(n2845), .Z(n44) );
  AND U2820 ( .A(n62), .B(n2846), .Z(n2845) );
  XOR U2821 ( .A(p_input[16]), .B(n2844), .Z(n2846) );
  XNOR U2822 ( .A(n2847), .B(n2848), .Z(n2844) );
  AND U2823 ( .A(n66), .B(n2843), .Z(n2848) );
  XNOR U2824 ( .A(n2847), .B(n2841), .Z(n2843) );
  XOR U2825 ( .A(n2849), .B(n2850), .Z(n2841) );
  AND U2826 ( .A(n82), .B(n2851), .Z(n2850) );
  XNOR U2827 ( .A(n2852), .B(n2853), .Z(n2847) );
  AND U2828 ( .A(n74), .B(n2854), .Z(n2853) );
  XOR U2829 ( .A(p_input[48]), .B(n2852), .Z(n2854) );
  XNOR U2830 ( .A(n2855), .B(n2856), .Z(n2852) );
  AND U2831 ( .A(n78), .B(n2851), .Z(n2856) );
  XNOR U2832 ( .A(n2855), .B(n2849), .Z(n2851) );
  XOR U2833 ( .A(n2857), .B(n2858), .Z(n2849) );
  AND U2834 ( .A(n93), .B(n2859), .Z(n2858) );
  XNOR U2835 ( .A(n2860), .B(n2861), .Z(n2855) );
  AND U2836 ( .A(n85), .B(n2862), .Z(n2861) );
  XOR U2837 ( .A(p_input[80]), .B(n2860), .Z(n2862) );
  XNOR U2838 ( .A(n2863), .B(n2864), .Z(n2860) );
  AND U2839 ( .A(n89), .B(n2859), .Z(n2864) );
  XNOR U2840 ( .A(n2863), .B(n2857), .Z(n2859) );
  XOR U2841 ( .A(n2865), .B(n2866), .Z(n2857) );
  AND U2842 ( .A(n104), .B(n2867), .Z(n2866) );
  XNOR U2843 ( .A(n2868), .B(n2869), .Z(n2863) );
  AND U2844 ( .A(n96), .B(n2870), .Z(n2869) );
  XOR U2845 ( .A(p_input[112]), .B(n2868), .Z(n2870) );
  XNOR U2846 ( .A(n2871), .B(n2872), .Z(n2868) );
  AND U2847 ( .A(n100), .B(n2867), .Z(n2872) );
  XNOR U2848 ( .A(n2871), .B(n2865), .Z(n2867) );
  XOR U2849 ( .A(n2873), .B(n2874), .Z(n2865) );
  AND U2850 ( .A(n115), .B(n2875), .Z(n2874) );
  XNOR U2851 ( .A(n2876), .B(n2877), .Z(n2871) );
  AND U2852 ( .A(n107), .B(n2878), .Z(n2877) );
  XOR U2853 ( .A(p_input[144]), .B(n2876), .Z(n2878) );
  XNOR U2854 ( .A(n2879), .B(n2880), .Z(n2876) );
  AND U2855 ( .A(n111), .B(n2875), .Z(n2880) );
  XNOR U2856 ( .A(n2879), .B(n2873), .Z(n2875) );
  XOR U2857 ( .A(n2881), .B(n2882), .Z(n2873) );
  AND U2858 ( .A(n126), .B(n2883), .Z(n2882) );
  XNOR U2859 ( .A(n2884), .B(n2885), .Z(n2879) );
  AND U2860 ( .A(n118), .B(n2886), .Z(n2885) );
  XOR U2861 ( .A(p_input[176]), .B(n2884), .Z(n2886) );
  XNOR U2862 ( .A(n2887), .B(n2888), .Z(n2884) );
  AND U2863 ( .A(n122), .B(n2883), .Z(n2888) );
  XNOR U2864 ( .A(n2887), .B(n2881), .Z(n2883) );
  XOR U2865 ( .A(n2889), .B(n2890), .Z(n2881) );
  AND U2866 ( .A(n137), .B(n2891), .Z(n2890) );
  XNOR U2867 ( .A(n2892), .B(n2893), .Z(n2887) );
  AND U2868 ( .A(n129), .B(n2894), .Z(n2893) );
  XOR U2869 ( .A(p_input[208]), .B(n2892), .Z(n2894) );
  XNOR U2870 ( .A(n2895), .B(n2896), .Z(n2892) );
  AND U2871 ( .A(n133), .B(n2891), .Z(n2896) );
  XNOR U2872 ( .A(n2895), .B(n2889), .Z(n2891) );
  XOR U2873 ( .A(n2897), .B(n2898), .Z(n2889) );
  AND U2874 ( .A(n148), .B(n2899), .Z(n2898) );
  XNOR U2875 ( .A(n2900), .B(n2901), .Z(n2895) );
  AND U2876 ( .A(n140), .B(n2902), .Z(n2901) );
  XOR U2877 ( .A(p_input[240]), .B(n2900), .Z(n2902) );
  XNOR U2878 ( .A(n2903), .B(n2904), .Z(n2900) );
  AND U2879 ( .A(n144), .B(n2899), .Z(n2904) );
  XNOR U2880 ( .A(n2903), .B(n2897), .Z(n2899) );
  XOR U2881 ( .A(n2905), .B(n2906), .Z(n2897) );
  AND U2882 ( .A(n159), .B(n2907), .Z(n2906) );
  XNOR U2883 ( .A(n2908), .B(n2909), .Z(n2903) );
  AND U2884 ( .A(n151), .B(n2910), .Z(n2909) );
  XOR U2885 ( .A(p_input[272]), .B(n2908), .Z(n2910) );
  XNOR U2886 ( .A(n2911), .B(n2912), .Z(n2908) );
  AND U2887 ( .A(n155), .B(n2907), .Z(n2912) );
  XNOR U2888 ( .A(n2911), .B(n2905), .Z(n2907) );
  XOR U2889 ( .A(n2913), .B(n2914), .Z(n2905) );
  AND U2890 ( .A(n170), .B(n2915), .Z(n2914) );
  XNOR U2891 ( .A(n2916), .B(n2917), .Z(n2911) );
  AND U2892 ( .A(n162), .B(n2918), .Z(n2917) );
  XOR U2893 ( .A(p_input[304]), .B(n2916), .Z(n2918) );
  XNOR U2894 ( .A(n2919), .B(n2920), .Z(n2916) );
  AND U2895 ( .A(n166), .B(n2915), .Z(n2920) );
  XNOR U2896 ( .A(n2919), .B(n2913), .Z(n2915) );
  XOR U2897 ( .A(n2921), .B(n2922), .Z(n2913) );
  AND U2898 ( .A(n181), .B(n2923), .Z(n2922) );
  XNOR U2899 ( .A(n2924), .B(n2925), .Z(n2919) );
  AND U2900 ( .A(n173), .B(n2926), .Z(n2925) );
  XOR U2901 ( .A(p_input[336]), .B(n2924), .Z(n2926) );
  XNOR U2902 ( .A(n2927), .B(n2928), .Z(n2924) );
  AND U2903 ( .A(n177), .B(n2923), .Z(n2928) );
  XNOR U2904 ( .A(n2927), .B(n2921), .Z(n2923) );
  XOR U2905 ( .A(n2929), .B(n2930), .Z(n2921) );
  AND U2906 ( .A(n192), .B(n2931), .Z(n2930) );
  XNOR U2907 ( .A(n2932), .B(n2933), .Z(n2927) );
  AND U2908 ( .A(n184), .B(n2934), .Z(n2933) );
  XOR U2909 ( .A(p_input[368]), .B(n2932), .Z(n2934) );
  XNOR U2910 ( .A(n2935), .B(n2936), .Z(n2932) );
  AND U2911 ( .A(n188), .B(n2931), .Z(n2936) );
  XNOR U2912 ( .A(n2935), .B(n2929), .Z(n2931) );
  XOR U2913 ( .A(n2937), .B(n2938), .Z(n2929) );
  AND U2914 ( .A(n203), .B(n2939), .Z(n2938) );
  XNOR U2915 ( .A(n2940), .B(n2941), .Z(n2935) );
  AND U2916 ( .A(n195), .B(n2942), .Z(n2941) );
  XOR U2917 ( .A(p_input[400]), .B(n2940), .Z(n2942) );
  XNOR U2918 ( .A(n2943), .B(n2944), .Z(n2940) );
  AND U2919 ( .A(n199), .B(n2939), .Z(n2944) );
  XNOR U2920 ( .A(n2943), .B(n2937), .Z(n2939) );
  XOR U2921 ( .A(\knn_comb_/min_val_out[0][16] ), .B(n2945), .Z(n2937) );
  AND U2922 ( .A(n213), .B(n2946), .Z(n2945) );
  XNOR U2923 ( .A(n2947), .B(n2948), .Z(n2943) );
  AND U2924 ( .A(n206), .B(n2949), .Z(n2948) );
  XOR U2925 ( .A(p_input[432]), .B(n2947), .Z(n2949) );
  XNOR U2926 ( .A(n2950), .B(n2951), .Z(n2947) );
  AND U2927 ( .A(n210), .B(n2946), .Z(n2951) );
  XOR U2928 ( .A(n2952), .B(n2950), .Z(n2946) );
  IV U2929 ( .A(\knn_comb_/min_val_out[0][16] ), .Z(n2952) );
  IV U2930 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .Z(n2950) );
  XOR U2931 ( .A(n45), .B(n2953), .Z(o[15]) );
  AND U2932 ( .A(n58), .B(n2954), .Z(n45) );
  XOR U2933 ( .A(n46), .B(n2953), .Z(n2954) );
  XOR U2934 ( .A(n2955), .B(n2956), .Z(n2953) );
  AND U2935 ( .A(n70), .B(n2957), .Z(n2956) );
  XOR U2936 ( .A(n2958), .B(n2959), .Z(n46) );
  AND U2937 ( .A(n62), .B(n2960), .Z(n2959) );
  XOR U2938 ( .A(p_input[15]), .B(n2958), .Z(n2960) );
  XNOR U2939 ( .A(n2961), .B(n2962), .Z(n2958) );
  AND U2940 ( .A(n66), .B(n2957), .Z(n2962) );
  XNOR U2941 ( .A(n2961), .B(n2955), .Z(n2957) );
  XOR U2942 ( .A(n2963), .B(n2964), .Z(n2955) );
  AND U2943 ( .A(n82), .B(n2965), .Z(n2964) );
  XNOR U2944 ( .A(n2966), .B(n2967), .Z(n2961) );
  AND U2945 ( .A(n74), .B(n2968), .Z(n2967) );
  XOR U2946 ( .A(p_input[47]), .B(n2966), .Z(n2968) );
  XNOR U2947 ( .A(n2969), .B(n2970), .Z(n2966) );
  AND U2948 ( .A(n78), .B(n2965), .Z(n2970) );
  XNOR U2949 ( .A(n2969), .B(n2963), .Z(n2965) );
  XOR U2950 ( .A(n2971), .B(n2972), .Z(n2963) );
  AND U2951 ( .A(n93), .B(n2973), .Z(n2972) );
  XNOR U2952 ( .A(n2974), .B(n2975), .Z(n2969) );
  AND U2953 ( .A(n85), .B(n2976), .Z(n2975) );
  XOR U2954 ( .A(p_input[79]), .B(n2974), .Z(n2976) );
  XNOR U2955 ( .A(n2977), .B(n2978), .Z(n2974) );
  AND U2956 ( .A(n89), .B(n2973), .Z(n2978) );
  XNOR U2957 ( .A(n2977), .B(n2971), .Z(n2973) );
  XOR U2958 ( .A(n2979), .B(n2980), .Z(n2971) );
  AND U2959 ( .A(n104), .B(n2981), .Z(n2980) );
  XNOR U2960 ( .A(n2982), .B(n2983), .Z(n2977) );
  AND U2961 ( .A(n96), .B(n2984), .Z(n2983) );
  XOR U2962 ( .A(p_input[111]), .B(n2982), .Z(n2984) );
  XNOR U2963 ( .A(n2985), .B(n2986), .Z(n2982) );
  AND U2964 ( .A(n100), .B(n2981), .Z(n2986) );
  XNOR U2965 ( .A(n2985), .B(n2979), .Z(n2981) );
  XOR U2966 ( .A(n2987), .B(n2988), .Z(n2979) );
  AND U2967 ( .A(n115), .B(n2989), .Z(n2988) );
  XNOR U2968 ( .A(n2990), .B(n2991), .Z(n2985) );
  AND U2969 ( .A(n107), .B(n2992), .Z(n2991) );
  XOR U2970 ( .A(p_input[143]), .B(n2990), .Z(n2992) );
  XNOR U2971 ( .A(n2993), .B(n2994), .Z(n2990) );
  AND U2972 ( .A(n111), .B(n2989), .Z(n2994) );
  XNOR U2973 ( .A(n2993), .B(n2987), .Z(n2989) );
  XOR U2974 ( .A(n2995), .B(n2996), .Z(n2987) );
  AND U2975 ( .A(n126), .B(n2997), .Z(n2996) );
  XNOR U2976 ( .A(n2998), .B(n2999), .Z(n2993) );
  AND U2977 ( .A(n118), .B(n3000), .Z(n2999) );
  XOR U2978 ( .A(p_input[175]), .B(n2998), .Z(n3000) );
  XNOR U2979 ( .A(n3001), .B(n3002), .Z(n2998) );
  AND U2980 ( .A(n122), .B(n2997), .Z(n3002) );
  XNOR U2981 ( .A(n3001), .B(n2995), .Z(n2997) );
  XOR U2982 ( .A(n3003), .B(n3004), .Z(n2995) );
  AND U2983 ( .A(n137), .B(n3005), .Z(n3004) );
  XNOR U2984 ( .A(n3006), .B(n3007), .Z(n3001) );
  AND U2985 ( .A(n129), .B(n3008), .Z(n3007) );
  XOR U2986 ( .A(p_input[207]), .B(n3006), .Z(n3008) );
  XNOR U2987 ( .A(n3009), .B(n3010), .Z(n3006) );
  AND U2988 ( .A(n133), .B(n3005), .Z(n3010) );
  XNOR U2989 ( .A(n3009), .B(n3003), .Z(n3005) );
  XOR U2990 ( .A(n3011), .B(n3012), .Z(n3003) );
  AND U2991 ( .A(n148), .B(n3013), .Z(n3012) );
  XNOR U2992 ( .A(n3014), .B(n3015), .Z(n3009) );
  AND U2993 ( .A(n140), .B(n3016), .Z(n3015) );
  XOR U2994 ( .A(p_input[239]), .B(n3014), .Z(n3016) );
  XNOR U2995 ( .A(n3017), .B(n3018), .Z(n3014) );
  AND U2996 ( .A(n144), .B(n3013), .Z(n3018) );
  XNOR U2997 ( .A(n3017), .B(n3011), .Z(n3013) );
  XOR U2998 ( .A(n3019), .B(n3020), .Z(n3011) );
  AND U2999 ( .A(n159), .B(n3021), .Z(n3020) );
  XNOR U3000 ( .A(n3022), .B(n3023), .Z(n3017) );
  AND U3001 ( .A(n151), .B(n3024), .Z(n3023) );
  XOR U3002 ( .A(p_input[271]), .B(n3022), .Z(n3024) );
  XNOR U3003 ( .A(n3025), .B(n3026), .Z(n3022) );
  AND U3004 ( .A(n155), .B(n3021), .Z(n3026) );
  XNOR U3005 ( .A(n3025), .B(n3019), .Z(n3021) );
  XOR U3006 ( .A(n3027), .B(n3028), .Z(n3019) );
  AND U3007 ( .A(n170), .B(n3029), .Z(n3028) );
  XNOR U3008 ( .A(n3030), .B(n3031), .Z(n3025) );
  AND U3009 ( .A(n162), .B(n3032), .Z(n3031) );
  XOR U3010 ( .A(p_input[303]), .B(n3030), .Z(n3032) );
  XNOR U3011 ( .A(n3033), .B(n3034), .Z(n3030) );
  AND U3012 ( .A(n166), .B(n3029), .Z(n3034) );
  XNOR U3013 ( .A(n3033), .B(n3027), .Z(n3029) );
  XOR U3014 ( .A(n3035), .B(n3036), .Z(n3027) );
  AND U3015 ( .A(n181), .B(n3037), .Z(n3036) );
  XNOR U3016 ( .A(n3038), .B(n3039), .Z(n3033) );
  AND U3017 ( .A(n173), .B(n3040), .Z(n3039) );
  XOR U3018 ( .A(p_input[335]), .B(n3038), .Z(n3040) );
  XNOR U3019 ( .A(n3041), .B(n3042), .Z(n3038) );
  AND U3020 ( .A(n177), .B(n3037), .Z(n3042) );
  XNOR U3021 ( .A(n3041), .B(n3035), .Z(n3037) );
  XOR U3022 ( .A(n3043), .B(n3044), .Z(n3035) );
  AND U3023 ( .A(n192), .B(n3045), .Z(n3044) );
  XNOR U3024 ( .A(n3046), .B(n3047), .Z(n3041) );
  AND U3025 ( .A(n184), .B(n3048), .Z(n3047) );
  XOR U3026 ( .A(p_input[367]), .B(n3046), .Z(n3048) );
  XNOR U3027 ( .A(n3049), .B(n3050), .Z(n3046) );
  AND U3028 ( .A(n188), .B(n3045), .Z(n3050) );
  XNOR U3029 ( .A(n3049), .B(n3043), .Z(n3045) );
  XOR U3030 ( .A(n3051), .B(n3052), .Z(n3043) );
  AND U3031 ( .A(n203), .B(n3053), .Z(n3052) );
  XNOR U3032 ( .A(n3054), .B(n3055), .Z(n3049) );
  AND U3033 ( .A(n195), .B(n3056), .Z(n3055) );
  XOR U3034 ( .A(p_input[399]), .B(n3054), .Z(n3056) );
  XNOR U3035 ( .A(n3057), .B(n3058), .Z(n3054) );
  AND U3036 ( .A(n199), .B(n3053), .Z(n3058) );
  XNOR U3037 ( .A(n3057), .B(n3051), .Z(n3053) );
  XOR U3038 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n3059), .Z(n3051) );
  AND U3039 ( .A(n213), .B(n3060), .Z(n3059) );
  XNOR U3040 ( .A(n3061), .B(n3062), .Z(n3057) );
  AND U3041 ( .A(n206), .B(n3063), .Z(n3062) );
  XOR U3042 ( .A(p_input[431]), .B(n3061), .Z(n3063) );
  XNOR U3043 ( .A(n3064), .B(n3065), .Z(n3061) );
  AND U3044 ( .A(n210), .B(n3060), .Z(n3065) );
  XOR U3045 ( .A(n3066), .B(n3064), .Z(n3060) );
  IV U3046 ( .A(\knn_comb_/min_val_out[0][15] ), .Z(n3066) );
  IV U3047 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .Z(n3064) );
  XOR U3048 ( .A(n47), .B(n3067), .Z(o[14]) );
  AND U3049 ( .A(n58), .B(n3068), .Z(n47) );
  XOR U3050 ( .A(n48), .B(n3067), .Z(n3068) );
  XOR U3051 ( .A(n3069), .B(n3070), .Z(n3067) );
  AND U3052 ( .A(n70), .B(n3071), .Z(n3070) );
  XOR U3053 ( .A(n3072), .B(n3073), .Z(n48) );
  AND U3054 ( .A(n62), .B(n3074), .Z(n3073) );
  XOR U3055 ( .A(p_input[14]), .B(n3072), .Z(n3074) );
  XNOR U3056 ( .A(n3075), .B(n3076), .Z(n3072) );
  AND U3057 ( .A(n66), .B(n3071), .Z(n3076) );
  XNOR U3058 ( .A(n3075), .B(n3069), .Z(n3071) );
  XOR U3059 ( .A(n3077), .B(n3078), .Z(n3069) );
  AND U3060 ( .A(n82), .B(n3079), .Z(n3078) );
  XNOR U3061 ( .A(n3080), .B(n3081), .Z(n3075) );
  AND U3062 ( .A(n74), .B(n3082), .Z(n3081) );
  XOR U3063 ( .A(p_input[46]), .B(n3080), .Z(n3082) );
  XNOR U3064 ( .A(n3083), .B(n3084), .Z(n3080) );
  AND U3065 ( .A(n78), .B(n3079), .Z(n3084) );
  XNOR U3066 ( .A(n3083), .B(n3077), .Z(n3079) );
  XOR U3067 ( .A(n3085), .B(n3086), .Z(n3077) );
  AND U3068 ( .A(n93), .B(n3087), .Z(n3086) );
  XNOR U3069 ( .A(n3088), .B(n3089), .Z(n3083) );
  AND U3070 ( .A(n85), .B(n3090), .Z(n3089) );
  XOR U3071 ( .A(p_input[78]), .B(n3088), .Z(n3090) );
  XNOR U3072 ( .A(n3091), .B(n3092), .Z(n3088) );
  AND U3073 ( .A(n89), .B(n3087), .Z(n3092) );
  XNOR U3074 ( .A(n3091), .B(n3085), .Z(n3087) );
  XOR U3075 ( .A(n3093), .B(n3094), .Z(n3085) );
  AND U3076 ( .A(n104), .B(n3095), .Z(n3094) );
  XNOR U3077 ( .A(n3096), .B(n3097), .Z(n3091) );
  AND U3078 ( .A(n96), .B(n3098), .Z(n3097) );
  XOR U3079 ( .A(p_input[110]), .B(n3096), .Z(n3098) );
  XNOR U3080 ( .A(n3099), .B(n3100), .Z(n3096) );
  AND U3081 ( .A(n100), .B(n3095), .Z(n3100) );
  XNOR U3082 ( .A(n3099), .B(n3093), .Z(n3095) );
  XOR U3083 ( .A(n3101), .B(n3102), .Z(n3093) );
  AND U3084 ( .A(n115), .B(n3103), .Z(n3102) );
  XNOR U3085 ( .A(n3104), .B(n3105), .Z(n3099) );
  AND U3086 ( .A(n107), .B(n3106), .Z(n3105) );
  XOR U3087 ( .A(p_input[142]), .B(n3104), .Z(n3106) );
  XNOR U3088 ( .A(n3107), .B(n3108), .Z(n3104) );
  AND U3089 ( .A(n111), .B(n3103), .Z(n3108) );
  XNOR U3090 ( .A(n3107), .B(n3101), .Z(n3103) );
  XOR U3091 ( .A(n3109), .B(n3110), .Z(n3101) );
  AND U3092 ( .A(n126), .B(n3111), .Z(n3110) );
  XNOR U3093 ( .A(n3112), .B(n3113), .Z(n3107) );
  AND U3094 ( .A(n118), .B(n3114), .Z(n3113) );
  XOR U3095 ( .A(p_input[174]), .B(n3112), .Z(n3114) );
  XNOR U3096 ( .A(n3115), .B(n3116), .Z(n3112) );
  AND U3097 ( .A(n122), .B(n3111), .Z(n3116) );
  XNOR U3098 ( .A(n3115), .B(n3109), .Z(n3111) );
  XOR U3099 ( .A(n3117), .B(n3118), .Z(n3109) );
  AND U3100 ( .A(n137), .B(n3119), .Z(n3118) );
  XNOR U3101 ( .A(n3120), .B(n3121), .Z(n3115) );
  AND U3102 ( .A(n129), .B(n3122), .Z(n3121) );
  XOR U3103 ( .A(p_input[206]), .B(n3120), .Z(n3122) );
  XNOR U3104 ( .A(n3123), .B(n3124), .Z(n3120) );
  AND U3105 ( .A(n133), .B(n3119), .Z(n3124) );
  XNOR U3106 ( .A(n3123), .B(n3117), .Z(n3119) );
  XOR U3107 ( .A(n3125), .B(n3126), .Z(n3117) );
  AND U3108 ( .A(n148), .B(n3127), .Z(n3126) );
  XNOR U3109 ( .A(n3128), .B(n3129), .Z(n3123) );
  AND U3110 ( .A(n140), .B(n3130), .Z(n3129) );
  XOR U3111 ( .A(p_input[238]), .B(n3128), .Z(n3130) );
  XNOR U3112 ( .A(n3131), .B(n3132), .Z(n3128) );
  AND U3113 ( .A(n144), .B(n3127), .Z(n3132) );
  XNOR U3114 ( .A(n3131), .B(n3125), .Z(n3127) );
  XOR U3115 ( .A(n3133), .B(n3134), .Z(n3125) );
  AND U3116 ( .A(n159), .B(n3135), .Z(n3134) );
  XNOR U3117 ( .A(n3136), .B(n3137), .Z(n3131) );
  AND U3118 ( .A(n151), .B(n3138), .Z(n3137) );
  XOR U3119 ( .A(p_input[270]), .B(n3136), .Z(n3138) );
  XNOR U3120 ( .A(n3139), .B(n3140), .Z(n3136) );
  AND U3121 ( .A(n155), .B(n3135), .Z(n3140) );
  XNOR U3122 ( .A(n3139), .B(n3133), .Z(n3135) );
  XOR U3123 ( .A(n3141), .B(n3142), .Z(n3133) );
  AND U3124 ( .A(n170), .B(n3143), .Z(n3142) );
  XNOR U3125 ( .A(n3144), .B(n3145), .Z(n3139) );
  AND U3126 ( .A(n162), .B(n3146), .Z(n3145) );
  XOR U3127 ( .A(p_input[302]), .B(n3144), .Z(n3146) );
  XNOR U3128 ( .A(n3147), .B(n3148), .Z(n3144) );
  AND U3129 ( .A(n166), .B(n3143), .Z(n3148) );
  XNOR U3130 ( .A(n3147), .B(n3141), .Z(n3143) );
  XOR U3131 ( .A(n3149), .B(n3150), .Z(n3141) );
  AND U3132 ( .A(n181), .B(n3151), .Z(n3150) );
  XNOR U3133 ( .A(n3152), .B(n3153), .Z(n3147) );
  AND U3134 ( .A(n173), .B(n3154), .Z(n3153) );
  XOR U3135 ( .A(p_input[334]), .B(n3152), .Z(n3154) );
  XNOR U3136 ( .A(n3155), .B(n3156), .Z(n3152) );
  AND U3137 ( .A(n177), .B(n3151), .Z(n3156) );
  XNOR U3138 ( .A(n3155), .B(n3149), .Z(n3151) );
  XOR U3139 ( .A(n3157), .B(n3158), .Z(n3149) );
  AND U3140 ( .A(n192), .B(n3159), .Z(n3158) );
  XNOR U3141 ( .A(n3160), .B(n3161), .Z(n3155) );
  AND U3142 ( .A(n184), .B(n3162), .Z(n3161) );
  XOR U3143 ( .A(p_input[366]), .B(n3160), .Z(n3162) );
  XNOR U3144 ( .A(n3163), .B(n3164), .Z(n3160) );
  AND U3145 ( .A(n188), .B(n3159), .Z(n3164) );
  XNOR U3146 ( .A(n3163), .B(n3157), .Z(n3159) );
  XOR U3147 ( .A(n3165), .B(n3166), .Z(n3157) );
  AND U3148 ( .A(n203), .B(n3167), .Z(n3166) );
  XNOR U3149 ( .A(n3168), .B(n3169), .Z(n3163) );
  AND U3150 ( .A(n195), .B(n3170), .Z(n3169) );
  XOR U3151 ( .A(p_input[398]), .B(n3168), .Z(n3170) );
  XNOR U3152 ( .A(n3171), .B(n3172), .Z(n3168) );
  AND U3153 ( .A(n199), .B(n3167), .Z(n3172) );
  XNOR U3154 ( .A(n3171), .B(n3165), .Z(n3167) );
  XOR U3155 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n3173), .Z(n3165) );
  AND U3156 ( .A(n213), .B(n3174), .Z(n3173) );
  XNOR U3157 ( .A(n3175), .B(n3176), .Z(n3171) );
  AND U3158 ( .A(n206), .B(n3177), .Z(n3176) );
  XOR U3159 ( .A(p_input[430]), .B(n3175), .Z(n3177) );
  XNOR U3160 ( .A(n3178), .B(n3179), .Z(n3175) );
  AND U3161 ( .A(n210), .B(n3174), .Z(n3179) );
  XOR U3162 ( .A(\knn_comb_/min_val_out[0][14] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n3174) );
  XOR U3163 ( .A(n49), .B(n3180), .Z(o[13]) );
  AND U3164 ( .A(n58), .B(n3181), .Z(n49) );
  XOR U3165 ( .A(n50), .B(n3180), .Z(n3181) );
  XOR U3166 ( .A(n3182), .B(n3183), .Z(n3180) );
  AND U3167 ( .A(n70), .B(n3184), .Z(n3183) );
  XOR U3168 ( .A(n3185), .B(n3186), .Z(n50) );
  AND U3169 ( .A(n62), .B(n3187), .Z(n3186) );
  XOR U3170 ( .A(p_input[13]), .B(n3185), .Z(n3187) );
  XNOR U3171 ( .A(n3188), .B(n3189), .Z(n3185) );
  AND U3172 ( .A(n66), .B(n3184), .Z(n3189) );
  XNOR U3173 ( .A(n3188), .B(n3182), .Z(n3184) );
  XOR U3174 ( .A(n3190), .B(n3191), .Z(n3182) );
  AND U3175 ( .A(n82), .B(n3192), .Z(n3191) );
  XNOR U3176 ( .A(n3193), .B(n3194), .Z(n3188) );
  AND U3177 ( .A(n74), .B(n3195), .Z(n3194) );
  XOR U3178 ( .A(p_input[45]), .B(n3193), .Z(n3195) );
  XNOR U3179 ( .A(n3196), .B(n3197), .Z(n3193) );
  AND U3180 ( .A(n78), .B(n3192), .Z(n3197) );
  XNOR U3181 ( .A(n3196), .B(n3190), .Z(n3192) );
  XOR U3182 ( .A(n3198), .B(n3199), .Z(n3190) );
  AND U3183 ( .A(n93), .B(n3200), .Z(n3199) );
  XNOR U3184 ( .A(n3201), .B(n3202), .Z(n3196) );
  AND U3185 ( .A(n85), .B(n3203), .Z(n3202) );
  XOR U3186 ( .A(p_input[77]), .B(n3201), .Z(n3203) );
  XNOR U3187 ( .A(n3204), .B(n3205), .Z(n3201) );
  AND U3188 ( .A(n89), .B(n3200), .Z(n3205) );
  XNOR U3189 ( .A(n3204), .B(n3198), .Z(n3200) );
  XOR U3190 ( .A(n3206), .B(n3207), .Z(n3198) );
  AND U3191 ( .A(n104), .B(n3208), .Z(n3207) );
  XNOR U3192 ( .A(n3209), .B(n3210), .Z(n3204) );
  AND U3193 ( .A(n96), .B(n3211), .Z(n3210) );
  XOR U3194 ( .A(p_input[109]), .B(n3209), .Z(n3211) );
  XNOR U3195 ( .A(n3212), .B(n3213), .Z(n3209) );
  AND U3196 ( .A(n100), .B(n3208), .Z(n3213) );
  XNOR U3197 ( .A(n3212), .B(n3206), .Z(n3208) );
  XOR U3198 ( .A(n3214), .B(n3215), .Z(n3206) );
  AND U3199 ( .A(n115), .B(n3216), .Z(n3215) );
  XNOR U3200 ( .A(n3217), .B(n3218), .Z(n3212) );
  AND U3201 ( .A(n107), .B(n3219), .Z(n3218) );
  XOR U3202 ( .A(p_input[141]), .B(n3217), .Z(n3219) );
  XNOR U3203 ( .A(n3220), .B(n3221), .Z(n3217) );
  AND U3204 ( .A(n111), .B(n3216), .Z(n3221) );
  XNOR U3205 ( .A(n3220), .B(n3214), .Z(n3216) );
  XOR U3206 ( .A(n3222), .B(n3223), .Z(n3214) );
  AND U3207 ( .A(n126), .B(n3224), .Z(n3223) );
  XNOR U3208 ( .A(n3225), .B(n3226), .Z(n3220) );
  AND U3209 ( .A(n118), .B(n3227), .Z(n3226) );
  XOR U3210 ( .A(p_input[173]), .B(n3225), .Z(n3227) );
  XNOR U3211 ( .A(n3228), .B(n3229), .Z(n3225) );
  AND U3212 ( .A(n122), .B(n3224), .Z(n3229) );
  XNOR U3213 ( .A(n3228), .B(n3222), .Z(n3224) );
  XOR U3214 ( .A(n3230), .B(n3231), .Z(n3222) );
  AND U3215 ( .A(n137), .B(n3232), .Z(n3231) );
  XNOR U3216 ( .A(n3233), .B(n3234), .Z(n3228) );
  AND U3217 ( .A(n129), .B(n3235), .Z(n3234) );
  XOR U3218 ( .A(p_input[205]), .B(n3233), .Z(n3235) );
  XNOR U3219 ( .A(n3236), .B(n3237), .Z(n3233) );
  AND U3220 ( .A(n133), .B(n3232), .Z(n3237) );
  XNOR U3221 ( .A(n3236), .B(n3230), .Z(n3232) );
  XOR U3222 ( .A(n3238), .B(n3239), .Z(n3230) );
  AND U3223 ( .A(n148), .B(n3240), .Z(n3239) );
  XNOR U3224 ( .A(n3241), .B(n3242), .Z(n3236) );
  AND U3225 ( .A(n140), .B(n3243), .Z(n3242) );
  XOR U3226 ( .A(p_input[237]), .B(n3241), .Z(n3243) );
  XNOR U3227 ( .A(n3244), .B(n3245), .Z(n3241) );
  AND U3228 ( .A(n144), .B(n3240), .Z(n3245) );
  XNOR U3229 ( .A(n3244), .B(n3238), .Z(n3240) );
  XOR U3230 ( .A(n3246), .B(n3247), .Z(n3238) );
  AND U3231 ( .A(n159), .B(n3248), .Z(n3247) );
  XNOR U3232 ( .A(n3249), .B(n3250), .Z(n3244) );
  AND U3233 ( .A(n151), .B(n3251), .Z(n3250) );
  XOR U3234 ( .A(p_input[269]), .B(n3249), .Z(n3251) );
  XNOR U3235 ( .A(n3252), .B(n3253), .Z(n3249) );
  AND U3236 ( .A(n155), .B(n3248), .Z(n3253) );
  XNOR U3237 ( .A(n3252), .B(n3246), .Z(n3248) );
  XOR U3238 ( .A(n3254), .B(n3255), .Z(n3246) );
  AND U3239 ( .A(n170), .B(n3256), .Z(n3255) );
  XNOR U3240 ( .A(n3257), .B(n3258), .Z(n3252) );
  AND U3241 ( .A(n162), .B(n3259), .Z(n3258) );
  XOR U3242 ( .A(p_input[301]), .B(n3257), .Z(n3259) );
  XNOR U3243 ( .A(n3260), .B(n3261), .Z(n3257) );
  AND U3244 ( .A(n166), .B(n3256), .Z(n3261) );
  XNOR U3245 ( .A(n3260), .B(n3254), .Z(n3256) );
  XOR U3246 ( .A(n3262), .B(n3263), .Z(n3254) );
  AND U3247 ( .A(n181), .B(n3264), .Z(n3263) );
  XNOR U3248 ( .A(n3265), .B(n3266), .Z(n3260) );
  AND U3249 ( .A(n173), .B(n3267), .Z(n3266) );
  XOR U3250 ( .A(p_input[333]), .B(n3265), .Z(n3267) );
  XNOR U3251 ( .A(n3268), .B(n3269), .Z(n3265) );
  AND U3252 ( .A(n177), .B(n3264), .Z(n3269) );
  XNOR U3253 ( .A(n3268), .B(n3262), .Z(n3264) );
  XOR U3254 ( .A(n3270), .B(n3271), .Z(n3262) );
  AND U3255 ( .A(n192), .B(n3272), .Z(n3271) );
  XNOR U3256 ( .A(n3273), .B(n3274), .Z(n3268) );
  AND U3257 ( .A(n184), .B(n3275), .Z(n3274) );
  XOR U3258 ( .A(p_input[365]), .B(n3273), .Z(n3275) );
  XNOR U3259 ( .A(n3276), .B(n3277), .Z(n3273) );
  AND U3260 ( .A(n188), .B(n3272), .Z(n3277) );
  XNOR U3261 ( .A(n3276), .B(n3270), .Z(n3272) );
  XOR U3262 ( .A(n3278), .B(n3279), .Z(n3270) );
  AND U3263 ( .A(n203), .B(n3280), .Z(n3279) );
  XNOR U3264 ( .A(n3281), .B(n3282), .Z(n3276) );
  AND U3265 ( .A(n195), .B(n3283), .Z(n3282) );
  XOR U3266 ( .A(p_input[397]), .B(n3281), .Z(n3283) );
  XNOR U3267 ( .A(n3284), .B(n3285), .Z(n3281) );
  AND U3268 ( .A(n199), .B(n3280), .Z(n3285) );
  XNOR U3269 ( .A(n3284), .B(n3278), .Z(n3280) );
  XOR U3270 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n3286), .Z(n3278) );
  AND U3271 ( .A(n213), .B(n3287), .Z(n3286) );
  XNOR U3272 ( .A(n3288), .B(n3289), .Z(n3284) );
  AND U3273 ( .A(n206), .B(n3290), .Z(n3289) );
  XOR U3274 ( .A(p_input[429]), .B(n3288), .Z(n3290) );
  XNOR U3275 ( .A(n3291), .B(n3292), .Z(n3288) );
  AND U3276 ( .A(n210), .B(n3287), .Z(n3292) );
  XOR U3277 ( .A(\knn_comb_/min_val_out[0][13] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n3287) );
  XOR U3278 ( .A(n51), .B(n3293), .Z(o[12]) );
  AND U3279 ( .A(n58), .B(n3294), .Z(n51) );
  XOR U3280 ( .A(n52), .B(n3293), .Z(n3294) );
  XOR U3281 ( .A(n3295), .B(n3296), .Z(n3293) );
  AND U3282 ( .A(n70), .B(n3297), .Z(n3296) );
  XOR U3283 ( .A(n3298), .B(n3299), .Z(n52) );
  AND U3284 ( .A(n62), .B(n3300), .Z(n3299) );
  XOR U3285 ( .A(p_input[12]), .B(n3298), .Z(n3300) );
  XNOR U3286 ( .A(n3301), .B(n3302), .Z(n3298) );
  AND U3287 ( .A(n66), .B(n3297), .Z(n3302) );
  XNOR U3288 ( .A(n3301), .B(n3295), .Z(n3297) );
  XOR U3289 ( .A(n3303), .B(n3304), .Z(n3295) );
  AND U3290 ( .A(n82), .B(n3305), .Z(n3304) );
  XNOR U3291 ( .A(n3306), .B(n3307), .Z(n3301) );
  AND U3292 ( .A(n74), .B(n3308), .Z(n3307) );
  XOR U3293 ( .A(p_input[44]), .B(n3306), .Z(n3308) );
  XNOR U3294 ( .A(n3309), .B(n3310), .Z(n3306) );
  AND U3295 ( .A(n78), .B(n3305), .Z(n3310) );
  XNOR U3296 ( .A(n3309), .B(n3303), .Z(n3305) );
  XOR U3297 ( .A(n3311), .B(n3312), .Z(n3303) );
  AND U3298 ( .A(n93), .B(n3313), .Z(n3312) );
  XNOR U3299 ( .A(n3314), .B(n3315), .Z(n3309) );
  AND U3300 ( .A(n85), .B(n3316), .Z(n3315) );
  XOR U3301 ( .A(p_input[76]), .B(n3314), .Z(n3316) );
  XNOR U3302 ( .A(n3317), .B(n3318), .Z(n3314) );
  AND U3303 ( .A(n89), .B(n3313), .Z(n3318) );
  XNOR U3304 ( .A(n3317), .B(n3311), .Z(n3313) );
  XOR U3305 ( .A(n3319), .B(n3320), .Z(n3311) );
  AND U3306 ( .A(n104), .B(n3321), .Z(n3320) );
  XNOR U3307 ( .A(n3322), .B(n3323), .Z(n3317) );
  AND U3308 ( .A(n96), .B(n3324), .Z(n3323) );
  XOR U3309 ( .A(p_input[108]), .B(n3322), .Z(n3324) );
  XNOR U3310 ( .A(n3325), .B(n3326), .Z(n3322) );
  AND U3311 ( .A(n100), .B(n3321), .Z(n3326) );
  XNOR U3312 ( .A(n3325), .B(n3319), .Z(n3321) );
  XOR U3313 ( .A(n3327), .B(n3328), .Z(n3319) );
  AND U3314 ( .A(n115), .B(n3329), .Z(n3328) );
  XNOR U3315 ( .A(n3330), .B(n3331), .Z(n3325) );
  AND U3316 ( .A(n107), .B(n3332), .Z(n3331) );
  XOR U3317 ( .A(p_input[140]), .B(n3330), .Z(n3332) );
  XNOR U3318 ( .A(n3333), .B(n3334), .Z(n3330) );
  AND U3319 ( .A(n111), .B(n3329), .Z(n3334) );
  XNOR U3320 ( .A(n3333), .B(n3327), .Z(n3329) );
  XOR U3321 ( .A(n3335), .B(n3336), .Z(n3327) );
  AND U3322 ( .A(n126), .B(n3337), .Z(n3336) );
  XNOR U3323 ( .A(n3338), .B(n3339), .Z(n3333) );
  AND U3324 ( .A(n118), .B(n3340), .Z(n3339) );
  XOR U3325 ( .A(p_input[172]), .B(n3338), .Z(n3340) );
  XNOR U3326 ( .A(n3341), .B(n3342), .Z(n3338) );
  AND U3327 ( .A(n122), .B(n3337), .Z(n3342) );
  XNOR U3328 ( .A(n3341), .B(n3335), .Z(n3337) );
  XOR U3329 ( .A(n3343), .B(n3344), .Z(n3335) );
  AND U3330 ( .A(n137), .B(n3345), .Z(n3344) );
  XNOR U3331 ( .A(n3346), .B(n3347), .Z(n3341) );
  AND U3332 ( .A(n129), .B(n3348), .Z(n3347) );
  XOR U3333 ( .A(p_input[204]), .B(n3346), .Z(n3348) );
  XNOR U3334 ( .A(n3349), .B(n3350), .Z(n3346) );
  AND U3335 ( .A(n133), .B(n3345), .Z(n3350) );
  XNOR U3336 ( .A(n3349), .B(n3343), .Z(n3345) );
  XOR U3337 ( .A(n3351), .B(n3352), .Z(n3343) );
  AND U3338 ( .A(n148), .B(n3353), .Z(n3352) );
  XNOR U3339 ( .A(n3354), .B(n3355), .Z(n3349) );
  AND U3340 ( .A(n140), .B(n3356), .Z(n3355) );
  XOR U3341 ( .A(p_input[236]), .B(n3354), .Z(n3356) );
  XNOR U3342 ( .A(n3357), .B(n3358), .Z(n3354) );
  AND U3343 ( .A(n144), .B(n3353), .Z(n3358) );
  XNOR U3344 ( .A(n3357), .B(n3351), .Z(n3353) );
  XOR U3345 ( .A(n3359), .B(n3360), .Z(n3351) );
  AND U3346 ( .A(n159), .B(n3361), .Z(n3360) );
  XNOR U3347 ( .A(n3362), .B(n3363), .Z(n3357) );
  AND U3348 ( .A(n151), .B(n3364), .Z(n3363) );
  XOR U3349 ( .A(p_input[268]), .B(n3362), .Z(n3364) );
  XNOR U3350 ( .A(n3365), .B(n3366), .Z(n3362) );
  AND U3351 ( .A(n155), .B(n3361), .Z(n3366) );
  XNOR U3352 ( .A(n3365), .B(n3359), .Z(n3361) );
  XOR U3353 ( .A(n3367), .B(n3368), .Z(n3359) );
  AND U3354 ( .A(n170), .B(n3369), .Z(n3368) );
  XNOR U3355 ( .A(n3370), .B(n3371), .Z(n3365) );
  AND U3356 ( .A(n162), .B(n3372), .Z(n3371) );
  XOR U3357 ( .A(p_input[300]), .B(n3370), .Z(n3372) );
  XNOR U3358 ( .A(n3373), .B(n3374), .Z(n3370) );
  AND U3359 ( .A(n166), .B(n3369), .Z(n3374) );
  XNOR U3360 ( .A(n3373), .B(n3367), .Z(n3369) );
  XOR U3361 ( .A(n3375), .B(n3376), .Z(n3367) );
  AND U3362 ( .A(n181), .B(n3377), .Z(n3376) );
  XNOR U3363 ( .A(n3378), .B(n3379), .Z(n3373) );
  AND U3364 ( .A(n173), .B(n3380), .Z(n3379) );
  XOR U3365 ( .A(p_input[332]), .B(n3378), .Z(n3380) );
  XNOR U3366 ( .A(n3381), .B(n3382), .Z(n3378) );
  AND U3367 ( .A(n177), .B(n3377), .Z(n3382) );
  XNOR U3368 ( .A(n3381), .B(n3375), .Z(n3377) );
  XOR U3369 ( .A(n3383), .B(n3384), .Z(n3375) );
  AND U3370 ( .A(n192), .B(n3385), .Z(n3384) );
  XNOR U3371 ( .A(n3386), .B(n3387), .Z(n3381) );
  AND U3372 ( .A(n184), .B(n3388), .Z(n3387) );
  XOR U3373 ( .A(p_input[364]), .B(n3386), .Z(n3388) );
  XNOR U3374 ( .A(n3389), .B(n3390), .Z(n3386) );
  AND U3375 ( .A(n188), .B(n3385), .Z(n3390) );
  XNOR U3376 ( .A(n3389), .B(n3383), .Z(n3385) );
  XOR U3377 ( .A(n3391), .B(n3392), .Z(n3383) );
  AND U3378 ( .A(n203), .B(n3393), .Z(n3392) );
  XNOR U3379 ( .A(n3394), .B(n3395), .Z(n3389) );
  AND U3380 ( .A(n195), .B(n3396), .Z(n3395) );
  XOR U3381 ( .A(p_input[396]), .B(n3394), .Z(n3396) );
  XNOR U3382 ( .A(n3397), .B(n3398), .Z(n3394) );
  AND U3383 ( .A(n199), .B(n3393), .Z(n3398) );
  XNOR U3384 ( .A(n3397), .B(n3391), .Z(n3393) );
  XOR U3385 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n3399), .Z(n3391) );
  AND U3386 ( .A(n213), .B(n3400), .Z(n3399) );
  XNOR U3387 ( .A(n3401), .B(n3402), .Z(n3397) );
  AND U3388 ( .A(n206), .B(n3403), .Z(n3402) );
  XOR U3389 ( .A(p_input[428]), .B(n3401), .Z(n3403) );
  XNOR U3390 ( .A(n3404), .B(n3405), .Z(n3401) );
  AND U3391 ( .A(n210), .B(n3400), .Z(n3405) );
  XOR U3392 ( .A(n3406), .B(n3404), .Z(n3400) );
  IV U3393 ( .A(\knn_comb_/min_val_out[0][12] ), .Z(n3406) );
  IV U3394 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n3404) );
  XOR U3395 ( .A(n53), .B(n3407), .Z(o[11]) );
  AND U3396 ( .A(n58), .B(n3408), .Z(n53) );
  XOR U3397 ( .A(n54), .B(n3407), .Z(n3408) );
  XOR U3398 ( .A(n3409), .B(n3410), .Z(n3407) );
  AND U3399 ( .A(n70), .B(n3411), .Z(n3410) );
  XOR U3400 ( .A(n3412), .B(n3413), .Z(n54) );
  AND U3401 ( .A(n62), .B(n3414), .Z(n3413) );
  XOR U3402 ( .A(p_input[11]), .B(n3412), .Z(n3414) );
  XNOR U3403 ( .A(n3415), .B(n3416), .Z(n3412) );
  AND U3404 ( .A(n66), .B(n3411), .Z(n3416) );
  XNOR U3405 ( .A(n3415), .B(n3409), .Z(n3411) );
  XOR U3406 ( .A(n3417), .B(n3418), .Z(n3409) );
  AND U3407 ( .A(n82), .B(n3419), .Z(n3418) );
  XNOR U3408 ( .A(n3420), .B(n3421), .Z(n3415) );
  AND U3409 ( .A(n74), .B(n3422), .Z(n3421) );
  XOR U3410 ( .A(p_input[43]), .B(n3420), .Z(n3422) );
  XNOR U3411 ( .A(n3423), .B(n3424), .Z(n3420) );
  AND U3412 ( .A(n78), .B(n3419), .Z(n3424) );
  XNOR U3413 ( .A(n3423), .B(n3417), .Z(n3419) );
  XOR U3414 ( .A(n3425), .B(n3426), .Z(n3417) );
  AND U3415 ( .A(n93), .B(n3427), .Z(n3426) );
  XNOR U3416 ( .A(n3428), .B(n3429), .Z(n3423) );
  AND U3417 ( .A(n85), .B(n3430), .Z(n3429) );
  XOR U3418 ( .A(p_input[75]), .B(n3428), .Z(n3430) );
  XNOR U3419 ( .A(n3431), .B(n3432), .Z(n3428) );
  AND U3420 ( .A(n89), .B(n3427), .Z(n3432) );
  XNOR U3421 ( .A(n3431), .B(n3425), .Z(n3427) );
  XOR U3422 ( .A(n3433), .B(n3434), .Z(n3425) );
  AND U3423 ( .A(n104), .B(n3435), .Z(n3434) );
  XNOR U3424 ( .A(n3436), .B(n3437), .Z(n3431) );
  AND U3425 ( .A(n96), .B(n3438), .Z(n3437) );
  XOR U3426 ( .A(p_input[107]), .B(n3436), .Z(n3438) );
  XNOR U3427 ( .A(n3439), .B(n3440), .Z(n3436) );
  AND U3428 ( .A(n100), .B(n3435), .Z(n3440) );
  XNOR U3429 ( .A(n3439), .B(n3433), .Z(n3435) );
  XOR U3430 ( .A(n3441), .B(n3442), .Z(n3433) );
  AND U3431 ( .A(n115), .B(n3443), .Z(n3442) );
  XNOR U3432 ( .A(n3444), .B(n3445), .Z(n3439) );
  AND U3433 ( .A(n107), .B(n3446), .Z(n3445) );
  XOR U3434 ( .A(p_input[139]), .B(n3444), .Z(n3446) );
  XNOR U3435 ( .A(n3447), .B(n3448), .Z(n3444) );
  AND U3436 ( .A(n111), .B(n3443), .Z(n3448) );
  XNOR U3437 ( .A(n3447), .B(n3441), .Z(n3443) );
  XOR U3438 ( .A(n3449), .B(n3450), .Z(n3441) );
  AND U3439 ( .A(n126), .B(n3451), .Z(n3450) );
  XNOR U3440 ( .A(n3452), .B(n3453), .Z(n3447) );
  AND U3441 ( .A(n118), .B(n3454), .Z(n3453) );
  XOR U3442 ( .A(p_input[171]), .B(n3452), .Z(n3454) );
  XNOR U3443 ( .A(n3455), .B(n3456), .Z(n3452) );
  AND U3444 ( .A(n122), .B(n3451), .Z(n3456) );
  XNOR U3445 ( .A(n3455), .B(n3449), .Z(n3451) );
  XOR U3446 ( .A(n3457), .B(n3458), .Z(n3449) );
  AND U3447 ( .A(n137), .B(n3459), .Z(n3458) );
  XNOR U3448 ( .A(n3460), .B(n3461), .Z(n3455) );
  AND U3449 ( .A(n129), .B(n3462), .Z(n3461) );
  XOR U3450 ( .A(p_input[203]), .B(n3460), .Z(n3462) );
  XNOR U3451 ( .A(n3463), .B(n3464), .Z(n3460) );
  AND U3452 ( .A(n133), .B(n3459), .Z(n3464) );
  XNOR U3453 ( .A(n3463), .B(n3457), .Z(n3459) );
  XOR U3454 ( .A(n3465), .B(n3466), .Z(n3457) );
  AND U3455 ( .A(n148), .B(n3467), .Z(n3466) );
  XNOR U3456 ( .A(n3468), .B(n3469), .Z(n3463) );
  AND U3457 ( .A(n140), .B(n3470), .Z(n3469) );
  XOR U3458 ( .A(p_input[235]), .B(n3468), .Z(n3470) );
  XNOR U3459 ( .A(n3471), .B(n3472), .Z(n3468) );
  AND U3460 ( .A(n144), .B(n3467), .Z(n3472) );
  XNOR U3461 ( .A(n3471), .B(n3465), .Z(n3467) );
  XOR U3462 ( .A(n3473), .B(n3474), .Z(n3465) );
  AND U3463 ( .A(n159), .B(n3475), .Z(n3474) );
  XNOR U3464 ( .A(n3476), .B(n3477), .Z(n3471) );
  AND U3465 ( .A(n151), .B(n3478), .Z(n3477) );
  XOR U3466 ( .A(p_input[267]), .B(n3476), .Z(n3478) );
  XNOR U3467 ( .A(n3479), .B(n3480), .Z(n3476) );
  AND U3468 ( .A(n155), .B(n3475), .Z(n3480) );
  XNOR U3469 ( .A(n3479), .B(n3473), .Z(n3475) );
  XOR U3470 ( .A(n3481), .B(n3482), .Z(n3473) );
  AND U3471 ( .A(n170), .B(n3483), .Z(n3482) );
  XNOR U3472 ( .A(n3484), .B(n3485), .Z(n3479) );
  AND U3473 ( .A(n162), .B(n3486), .Z(n3485) );
  XOR U3474 ( .A(p_input[299]), .B(n3484), .Z(n3486) );
  XNOR U3475 ( .A(n3487), .B(n3488), .Z(n3484) );
  AND U3476 ( .A(n166), .B(n3483), .Z(n3488) );
  XNOR U3477 ( .A(n3487), .B(n3481), .Z(n3483) );
  XOR U3478 ( .A(n3489), .B(n3490), .Z(n3481) );
  AND U3479 ( .A(n181), .B(n3491), .Z(n3490) );
  XNOR U3480 ( .A(n3492), .B(n3493), .Z(n3487) );
  AND U3481 ( .A(n173), .B(n3494), .Z(n3493) );
  XOR U3482 ( .A(p_input[331]), .B(n3492), .Z(n3494) );
  XNOR U3483 ( .A(n3495), .B(n3496), .Z(n3492) );
  AND U3484 ( .A(n177), .B(n3491), .Z(n3496) );
  XNOR U3485 ( .A(n3495), .B(n3489), .Z(n3491) );
  XOR U3486 ( .A(n3497), .B(n3498), .Z(n3489) );
  AND U3487 ( .A(n192), .B(n3499), .Z(n3498) );
  XNOR U3488 ( .A(n3500), .B(n3501), .Z(n3495) );
  AND U3489 ( .A(n184), .B(n3502), .Z(n3501) );
  XOR U3490 ( .A(p_input[363]), .B(n3500), .Z(n3502) );
  XNOR U3491 ( .A(n3503), .B(n3504), .Z(n3500) );
  AND U3492 ( .A(n188), .B(n3499), .Z(n3504) );
  XNOR U3493 ( .A(n3503), .B(n3497), .Z(n3499) );
  XOR U3494 ( .A(n3505), .B(n3506), .Z(n3497) );
  AND U3495 ( .A(n203), .B(n3507), .Z(n3506) );
  XNOR U3496 ( .A(n3508), .B(n3509), .Z(n3503) );
  AND U3497 ( .A(n195), .B(n3510), .Z(n3509) );
  XOR U3498 ( .A(p_input[395]), .B(n3508), .Z(n3510) );
  XNOR U3499 ( .A(n3511), .B(n3512), .Z(n3508) );
  AND U3500 ( .A(n199), .B(n3507), .Z(n3512) );
  XNOR U3501 ( .A(n3511), .B(n3505), .Z(n3507) );
  XOR U3502 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n3513), .Z(n3505) );
  AND U3503 ( .A(n213), .B(n3514), .Z(n3513) );
  XNOR U3504 ( .A(n3515), .B(n3516), .Z(n3511) );
  AND U3505 ( .A(n206), .B(n3517), .Z(n3516) );
  XOR U3506 ( .A(p_input[427]), .B(n3515), .Z(n3517) );
  XNOR U3507 ( .A(n3518), .B(n3519), .Z(n3515) );
  AND U3508 ( .A(n210), .B(n3514), .Z(n3519) );
  XOR U3509 ( .A(\knn_comb_/min_val_out[0][11] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n3514) );
  XOR U3510 ( .A(n55), .B(n3520), .Z(o[10]) );
  AND U3511 ( .A(n58), .B(n3521), .Z(n55) );
  XOR U3512 ( .A(n56), .B(n3520), .Z(n3521) );
  XOR U3513 ( .A(n3522), .B(n3523), .Z(n3520) );
  AND U3514 ( .A(n70), .B(n3524), .Z(n3523) );
  XOR U3515 ( .A(n3525), .B(n3526), .Z(n56) );
  AND U3516 ( .A(n62), .B(n3527), .Z(n3526) );
  XOR U3517 ( .A(p_input[10]), .B(n3525), .Z(n3527) );
  XNOR U3518 ( .A(n3528), .B(n3529), .Z(n3525) );
  AND U3519 ( .A(n66), .B(n3524), .Z(n3529) );
  XNOR U3520 ( .A(n3528), .B(n3522), .Z(n3524) );
  XOR U3521 ( .A(n3530), .B(n3531), .Z(n3522) );
  AND U3522 ( .A(n82), .B(n3532), .Z(n3531) );
  XNOR U3523 ( .A(n3533), .B(n3534), .Z(n3528) );
  AND U3524 ( .A(n74), .B(n3535), .Z(n3534) );
  XOR U3525 ( .A(p_input[42]), .B(n3533), .Z(n3535) );
  XNOR U3526 ( .A(n3536), .B(n3537), .Z(n3533) );
  AND U3527 ( .A(n78), .B(n3532), .Z(n3537) );
  XNOR U3528 ( .A(n3536), .B(n3530), .Z(n3532) );
  XOR U3529 ( .A(n3538), .B(n3539), .Z(n3530) );
  AND U3530 ( .A(n93), .B(n3540), .Z(n3539) );
  XNOR U3531 ( .A(n3541), .B(n3542), .Z(n3536) );
  AND U3532 ( .A(n85), .B(n3543), .Z(n3542) );
  XOR U3533 ( .A(p_input[74]), .B(n3541), .Z(n3543) );
  XNOR U3534 ( .A(n3544), .B(n3545), .Z(n3541) );
  AND U3535 ( .A(n89), .B(n3540), .Z(n3545) );
  XNOR U3536 ( .A(n3544), .B(n3538), .Z(n3540) );
  XOR U3537 ( .A(n3546), .B(n3547), .Z(n3538) );
  AND U3538 ( .A(n104), .B(n3548), .Z(n3547) );
  XNOR U3539 ( .A(n3549), .B(n3550), .Z(n3544) );
  AND U3540 ( .A(n96), .B(n3551), .Z(n3550) );
  XOR U3541 ( .A(p_input[106]), .B(n3549), .Z(n3551) );
  XNOR U3542 ( .A(n3552), .B(n3553), .Z(n3549) );
  AND U3543 ( .A(n100), .B(n3548), .Z(n3553) );
  XNOR U3544 ( .A(n3552), .B(n3546), .Z(n3548) );
  XOR U3545 ( .A(n3554), .B(n3555), .Z(n3546) );
  AND U3546 ( .A(n115), .B(n3556), .Z(n3555) );
  XNOR U3547 ( .A(n3557), .B(n3558), .Z(n3552) );
  AND U3548 ( .A(n107), .B(n3559), .Z(n3558) );
  XOR U3549 ( .A(p_input[138]), .B(n3557), .Z(n3559) );
  XNOR U3550 ( .A(n3560), .B(n3561), .Z(n3557) );
  AND U3551 ( .A(n111), .B(n3556), .Z(n3561) );
  XNOR U3552 ( .A(n3560), .B(n3554), .Z(n3556) );
  XOR U3553 ( .A(n3562), .B(n3563), .Z(n3554) );
  AND U3554 ( .A(n126), .B(n3564), .Z(n3563) );
  XNOR U3555 ( .A(n3565), .B(n3566), .Z(n3560) );
  AND U3556 ( .A(n118), .B(n3567), .Z(n3566) );
  XOR U3557 ( .A(p_input[170]), .B(n3565), .Z(n3567) );
  XNOR U3558 ( .A(n3568), .B(n3569), .Z(n3565) );
  AND U3559 ( .A(n122), .B(n3564), .Z(n3569) );
  XNOR U3560 ( .A(n3568), .B(n3562), .Z(n3564) );
  XOR U3561 ( .A(n3570), .B(n3571), .Z(n3562) );
  AND U3562 ( .A(n137), .B(n3572), .Z(n3571) );
  XNOR U3563 ( .A(n3573), .B(n3574), .Z(n3568) );
  AND U3564 ( .A(n129), .B(n3575), .Z(n3574) );
  XOR U3565 ( .A(p_input[202]), .B(n3573), .Z(n3575) );
  XNOR U3566 ( .A(n3576), .B(n3577), .Z(n3573) );
  AND U3567 ( .A(n133), .B(n3572), .Z(n3577) );
  XNOR U3568 ( .A(n3576), .B(n3570), .Z(n3572) );
  XOR U3569 ( .A(n3578), .B(n3579), .Z(n3570) );
  AND U3570 ( .A(n148), .B(n3580), .Z(n3579) );
  XNOR U3571 ( .A(n3581), .B(n3582), .Z(n3576) );
  AND U3572 ( .A(n140), .B(n3583), .Z(n3582) );
  XOR U3573 ( .A(p_input[234]), .B(n3581), .Z(n3583) );
  XNOR U3574 ( .A(n3584), .B(n3585), .Z(n3581) );
  AND U3575 ( .A(n144), .B(n3580), .Z(n3585) );
  XNOR U3576 ( .A(n3584), .B(n3578), .Z(n3580) );
  XOR U3577 ( .A(n3586), .B(n3587), .Z(n3578) );
  AND U3578 ( .A(n159), .B(n3588), .Z(n3587) );
  XNOR U3579 ( .A(n3589), .B(n3590), .Z(n3584) );
  AND U3580 ( .A(n151), .B(n3591), .Z(n3590) );
  XOR U3581 ( .A(p_input[266]), .B(n3589), .Z(n3591) );
  XNOR U3582 ( .A(n3592), .B(n3593), .Z(n3589) );
  AND U3583 ( .A(n155), .B(n3588), .Z(n3593) );
  XNOR U3584 ( .A(n3592), .B(n3586), .Z(n3588) );
  XOR U3585 ( .A(n3594), .B(n3595), .Z(n3586) );
  AND U3586 ( .A(n170), .B(n3596), .Z(n3595) );
  XNOR U3587 ( .A(n3597), .B(n3598), .Z(n3592) );
  AND U3588 ( .A(n162), .B(n3599), .Z(n3598) );
  XOR U3589 ( .A(p_input[298]), .B(n3597), .Z(n3599) );
  XNOR U3590 ( .A(n3600), .B(n3601), .Z(n3597) );
  AND U3591 ( .A(n166), .B(n3596), .Z(n3601) );
  XNOR U3592 ( .A(n3600), .B(n3594), .Z(n3596) );
  XOR U3593 ( .A(n3602), .B(n3603), .Z(n3594) );
  AND U3594 ( .A(n181), .B(n3604), .Z(n3603) );
  XNOR U3595 ( .A(n3605), .B(n3606), .Z(n3600) );
  AND U3596 ( .A(n173), .B(n3607), .Z(n3606) );
  XOR U3597 ( .A(p_input[330]), .B(n3605), .Z(n3607) );
  XNOR U3598 ( .A(n3608), .B(n3609), .Z(n3605) );
  AND U3599 ( .A(n177), .B(n3604), .Z(n3609) );
  XNOR U3600 ( .A(n3608), .B(n3602), .Z(n3604) );
  XOR U3601 ( .A(n3610), .B(n3611), .Z(n3602) );
  AND U3602 ( .A(n192), .B(n3612), .Z(n3611) );
  XNOR U3603 ( .A(n3613), .B(n3614), .Z(n3608) );
  AND U3604 ( .A(n184), .B(n3615), .Z(n3614) );
  XOR U3605 ( .A(p_input[362]), .B(n3613), .Z(n3615) );
  XNOR U3606 ( .A(n3616), .B(n3617), .Z(n3613) );
  AND U3607 ( .A(n188), .B(n3612), .Z(n3617) );
  XNOR U3608 ( .A(n3616), .B(n3610), .Z(n3612) );
  XOR U3609 ( .A(n3618), .B(n3619), .Z(n3610) );
  AND U3610 ( .A(n203), .B(n3620), .Z(n3619) );
  XNOR U3611 ( .A(n3621), .B(n3622), .Z(n3616) );
  AND U3612 ( .A(n195), .B(n3623), .Z(n3622) );
  XOR U3613 ( .A(p_input[394]), .B(n3621), .Z(n3623) );
  XNOR U3614 ( .A(n3624), .B(n3625), .Z(n3621) );
  AND U3615 ( .A(n199), .B(n3620), .Z(n3625) );
  XNOR U3616 ( .A(n3624), .B(n3618), .Z(n3620) );
  XOR U3617 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n3626), .Z(n3618) );
  AND U3618 ( .A(n213), .B(n3627), .Z(n3626) );
  XNOR U3619 ( .A(n3628), .B(n3629), .Z(n3624) );
  AND U3620 ( .A(n206), .B(n3630), .Z(n3629) );
  XOR U3621 ( .A(p_input[426]), .B(n3628), .Z(n3630) );
  XNOR U3622 ( .A(n3631), .B(n3632), .Z(n3628) );
  AND U3623 ( .A(n210), .B(n3627), .Z(n3632) );
  XOR U3624 ( .A(\knn_comb_/min_val_out[0][10] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n3627) );
  XOR U3625 ( .A(n911), .B(n3633), .Z(o[0]) );
  AND U3626 ( .A(n58), .B(n3634), .Z(n911) );
  XOR U3627 ( .A(n912), .B(n3633), .Z(n3634) );
  XOR U3628 ( .A(n3635), .B(n3636), .Z(n3633) );
  AND U3629 ( .A(n70), .B(n3637), .Z(n3636) );
  XOR U3630 ( .A(n3638), .B(n3639), .Z(n912) );
  AND U3631 ( .A(n62), .B(n3640), .Z(n3639) );
  XOR U3632 ( .A(p_input[0]), .B(n3638), .Z(n3640) );
  XNOR U3633 ( .A(n3641), .B(n3642), .Z(n3638) );
  AND U3634 ( .A(n66), .B(n3637), .Z(n3642) );
  XNOR U3635 ( .A(n3641), .B(n3635), .Z(n3637) );
  XOR U3636 ( .A(n3643), .B(n3644), .Z(n3635) );
  AND U3637 ( .A(n82), .B(n3645), .Z(n3644) );
  XNOR U3638 ( .A(n3646), .B(n3647), .Z(n3641) );
  AND U3639 ( .A(n74), .B(n3648), .Z(n3647) );
  XOR U3640 ( .A(p_input[32]), .B(n3646), .Z(n3648) );
  XNOR U3641 ( .A(n3649), .B(n3650), .Z(n3646) );
  AND U3642 ( .A(n78), .B(n3645), .Z(n3650) );
  XNOR U3643 ( .A(n3649), .B(n3643), .Z(n3645) );
  XOR U3644 ( .A(n3651), .B(n3652), .Z(n3643) );
  AND U3645 ( .A(n93), .B(n3653), .Z(n3652) );
  XNOR U3646 ( .A(n3654), .B(n3655), .Z(n3649) );
  AND U3647 ( .A(n85), .B(n3656), .Z(n3655) );
  XOR U3648 ( .A(p_input[64]), .B(n3654), .Z(n3656) );
  XNOR U3649 ( .A(n3657), .B(n3658), .Z(n3654) );
  AND U3650 ( .A(n89), .B(n3653), .Z(n3658) );
  XNOR U3651 ( .A(n3657), .B(n3651), .Z(n3653) );
  XOR U3652 ( .A(n3659), .B(n3660), .Z(n3651) );
  AND U3653 ( .A(n104), .B(n3661), .Z(n3660) );
  XNOR U3654 ( .A(n3662), .B(n3663), .Z(n3657) );
  AND U3655 ( .A(n96), .B(n3664), .Z(n3663) );
  XOR U3656 ( .A(p_input[96]), .B(n3662), .Z(n3664) );
  XNOR U3657 ( .A(n3665), .B(n3666), .Z(n3662) );
  AND U3658 ( .A(n100), .B(n3661), .Z(n3666) );
  XNOR U3659 ( .A(n3665), .B(n3659), .Z(n3661) );
  XOR U3660 ( .A(n3667), .B(n3668), .Z(n3659) );
  AND U3661 ( .A(n115), .B(n3669), .Z(n3668) );
  XNOR U3662 ( .A(n3670), .B(n3671), .Z(n3665) );
  AND U3663 ( .A(n107), .B(n3672), .Z(n3671) );
  XOR U3664 ( .A(p_input[128]), .B(n3670), .Z(n3672) );
  XNOR U3665 ( .A(n3673), .B(n3674), .Z(n3670) );
  AND U3666 ( .A(n111), .B(n3669), .Z(n3674) );
  XNOR U3667 ( .A(n3673), .B(n3667), .Z(n3669) );
  XOR U3668 ( .A(n3675), .B(n3676), .Z(n3667) );
  AND U3669 ( .A(n126), .B(n3677), .Z(n3676) );
  XNOR U3670 ( .A(n3678), .B(n3679), .Z(n3673) );
  AND U3671 ( .A(n118), .B(n3680), .Z(n3679) );
  XOR U3672 ( .A(p_input[160]), .B(n3678), .Z(n3680) );
  XNOR U3673 ( .A(n3681), .B(n3682), .Z(n3678) );
  AND U3674 ( .A(n122), .B(n3677), .Z(n3682) );
  XNOR U3675 ( .A(n3681), .B(n3675), .Z(n3677) );
  XOR U3676 ( .A(n3683), .B(n3684), .Z(n3675) );
  AND U3677 ( .A(n137), .B(n3685), .Z(n3684) );
  XNOR U3678 ( .A(n3686), .B(n3687), .Z(n3681) );
  AND U3679 ( .A(n129), .B(n3688), .Z(n3687) );
  XOR U3680 ( .A(p_input[192]), .B(n3686), .Z(n3688) );
  XNOR U3681 ( .A(n3689), .B(n3690), .Z(n3686) );
  AND U3682 ( .A(n133), .B(n3685), .Z(n3690) );
  XNOR U3683 ( .A(n3689), .B(n3683), .Z(n3685) );
  XOR U3684 ( .A(n3691), .B(n3692), .Z(n3683) );
  AND U3685 ( .A(n148), .B(n3693), .Z(n3692) );
  XNOR U3686 ( .A(n3694), .B(n3695), .Z(n3689) );
  AND U3687 ( .A(n140), .B(n3696), .Z(n3695) );
  XOR U3688 ( .A(p_input[224]), .B(n3694), .Z(n3696) );
  XNOR U3689 ( .A(n3697), .B(n3698), .Z(n3694) );
  AND U3690 ( .A(n144), .B(n3693), .Z(n3698) );
  XNOR U3691 ( .A(n3697), .B(n3691), .Z(n3693) );
  XOR U3692 ( .A(n3699), .B(n3700), .Z(n3691) );
  AND U3693 ( .A(n159), .B(n3701), .Z(n3700) );
  XNOR U3694 ( .A(n3702), .B(n3703), .Z(n3697) );
  AND U3695 ( .A(n151), .B(n3704), .Z(n3703) );
  XOR U3696 ( .A(p_input[256]), .B(n3702), .Z(n3704) );
  XNOR U3697 ( .A(n3705), .B(n3706), .Z(n3702) );
  AND U3698 ( .A(n155), .B(n3701), .Z(n3706) );
  XNOR U3699 ( .A(n3705), .B(n3699), .Z(n3701) );
  XOR U3700 ( .A(n3707), .B(n3708), .Z(n3699) );
  AND U3701 ( .A(n170), .B(n3709), .Z(n3708) );
  XNOR U3702 ( .A(n3710), .B(n3711), .Z(n3705) );
  AND U3703 ( .A(n162), .B(n3712), .Z(n3711) );
  XOR U3704 ( .A(p_input[288]), .B(n3710), .Z(n3712) );
  XNOR U3705 ( .A(n3713), .B(n3714), .Z(n3710) );
  AND U3706 ( .A(n166), .B(n3709), .Z(n3714) );
  XNOR U3707 ( .A(n3713), .B(n3707), .Z(n3709) );
  XOR U3708 ( .A(n3715), .B(n3716), .Z(n3707) );
  AND U3709 ( .A(n181), .B(n3717), .Z(n3716) );
  XNOR U3710 ( .A(n3718), .B(n3719), .Z(n3713) );
  AND U3711 ( .A(n173), .B(n3720), .Z(n3719) );
  XOR U3712 ( .A(p_input[320]), .B(n3718), .Z(n3720) );
  XNOR U3713 ( .A(n3721), .B(n3722), .Z(n3718) );
  AND U3714 ( .A(n177), .B(n3717), .Z(n3722) );
  XNOR U3715 ( .A(n3721), .B(n3715), .Z(n3717) );
  XOR U3716 ( .A(n3723), .B(n3724), .Z(n3715) );
  AND U3717 ( .A(n192), .B(n3725), .Z(n3724) );
  XNOR U3718 ( .A(n3726), .B(n3727), .Z(n3721) );
  AND U3719 ( .A(n184), .B(n3728), .Z(n3727) );
  XOR U3720 ( .A(p_input[352]), .B(n3726), .Z(n3728) );
  XNOR U3721 ( .A(n3729), .B(n3730), .Z(n3726) );
  AND U3722 ( .A(n188), .B(n3725), .Z(n3730) );
  XNOR U3723 ( .A(n3729), .B(n3723), .Z(n3725) );
  XOR U3724 ( .A(n3731), .B(n3732), .Z(n3723) );
  AND U3725 ( .A(n203), .B(n3733), .Z(n3732) );
  XNOR U3726 ( .A(n3734), .B(n3735), .Z(n3729) );
  AND U3727 ( .A(n195), .B(n3736), .Z(n3735) );
  XOR U3728 ( .A(p_input[384]), .B(n3734), .Z(n3736) );
  XNOR U3729 ( .A(n3737), .B(n3738), .Z(n3734) );
  AND U3730 ( .A(n199), .B(n3733), .Z(n3738) );
  XNOR U3731 ( .A(n3737), .B(n3731), .Z(n3733) );
  XOR U3732 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n3739), .Z(n3731) );
  AND U3733 ( .A(n213), .B(n3740), .Z(n3739) );
  XNOR U3734 ( .A(n3741), .B(n3742), .Z(n3737) );
  AND U3735 ( .A(n206), .B(n3743), .Z(n3742) );
  XOR U3736 ( .A(p_input[416]), .B(n3741), .Z(n3743) );
  XNOR U3737 ( .A(n3744), .B(n3745), .Z(n3741) );
  AND U3738 ( .A(n210), .B(n3740), .Z(n3745) );
  XOR U3739 ( .A(\knn_comb_/min_val_out[0][0] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n3740) );
  IV U3740 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n3744) );
  XNOR U3741 ( .A(n3746), .B(n3747), .Z(n58) );
  AND U3742 ( .A(n3748), .B(n3749), .Z(n3747) );
  XNOR U3743 ( .A(n3746), .B(n3750), .Z(n3749) );
  XOR U3744 ( .A(n3751), .B(n3752), .Z(n3750) );
  AND U3745 ( .A(n62), .B(n3753), .Z(n3752) );
  XNOR U3746 ( .A(n3751), .B(n3754), .Z(n3753) );
  XNOR U3747 ( .A(n3746), .B(n3755), .Z(n3748) );
  XOR U3748 ( .A(n3756), .B(n3757), .Z(n3755) );
  AND U3749 ( .A(n70), .B(n3758), .Z(n3757) );
  XOR U3750 ( .A(n3759), .B(n3760), .Z(n3746) );
  AND U3751 ( .A(n3761), .B(n3762), .Z(n3760) );
  XOR U3752 ( .A(n3763), .B(n3759), .Z(n3762) );
  XOR U3753 ( .A(n3764), .B(n3765), .Z(n3763) );
  AND U3754 ( .A(n62), .B(n3766), .Z(n3765) );
  XOR U3755 ( .A(n3767), .B(n3764), .Z(n3766) );
  XNOR U3756 ( .A(n3759), .B(n3768), .Z(n3761) );
  XOR U3757 ( .A(n3769), .B(n3770), .Z(n3768) );
  AND U3758 ( .A(n70), .B(n3771), .Z(n3770) );
  XOR U3759 ( .A(n3772), .B(n3773), .Z(n3759) );
  AND U3760 ( .A(n3774), .B(n3775), .Z(n3773) );
  XOR U3761 ( .A(n3776), .B(n3772), .Z(n3775) );
  XOR U3762 ( .A(n3777), .B(n3778), .Z(n3776) );
  AND U3763 ( .A(n62), .B(n3779), .Z(n3778) );
  XNOR U3764 ( .A(n3780), .B(n3777), .Z(n3779) );
  XNOR U3765 ( .A(n3772), .B(n3781), .Z(n3774) );
  XOR U3766 ( .A(n3782), .B(n3783), .Z(n3781) );
  AND U3767 ( .A(n70), .B(n3784), .Z(n3783) );
  XOR U3768 ( .A(n3785), .B(n3786), .Z(n3772) );
  AND U3769 ( .A(n3787), .B(n3788), .Z(n3786) );
  XOR U3770 ( .A(n3789), .B(n3785), .Z(n3788) );
  XOR U3771 ( .A(n3790), .B(n3791), .Z(n3789) );
  AND U3772 ( .A(n62), .B(n3792), .Z(n3791) );
  XOR U3773 ( .A(n3793), .B(n3790), .Z(n3792) );
  XNOR U3774 ( .A(n3785), .B(n3794), .Z(n3787) );
  XOR U3775 ( .A(n3795), .B(n3796), .Z(n3794) );
  AND U3776 ( .A(n70), .B(n3797), .Z(n3796) );
  XOR U3777 ( .A(n3798), .B(n3799), .Z(n3785) );
  AND U3778 ( .A(n3800), .B(n3801), .Z(n3799) );
  XOR U3779 ( .A(n3798), .B(n3802), .Z(n3801) );
  XOR U3780 ( .A(n3803), .B(n3804), .Z(n3802) );
  AND U3781 ( .A(n62), .B(n3805), .Z(n3804) );
  XNOR U3782 ( .A(n3806), .B(n3803), .Z(n3805) );
  XNOR U3783 ( .A(n3807), .B(n3798), .Z(n3800) );
  XNOR U3784 ( .A(n3808), .B(n3809), .Z(n3807) );
  AND U3785 ( .A(n70), .B(n3810), .Z(n3809) );
  AND U3786 ( .A(n3811), .B(n3812), .Z(n3798) );
  XNOR U3787 ( .A(n3813), .B(n3814), .Z(n3812) );
  AND U3788 ( .A(n62), .B(n3815), .Z(n3814) );
  XNOR U3789 ( .A(n3816), .B(n3813), .Z(n3815) );
  XNOR U3790 ( .A(n3817), .B(n3818), .Z(n62) );
  AND U3791 ( .A(n3819), .B(n3820), .Z(n3818) );
  XOR U3792 ( .A(n3754), .B(n3817), .Z(n3820) );
  AND U3793 ( .A(n3821), .B(n3822), .Z(n3754) );
  XOR U3794 ( .A(n3817), .B(n3751), .Z(n3819) );
  XNOR U3795 ( .A(n3823), .B(n3824), .Z(n3751) );
  AND U3796 ( .A(n66), .B(n3758), .Z(n3824) );
  XOR U3797 ( .A(n3756), .B(n3823), .Z(n3758) );
  XOR U3798 ( .A(n3825), .B(n3826), .Z(n3817) );
  AND U3799 ( .A(n3827), .B(n3828), .Z(n3826) );
  XNOR U3800 ( .A(n3825), .B(n3821), .Z(n3828) );
  IV U3801 ( .A(n3767), .Z(n3821) );
  XOR U3802 ( .A(n3829), .B(n3830), .Z(n3767) );
  XOR U3803 ( .A(n3831), .B(n3822), .Z(n3830) );
  AND U3804 ( .A(n3780), .B(n3832), .Z(n3822) );
  AND U3805 ( .A(n3833), .B(n3834), .Z(n3831) );
  XOR U3806 ( .A(n3835), .B(n3829), .Z(n3833) );
  XNOR U3807 ( .A(n3764), .B(n3825), .Z(n3827) );
  XNOR U3808 ( .A(n3836), .B(n3837), .Z(n3764) );
  AND U3809 ( .A(n66), .B(n3771), .Z(n3837) );
  XOR U3810 ( .A(n3836), .B(n3838), .Z(n3771) );
  XOR U3811 ( .A(n3839), .B(n3840), .Z(n3825) );
  AND U3812 ( .A(n3841), .B(n3842), .Z(n3840) );
  XNOR U3813 ( .A(n3839), .B(n3780), .Z(n3842) );
  XOR U3814 ( .A(n3843), .B(n3834), .Z(n3780) );
  XNOR U3815 ( .A(n3844), .B(n3829), .Z(n3834) );
  XOR U3816 ( .A(n3845), .B(n3846), .Z(n3829) );
  AND U3817 ( .A(n3847), .B(n3848), .Z(n3846) );
  XOR U3818 ( .A(n3849), .B(n3845), .Z(n3847) );
  XNOR U3819 ( .A(n3850), .B(n3851), .Z(n3844) );
  AND U3820 ( .A(n3852), .B(n3853), .Z(n3851) );
  XOR U3821 ( .A(n3850), .B(n3854), .Z(n3852) );
  XNOR U3822 ( .A(n3835), .B(n3832), .Z(n3843) );
  AND U3823 ( .A(n3855), .B(n3856), .Z(n3832) );
  XOR U3824 ( .A(n3857), .B(n3858), .Z(n3835) );
  AND U3825 ( .A(n3859), .B(n3860), .Z(n3858) );
  XOR U3826 ( .A(n3857), .B(n3861), .Z(n3859) );
  XNOR U3827 ( .A(n3777), .B(n3839), .Z(n3841) );
  XNOR U3828 ( .A(n3862), .B(n3863), .Z(n3777) );
  AND U3829 ( .A(n66), .B(n3784), .Z(n3863) );
  XOR U3830 ( .A(n3862), .B(n3864), .Z(n3784) );
  XOR U3831 ( .A(n3865), .B(n3866), .Z(n3839) );
  AND U3832 ( .A(n3867), .B(n3868), .Z(n3866) );
  XNOR U3833 ( .A(n3865), .B(n3855), .Z(n3868) );
  IV U3834 ( .A(n3793), .Z(n3855) );
  XNOR U3835 ( .A(n3869), .B(n3848), .Z(n3793) );
  XNOR U3836 ( .A(n3870), .B(n3854), .Z(n3848) );
  XOR U3837 ( .A(n3871), .B(n3872), .Z(n3854) );
  AND U3838 ( .A(n3873), .B(n3874), .Z(n3872) );
  XOR U3839 ( .A(n3871), .B(n3875), .Z(n3873) );
  XNOR U3840 ( .A(n3853), .B(n3845), .Z(n3870) );
  XOR U3841 ( .A(n3876), .B(n3877), .Z(n3845) );
  AND U3842 ( .A(n3878), .B(n3879), .Z(n3877) );
  XNOR U3843 ( .A(n3880), .B(n3876), .Z(n3878) );
  XNOR U3844 ( .A(n3881), .B(n3850), .Z(n3853) );
  XOR U3845 ( .A(n3882), .B(n3883), .Z(n3850) );
  AND U3846 ( .A(n3884), .B(n3885), .Z(n3883) );
  XOR U3847 ( .A(n3882), .B(n3886), .Z(n3884) );
  XNOR U3848 ( .A(n3887), .B(n3888), .Z(n3881) );
  AND U3849 ( .A(n3889), .B(n3890), .Z(n3888) );
  XNOR U3850 ( .A(n3887), .B(n3891), .Z(n3889) );
  XNOR U3851 ( .A(n3849), .B(n3856), .Z(n3869) );
  AND U3852 ( .A(n3806), .B(n3892), .Z(n3856) );
  XOR U3853 ( .A(n3861), .B(n3860), .Z(n3849) );
  XNOR U3854 ( .A(n3893), .B(n3857), .Z(n3860) );
  XOR U3855 ( .A(n3894), .B(n3895), .Z(n3857) );
  AND U3856 ( .A(n3896), .B(n3897), .Z(n3895) );
  XOR U3857 ( .A(n3894), .B(n3898), .Z(n3896) );
  XNOR U3858 ( .A(n3899), .B(n3900), .Z(n3893) );
  AND U3859 ( .A(n3901), .B(n3902), .Z(n3900) );
  XOR U3860 ( .A(n3899), .B(n3903), .Z(n3901) );
  XOR U3861 ( .A(n3904), .B(n3905), .Z(n3861) );
  AND U3862 ( .A(n3906), .B(n3907), .Z(n3905) );
  XOR U3863 ( .A(n3904), .B(n3908), .Z(n3906) );
  XNOR U3864 ( .A(n3790), .B(n3865), .Z(n3867) );
  XNOR U3865 ( .A(n3909), .B(n3910), .Z(n3790) );
  AND U3866 ( .A(n66), .B(n3797), .Z(n3910) );
  XOR U3867 ( .A(n3909), .B(n3911), .Z(n3797) );
  XOR U3868 ( .A(n3912), .B(n3913), .Z(n3865) );
  AND U3869 ( .A(n3914), .B(n3915), .Z(n3913) );
  XNOR U3870 ( .A(n3912), .B(n3806), .Z(n3915) );
  XOR U3871 ( .A(n3916), .B(n3879), .Z(n3806) );
  XNOR U3872 ( .A(n3917), .B(n3886), .Z(n3879) );
  XOR U3873 ( .A(n3875), .B(n3874), .Z(n3886) );
  XNOR U3874 ( .A(n3918), .B(n3871), .Z(n3874) );
  XOR U3875 ( .A(n3919), .B(n3920), .Z(n3871) );
  AND U3876 ( .A(n3921), .B(n3922), .Z(n3920) );
  XNOR U3877 ( .A(n3923), .B(n3924), .Z(n3921) );
  IV U3878 ( .A(n3919), .Z(n3923) );
  XNOR U3879 ( .A(n3925), .B(n3926), .Z(n3918) );
  NOR U3880 ( .A(n3927), .B(n3928), .Z(n3926) );
  XNOR U3881 ( .A(n3925), .B(n3929), .Z(n3927) );
  XOR U3882 ( .A(n3930), .B(n3931), .Z(n3875) );
  NOR U3883 ( .A(n3932), .B(n3933), .Z(n3931) );
  XNOR U3884 ( .A(n3930), .B(n3934), .Z(n3932) );
  XNOR U3885 ( .A(n3885), .B(n3876), .Z(n3917) );
  XOR U3886 ( .A(n3935), .B(n3936), .Z(n3876) );
  AND U3887 ( .A(n3937), .B(n3938), .Z(n3936) );
  XOR U3888 ( .A(n3935), .B(n3939), .Z(n3937) );
  XOR U3889 ( .A(n3940), .B(n3891), .Z(n3885) );
  XOR U3890 ( .A(n3941), .B(n3942), .Z(n3891) );
  NOR U3891 ( .A(n3943), .B(n3944), .Z(n3942) );
  XOR U3892 ( .A(n3941), .B(n3945), .Z(n3943) );
  XNOR U3893 ( .A(n3890), .B(n3882), .Z(n3940) );
  XOR U3894 ( .A(n3946), .B(n3947), .Z(n3882) );
  AND U3895 ( .A(n3948), .B(n3949), .Z(n3947) );
  XOR U3896 ( .A(n3946), .B(n3950), .Z(n3948) );
  XNOR U3897 ( .A(n3951), .B(n3887), .Z(n3890) );
  XOR U3898 ( .A(n3952), .B(n3953), .Z(n3887) );
  AND U3899 ( .A(n3954), .B(n3955), .Z(n3953) );
  XNOR U3900 ( .A(n3956), .B(n3957), .Z(n3954) );
  IV U3901 ( .A(n3952), .Z(n3956) );
  XNOR U3902 ( .A(n3958), .B(n3959), .Z(n3951) );
  NOR U3903 ( .A(n3960), .B(n3961), .Z(n3959) );
  XNOR U3904 ( .A(n3958), .B(n3962), .Z(n3960) );
  XOR U3905 ( .A(n3880), .B(n3892), .Z(n3916) );
  NOR U3906 ( .A(n3816), .B(n3963), .Z(n3892) );
  XNOR U3907 ( .A(n3898), .B(n3897), .Z(n3880) );
  XNOR U3908 ( .A(n3964), .B(n3903), .Z(n3897) );
  XNOR U3909 ( .A(n3965), .B(n3966), .Z(n3903) );
  NOR U3910 ( .A(n3967), .B(n3968), .Z(n3966) );
  XOR U3911 ( .A(n3965), .B(n3969), .Z(n3967) );
  XNOR U3912 ( .A(n3902), .B(n3894), .Z(n3964) );
  XOR U3913 ( .A(n3970), .B(n3971), .Z(n3894) );
  AND U3914 ( .A(n3972), .B(n3973), .Z(n3971) );
  XNOR U3915 ( .A(n3970), .B(n3974), .Z(n3972) );
  XNOR U3916 ( .A(n3975), .B(n3899), .Z(n3902) );
  XOR U3917 ( .A(n3976), .B(n3977), .Z(n3899) );
  AND U3918 ( .A(n3978), .B(n3979), .Z(n3977) );
  XNOR U3919 ( .A(n3980), .B(n3981), .Z(n3978) );
  IV U3920 ( .A(n3976), .Z(n3980) );
  XNOR U3921 ( .A(n3982), .B(n3983), .Z(n3975) );
  NOR U3922 ( .A(n3984), .B(n3985), .Z(n3983) );
  XNOR U3923 ( .A(n3982), .B(n3986), .Z(n3984) );
  XOR U3924 ( .A(n3908), .B(n3907), .Z(n3898) );
  XNOR U3925 ( .A(n3987), .B(n3904), .Z(n3907) );
  XOR U3926 ( .A(n3988), .B(n3989), .Z(n3904) );
  AND U3927 ( .A(n3990), .B(n3991), .Z(n3989) );
  XNOR U3928 ( .A(n3992), .B(n3993), .Z(n3990) );
  IV U3929 ( .A(n3988), .Z(n3992) );
  XNOR U3930 ( .A(n3994), .B(n3995), .Z(n3987) );
  NOR U3931 ( .A(n3996), .B(n3997), .Z(n3995) );
  XNOR U3932 ( .A(n3994), .B(n3998), .Z(n3996) );
  XOR U3933 ( .A(n3999), .B(n4000), .Z(n3908) );
  NOR U3934 ( .A(n4001), .B(n4002), .Z(n4000) );
  XNOR U3935 ( .A(n3999), .B(n4003), .Z(n4001) );
  XNOR U3936 ( .A(n3803), .B(n3912), .Z(n3914) );
  XNOR U3937 ( .A(n4004), .B(n4005), .Z(n3803) );
  AND U3938 ( .A(n66), .B(n3810), .Z(n4005) );
  XOR U3939 ( .A(n4004), .B(n3808), .Z(n3810) );
  AND U3940 ( .A(n3813), .B(n3816), .Z(n3912) );
  XOR U3941 ( .A(n4006), .B(n3963), .Z(n3816) );
  XNOR U3942 ( .A(p_input[0]), .B(p_input[512]), .Z(n3963) );
  XNOR U3943 ( .A(n3939), .B(n3938), .Z(n4006) );
  XNOR U3944 ( .A(n4007), .B(n3950), .Z(n3938) );
  XOR U3945 ( .A(n3924), .B(n3922), .Z(n3950) );
  XNOR U3946 ( .A(n4008), .B(n3929), .Z(n3922) );
  XOR U3947 ( .A(p_input[24]), .B(p_input[536]), .Z(n3929) );
  XOR U3948 ( .A(n3919), .B(n3928), .Z(n4008) );
  XOR U3949 ( .A(n4009), .B(n3925), .Z(n3928) );
  XOR U3950 ( .A(p_input[22]), .B(p_input[534]), .Z(n3925) );
  XOR U3951 ( .A(p_input[23]), .B(n4010), .Z(n4009) );
  XOR U3952 ( .A(p_input[18]), .B(p_input[530]), .Z(n3919) );
  XNOR U3953 ( .A(n3934), .B(n3933), .Z(n3924) );
  XOR U3954 ( .A(n4011), .B(n3930), .Z(n3933) );
  XOR U3955 ( .A(p_input[19]), .B(p_input[531]), .Z(n3930) );
  XOR U3956 ( .A(p_input[20]), .B(n4012), .Z(n4011) );
  XOR U3957 ( .A(p_input[21]), .B(p_input[533]), .Z(n3934) );
  XOR U3958 ( .A(n3949), .B(n4013), .Z(n4007) );
  IV U3959 ( .A(n3935), .Z(n4013) );
  XOR U3960 ( .A(p_input[1]), .B(p_input[513]), .Z(n3935) );
  XNOR U3961 ( .A(n4014), .B(n3957), .Z(n3949) );
  XNOR U3962 ( .A(n3945), .B(n3944), .Z(n3957) );
  XNOR U3963 ( .A(n4015), .B(n3941), .Z(n3944) );
  XNOR U3964 ( .A(p_input[26]), .B(p_input[538]), .Z(n3941) );
  XOR U3965 ( .A(p_input[27]), .B(n4016), .Z(n4015) );
  XOR U3966 ( .A(p_input[28]), .B(p_input[540]), .Z(n3945) );
  XOR U3967 ( .A(n3955), .B(n4017), .Z(n4014) );
  IV U3968 ( .A(n3946), .Z(n4017) );
  XOR U3969 ( .A(p_input[17]), .B(p_input[529]), .Z(n3946) );
  XNOR U3970 ( .A(n4018), .B(n3962), .Z(n3955) );
  XNOR U3971 ( .A(p_input[31]), .B(n4019), .Z(n3962) );
  XOR U3972 ( .A(n3952), .B(n3961), .Z(n4018) );
  XOR U3973 ( .A(n4020), .B(n3958), .Z(n3961) );
  XOR U3974 ( .A(p_input[29]), .B(p_input[541]), .Z(n3958) );
  XOR U3975 ( .A(p_input[30]), .B(n4021), .Z(n4020) );
  XOR U3976 ( .A(p_input[25]), .B(p_input[537]), .Z(n3952) );
  XNOR U3977 ( .A(n3974), .B(n3973), .Z(n3939) );
  XNOR U3978 ( .A(n4022), .B(n3981), .Z(n3973) );
  XNOR U3979 ( .A(n3969), .B(n3968), .Z(n3981) );
  XNOR U3980 ( .A(n4023), .B(n3965), .Z(n3968) );
  XNOR U3981 ( .A(p_input[11]), .B(p_input[523]), .Z(n3965) );
  XOR U3982 ( .A(p_input[12]), .B(n4024), .Z(n4023) );
  XOR U3983 ( .A(p_input[13]), .B(p_input[525]), .Z(n3969) );
  XOR U3984 ( .A(n3979), .B(n4025), .Z(n4022) );
  IV U3985 ( .A(n3970), .Z(n4025) );
  XOR U3986 ( .A(p_input[2]), .B(p_input[514]), .Z(n3970) );
  XNOR U3987 ( .A(n4026), .B(n3986), .Z(n3979) );
  XNOR U3988 ( .A(p_input[16]), .B(n4027), .Z(n3986) );
  XOR U3989 ( .A(n3976), .B(n3985), .Z(n4026) );
  XOR U3990 ( .A(n4028), .B(n3982), .Z(n3985) );
  XOR U3991 ( .A(p_input[14]), .B(p_input[526]), .Z(n3982) );
  XOR U3992 ( .A(p_input[15]), .B(n4029), .Z(n4028) );
  XOR U3993 ( .A(p_input[10]), .B(p_input[522]), .Z(n3976) );
  XNOR U3994 ( .A(n3993), .B(n3991), .Z(n3974) );
  XNOR U3995 ( .A(n4030), .B(n3998), .Z(n3991) );
  XOR U3996 ( .A(p_input[521]), .B(p_input[9]), .Z(n3998) );
  XOR U3997 ( .A(n3988), .B(n3997), .Z(n4030) );
  XOR U3998 ( .A(n4031), .B(n3994), .Z(n3997) );
  XOR U3999 ( .A(p_input[519]), .B(p_input[7]), .Z(n3994) );
  XNOR U4000 ( .A(p_input[520]), .B(p_input[8]), .Z(n4031) );
  XOR U4001 ( .A(p_input[3]), .B(p_input[515]), .Z(n3988) );
  XNOR U4002 ( .A(n4003), .B(n4002), .Z(n3993) );
  XOR U4003 ( .A(n4032), .B(n3999), .Z(n4002) );
  XOR U4004 ( .A(p_input[4]), .B(p_input[516]), .Z(n3999) );
  XNOR U4005 ( .A(p_input[517]), .B(p_input[5]), .Z(n4032) );
  XOR U4006 ( .A(p_input[518]), .B(p_input[6]), .Z(n4003) );
  XNOR U4007 ( .A(n4033), .B(n4034), .Z(n3813) );
  AND U4008 ( .A(n66), .B(n4035), .Z(n4034) );
  XNOR U4009 ( .A(n4036), .B(n4037), .Z(n66) );
  AND U4010 ( .A(n4038), .B(n4039), .Z(n4037) );
  XOR U4011 ( .A(n4036), .B(n3823), .Z(n4039) );
  XNOR U4012 ( .A(n4036), .B(n3756), .Z(n4038) );
  XOR U4013 ( .A(n4040), .B(n4041), .Z(n4036) );
  AND U4014 ( .A(n4042), .B(n4043), .Z(n4041) );
  XNOR U4015 ( .A(n3836), .B(n4040), .Z(n4043) );
  XOR U4016 ( .A(n4040), .B(n3838), .Z(n4042) );
  XOR U4017 ( .A(n4044), .B(n4045), .Z(n4040) );
  AND U4018 ( .A(n4046), .B(n4047), .Z(n4045) );
  XNOR U4019 ( .A(n3862), .B(n4044), .Z(n4047) );
  XOR U4020 ( .A(n4044), .B(n3864), .Z(n4046) );
  IV U4021 ( .A(n3782), .Z(n3864) );
  XOR U4022 ( .A(n4048), .B(n4049), .Z(n4044) );
  AND U4023 ( .A(n4050), .B(n4051), .Z(n4049) );
  XOR U4024 ( .A(n4048), .B(n3911), .Z(n4050) );
  XOR U4025 ( .A(n4052), .B(n4053), .Z(n3811) );
  AND U4026 ( .A(n70), .B(n4035), .Z(n4053) );
  XNOR U4027 ( .A(n4033), .B(n4052), .Z(n4035) );
  XNOR U4028 ( .A(n4054), .B(n4055), .Z(n70) );
  AND U4029 ( .A(n4056), .B(n4057), .Z(n4055) );
  XNOR U4030 ( .A(n4058), .B(n4054), .Z(n4057) );
  IV U4031 ( .A(n3823), .Z(n4058) );
  XNOR U4032 ( .A(n4059), .B(n4060), .Z(n3823) );
  AND U4033 ( .A(n74), .B(n4061), .Z(n4060) );
  XNOR U4034 ( .A(n4059), .B(n4062), .Z(n4061) );
  XNOR U4035 ( .A(n3756), .B(n4054), .Z(n4056) );
  XOR U4036 ( .A(n4063), .B(n4064), .Z(n3756) );
  AND U4037 ( .A(n82), .B(n4065), .Z(n4064) );
  XOR U4038 ( .A(n4066), .B(n4067), .Z(n4054) );
  AND U4039 ( .A(n4068), .B(n4069), .Z(n4067) );
  XNOR U4040 ( .A(n4066), .B(n3836), .Z(n4069) );
  XNOR U4041 ( .A(n4070), .B(n4071), .Z(n3836) );
  AND U4042 ( .A(n74), .B(n4072), .Z(n4071) );
  XOR U4043 ( .A(n4073), .B(n4070), .Z(n4072) );
  XNOR U4044 ( .A(n3769), .B(n4066), .Z(n4068) );
  IV U4045 ( .A(n3838), .Z(n3769) );
  XOR U4046 ( .A(n4074), .B(n4075), .Z(n3838) );
  AND U4047 ( .A(n82), .B(n4076), .Z(n4075) );
  XOR U4048 ( .A(n4077), .B(n4078), .Z(n4066) );
  AND U4049 ( .A(n4079), .B(n4080), .Z(n4078) );
  XNOR U4050 ( .A(n4077), .B(n3862), .Z(n4080) );
  XNOR U4051 ( .A(n4081), .B(n4082), .Z(n3862) );
  AND U4052 ( .A(n74), .B(n4083), .Z(n4082) );
  XNOR U4053 ( .A(n4084), .B(n4081), .Z(n4083) );
  XNOR U4054 ( .A(n3782), .B(n4077), .Z(n4079) );
  XNOR U4055 ( .A(n4085), .B(n4086), .Z(n3782) );
  AND U4056 ( .A(n82), .B(n4087), .Z(n4086) );
  XOR U4057 ( .A(n4048), .B(n4088), .Z(n4077) );
  AND U4058 ( .A(n4089), .B(n4051), .Z(n4088) );
  XNOR U4059 ( .A(n3909), .B(n4048), .Z(n4051) );
  XNOR U4060 ( .A(n4090), .B(n4091), .Z(n3909) );
  AND U4061 ( .A(n74), .B(n4092), .Z(n4091) );
  XOR U4062 ( .A(n4093), .B(n4090), .Z(n4092) );
  XNOR U4063 ( .A(n3795), .B(n4048), .Z(n4089) );
  IV U4064 ( .A(n3911), .Z(n3795) );
  XOR U4065 ( .A(n4094), .B(n4095), .Z(n3911) );
  AND U4066 ( .A(n82), .B(n4096), .Z(n4095) );
  XOR U4067 ( .A(n4097), .B(n4098), .Z(n4048) );
  AND U4068 ( .A(n4099), .B(n4100), .Z(n4098) );
  XNOR U4069 ( .A(n4097), .B(n4004), .Z(n4100) );
  XNOR U4070 ( .A(n4101), .B(n4102), .Z(n4004) );
  AND U4071 ( .A(n74), .B(n4103), .Z(n4102) );
  XNOR U4072 ( .A(n4104), .B(n4101), .Z(n4103) );
  XNOR U4073 ( .A(n4105), .B(n4097), .Z(n4099) );
  IV U4074 ( .A(n3808), .Z(n4105) );
  XOR U4075 ( .A(n4106), .B(n4107), .Z(n3808) );
  AND U4076 ( .A(n82), .B(n4108), .Z(n4107) );
  AND U4077 ( .A(n4052), .B(n4033), .Z(n4097) );
  XNOR U4078 ( .A(n4109), .B(n4110), .Z(n4033) );
  AND U4079 ( .A(n74), .B(n4111), .Z(n4110) );
  XNOR U4080 ( .A(n4112), .B(n4109), .Z(n4111) );
  XNOR U4081 ( .A(n4113), .B(n4114), .Z(n74) );
  AND U4082 ( .A(n4115), .B(n4116), .Z(n4114) );
  XOR U4083 ( .A(n4062), .B(n4113), .Z(n4116) );
  AND U4084 ( .A(n4117), .B(n4118), .Z(n4062) );
  XOR U4085 ( .A(n4113), .B(n4059), .Z(n4115) );
  XNOR U4086 ( .A(n4119), .B(n4120), .Z(n4059) );
  AND U4087 ( .A(n78), .B(n4065), .Z(n4120) );
  XOR U4088 ( .A(n4063), .B(n4119), .Z(n4065) );
  XOR U4089 ( .A(n4121), .B(n4122), .Z(n4113) );
  AND U4090 ( .A(n4123), .B(n4124), .Z(n4122) );
  XNOR U4091 ( .A(n4121), .B(n4117), .Z(n4124) );
  IV U4092 ( .A(n4073), .Z(n4117) );
  XOR U4093 ( .A(n4125), .B(n4126), .Z(n4073) );
  XOR U4094 ( .A(n4127), .B(n4118), .Z(n4126) );
  AND U4095 ( .A(n4084), .B(n4128), .Z(n4118) );
  AND U4096 ( .A(n4129), .B(n4130), .Z(n4127) );
  XOR U4097 ( .A(n4131), .B(n4125), .Z(n4129) );
  XNOR U4098 ( .A(n4070), .B(n4121), .Z(n4123) );
  XNOR U4099 ( .A(n4132), .B(n4133), .Z(n4070) );
  AND U4100 ( .A(n78), .B(n4076), .Z(n4133) );
  XOR U4101 ( .A(n4132), .B(n4074), .Z(n4076) );
  XOR U4102 ( .A(n4134), .B(n4135), .Z(n4121) );
  AND U4103 ( .A(n4136), .B(n4137), .Z(n4135) );
  XNOR U4104 ( .A(n4134), .B(n4084), .Z(n4137) );
  XOR U4105 ( .A(n4138), .B(n4130), .Z(n4084) );
  XNOR U4106 ( .A(n4139), .B(n4125), .Z(n4130) );
  XOR U4107 ( .A(n4140), .B(n4141), .Z(n4125) );
  AND U4108 ( .A(n4142), .B(n4143), .Z(n4141) );
  XOR U4109 ( .A(n4144), .B(n4140), .Z(n4142) );
  XNOR U4110 ( .A(n4145), .B(n4146), .Z(n4139) );
  AND U4111 ( .A(n4147), .B(n4148), .Z(n4146) );
  XOR U4112 ( .A(n4145), .B(n4149), .Z(n4147) );
  XNOR U4113 ( .A(n4131), .B(n4128), .Z(n4138) );
  AND U4114 ( .A(n4150), .B(n4151), .Z(n4128) );
  XOR U4115 ( .A(n4152), .B(n4153), .Z(n4131) );
  AND U4116 ( .A(n4154), .B(n4155), .Z(n4153) );
  XOR U4117 ( .A(n4152), .B(n4156), .Z(n4154) );
  XNOR U4118 ( .A(n4081), .B(n4134), .Z(n4136) );
  XNOR U4119 ( .A(n4157), .B(n4158), .Z(n4081) );
  AND U4120 ( .A(n78), .B(n4087), .Z(n4158) );
  XOR U4121 ( .A(n4157), .B(n4085), .Z(n4087) );
  XOR U4122 ( .A(n4159), .B(n4160), .Z(n4134) );
  AND U4123 ( .A(n4161), .B(n4162), .Z(n4160) );
  XNOR U4124 ( .A(n4159), .B(n4150), .Z(n4162) );
  IV U4125 ( .A(n4093), .Z(n4150) );
  XNOR U4126 ( .A(n4163), .B(n4143), .Z(n4093) );
  XNOR U4127 ( .A(n4164), .B(n4149), .Z(n4143) );
  XOR U4128 ( .A(n4165), .B(n4166), .Z(n4149) );
  AND U4129 ( .A(n4167), .B(n4168), .Z(n4166) );
  XOR U4130 ( .A(n4165), .B(n4169), .Z(n4167) );
  XNOR U4131 ( .A(n4148), .B(n4140), .Z(n4164) );
  XOR U4132 ( .A(n4170), .B(n4171), .Z(n4140) );
  AND U4133 ( .A(n4172), .B(n4173), .Z(n4171) );
  XNOR U4134 ( .A(n4174), .B(n4170), .Z(n4172) );
  XNOR U4135 ( .A(n4175), .B(n4145), .Z(n4148) );
  XOR U4136 ( .A(n4176), .B(n4177), .Z(n4145) );
  AND U4137 ( .A(n4178), .B(n4179), .Z(n4177) );
  XOR U4138 ( .A(n4176), .B(n4180), .Z(n4178) );
  XNOR U4139 ( .A(n4181), .B(n4182), .Z(n4175) );
  AND U4140 ( .A(n4183), .B(n4184), .Z(n4182) );
  XNOR U4141 ( .A(n4181), .B(n4185), .Z(n4183) );
  XNOR U4142 ( .A(n4144), .B(n4151), .Z(n4163) );
  AND U4143 ( .A(n4104), .B(n4186), .Z(n4151) );
  XOR U4144 ( .A(n4156), .B(n4155), .Z(n4144) );
  XNOR U4145 ( .A(n4187), .B(n4152), .Z(n4155) );
  XOR U4146 ( .A(n4188), .B(n4189), .Z(n4152) );
  AND U4147 ( .A(n4190), .B(n4191), .Z(n4189) );
  XOR U4148 ( .A(n4188), .B(n4192), .Z(n4190) );
  XNOR U4149 ( .A(n4193), .B(n4194), .Z(n4187) );
  AND U4150 ( .A(n4195), .B(n4196), .Z(n4194) );
  XOR U4151 ( .A(n4193), .B(n4197), .Z(n4195) );
  XOR U4152 ( .A(n4198), .B(n4199), .Z(n4156) );
  AND U4153 ( .A(n4200), .B(n4201), .Z(n4199) );
  XOR U4154 ( .A(n4198), .B(n4202), .Z(n4200) );
  XNOR U4155 ( .A(n4090), .B(n4159), .Z(n4161) );
  XNOR U4156 ( .A(n4203), .B(n4204), .Z(n4090) );
  AND U4157 ( .A(n78), .B(n4096), .Z(n4204) );
  XOR U4158 ( .A(n4203), .B(n4094), .Z(n4096) );
  XOR U4159 ( .A(n4205), .B(n4206), .Z(n4159) );
  AND U4160 ( .A(n4207), .B(n4208), .Z(n4206) );
  XNOR U4161 ( .A(n4205), .B(n4104), .Z(n4208) );
  XOR U4162 ( .A(n4209), .B(n4173), .Z(n4104) );
  XNOR U4163 ( .A(n4210), .B(n4180), .Z(n4173) );
  XOR U4164 ( .A(n4169), .B(n4168), .Z(n4180) );
  XNOR U4165 ( .A(n4211), .B(n4165), .Z(n4168) );
  XOR U4166 ( .A(n4212), .B(n4213), .Z(n4165) );
  AND U4167 ( .A(n4214), .B(n4215), .Z(n4213) );
  XNOR U4168 ( .A(n4216), .B(n4217), .Z(n4214) );
  IV U4169 ( .A(n4212), .Z(n4216) );
  XNOR U4170 ( .A(n4218), .B(n4219), .Z(n4211) );
  NOR U4171 ( .A(n4220), .B(n4221), .Z(n4219) );
  XNOR U4172 ( .A(n4218), .B(n4222), .Z(n4220) );
  XOR U4173 ( .A(n4223), .B(n4224), .Z(n4169) );
  NOR U4174 ( .A(n4225), .B(n4226), .Z(n4224) );
  XNOR U4175 ( .A(n4223), .B(n4227), .Z(n4225) );
  XNOR U4176 ( .A(n4179), .B(n4170), .Z(n4210) );
  XOR U4177 ( .A(n4228), .B(n4229), .Z(n4170) );
  NOR U4178 ( .A(n4230), .B(n4231), .Z(n4229) );
  XOR U4179 ( .A(n4232), .B(n4233), .Z(n4230) );
  XOR U4180 ( .A(n4234), .B(n4185), .Z(n4179) );
  XNOR U4181 ( .A(n4235), .B(n4236), .Z(n4185) );
  NOR U4182 ( .A(n4237), .B(n4238), .Z(n4236) );
  XNOR U4183 ( .A(n4235), .B(n4239), .Z(n4237) );
  XNOR U4184 ( .A(n4184), .B(n4176), .Z(n4234) );
  XOR U4185 ( .A(n4240), .B(n4241), .Z(n4176) );
  AND U4186 ( .A(n4242), .B(n4243), .Z(n4241) );
  XOR U4187 ( .A(n4240), .B(n4244), .Z(n4242) );
  XNOR U4188 ( .A(n4245), .B(n4181), .Z(n4184) );
  XOR U4189 ( .A(n4246), .B(n4247), .Z(n4181) );
  AND U4190 ( .A(n4248), .B(n4249), .Z(n4247) );
  XOR U4191 ( .A(n4246), .B(n4250), .Z(n4248) );
  XNOR U4192 ( .A(n4251), .B(n4252), .Z(n4245) );
  NOR U4193 ( .A(n4253), .B(n4254), .Z(n4252) );
  XOR U4194 ( .A(n4251), .B(n4255), .Z(n4253) );
  XOR U4195 ( .A(n4174), .B(n4186), .Z(n4209) );
  NOR U4196 ( .A(n4112), .B(n4256), .Z(n4186) );
  XNOR U4197 ( .A(n4192), .B(n4191), .Z(n4174) );
  XNOR U4198 ( .A(n4257), .B(n4197), .Z(n4191) );
  XNOR U4199 ( .A(n4258), .B(n4259), .Z(n4197) );
  NOR U4200 ( .A(n4260), .B(n4261), .Z(n4259) );
  XOR U4201 ( .A(n4258), .B(n4262), .Z(n4260) );
  XNOR U4202 ( .A(n4196), .B(n4188), .Z(n4257) );
  XOR U4203 ( .A(n4263), .B(n4264), .Z(n4188) );
  AND U4204 ( .A(n4265), .B(n4266), .Z(n4264) );
  XOR U4205 ( .A(n4263), .B(n4267), .Z(n4265) );
  XNOR U4206 ( .A(n4268), .B(n4193), .Z(n4196) );
  XOR U4207 ( .A(n4269), .B(n4270), .Z(n4193) );
  AND U4208 ( .A(n4271), .B(n4272), .Z(n4270) );
  XNOR U4209 ( .A(n4273), .B(n4274), .Z(n4271) );
  IV U4210 ( .A(n4269), .Z(n4273) );
  XNOR U4211 ( .A(n4275), .B(n4276), .Z(n4268) );
  NOR U4212 ( .A(n4277), .B(n4278), .Z(n4276) );
  XNOR U4213 ( .A(n4275), .B(n4279), .Z(n4277) );
  XOR U4214 ( .A(n4202), .B(n4201), .Z(n4192) );
  XNOR U4215 ( .A(n4280), .B(n4198), .Z(n4201) );
  XOR U4216 ( .A(n4281), .B(n4282), .Z(n4198) );
  AND U4217 ( .A(n4283), .B(n4284), .Z(n4282) );
  XNOR U4218 ( .A(n4285), .B(n4286), .Z(n4283) );
  IV U4219 ( .A(n4281), .Z(n4285) );
  XNOR U4220 ( .A(n4287), .B(n4288), .Z(n4280) );
  NOR U4221 ( .A(n4289), .B(n4290), .Z(n4288) );
  XNOR U4222 ( .A(n4287), .B(n4291), .Z(n4289) );
  XOR U4223 ( .A(n4292), .B(n4293), .Z(n4202) );
  NOR U4224 ( .A(n4294), .B(n4295), .Z(n4293) );
  XNOR U4225 ( .A(n4292), .B(n4296), .Z(n4294) );
  XNOR U4226 ( .A(n4101), .B(n4205), .Z(n4207) );
  XNOR U4227 ( .A(n4297), .B(n4298), .Z(n4101) );
  AND U4228 ( .A(n78), .B(n4108), .Z(n4298) );
  XOR U4229 ( .A(n4297), .B(n4106), .Z(n4108) );
  AND U4230 ( .A(n4109), .B(n4112), .Z(n4205) );
  XOR U4231 ( .A(n4299), .B(n4256), .Z(n4112) );
  XNOR U4232 ( .A(p_input[32]), .B(p_input[512]), .Z(n4256) );
  XOR U4233 ( .A(n4233), .B(n4231), .Z(n4299) );
  XOR U4234 ( .A(n4300), .B(n4244), .Z(n4231) );
  XOR U4235 ( .A(n4217), .B(n4215), .Z(n4244) );
  XNOR U4236 ( .A(n4301), .B(n4222), .Z(n4215) );
  XOR U4237 ( .A(p_input[536]), .B(p_input[56]), .Z(n4222) );
  XOR U4238 ( .A(n4212), .B(n4221), .Z(n4301) );
  XOR U4239 ( .A(n4302), .B(n4218), .Z(n4221) );
  XOR U4240 ( .A(p_input[534]), .B(p_input[54]), .Z(n4218) );
  XNOR U4241 ( .A(p_input[535]), .B(p_input[55]), .Z(n4302) );
  XOR U4242 ( .A(p_input[50]), .B(p_input[530]), .Z(n4212) );
  XNOR U4243 ( .A(n4227), .B(n4226), .Z(n4217) );
  XOR U4244 ( .A(n4303), .B(n4223), .Z(n4226) );
  XOR U4245 ( .A(p_input[51]), .B(p_input[531]), .Z(n4223) );
  XOR U4246 ( .A(p_input[52]), .B(n4012), .Z(n4303) );
  XOR U4247 ( .A(p_input[533]), .B(p_input[53]), .Z(n4227) );
  XOR U4248 ( .A(n4243), .B(n4232), .Z(n4300) );
  IV U4249 ( .A(n4228), .Z(n4232) );
  XOR U4250 ( .A(p_input[33]), .B(p_input[513]), .Z(n4228) );
  XNOR U4251 ( .A(n4304), .B(n4250), .Z(n4243) );
  XNOR U4252 ( .A(n4239), .B(n4238), .Z(n4250) );
  XOR U4253 ( .A(n4305), .B(n4235), .Z(n4238) );
  XNOR U4254 ( .A(n4306), .B(p_input[58]), .Z(n4235) );
  XNOR U4255 ( .A(p_input[539]), .B(p_input[59]), .Z(n4305) );
  XOR U4256 ( .A(p_input[540]), .B(p_input[60]), .Z(n4239) );
  XOR U4257 ( .A(n4249), .B(n4307), .Z(n4304) );
  IV U4258 ( .A(n4240), .Z(n4307) );
  XOR U4259 ( .A(p_input[49]), .B(p_input[529]), .Z(n4240) );
  XOR U4260 ( .A(n4308), .B(n4255), .Z(n4249) );
  XNOR U4261 ( .A(p_input[543]), .B(p_input[63]), .Z(n4255) );
  XOR U4262 ( .A(n4246), .B(n4254), .Z(n4308) );
  XOR U4263 ( .A(n4309), .B(n4251), .Z(n4254) );
  XOR U4264 ( .A(p_input[541]), .B(p_input[61]), .Z(n4251) );
  XNOR U4265 ( .A(p_input[542]), .B(p_input[62]), .Z(n4309) );
  XNOR U4266 ( .A(n4310), .B(p_input[57]), .Z(n4246) );
  XOR U4267 ( .A(n4267), .B(n4266), .Z(n4233) );
  XNOR U4268 ( .A(n4311), .B(n4274), .Z(n4266) );
  XNOR U4269 ( .A(n4262), .B(n4261), .Z(n4274) );
  XNOR U4270 ( .A(n4312), .B(n4258), .Z(n4261) );
  XNOR U4271 ( .A(p_input[43]), .B(p_input[523]), .Z(n4258) );
  XOR U4272 ( .A(p_input[44]), .B(n4024), .Z(n4312) );
  XOR U4273 ( .A(p_input[45]), .B(p_input[525]), .Z(n4262) );
  XOR U4274 ( .A(n4272), .B(n4313), .Z(n4311) );
  IV U4275 ( .A(n4263), .Z(n4313) );
  XOR U4276 ( .A(p_input[34]), .B(p_input[514]), .Z(n4263) );
  XNOR U4277 ( .A(n4314), .B(n4279), .Z(n4272) );
  XNOR U4278 ( .A(p_input[48]), .B(n4027), .Z(n4279) );
  XOR U4279 ( .A(n4269), .B(n4278), .Z(n4314) );
  XOR U4280 ( .A(n4315), .B(n4275), .Z(n4278) );
  XOR U4281 ( .A(p_input[46]), .B(p_input[526]), .Z(n4275) );
  XOR U4282 ( .A(p_input[47]), .B(n4029), .Z(n4315) );
  XOR U4283 ( .A(p_input[42]), .B(p_input[522]), .Z(n4269) );
  XOR U4284 ( .A(n4286), .B(n4284), .Z(n4267) );
  XNOR U4285 ( .A(n4316), .B(n4291), .Z(n4284) );
  XOR U4286 ( .A(p_input[41]), .B(p_input[521]), .Z(n4291) );
  XOR U4287 ( .A(n4281), .B(n4290), .Z(n4316) );
  XOR U4288 ( .A(n4317), .B(n4287), .Z(n4290) );
  XOR U4289 ( .A(p_input[39]), .B(p_input[519]), .Z(n4287) );
  XOR U4290 ( .A(p_input[40]), .B(n4318), .Z(n4317) );
  XOR U4291 ( .A(p_input[35]), .B(p_input[515]), .Z(n4281) );
  XNOR U4292 ( .A(n4296), .B(n4295), .Z(n4286) );
  XOR U4293 ( .A(n4319), .B(n4292), .Z(n4295) );
  XOR U4294 ( .A(p_input[36]), .B(p_input[516]), .Z(n4292) );
  XOR U4295 ( .A(p_input[37]), .B(n4320), .Z(n4319) );
  XOR U4296 ( .A(p_input[38]), .B(p_input[518]), .Z(n4296) );
  XNOR U4297 ( .A(n4321), .B(n4322), .Z(n4109) );
  AND U4298 ( .A(n78), .B(n4323), .Z(n4322) );
  XNOR U4299 ( .A(n4324), .B(n4325), .Z(n78) );
  AND U4300 ( .A(n4326), .B(n4327), .Z(n4325) );
  XOR U4301 ( .A(n4324), .B(n4119), .Z(n4327) );
  XNOR U4302 ( .A(n4324), .B(n4063), .Z(n4326) );
  XOR U4303 ( .A(n4328), .B(n4329), .Z(n4324) );
  AND U4304 ( .A(n4330), .B(n4331), .Z(n4329) );
  XNOR U4305 ( .A(n4132), .B(n4328), .Z(n4331) );
  XOR U4306 ( .A(n4328), .B(n4074), .Z(n4330) );
  XOR U4307 ( .A(n4332), .B(n4333), .Z(n4328) );
  AND U4308 ( .A(n4334), .B(n4335), .Z(n4333) );
  XNOR U4309 ( .A(n4157), .B(n4332), .Z(n4335) );
  XOR U4310 ( .A(n4332), .B(n4085), .Z(n4334) );
  XOR U4311 ( .A(n4336), .B(n4337), .Z(n4332) );
  AND U4312 ( .A(n4338), .B(n4339), .Z(n4337) );
  XOR U4313 ( .A(n4336), .B(n4094), .Z(n4338) );
  XOR U4314 ( .A(n4340), .B(n4341), .Z(n4052) );
  AND U4315 ( .A(n82), .B(n4323), .Z(n4341) );
  XNOR U4316 ( .A(n4321), .B(n4340), .Z(n4323) );
  XNOR U4317 ( .A(n4342), .B(n4343), .Z(n82) );
  AND U4318 ( .A(n4344), .B(n4345), .Z(n4343) );
  XNOR U4319 ( .A(n4346), .B(n4342), .Z(n4345) );
  IV U4320 ( .A(n4119), .Z(n4346) );
  XNOR U4321 ( .A(n4347), .B(n4348), .Z(n4119) );
  AND U4322 ( .A(n85), .B(n4349), .Z(n4348) );
  XNOR U4323 ( .A(n4347), .B(n4350), .Z(n4349) );
  XNOR U4324 ( .A(n4063), .B(n4342), .Z(n4344) );
  XOR U4325 ( .A(n4351), .B(n4352), .Z(n4063) );
  AND U4326 ( .A(n93), .B(n4353), .Z(n4352) );
  XOR U4327 ( .A(n4354), .B(n4355), .Z(n4342) );
  AND U4328 ( .A(n4356), .B(n4357), .Z(n4355) );
  XNOR U4329 ( .A(n4354), .B(n4132), .Z(n4357) );
  XNOR U4330 ( .A(n4358), .B(n4359), .Z(n4132) );
  AND U4331 ( .A(n85), .B(n4360), .Z(n4359) );
  XOR U4332 ( .A(n4361), .B(n4358), .Z(n4360) );
  XNOR U4333 ( .A(n4362), .B(n4354), .Z(n4356) );
  IV U4334 ( .A(n4074), .Z(n4362) );
  XOR U4335 ( .A(n4363), .B(n4364), .Z(n4074) );
  AND U4336 ( .A(n93), .B(n4365), .Z(n4364) );
  XOR U4337 ( .A(n4366), .B(n4367), .Z(n4354) );
  AND U4338 ( .A(n4368), .B(n4369), .Z(n4367) );
  XNOR U4339 ( .A(n4366), .B(n4157), .Z(n4369) );
  XNOR U4340 ( .A(n4370), .B(n4371), .Z(n4157) );
  AND U4341 ( .A(n85), .B(n4372), .Z(n4371) );
  XNOR U4342 ( .A(n4373), .B(n4370), .Z(n4372) );
  XOR U4343 ( .A(n4085), .B(n4366), .Z(n4368) );
  XOR U4344 ( .A(n4374), .B(n4375), .Z(n4085) );
  AND U4345 ( .A(n93), .B(n4376), .Z(n4375) );
  XOR U4346 ( .A(n4336), .B(n4377), .Z(n4366) );
  AND U4347 ( .A(n4378), .B(n4339), .Z(n4377) );
  XNOR U4348 ( .A(n4203), .B(n4336), .Z(n4339) );
  XNOR U4349 ( .A(n4379), .B(n4380), .Z(n4203) );
  AND U4350 ( .A(n85), .B(n4381), .Z(n4380) );
  XOR U4351 ( .A(n4382), .B(n4379), .Z(n4381) );
  XNOR U4352 ( .A(n4383), .B(n4336), .Z(n4378) );
  IV U4353 ( .A(n4094), .Z(n4383) );
  XOR U4354 ( .A(n4384), .B(n4385), .Z(n4094) );
  AND U4355 ( .A(n93), .B(n4386), .Z(n4385) );
  XOR U4356 ( .A(n4387), .B(n4388), .Z(n4336) );
  AND U4357 ( .A(n4389), .B(n4390), .Z(n4388) );
  XNOR U4358 ( .A(n4387), .B(n4297), .Z(n4390) );
  XNOR U4359 ( .A(n4391), .B(n4392), .Z(n4297) );
  AND U4360 ( .A(n85), .B(n4393), .Z(n4392) );
  XNOR U4361 ( .A(n4394), .B(n4391), .Z(n4393) );
  XNOR U4362 ( .A(n4395), .B(n4387), .Z(n4389) );
  IV U4363 ( .A(n4106), .Z(n4395) );
  XOR U4364 ( .A(n4396), .B(n4397), .Z(n4106) );
  AND U4365 ( .A(n93), .B(n4398), .Z(n4397) );
  AND U4366 ( .A(n4340), .B(n4321), .Z(n4387) );
  XNOR U4367 ( .A(n4399), .B(n4400), .Z(n4321) );
  AND U4368 ( .A(n85), .B(n4401), .Z(n4400) );
  XNOR U4369 ( .A(n4402), .B(n4399), .Z(n4401) );
  XNOR U4370 ( .A(n4403), .B(n4404), .Z(n85) );
  AND U4371 ( .A(n4405), .B(n4406), .Z(n4404) );
  XOR U4372 ( .A(n4350), .B(n4403), .Z(n4406) );
  AND U4373 ( .A(n4407), .B(n4408), .Z(n4350) );
  XOR U4374 ( .A(n4403), .B(n4347), .Z(n4405) );
  XNOR U4375 ( .A(n4409), .B(n4410), .Z(n4347) );
  AND U4376 ( .A(n89), .B(n4353), .Z(n4410) );
  XOR U4377 ( .A(n4351), .B(n4409), .Z(n4353) );
  XOR U4378 ( .A(n4411), .B(n4412), .Z(n4403) );
  AND U4379 ( .A(n4413), .B(n4414), .Z(n4412) );
  XNOR U4380 ( .A(n4411), .B(n4407), .Z(n4414) );
  IV U4381 ( .A(n4361), .Z(n4407) );
  XOR U4382 ( .A(n4415), .B(n4416), .Z(n4361) );
  XOR U4383 ( .A(n4417), .B(n4408), .Z(n4416) );
  AND U4384 ( .A(n4373), .B(n4418), .Z(n4408) );
  AND U4385 ( .A(n4419), .B(n4420), .Z(n4417) );
  XOR U4386 ( .A(n4421), .B(n4415), .Z(n4419) );
  XNOR U4387 ( .A(n4358), .B(n4411), .Z(n4413) );
  XNOR U4388 ( .A(n4422), .B(n4423), .Z(n4358) );
  AND U4389 ( .A(n89), .B(n4365), .Z(n4423) );
  XOR U4390 ( .A(n4422), .B(n4363), .Z(n4365) );
  XOR U4391 ( .A(n4424), .B(n4425), .Z(n4411) );
  AND U4392 ( .A(n4426), .B(n4427), .Z(n4425) );
  XNOR U4393 ( .A(n4424), .B(n4373), .Z(n4427) );
  XOR U4394 ( .A(n4428), .B(n4420), .Z(n4373) );
  XNOR U4395 ( .A(n4429), .B(n4415), .Z(n4420) );
  XOR U4396 ( .A(n4430), .B(n4431), .Z(n4415) );
  AND U4397 ( .A(n4432), .B(n4433), .Z(n4431) );
  XOR U4398 ( .A(n4434), .B(n4430), .Z(n4432) );
  XNOR U4399 ( .A(n4435), .B(n4436), .Z(n4429) );
  AND U4400 ( .A(n4437), .B(n4438), .Z(n4436) );
  XOR U4401 ( .A(n4435), .B(n4439), .Z(n4437) );
  XNOR U4402 ( .A(n4421), .B(n4418), .Z(n4428) );
  AND U4403 ( .A(n4440), .B(n4441), .Z(n4418) );
  XOR U4404 ( .A(n4442), .B(n4443), .Z(n4421) );
  AND U4405 ( .A(n4444), .B(n4445), .Z(n4443) );
  XOR U4406 ( .A(n4442), .B(n4446), .Z(n4444) );
  XNOR U4407 ( .A(n4370), .B(n4424), .Z(n4426) );
  XNOR U4408 ( .A(n4447), .B(n4448), .Z(n4370) );
  AND U4409 ( .A(n89), .B(n4376), .Z(n4448) );
  XOR U4410 ( .A(n4447), .B(n4374), .Z(n4376) );
  XOR U4411 ( .A(n4449), .B(n4450), .Z(n4424) );
  AND U4412 ( .A(n4451), .B(n4452), .Z(n4450) );
  XNOR U4413 ( .A(n4449), .B(n4440), .Z(n4452) );
  IV U4414 ( .A(n4382), .Z(n4440) );
  XNOR U4415 ( .A(n4453), .B(n4433), .Z(n4382) );
  XNOR U4416 ( .A(n4454), .B(n4439), .Z(n4433) );
  XOR U4417 ( .A(n4455), .B(n4456), .Z(n4439) );
  AND U4418 ( .A(n4457), .B(n4458), .Z(n4456) );
  XOR U4419 ( .A(n4455), .B(n4459), .Z(n4457) );
  XNOR U4420 ( .A(n4438), .B(n4430), .Z(n4454) );
  XOR U4421 ( .A(n4460), .B(n4461), .Z(n4430) );
  AND U4422 ( .A(n4462), .B(n4463), .Z(n4461) );
  XNOR U4423 ( .A(n4464), .B(n4460), .Z(n4462) );
  XNOR U4424 ( .A(n4465), .B(n4435), .Z(n4438) );
  XOR U4425 ( .A(n4466), .B(n4467), .Z(n4435) );
  AND U4426 ( .A(n4468), .B(n4469), .Z(n4467) );
  XOR U4427 ( .A(n4466), .B(n4470), .Z(n4468) );
  XNOR U4428 ( .A(n4471), .B(n4472), .Z(n4465) );
  AND U4429 ( .A(n4473), .B(n4474), .Z(n4472) );
  XNOR U4430 ( .A(n4471), .B(n4475), .Z(n4473) );
  XNOR U4431 ( .A(n4434), .B(n4441), .Z(n4453) );
  AND U4432 ( .A(n4394), .B(n4476), .Z(n4441) );
  XOR U4433 ( .A(n4446), .B(n4445), .Z(n4434) );
  XNOR U4434 ( .A(n4477), .B(n4442), .Z(n4445) );
  XOR U4435 ( .A(n4478), .B(n4479), .Z(n4442) );
  AND U4436 ( .A(n4480), .B(n4481), .Z(n4479) );
  XOR U4437 ( .A(n4478), .B(n4482), .Z(n4480) );
  XNOR U4438 ( .A(n4483), .B(n4484), .Z(n4477) );
  AND U4439 ( .A(n4485), .B(n4486), .Z(n4484) );
  XOR U4440 ( .A(n4483), .B(n4487), .Z(n4485) );
  XOR U4441 ( .A(n4488), .B(n4489), .Z(n4446) );
  AND U4442 ( .A(n4490), .B(n4491), .Z(n4489) );
  XOR U4443 ( .A(n4488), .B(n4492), .Z(n4490) );
  XNOR U4444 ( .A(n4379), .B(n4449), .Z(n4451) );
  XNOR U4445 ( .A(n4493), .B(n4494), .Z(n4379) );
  AND U4446 ( .A(n89), .B(n4386), .Z(n4494) );
  XOR U4447 ( .A(n4493), .B(n4384), .Z(n4386) );
  XOR U4448 ( .A(n4495), .B(n4496), .Z(n4449) );
  AND U4449 ( .A(n4497), .B(n4498), .Z(n4496) );
  XNOR U4450 ( .A(n4495), .B(n4394), .Z(n4498) );
  XOR U4451 ( .A(n4499), .B(n4463), .Z(n4394) );
  XNOR U4452 ( .A(n4500), .B(n4470), .Z(n4463) );
  XOR U4453 ( .A(n4459), .B(n4458), .Z(n4470) );
  XNOR U4454 ( .A(n4501), .B(n4455), .Z(n4458) );
  XOR U4455 ( .A(n4502), .B(n4503), .Z(n4455) );
  AND U4456 ( .A(n4504), .B(n4505), .Z(n4503) );
  XOR U4457 ( .A(n4502), .B(n4506), .Z(n4504) );
  XNOR U4458 ( .A(n4507), .B(n4508), .Z(n4501) );
  NOR U4459 ( .A(n4509), .B(n4510), .Z(n4508) );
  XNOR U4460 ( .A(n4507), .B(n4511), .Z(n4509) );
  XOR U4461 ( .A(n4512), .B(n4513), .Z(n4459) );
  NOR U4462 ( .A(n4514), .B(n4515), .Z(n4513) );
  XNOR U4463 ( .A(n4512), .B(n4516), .Z(n4514) );
  XNOR U4464 ( .A(n4469), .B(n4460), .Z(n4500) );
  XOR U4465 ( .A(n4517), .B(n4518), .Z(n4460) );
  NOR U4466 ( .A(n4519), .B(n4520), .Z(n4518) );
  XNOR U4467 ( .A(n4517), .B(n4521), .Z(n4519) );
  XOR U4468 ( .A(n4522), .B(n4475), .Z(n4469) );
  XNOR U4469 ( .A(n4523), .B(n4524), .Z(n4475) );
  NOR U4470 ( .A(n4525), .B(n4526), .Z(n4524) );
  XNOR U4471 ( .A(n4523), .B(n4527), .Z(n4525) );
  XNOR U4472 ( .A(n4474), .B(n4466), .Z(n4522) );
  XOR U4473 ( .A(n4528), .B(n4529), .Z(n4466) );
  AND U4474 ( .A(n4530), .B(n4531), .Z(n4529) );
  XOR U4475 ( .A(n4528), .B(n4532), .Z(n4530) );
  XNOR U4476 ( .A(n4533), .B(n4471), .Z(n4474) );
  XOR U4477 ( .A(n4534), .B(n4535), .Z(n4471) );
  AND U4478 ( .A(n4536), .B(n4537), .Z(n4535) );
  XOR U4479 ( .A(n4534), .B(n4538), .Z(n4536) );
  XNOR U4480 ( .A(n4539), .B(n4540), .Z(n4533) );
  NOR U4481 ( .A(n4541), .B(n4542), .Z(n4540) );
  XOR U4482 ( .A(n4539), .B(n4543), .Z(n4541) );
  XOR U4483 ( .A(n4464), .B(n4476), .Z(n4499) );
  NOR U4484 ( .A(n4402), .B(n4544), .Z(n4476) );
  XNOR U4485 ( .A(n4482), .B(n4481), .Z(n4464) );
  XNOR U4486 ( .A(n4545), .B(n4487), .Z(n4481) );
  XOR U4487 ( .A(n4546), .B(n4547), .Z(n4487) );
  NOR U4488 ( .A(n4548), .B(n4549), .Z(n4547) );
  XNOR U4489 ( .A(n4546), .B(n4550), .Z(n4548) );
  XNOR U4490 ( .A(n4486), .B(n4478), .Z(n4545) );
  XOR U4491 ( .A(n4551), .B(n4552), .Z(n4478) );
  AND U4492 ( .A(n4553), .B(n4554), .Z(n4552) );
  XNOR U4493 ( .A(n4551), .B(n4555), .Z(n4553) );
  XNOR U4494 ( .A(n4556), .B(n4483), .Z(n4486) );
  XOR U4495 ( .A(n4557), .B(n4558), .Z(n4483) );
  AND U4496 ( .A(n4559), .B(n4560), .Z(n4558) );
  XOR U4497 ( .A(n4557), .B(n4561), .Z(n4559) );
  XNOR U4498 ( .A(n4562), .B(n4563), .Z(n4556) );
  NOR U4499 ( .A(n4564), .B(n4565), .Z(n4563) );
  XOR U4500 ( .A(n4562), .B(n4566), .Z(n4564) );
  XOR U4501 ( .A(n4492), .B(n4491), .Z(n4482) );
  XNOR U4502 ( .A(n4567), .B(n4488), .Z(n4491) );
  XOR U4503 ( .A(n4568), .B(n4569), .Z(n4488) );
  AND U4504 ( .A(n4570), .B(n4571), .Z(n4569) );
  XOR U4505 ( .A(n4568), .B(n4572), .Z(n4570) );
  XNOR U4506 ( .A(n4573), .B(n4574), .Z(n4567) );
  NOR U4507 ( .A(n4575), .B(n4576), .Z(n4574) );
  XNOR U4508 ( .A(n4573), .B(n4577), .Z(n4575) );
  XOR U4509 ( .A(n4578), .B(n4579), .Z(n4492) );
  NOR U4510 ( .A(n4580), .B(n4581), .Z(n4579) );
  XNOR U4511 ( .A(n4578), .B(n4582), .Z(n4580) );
  XNOR U4512 ( .A(n4391), .B(n4495), .Z(n4497) );
  XNOR U4513 ( .A(n4583), .B(n4584), .Z(n4391) );
  AND U4514 ( .A(n89), .B(n4398), .Z(n4584) );
  XOR U4515 ( .A(n4583), .B(n4396), .Z(n4398) );
  AND U4516 ( .A(n4399), .B(n4402), .Z(n4495) );
  XOR U4517 ( .A(n4585), .B(n4544), .Z(n4402) );
  XNOR U4518 ( .A(p_input[512]), .B(p_input[64]), .Z(n4544) );
  XOR U4519 ( .A(n4521), .B(n4520), .Z(n4585) );
  XOR U4520 ( .A(n4586), .B(n4532), .Z(n4520) );
  XOR U4521 ( .A(n4506), .B(n4505), .Z(n4532) );
  XNOR U4522 ( .A(n4587), .B(n4511), .Z(n4505) );
  XOR U4523 ( .A(p_input[536]), .B(p_input[88]), .Z(n4511) );
  XOR U4524 ( .A(n4502), .B(n4510), .Z(n4587) );
  XOR U4525 ( .A(n4588), .B(n4507), .Z(n4510) );
  XOR U4526 ( .A(p_input[534]), .B(p_input[86]), .Z(n4507) );
  XNOR U4527 ( .A(p_input[535]), .B(p_input[87]), .Z(n4588) );
  XNOR U4528 ( .A(n4589), .B(p_input[82]), .Z(n4502) );
  XNOR U4529 ( .A(n4516), .B(n4515), .Z(n4506) );
  XOR U4530 ( .A(n4590), .B(n4512), .Z(n4515) );
  XOR U4531 ( .A(p_input[531]), .B(p_input[83]), .Z(n4512) );
  XNOR U4532 ( .A(p_input[532]), .B(p_input[84]), .Z(n4590) );
  XOR U4533 ( .A(p_input[533]), .B(p_input[85]), .Z(n4516) );
  XNOR U4534 ( .A(n4531), .B(n4517), .Z(n4586) );
  XNOR U4535 ( .A(n4591), .B(p_input[65]), .Z(n4517) );
  XNOR U4536 ( .A(n4592), .B(n4538), .Z(n4531) );
  XNOR U4537 ( .A(n4527), .B(n4526), .Z(n4538) );
  XOR U4538 ( .A(n4593), .B(n4523), .Z(n4526) );
  XNOR U4539 ( .A(n4306), .B(p_input[90]), .Z(n4523) );
  XNOR U4540 ( .A(p_input[539]), .B(p_input[91]), .Z(n4593) );
  XOR U4541 ( .A(p_input[540]), .B(p_input[92]), .Z(n4527) );
  XNOR U4542 ( .A(n4537), .B(n4528), .Z(n4592) );
  XNOR U4543 ( .A(n4594), .B(p_input[81]), .Z(n4528) );
  XOR U4544 ( .A(n4595), .B(n4543), .Z(n4537) );
  XNOR U4545 ( .A(p_input[543]), .B(p_input[95]), .Z(n4543) );
  XOR U4546 ( .A(n4534), .B(n4542), .Z(n4595) );
  XOR U4547 ( .A(n4596), .B(n4539), .Z(n4542) );
  XOR U4548 ( .A(p_input[541]), .B(p_input[93]), .Z(n4539) );
  XNOR U4549 ( .A(p_input[542]), .B(p_input[94]), .Z(n4596) );
  XNOR U4550 ( .A(n4310), .B(p_input[89]), .Z(n4534) );
  XNOR U4551 ( .A(n4555), .B(n4554), .Z(n4521) );
  XNOR U4552 ( .A(n4597), .B(n4561), .Z(n4554) );
  XNOR U4553 ( .A(n4550), .B(n4549), .Z(n4561) );
  XOR U4554 ( .A(n4598), .B(n4546), .Z(n4549) );
  XNOR U4555 ( .A(n4599), .B(p_input[75]), .Z(n4546) );
  XNOR U4556 ( .A(p_input[524]), .B(p_input[76]), .Z(n4598) );
  XOR U4557 ( .A(p_input[525]), .B(p_input[77]), .Z(n4550) );
  XNOR U4558 ( .A(n4560), .B(n4551), .Z(n4597) );
  XNOR U4559 ( .A(n4600), .B(p_input[66]), .Z(n4551) );
  XOR U4560 ( .A(n4601), .B(n4566), .Z(n4560) );
  XNOR U4561 ( .A(p_input[528]), .B(p_input[80]), .Z(n4566) );
  XOR U4562 ( .A(n4557), .B(n4565), .Z(n4601) );
  XOR U4563 ( .A(n4602), .B(n4562), .Z(n4565) );
  XOR U4564 ( .A(p_input[526]), .B(p_input[78]), .Z(n4562) );
  XNOR U4565 ( .A(p_input[527]), .B(p_input[79]), .Z(n4602) );
  XNOR U4566 ( .A(n4603), .B(p_input[74]), .Z(n4557) );
  XNOR U4567 ( .A(n4572), .B(n4571), .Z(n4555) );
  XNOR U4568 ( .A(n4604), .B(n4577), .Z(n4571) );
  XOR U4569 ( .A(p_input[521]), .B(p_input[73]), .Z(n4577) );
  XOR U4570 ( .A(n4568), .B(n4576), .Z(n4604) );
  XOR U4571 ( .A(n4605), .B(n4573), .Z(n4576) );
  XOR U4572 ( .A(p_input[519]), .B(p_input[71]), .Z(n4573) );
  XNOR U4573 ( .A(p_input[520]), .B(p_input[72]), .Z(n4605) );
  XNOR U4574 ( .A(n4606), .B(p_input[67]), .Z(n4568) );
  XNOR U4575 ( .A(n4582), .B(n4581), .Z(n4572) );
  XOR U4576 ( .A(n4607), .B(n4578), .Z(n4581) );
  XOR U4577 ( .A(p_input[516]), .B(p_input[68]), .Z(n4578) );
  XNOR U4578 ( .A(p_input[517]), .B(p_input[69]), .Z(n4607) );
  XOR U4579 ( .A(p_input[518]), .B(p_input[70]), .Z(n4582) );
  XNOR U4580 ( .A(n4608), .B(n4609), .Z(n4399) );
  AND U4581 ( .A(n89), .B(n4610), .Z(n4609) );
  XNOR U4582 ( .A(n4611), .B(n4612), .Z(n89) );
  AND U4583 ( .A(n4613), .B(n4614), .Z(n4612) );
  XOR U4584 ( .A(n4611), .B(n4409), .Z(n4614) );
  XNOR U4585 ( .A(n4611), .B(n4351), .Z(n4613) );
  XOR U4586 ( .A(n4615), .B(n4616), .Z(n4611) );
  AND U4587 ( .A(n4617), .B(n4618), .Z(n4616) );
  XNOR U4588 ( .A(n4422), .B(n4615), .Z(n4618) );
  XOR U4589 ( .A(n4615), .B(n4363), .Z(n4617) );
  XOR U4590 ( .A(n4619), .B(n4620), .Z(n4615) );
  AND U4591 ( .A(n4621), .B(n4622), .Z(n4620) );
  XNOR U4592 ( .A(n4447), .B(n4619), .Z(n4622) );
  XOR U4593 ( .A(n4619), .B(n4374), .Z(n4621) );
  XOR U4594 ( .A(n4623), .B(n4624), .Z(n4619) );
  AND U4595 ( .A(n4625), .B(n4626), .Z(n4624) );
  XOR U4596 ( .A(n4623), .B(n4384), .Z(n4625) );
  XOR U4597 ( .A(n4627), .B(n4628), .Z(n4340) );
  AND U4598 ( .A(n93), .B(n4610), .Z(n4628) );
  XNOR U4599 ( .A(n4608), .B(n4627), .Z(n4610) );
  XNOR U4600 ( .A(n4629), .B(n4630), .Z(n93) );
  AND U4601 ( .A(n4631), .B(n4632), .Z(n4630) );
  XNOR U4602 ( .A(n4633), .B(n4629), .Z(n4632) );
  IV U4603 ( .A(n4409), .Z(n4633) );
  XNOR U4604 ( .A(n4634), .B(n4635), .Z(n4409) );
  AND U4605 ( .A(n96), .B(n4636), .Z(n4635) );
  XNOR U4606 ( .A(n4634), .B(n4637), .Z(n4636) );
  XNOR U4607 ( .A(n4351), .B(n4629), .Z(n4631) );
  XOR U4608 ( .A(n4638), .B(n4639), .Z(n4351) );
  AND U4609 ( .A(n104), .B(n4640), .Z(n4639) );
  XOR U4610 ( .A(n4641), .B(n4642), .Z(n4629) );
  AND U4611 ( .A(n4643), .B(n4644), .Z(n4642) );
  XNOR U4612 ( .A(n4641), .B(n4422), .Z(n4644) );
  XNOR U4613 ( .A(n4645), .B(n4646), .Z(n4422) );
  AND U4614 ( .A(n96), .B(n4647), .Z(n4646) );
  XOR U4615 ( .A(n4648), .B(n4645), .Z(n4647) );
  XNOR U4616 ( .A(n4649), .B(n4641), .Z(n4643) );
  IV U4617 ( .A(n4363), .Z(n4649) );
  XOR U4618 ( .A(n4650), .B(n4651), .Z(n4363) );
  AND U4619 ( .A(n104), .B(n4652), .Z(n4651) );
  XOR U4620 ( .A(n4653), .B(n4654), .Z(n4641) );
  AND U4621 ( .A(n4655), .B(n4656), .Z(n4654) );
  XNOR U4622 ( .A(n4653), .B(n4447), .Z(n4656) );
  XNOR U4623 ( .A(n4657), .B(n4658), .Z(n4447) );
  AND U4624 ( .A(n96), .B(n4659), .Z(n4658) );
  XNOR U4625 ( .A(n4660), .B(n4657), .Z(n4659) );
  XOR U4626 ( .A(n4374), .B(n4653), .Z(n4655) );
  XOR U4627 ( .A(n4661), .B(n4662), .Z(n4374) );
  AND U4628 ( .A(n104), .B(n4663), .Z(n4662) );
  XOR U4629 ( .A(n4623), .B(n4664), .Z(n4653) );
  AND U4630 ( .A(n4665), .B(n4626), .Z(n4664) );
  XNOR U4631 ( .A(n4493), .B(n4623), .Z(n4626) );
  XNOR U4632 ( .A(n4666), .B(n4667), .Z(n4493) );
  AND U4633 ( .A(n96), .B(n4668), .Z(n4667) );
  XOR U4634 ( .A(n4669), .B(n4666), .Z(n4668) );
  XNOR U4635 ( .A(n4670), .B(n4623), .Z(n4665) );
  IV U4636 ( .A(n4384), .Z(n4670) );
  XOR U4637 ( .A(n4671), .B(n4672), .Z(n4384) );
  AND U4638 ( .A(n104), .B(n4673), .Z(n4672) );
  XOR U4639 ( .A(n4674), .B(n4675), .Z(n4623) );
  AND U4640 ( .A(n4676), .B(n4677), .Z(n4675) );
  XNOR U4641 ( .A(n4674), .B(n4583), .Z(n4677) );
  XNOR U4642 ( .A(n4678), .B(n4679), .Z(n4583) );
  AND U4643 ( .A(n96), .B(n4680), .Z(n4679) );
  XNOR U4644 ( .A(n4681), .B(n4678), .Z(n4680) );
  XNOR U4645 ( .A(n4682), .B(n4674), .Z(n4676) );
  IV U4646 ( .A(n4396), .Z(n4682) );
  XOR U4647 ( .A(n4683), .B(n4684), .Z(n4396) );
  AND U4648 ( .A(n104), .B(n4685), .Z(n4684) );
  AND U4649 ( .A(n4627), .B(n4608), .Z(n4674) );
  XNOR U4650 ( .A(n4686), .B(n4687), .Z(n4608) );
  AND U4651 ( .A(n96), .B(n4688), .Z(n4687) );
  XNOR U4652 ( .A(n4689), .B(n4686), .Z(n4688) );
  XNOR U4653 ( .A(n4690), .B(n4691), .Z(n96) );
  AND U4654 ( .A(n4692), .B(n4693), .Z(n4691) );
  XOR U4655 ( .A(n4637), .B(n4690), .Z(n4693) );
  AND U4656 ( .A(n4694), .B(n4695), .Z(n4637) );
  XOR U4657 ( .A(n4690), .B(n4634), .Z(n4692) );
  XNOR U4658 ( .A(n4696), .B(n4697), .Z(n4634) );
  AND U4659 ( .A(n100), .B(n4640), .Z(n4697) );
  XOR U4660 ( .A(n4638), .B(n4696), .Z(n4640) );
  XOR U4661 ( .A(n4698), .B(n4699), .Z(n4690) );
  AND U4662 ( .A(n4700), .B(n4701), .Z(n4699) );
  XNOR U4663 ( .A(n4698), .B(n4694), .Z(n4701) );
  IV U4664 ( .A(n4648), .Z(n4694) );
  XOR U4665 ( .A(n4702), .B(n4703), .Z(n4648) );
  XOR U4666 ( .A(n4704), .B(n4695), .Z(n4703) );
  AND U4667 ( .A(n4660), .B(n4705), .Z(n4695) );
  AND U4668 ( .A(n4706), .B(n4707), .Z(n4704) );
  XOR U4669 ( .A(n4708), .B(n4702), .Z(n4706) );
  XNOR U4670 ( .A(n4645), .B(n4698), .Z(n4700) );
  XNOR U4671 ( .A(n4709), .B(n4710), .Z(n4645) );
  AND U4672 ( .A(n100), .B(n4652), .Z(n4710) );
  XOR U4673 ( .A(n4709), .B(n4650), .Z(n4652) );
  XOR U4674 ( .A(n4711), .B(n4712), .Z(n4698) );
  AND U4675 ( .A(n4713), .B(n4714), .Z(n4712) );
  XNOR U4676 ( .A(n4711), .B(n4660), .Z(n4714) );
  XOR U4677 ( .A(n4715), .B(n4707), .Z(n4660) );
  XNOR U4678 ( .A(n4716), .B(n4702), .Z(n4707) );
  XOR U4679 ( .A(n4717), .B(n4718), .Z(n4702) );
  AND U4680 ( .A(n4719), .B(n4720), .Z(n4718) );
  XOR U4681 ( .A(n4721), .B(n4717), .Z(n4719) );
  XNOR U4682 ( .A(n4722), .B(n4723), .Z(n4716) );
  AND U4683 ( .A(n4724), .B(n4725), .Z(n4723) );
  XOR U4684 ( .A(n4722), .B(n4726), .Z(n4724) );
  XNOR U4685 ( .A(n4708), .B(n4705), .Z(n4715) );
  AND U4686 ( .A(n4727), .B(n4728), .Z(n4705) );
  XOR U4687 ( .A(n4729), .B(n4730), .Z(n4708) );
  AND U4688 ( .A(n4731), .B(n4732), .Z(n4730) );
  XOR U4689 ( .A(n4729), .B(n4733), .Z(n4731) );
  XNOR U4690 ( .A(n4657), .B(n4711), .Z(n4713) );
  XNOR U4691 ( .A(n4734), .B(n4735), .Z(n4657) );
  AND U4692 ( .A(n100), .B(n4663), .Z(n4735) );
  XOR U4693 ( .A(n4734), .B(n4661), .Z(n4663) );
  XOR U4694 ( .A(n4736), .B(n4737), .Z(n4711) );
  AND U4695 ( .A(n4738), .B(n4739), .Z(n4737) );
  XNOR U4696 ( .A(n4736), .B(n4727), .Z(n4739) );
  IV U4697 ( .A(n4669), .Z(n4727) );
  XNOR U4698 ( .A(n4740), .B(n4720), .Z(n4669) );
  XNOR U4699 ( .A(n4741), .B(n4726), .Z(n4720) );
  XOR U4700 ( .A(n4742), .B(n4743), .Z(n4726) );
  AND U4701 ( .A(n4744), .B(n4745), .Z(n4743) );
  XOR U4702 ( .A(n4742), .B(n4746), .Z(n4744) );
  XNOR U4703 ( .A(n4725), .B(n4717), .Z(n4741) );
  XOR U4704 ( .A(n4747), .B(n4748), .Z(n4717) );
  AND U4705 ( .A(n4749), .B(n4750), .Z(n4748) );
  XNOR U4706 ( .A(n4751), .B(n4747), .Z(n4749) );
  XNOR U4707 ( .A(n4752), .B(n4722), .Z(n4725) );
  XOR U4708 ( .A(n4753), .B(n4754), .Z(n4722) );
  AND U4709 ( .A(n4755), .B(n4756), .Z(n4754) );
  XOR U4710 ( .A(n4753), .B(n4757), .Z(n4755) );
  XNOR U4711 ( .A(n4758), .B(n4759), .Z(n4752) );
  AND U4712 ( .A(n4760), .B(n4761), .Z(n4759) );
  XNOR U4713 ( .A(n4758), .B(n4762), .Z(n4760) );
  XNOR U4714 ( .A(n4721), .B(n4728), .Z(n4740) );
  AND U4715 ( .A(n4681), .B(n4763), .Z(n4728) );
  XOR U4716 ( .A(n4733), .B(n4732), .Z(n4721) );
  XNOR U4717 ( .A(n4764), .B(n4729), .Z(n4732) );
  XOR U4718 ( .A(n4765), .B(n4766), .Z(n4729) );
  AND U4719 ( .A(n4767), .B(n4768), .Z(n4766) );
  XOR U4720 ( .A(n4765), .B(n4769), .Z(n4767) );
  XNOR U4721 ( .A(n4770), .B(n4771), .Z(n4764) );
  AND U4722 ( .A(n4772), .B(n4773), .Z(n4771) );
  XOR U4723 ( .A(n4770), .B(n4774), .Z(n4772) );
  XOR U4724 ( .A(n4775), .B(n4776), .Z(n4733) );
  AND U4725 ( .A(n4777), .B(n4778), .Z(n4776) );
  XOR U4726 ( .A(n4775), .B(n4779), .Z(n4777) );
  XNOR U4727 ( .A(n4666), .B(n4736), .Z(n4738) );
  XNOR U4728 ( .A(n4780), .B(n4781), .Z(n4666) );
  AND U4729 ( .A(n100), .B(n4673), .Z(n4781) );
  XOR U4730 ( .A(n4780), .B(n4671), .Z(n4673) );
  XOR U4731 ( .A(n4782), .B(n4783), .Z(n4736) );
  AND U4732 ( .A(n4784), .B(n4785), .Z(n4783) );
  XNOR U4733 ( .A(n4782), .B(n4681), .Z(n4785) );
  XOR U4734 ( .A(n4786), .B(n4750), .Z(n4681) );
  XNOR U4735 ( .A(n4787), .B(n4757), .Z(n4750) );
  XOR U4736 ( .A(n4746), .B(n4745), .Z(n4757) );
  XNOR U4737 ( .A(n4788), .B(n4742), .Z(n4745) );
  XOR U4738 ( .A(n4789), .B(n4790), .Z(n4742) );
  AND U4739 ( .A(n4791), .B(n4792), .Z(n4790) );
  XNOR U4740 ( .A(n4793), .B(n4794), .Z(n4791) );
  IV U4741 ( .A(n4789), .Z(n4793) );
  XNOR U4742 ( .A(n4795), .B(n4796), .Z(n4788) );
  NOR U4743 ( .A(n4797), .B(n4798), .Z(n4796) );
  XNOR U4744 ( .A(n4795), .B(n4799), .Z(n4797) );
  XOR U4745 ( .A(n4800), .B(n4801), .Z(n4746) );
  NOR U4746 ( .A(n4802), .B(n4803), .Z(n4801) );
  XNOR U4747 ( .A(n4800), .B(n4804), .Z(n4802) );
  XNOR U4748 ( .A(n4756), .B(n4747), .Z(n4787) );
  XOR U4749 ( .A(n4805), .B(n4806), .Z(n4747) );
  AND U4750 ( .A(n4807), .B(n4808), .Z(n4806) );
  XOR U4751 ( .A(n4805), .B(n4809), .Z(n4807) );
  XOR U4752 ( .A(n4810), .B(n4762), .Z(n4756) );
  XOR U4753 ( .A(n4811), .B(n4812), .Z(n4762) );
  NOR U4754 ( .A(n4813), .B(n4814), .Z(n4812) );
  XOR U4755 ( .A(n4811), .B(n4815), .Z(n4813) );
  XNOR U4756 ( .A(n4761), .B(n4753), .Z(n4810) );
  XOR U4757 ( .A(n4816), .B(n4817), .Z(n4753) );
  AND U4758 ( .A(n4818), .B(n4819), .Z(n4817) );
  XOR U4759 ( .A(n4816), .B(n4820), .Z(n4818) );
  XNOR U4760 ( .A(n4821), .B(n4758), .Z(n4761) );
  XOR U4761 ( .A(n4822), .B(n4823), .Z(n4758) );
  AND U4762 ( .A(n4824), .B(n4825), .Z(n4823) );
  XNOR U4763 ( .A(n4826), .B(n4827), .Z(n4824) );
  IV U4764 ( .A(n4822), .Z(n4826) );
  XNOR U4765 ( .A(n4828), .B(n4829), .Z(n4821) );
  NOR U4766 ( .A(n4830), .B(n4831), .Z(n4829) );
  XNOR U4767 ( .A(n4828), .B(n4832), .Z(n4830) );
  XOR U4768 ( .A(n4751), .B(n4763), .Z(n4786) );
  NOR U4769 ( .A(n4689), .B(n4833), .Z(n4763) );
  XNOR U4770 ( .A(n4769), .B(n4768), .Z(n4751) );
  XNOR U4771 ( .A(n4834), .B(n4774), .Z(n4768) );
  XNOR U4772 ( .A(n4835), .B(n4836), .Z(n4774) );
  NOR U4773 ( .A(n4837), .B(n4838), .Z(n4836) );
  XOR U4774 ( .A(n4835), .B(n4839), .Z(n4837) );
  XNOR U4775 ( .A(n4773), .B(n4765), .Z(n4834) );
  XOR U4776 ( .A(n4840), .B(n4841), .Z(n4765) );
  AND U4777 ( .A(n4842), .B(n4843), .Z(n4841) );
  XOR U4778 ( .A(n4840), .B(n4844), .Z(n4842) );
  XNOR U4779 ( .A(n4845), .B(n4770), .Z(n4773) );
  XOR U4780 ( .A(n4846), .B(n4847), .Z(n4770) );
  AND U4781 ( .A(n4848), .B(n4849), .Z(n4847) );
  XNOR U4782 ( .A(n4850), .B(n4851), .Z(n4848) );
  IV U4783 ( .A(n4846), .Z(n4850) );
  XNOR U4784 ( .A(n4852), .B(n4853), .Z(n4845) );
  NOR U4785 ( .A(n4854), .B(n4855), .Z(n4853) );
  XNOR U4786 ( .A(n4852), .B(n4856), .Z(n4854) );
  XOR U4787 ( .A(n4779), .B(n4778), .Z(n4769) );
  XNOR U4788 ( .A(n4857), .B(n4775), .Z(n4778) );
  XOR U4789 ( .A(n4858), .B(n4859), .Z(n4775) );
  AND U4790 ( .A(n4860), .B(n4861), .Z(n4859) );
  XOR U4791 ( .A(n4858), .B(n4862), .Z(n4860) );
  XNOR U4792 ( .A(n4863), .B(n4864), .Z(n4857) );
  NOR U4793 ( .A(n4865), .B(n4866), .Z(n4864) );
  XNOR U4794 ( .A(n4863), .B(n4867), .Z(n4865) );
  XOR U4795 ( .A(n4868), .B(n4869), .Z(n4779) );
  NOR U4796 ( .A(n4870), .B(n4871), .Z(n4869) );
  XNOR U4797 ( .A(n4868), .B(n4872), .Z(n4870) );
  XNOR U4798 ( .A(n4678), .B(n4782), .Z(n4784) );
  XNOR U4799 ( .A(n4873), .B(n4874), .Z(n4678) );
  AND U4800 ( .A(n100), .B(n4685), .Z(n4874) );
  XOR U4801 ( .A(n4873), .B(n4683), .Z(n4685) );
  AND U4802 ( .A(n4686), .B(n4689), .Z(n4782) );
  XOR U4803 ( .A(n4875), .B(n4833), .Z(n4689) );
  XNOR U4804 ( .A(p_input[512]), .B(p_input[96]), .Z(n4833) );
  XNOR U4805 ( .A(n4809), .B(n4808), .Z(n4875) );
  XNOR U4806 ( .A(n4876), .B(n4820), .Z(n4808) );
  XOR U4807 ( .A(n4794), .B(n4792), .Z(n4820) );
  XNOR U4808 ( .A(n4877), .B(n4799), .Z(n4792) );
  XOR U4809 ( .A(p_input[120]), .B(p_input[536]), .Z(n4799) );
  XOR U4810 ( .A(n4789), .B(n4798), .Z(n4877) );
  XOR U4811 ( .A(n4878), .B(n4795), .Z(n4798) );
  XOR U4812 ( .A(p_input[118]), .B(p_input[534]), .Z(n4795) );
  XOR U4813 ( .A(p_input[119]), .B(n4010), .Z(n4878) );
  XOR U4814 ( .A(p_input[114]), .B(p_input[530]), .Z(n4789) );
  XNOR U4815 ( .A(n4804), .B(n4803), .Z(n4794) );
  XOR U4816 ( .A(n4879), .B(n4800), .Z(n4803) );
  XOR U4817 ( .A(p_input[115]), .B(p_input[531]), .Z(n4800) );
  XOR U4818 ( .A(p_input[116]), .B(n4012), .Z(n4879) );
  XOR U4819 ( .A(p_input[117]), .B(p_input[533]), .Z(n4804) );
  XNOR U4820 ( .A(n4819), .B(n4805), .Z(n4876) );
  XNOR U4821 ( .A(n4591), .B(p_input[97]), .Z(n4805) );
  XNOR U4822 ( .A(n4880), .B(n4827), .Z(n4819) );
  XNOR U4823 ( .A(n4815), .B(n4814), .Z(n4827) );
  XNOR U4824 ( .A(n4881), .B(n4811), .Z(n4814) );
  XNOR U4825 ( .A(p_input[122]), .B(p_input[538]), .Z(n4811) );
  XOR U4826 ( .A(p_input[123]), .B(n4016), .Z(n4881) );
  XOR U4827 ( .A(p_input[124]), .B(p_input[540]), .Z(n4815) );
  XOR U4828 ( .A(n4825), .B(n4882), .Z(n4880) );
  IV U4829 ( .A(n4816), .Z(n4882) );
  XOR U4830 ( .A(p_input[113]), .B(p_input[529]), .Z(n4816) );
  XNOR U4831 ( .A(n4883), .B(n4832), .Z(n4825) );
  XNOR U4832 ( .A(p_input[127]), .B(n4019), .Z(n4832) );
  XOR U4833 ( .A(n4822), .B(n4831), .Z(n4883) );
  XOR U4834 ( .A(n4884), .B(n4828), .Z(n4831) );
  XOR U4835 ( .A(p_input[125]), .B(p_input[541]), .Z(n4828) );
  XOR U4836 ( .A(p_input[126]), .B(n4021), .Z(n4884) );
  XOR U4837 ( .A(p_input[121]), .B(p_input[537]), .Z(n4822) );
  XOR U4838 ( .A(n4844), .B(n4843), .Z(n4809) );
  XNOR U4839 ( .A(n4885), .B(n4851), .Z(n4843) );
  XNOR U4840 ( .A(n4839), .B(n4838), .Z(n4851) );
  XNOR U4841 ( .A(n4886), .B(n4835), .Z(n4838) );
  XNOR U4842 ( .A(p_input[107]), .B(p_input[523]), .Z(n4835) );
  XOR U4843 ( .A(p_input[108]), .B(n4024), .Z(n4886) );
  XOR U4844 ( .A(p_input[109]), .B(p_input[525]), .Z(n4839) );
  XNOR U4845 ( .A(n4849), .B(n4840), .Z(n4885) );
  XNOR U4846 ( .A(n4600), .B(p_input[98]), .Z(n4840) );
  XNOR U4847 ( .A(n4887), .B(n4856), .Z(n4849) );
  XNOR U4848 ( .A(p_input[112]), .B(n4027), .Z(n4856) );
  XOR U4849 ( .A(n4846), .B(n4855), .Z(n4887) );
  XOR U4850 ( .A(n4888), .B(n4852), .Z(n4855) );
  XOR U4851 ( .A(p_input[110]), .B(p_input[526]), .Z(n4852) );
  XOR U4852 ( .A(p_input[111]), .B(n4029), .Z(n4888) );
  XOR U4853 ( .A(p_input[106]), .B(p_input[522]), .Z(n4846) );
  XOR U4854 ( .A(n4862), .B(n4861), .Z(n4844) );
  XNOR U4855 ( .A(n4889), .B(n4867), .Z(n4861) );
  XOR U4856 ( .A(p_input[105]), .B(p_input[521]), .Z(n4867) );
  XOR U4857 ( .A(n4858), .B(n4866), .Z(n4889) );
  XOR U4858 ( .A(n4890), .B(n4863), .Z(n4866) );
  XOR U4859 ( .A(p_input[103]), .B(p_input[519]), .Z(n4863) );
  XOR U4860 ( .A(p_input[104]), .B(n4318), .Z(n4890) );
  XNOR U4861 ( .A(n4606), .B(p_input[99]), .Z(n4858) );
  IV U4862 ( .A(p_input[515]), .Z(n4606) );
  XNOR U4863 ( .A(n4872), .B(n4871), .Z(n4862) );
  XOR U4864 ( .A(n4891), .B(n4868), .Z(n4871) );
  XOR U4865 ( .A(p_input[100]), .B(p_input[516]), .Z(n4868) );
  XOR U4866 ( .A(p_input[101]), .B(n4320), .Z(n4891) );
  XOR U4867 ( .A(p_input[102]), .B(p_input[518]), .Z(n4872) );
  XNOR U4868 ( .A(n4892), .B(n4893), .Z(n4686) );
  AND U4869 ( .A(n100), .B(n4894), .Z(n4893) );
  XNOR U4870 ( .A(n4895), .B(n4896), .Z(n100) );
  AND U4871 ( .A(n4897), .B(n4898), .Z(n4896) );
  XOR U4872 ( .A(n4895), .B(n4696), .Z(n4898) );
  XNOR U4873 ( .A(n4895), .B(n4638), .Z(n4897) );
  XOR U4874 ( .A(n4899), .B(n4900), .Z(n4895) );
  AND U4875 ( .A(n4901), .B(n4902), .Z(n4900) );
  XNOR U4876 ( .A(n4709), .B(n4899), .Z(n4902) );
  XOR U4877 ( .A(n4899), .B(n4650), .Z(n4901) );
  XOR U4878 ( .A(n4903), .B(n4904), .Z(n4899) );
  AND U4879 ( .A(n4905), .B(n4906), .Z(n4904) );
  XNOR U4880 ( .A(n4734), .B(n4903), .Z(n4906) );
  XOR U4881 ( .A(n4903), .B(n4661), .Z(n4905) );
  XOR U4882 ( .A(n4907), .B(n4908), .Z(n4903) );
  AND U4883 ( .A(n4909), .B(n4910), .Z(n4908) );
  XOR U4884 ( .A(n4907), .B(n4671), .Z(n4909) );
  XOR U4885 ( .A(n4911), .B(n4912), .Z(n4627) );
  AND U4886 ( .A(n104), .B(n4894), .Z(n4912) );
  XNOR U4887 ( .A(n4892), .B(n4911), .Z(n4894) );
  XNOR U4888 ( .A(n4913), .B(n4914), .Z(n104) );
  AND U4889 ( .A(n4915), .B(n4916), .Z(n4914) );
  XNOR U4890 ( .A(n4917), .B(n4913), .Z(n4916) );
  IV U4891 ( .A(n4696), .Z(n4917) );
  XNOR U4892 ( .A(n4918), .B(n4919), .Z(n4696) );
  AND U4893 ( .A(n107), .B(n4920), .Z(n4919) );
  XNOR U4894 ( .A(n4918), .B(n4921), .Z(n4920) );
  XNOR U4895 ( .A(n4638), .B(n4913), .Z(n4915) );
  XOR U4896 ( .A(n4922), .B(n4923), .Z(n4638) );
  AND U4897 ( .A(n115), .B(n4924), .Z(n4923) );
  XOR U4898 ( .A(n4925), .B(n4926), .Z(n4913) );
  AND U4899 ( .A(n4927), .B(n4928), .Z(n4926) );
  XNOR U4900 ( .A(n4925), .B(n4709), .Z(n4928) );
  XNOR U4901 ( .A(n4929), .B(n4930), .Z(n4709) );
  AND U4902 ( .A(n107), .B(n4931), .Z(n4930) );
  XOR U4903 ( .A(n4932), .B(n4929), .Z(n4931) );
  XNOR U4904 ( .A(n4933), .B(n4925), .Z(n4927) );
  IV U4905 ( .A(n4650), .Z(n4933) );
  XOR U4906 ( .A(n4934), .B(n4935), .Z(n4650) );
  AND U4907 ( .A(n115), .B(n4936), .Z(n4935) );
  XOR U4908 ( .A(n4937), .B(n4938), .Z(n4925) );
  AND U4909 ( .A(n4939), .B(n4940), .Z(n4938) );
  XNOR U4910 ( .A(n4937), .B(n4734), .Z(n4940) );
  XNOR U4911 ( .A(n4941), .B(n4942), .Z(n4734) );
  AND U4912 ( .A(n107), .B(n4943), .Z(n4942) );
  XNOR U4913 ( .A(n4944), .B(n4941), .Z(n4943) );
  XOR U4914 ( .A(n4661), .B(n4937), .Z(n4939) );
  XOR U4915 ( .A(n4945), .B(n4946), .Z(n4661) );
  AND U4916 ( .A(n115), .B(n4947), .Z(n4946) );
  XOR U4917 ( .A(n4907), .B(n4948), .Z(n4937) );
  AND U4918 ( .A(n4949), .B(n4910), .Z(n4948) );
  XNOR U4919 ( .A(n4780), .B(n4907), .Z(n4910) );
  XNOR U4920 ( .A(n4950), .B(n4951), .Z(n4780) );
  AND U4921 ( .A(n107), .B(n4952), .Z(n4951) );
  XOR U4922 ( .A(n4953), .B(n4950), .Z(n4952) );
  XNOR U4923 ( .A(n4954), .B(n4907), .Z(n4949) );
  IV U4924 ( .A(n4671), .Z(n4954) );
  XOR U4925 ( .A(n4955), .B(n4956), .Z(n4671) );
  AND U4926 ( .A(n115), .B(n4957), .Z(n4956) );
  XOR U4927 ( .A(n4958), .B(n4959), .Z(n4907) );
  AND U4928 ( .A(n4960), .B(n4961), .Z(n4959) );
  XNOR U4929 ( .A(n4958), .B(n4873), .Z(n4961) );
  XNOR U4930 ( .A(n4962), .B(n4963), .Z(n4873) );
  AND U4931 ( .A(n107), .B(n4964), .Z(n4963) );
  XNOR U4932 ( .A(n4965), .B(n4962), .Z(n4964) );
  XNOR U4933 ( .A(n4966), .B(n4958), .Z(n4960) );
  IV U4934 ( .A(n4683), .Z(n4966) );
  XOR U4935 ( .A(n4967), .B(n4968), .Z(n4683) );
  AND U4936 ( .A(n115), .B(n4969), .Z(n4968) );
  AND U4937 ( .A(n4911), .B(n4892), .Z(n4958) );
  XNOR U4938 ( .A(n4970), .B(n4971), .Z(n4892) );
  AND U4939 ( .A(n107), .B(n4972), .Z(n4971) );
  XNOR U4940 ( .A(n4973), .B(n4970), .Z(n4972) );
  XNOR U4941 ( .A(n4974), .B(n4975), .Z(n107) );
  AND U4942 ( .A(n4976), .B(n4977), .Z(n4975) );
  XOR U4943 ( .A(n4921), .B(n4974), .Z(n4977) );
  AND U4944 ( .A(n4978), .B(n4979), .Z(n4921) );
  XOR U4945 ( .A(n4974), .B(n4918), .Z(n4976) );
  XNOR U4946 ( .A(n4980), .B(n4981), .Z(n4918) );
  AND U4947 ( .A(n111), .B(n4924), .Z(n4981) );
  XOR U4948 ( .A(n4922), .B(n4980), .Z(n4924) );
  XOR U4949 ( .A(n4982), .B(n4983), .Z(n4974) );
  AND U4950 ( .A(n4984), .B(n4985), .Z(n4983) );
  XNOR U4951 ( .A(n4982), .B(n4978), .Z(n4985) );
  IV U4952 ( .A(n4932), .Z(n4978) );
  XOR U4953 ( .A(n4986), .B(n4987), .Z(n4932) );
  XOR U4954 ( .A(n4988), .B(n4979), .Z(n4987) );
  AND U4955 ( .A(n4944), .B(n4989), .Z(n4979) );
  AND U4956 ( .A(n4990), .B(n4991), .Z(n4988) );
  XOR U4957 ( .A(n4992), .B(n4986), .Z(n4990) );
  XNOR U4958 ( .A(n4929), .B(n4982), .Z(n4984) );
  XNOR U4959 ( .A(n4993), .B(n4994), .Z(n4929) );
  AND U4960 ( .A(n111), .B(n4936), .Z(n4994) );
  XOR U4961 ( .A(n4993), .B(n4934), .Z(n4936) );
  XOR U4962 ( .A(n4995), .B(n4996), .Z(n4982) );
  AND U4963 ( .A(n4997), .B(n4998), .Z(n4996) );
  XNOR U4964 ( .A(n4995), .B(n4944), .Z(n4998) );
  XOR U4965 ( .A(n4999), .B(n4991), .Z(n4944) );
  XNOR U4966 ( .A(n5000), .B(n4986), .Z(n4991) );
  XOR U4967 ( .A(n5001), .B(n5002), .Z(n4986) );
  AND U4968 ( .A(n5003), .B(n5004), .Z(n5002) );
  XOR U4969 ( .A(n5005), .B(n5001), .Z(n5003) );
  XNOR U4970 ( .A(n5006), .B(n5007), .Z(n5000) );
  AND U4971 ( .A(n5008), .B(n5009), .Z(n5007) );
  XOR U4972 ( .A(n5006), .B(n5010), .Z(n5008) );
  XNOR U4973 ( .A(n4992), .B(n4989), .Z(n4999) );
  AND U4974 ( .A(n5011), .B(n5012), .Z(n4989) );
  XOR U4975 ( .A(n5013), .B(n5014), .Z(n4992) );
  AND U4976 ( .A(n5015), .B(n5016), .Z(n5014) );
  XOR U4977 ( .A(n5013), .B(n5017), .Z(n5015) );
  XNOR U4978 ( .A(n4941), .B(n4995), .Z(n4997) );
  XNOR U4979 ( .A(n5018), .B(n5019), .Z(n4941) );
  AND U4980 ( .A(n111), .B(n4947), .Z(n5019) );
  XOR U4981 ( .A(n5018), .B(n4945), .Z(n4947) );
  XOR U4982 ( .A(n5020), .B(n5021), .Z(n4995) );
  AND U4983 ( .A(n5022), .B(n5023), .Z(n5021) );
  XNOR U4984 ( .A(n5020), .B(n5011), .Z(n5023) );
  IV U4985 ( .A(n4953), .Z(n5011) );
  XNOR U4986 ( .A(n5024), .B(n5004), .Z(n4953) );
  XNOR U4987 ( .A(n5025), .B(n5010), .Z(n5004) );
  XOR U4988 ( .A(n5026), .B(n5027), .Z(n5010) );
  AND U4989 ( .A(n5028), .B(n5029), .Z(n5027) );
  XOR U4990 ( .A(n5026), .B(n5030), .Z(n5028) );
  XNOR U4991 ( .A(n5009), .B(n5001), .Z(n5025) );
  XOR U4992 ( .A(n5031), .B(n5032), .Z(n5001) );
  AND U4993 ( .A(n5033), .B(n5034), .Z(n5032) );
  XNOR U4994 ( .A(n5035), .B(n5031), .Z(n5033) );
  XNOR U4995 ( .A(n5036), .B(n5006), .Z(n5009) );
  XOR U4996 ( .A(n5037), .B(n5038), .Z(n5006) );
  AND U4997 ( .A(n5039), .B(n5040), .Z(n5038) );
  XOR U4998 ( .A(n5037), .B(n5041), .Z(n5039) );
  XNOR U4999 ( .A(n5042), .B(n5043), .Z(n5036) );
  AND U5000 ( .A(n5044), .B(n5045), .Z(n5043) );
  XNOR U5001 ( .A(n5042), .B(n5046), .Z(n5044) );
  XNOR U5002 ( .A(n5005), .B(n5012), .Z(n5024) );
  AND U5003 ( .A(n4965), .B(n5047), .Z(n5012) );
  XOR U5004 ( .A(n5017), .B(n5016), .Z(n5005) );
  XNOR U5005 ( .A(n5048), .B(n5013), .Z(n5016) );
  XOR U5006 ( .A(n5049), .B(n5050), .Z(n5013) );
  AND U5007 ( .A(n5051), .B(n5052), .Z(n5050) );
  XOR U5008 ( .A(n5049), .B(n5053), .Z(n5051) );
  XNOR U5009 ( .A(n5054), .B(n5055), .Z(n5048) );
  AND U5010 ( .A(n5056), .B(n5057), .Z(n5055) );
  XOR U5011 ( .A(n5054), .B(n5058), .Z(n5056) );
  XOR U5012 ( .A(n5059), .B(n5060), .Z(n5017) );
  AND U5013 ( .A(n5061), .B(n5062), .Z(n5060) );
  XOR U5014 ( .A(n5059), .B(n5063), .Z(n5061) );
  XNOR U5015 ( .A(n4950), .B(n5020), .Z(n5022) );
  XNOR U5016 ( .A(n5064), .B(n5065), .Z(n4950) );
  AND U5017 ( .A(n111), .B(n4957), .Z(n5065) );
  XOR U5018 ( .A(n5064), .B(n4955), .Z(n4957) );
  XOR U5019 ( .A(n5066), .B(n5067), .Z(n5020) );
  AND U5020 ( .A(n5068), .B(n5069), .Z(n5067) );
  XNOR U5021 ( .A(n5066), .B(n4965), .Z(n5069) );
  XOR U5022 ( .A(n5070), .B(n5034), .Z(n4965) );
  XNOR U5023 ( .A(n5071), .B(n5041), .Z(n5034) );
  XOR U5024 ( .A(n5030), .B(n5029), .Z(n5041) );
  XNOR U5025 ( .A(n5072), .B(n5026), .Z(n5029) );
  XOR U5026 ( .A(n5073), .B(n5074), .Z(n5026) );
  AND U5027 ( .A(n5075), .B(n5076), .Z(n5074) );
  XNOR U5028 ( .A(n5077), .B(n5078), .Z(n5075) );
  IV U5029 ( .A(n5073), .Z(n5077) );
  XNOR U5030 ( .A(n5079), .B(n5080), .Z(n5072) );
  NOR U5031 ( .A(n5081), .B(n5082), .Z(n5080) );
  XNOR U5032 ( .A(n5079), .B(n5083), .Z(n5081) );
  XOR U5033 ( .A(n5084), .B(n5085), .Z(n5030) );
  NOR U5034 ( .A(n5086), .B(n5087), .Z(n5085) );
  XNOR U5035 ( .A(n5084), .B(n5088), .Z(n5086) );
  XNOR U5036 ( .A(n5040), .B(n5031), .Z(n5071) );
  XOR U5037 ( .A(n5089), .B(n5090), .Z(n5031) );
  AND U5038 ( .A(n5091), .B(n5092), .Z(n5090) );
  XOR U5039 ( .A(n5089), .B(n5093), .Z(n5091) );
  XOR U5040 ( .A(n5094), .B(n5046), .Z(n5040) );
  XOR U5041 ( .A(n5095), .B(n5096), .Z(n5046) );
  NOR U5042 ( .A(n5097), .B(n5098), .Z(n5096) );
  XOR U5043 ( .A(n5095), .B(n5099), .Z(n5097) );
  XNOR U5044 ( .A(n5045), .B(n5037), .Z(n5094) );
  XOR U5045 ( .A(n5100), .B(n5101), .Z(n5037) );
  AND U5046 ( .A(n5102), .B(n5103), .Z(n5101) );
  XOR U5047 ( .A(n5100), .B(n5104), .Z(n5102) );
  XNOR U5048 ( .A(n5105), .B(n5042), .Z(n5045) );
  XOR U5049 ( .A(n5106), .B(n5107), .Z(n5042) );
  AND U5050 ( .A(n5108), .B(n5109), .Z(n5107) );
  XNOR U5051 ( .A(n5110), .B(n5111), .Z(n5108) );
  IV U5052 ( .A(n5106), .Z(n5110) );
  XNOR U5053 ( .A(n5112), .B(n5113), .Z(n5105) );
  NOR U5054 ( .A(n5114), .B(n5115), .Z(n5113) );
  XNOR U5055 ( .A(n5112), .B(n5116), .Z(n5114) );
  XOR U5056 ( .A(n5035), .B(n5047), .Z(n5070) );
  NOR U5057 ( .A(n4973), .B(n5117), .Z(n5047) );
  XNOR U5058 ( .A(n5053), .B(n5052), .Z(n5035) );
  XNOR U5059 ( .A(n5118), .B(n5058), .Z(n5052) );
  XNOR U5060 ( .A(n5119), .B(n5120), .Z(n5058) );
  NOR U5061 ( .A(n5121), .B(n5122), .Z(n5120) );
  XOR U5062 ( .A(n5119), .B(n5123), .Z(n5121) );
  XNOR U5063 ( .A(n5057), .B(n5049), .Z(n5118) );
  XOR U5064 ( .A(n5124), .B(n5125), .Z(n5049) );
  AND U5065 ( .A(n5126), .B(n5127), .Z(n5125) );
  XOR U5066 ( .A(n5124), .B(n5128), .Z(n5126) );
  XNOR U5067 ( .A(n5129), .B(n5054), .Z(n5057) );
  XOR U5068 ( .A(n5130), .B(n5131), .Z(n5054) );
  AND U5069 ( .A(n5132), .B(n5133), .Z(n5131) );
  XNOR U5070 ( .A(n5134), .B(n5135), .Z(n5132) );
  IV U5071 ( .A(n5130), .Z(n5134) );
  XNOR U5072 ( .A(n5136), .B(n5137), .Z(n5129) );
  NOR U5073 ( .A(n5138), .B(n5139), .Z(n5137) );
  XNOR U5074 ( .A(n5136), .B(n5140), .Z(n5138) );
  XOR U5075 ( .A(n5063), .B(n5062), .Z(n5053) );
  XNOR U5076 ( .A(n5141), .B(n5059), .Z(n5062) );
  XOR U5077 ( .A(n5142), .B(n5143), .Z(n5059) );
  AND U5078 ( .A(n5144), .B(n5145), .Z(n5143) );
  XNOR U5079 ( .A(n5146), .B(n5147), .Z(n5144) );
  IV U5080 ( .A(n5142), .Z(n5146) );
  XNOR U5081 ( .A(n5148), .B(n5149), .Z(n5141) );
  NOR U5082 ( .A(n5150), .B(n5151), .Z(n5149) );
  XNOR U5083 ( .A(n5148), .B(n5152), .Z(n5150) );
  XOR U5084 ( .A(n5153), .B(n5154), .Z(n5063) );
  NOR U5085 ( .A(n5155), .B(n5156), .Z(n5154) );
  XNOR U5086 ( .A(n5153), .B(n5157), .Z(n5155) );
  XNOR U5087 ( .A(n4962), .B(n5066), .Z(n5068) );
  XNOR U5088 ( .A(n5158), .B(n5159), .Z(n4962) );
  AND U5089 ( .A(n111), .B(n4969), .Z(n5159) );
  XOR U5090 ( .A(n5158), .B(n4967), .Z(n4969) );
  AND U5091 ( .A(n4970), .B(n4973), .Z(n5066) );
  XOR U5092 ( .A(n5160), .B(n5117), .Z(n4973) );
  XNOR U5093 ( .A(p_input[128]), .B(p_input[512]), .Z(n5117) );
  XNOR U5094 ( .A(n5093), .B(n5092), .Z(n5160) );
  XNOR U5095 ( .A(n5161), .B(n5104), .Z(n5092) );
  XOR U5096 ( .A(n5078), .B(n5076), .Z(n5104) );
  XNOR U5097 ( .A(n5162), .B(n5083), .Z(n5076) );
  XOR U5098 ( .A(p_input[152]), .B(p_input[536]), .Z(n5083) );
  XOR U5099 ( .A(n5073), .B(n5082), .Z(n5162) );
  XOR U5100 ( .A(n5163), .B(n5079), .Z(n5082) );
  XOR U5101 ( .A(p_input[150]), .B(p_input[534]), .Z(n5079) );
  XOR U5102 ( .A(p_input[151]), .B(n4010), .Z(n5163) );
  XOR U5103 ( .A(p_input[146]), .B(p_input[530]), .Z(n5073) );
  XNOR U5104 ( .A(n5088), .B(n5087), .Z(n5078) );
  XOR U5105 ( .A(n5164), .B(n5084), .Z(n5087) );
  XOR U5106 ( .A(p_input[147]), .B(p_input[531]), .Z(n5084) );
  XOR U5107 ( .A(p_input[148]), .B(n4012), .Z(n5164) );
  XOR U5108 ( .A(p_input[149]), .B(p_input[533]), .Z(n5088) );
  XOR U5109 ( .A(n5103), .B(n5165), .Z(n5161) );
  IV U5110 ( .A(n5089), .Z(n5165) );
  XOR U5111 ( .A(p_input[129]), .B(p_input[513]), .Z(n5089) );
  XNOR U5112 ( .A(n5166), .B(n5111), .Z(n5103) );
  XNOR U5113 ( .A(n5099), .B(n5098), .Z(n5111) );
  XNOR U5114 ( .A(n5167), .B(n5095), .Z(n5098) );
  XNOR U5115 ( .A(p_input[154]), .B(p_input[538]), .Z(n5095) );
  XOR U5116 ( .A(p_input[155]), .B(n4016), .Z(n5167) );
  XOR U5117 ( .A(p_input[156]), .B(p_input[540]), .Z(n5099) );
  XOR U5118 ( .A(n5109), .B(n5168), .Z(n5166) );
  IV U5119 ( .A(n5100), .Z(n5168) );
  XOR U5120 ( .A(p_input[145]), .B(p_input[529]), .Z(n5100) );
  XNOR U5121 ( .A(n5169), .B(n5116), .Z(n5109) );
  XNOR U5122 ( .A(p_input[159]), .B(n4019), .Z(n5116) );
  XOR U5123 ( .A(n5106), .B(n5115), .Z(n5169) );
  XOR U5124 ( .A(n5170), .B(n5112), .Z(n5115) );
  XOR U5125 ( .A(p_input[157]), .B(p_input[541]), .Z(n5112) );
  XOR U5126 ( .A(p_input[158]), .B(n4021), .Z(n5170) );
  XOR U5127 ( .A(p_input[153]), .B(p_input[537]), .Z(n5106) );
  XOR U5128 ( .A(n5128), .B(n5127), .Z(n5093) );
  XNOR U5129 ( .A(n5171), .B(n5135), .Z(n5127) );
  XNOR U5130 ( .A(n5123), .B(n5122), .Z(n5135) );
  XNOR U5131 ( .A(n5172), .B(n5119), .Z(n5122) );
  XNOR U5132 ( .A(p_input[139]), .B(p_input[523]), .Z(n5119) );
  XOR U5133 ( .A(p_input[140]), .B(n4024), .Z(n5172) );
  XOR U5134 ( .A(p_input[141]), .B(p_input[525]), .Z(n5123) );
  XOR U5135 ( .A(n5133), .B(n5173), .Z(n5171) );
  IV U5136 ( .A(n5124), .Z(n5173) );
  XOR U5137 ( .A(p_input[130]), .B(p_input[514]), .Z(n5124) );
  XNOR U5138 ( .A(n5174), .B(n5140), .Z(n5133) );
  XNOR U5139 ( .A(p_input[144]), .B(n4027), .Z(n5140) );
  XOR U5140 ( .A(n5130), .B(n5139), .Z(n5174) );
  XOR U5141 ( .A(n5175), .B(n5136), .Z(n5139) );
  XOR U5142 ( .A(p_input[142]), .B(p_input[526]), .Z(n5136) );
  XOR U5143 ( .A(p_input[143]), .B(n4029), .Z(n5175) );
  XOR U5144 ( .A(p_input[138]), .B(p_input[522]), .Z(n5130) );
  XOR U5145 ( .A(n5147), .B(n5145), .Z(n5128) );
  XNOR U5146 ( .A(n5176), .B(n5152), .Z(n5145) );
  XOR U5147 ( .A(p_input[137]), .B(p_input[521]), .Z(n5152) );
  XOR U5148 ( .A(n5142), .B(n5151), .Z(n5176) );
  XOR U5149 ( .A(n5177), .B(n5148), .Z(n5151) );
  XOR U5150 ( .A(p_input[135]), .B(p_input[519]), .Z(n5148) );
  XOR U5151 ( .A(p_input[136]), .B(n4318), .Z(n5177) );
  XOR U5152 ( .A(p_input[131]), .B(p_input[515]), .Z(n5142) );
  XNOR U5153 ( .A(n5157), .B(n5156), .Z(n5147) );
  XOR U5154 ( .A(n5178), .B(n5153), .Z(n5156) );
  XOR U5155 ( .A(p_input[132]), .B(p_input[516]), .Z(n5153) );
  XOR U5156 ( .A(p_input[133]), .B(n4320), .Z(n5178) );
  XOR U5157 ( .A(p_input[134]), .B(p_input[518]), .Z(n5157) );
  XNOR U5158 ( .A(n5179), .B(n5180), .Z(n4970) );
  AND U5159 ( .A(n111), .B(n5181), .Z(n5180) );
  XNOR U5160 ( .A(n5182), .B(n5183), .Z(n111) );
  AND U5161 ( .A(n5184), .B(n5185), .Z(n5183) );
  XOR U5162 ( .A(n5182), .B(n4980), .Z(n5185) );
  XNOR U5163 ( .A(n5182), .B(n4922), .Z(n5184) );
  XOR U5164 ( .A(n5186), .B(n5187), .Z(n5182) );
  AND U5165 ( .A(n5188), .B(n5189), .Z(n5187) );
  XNOR U5166 ( .A(n4993), .B(n5186), .Z(n5189) );
  XOR U5167 ( .A(n5186), .B(n4934), .Z(n5188) );
  XOR U5168 ( .A(n5190), .B(n5191), .Z(n5186) );
  AND U5169 ( .A(n5192), .B(n5193), .Z(n5191) );
  XNOR U5170 ( .A(n5018), .B(n5190), .Z(n5193) );
  XOR U5171 ( .A(n5190), .B(n4945), .Z(n5192) );
  XOR U5172 ( .A(n5194), .B(n5195), .Z(n5190) );
  AND U5173 ( .A(n5196), .B(n5197), .Z(n5195) );
  XOR U5174 ( .A(n5194), .B(n4955), .Z(n5196) );
  XOR U5175 ( .A(n5198), .B(n5199), .Z(n4911) );
  AND U5176 ( .A(n115), .B(n5181), .Z(n5199) );
  XNOR U5177 ( .A(n5179), .B(n5198), .Z(n5181) );
  XNOR U5178 ( .A(n5200), .B(n5201), .Z(n115) );
  AND U5179 ( .A(n5202), .B(n5203), .Z(n5201) );
  XNOR U5180 ( .A(n5204), .B(n5200), .Z(n5203) );
  IV U5181 ( .A(n4980), .Z(n5204) );
  XNOR U5182 ( .A(n5205), .B(n5206), .Z(n4980) );
  AND U5183 ( .A(n118), .B(n5207), .Z(n5206) );
  XNOR U5184 ( .A(n5205), .B(n5208), .Z(n5207) );
  XNOR U5185 ( .A(n4922), .B(n5200), .Z(n5202) );
  XOR U5186 ( .A(n5209), .B(n5210), .Z(n4922) );
  AND U5187 ( .A(n126), .B(n5211), .Z(n5210) );
  XOR U5188 ( .A(n5212), .B(n5213), .Z(n5200) );
  AND U5189 ( .A(n5214), .B(n5215), .Z(n5213) );
  XNOR U5190 ( .A(n5212), .B(n4993), .Z(n5215) );
  XNOR U5191 ( .A(n5216), .B(n5217), .Z(n4993) );
  AND U5192 ( .A(n118), .B(n5218), .Z(n5217) );
  XOR U5193 ( .A(n5219), .B(n5216), .Z(n5218) );
  XNOR U5194 ( .A(n5220), .B(n5212), .Z(n5214) );
  IV U5195 ( .A(n4934), .Z(n5220) );
  XOR U5196 ( .A(n5221), .B(n5222), .Z(n4934) );
  AND U5197 ( .A(n126), .B(n5223), .Z(n5222) );
  XOR U5198 ( .A(n5224), .B(n5225), .Z(n5212) );
  AND U5199 ( .A(n5226), .B(n5227), .Z(n5225) );
  XNOR U5200 ( .A(n5224), .B(n5018), .Z(n5227) );
  XNOR U5201 ( .A(n5228), .B(n5229), .Z(n5018) );
  AND U5202 ( .A(n118), .B(n5230), .Z(n5229) );
  XNOR U5203 ( .A(n5231), .B(n5228), .Z(n5230) );
  XOR U5204 ( .A(n4945), .B(n5224), .Z(n5226) );
  XOR U5205 ( .A(n5232), .B(n5233), .Z(n4945) );
  AND U5206 ( .A(n126), .B(n5234), .Z(n5233) );
  XOR U5207 ( .A(n5194), .B(n5235), .Z(n5224) );
  AND U5208 ( .A(n5236), .B(n5197), .Z(n5235) );
  XNOR U5209 ( .A(n5064), .B(n5194), .Z(n5197) );
  XNOR U5210 ( .A(n5237), .B(n5238), .Z(n5064) );
  AND U5211 ( .A(n118), .B(n5239), .Z(n5238) );
  XOR U5212 ( .A(n5240), .B(n5237), .Z(n5239) );
  XNOR U5213 ( .A(n5241), .B(n5194), .Z(n5236) );
  IV U5214 ( .A(n4955), .Z(n5241) );
  XOR U5215 ( .A(n5242), .B(n5243), .Z(n4955) );
  AND U5216 ( .A(n126), .B(n5244), .Z(n5243) );
  XOR U5217 ( .A(n5245), .B(n5246), .Z(n5194) );
  AND U5218 ( .A(n5247), .B(n5248), .Z(n5246) );
  XNOR U5219 ( .A(n5245), .B(n5158), .Z(n5248) );
  XNOR U5220 ( .A(n5249), .B(n5250), .Z(n5158) );
  AND U5221 ( .A(n118), .B(n5251), .Z(n5250) );
  XNOR U5222 ( .A(n5252), .B(n5249), .Z(n5251) );
  XNOR U5223 ( .A(n5253), .B(n5245), .Z(n5247) );
  IV U5224 ( .A(n4967), .Z(n5253) );
  XOR U5225 ( .A(n5254), .B(n5255), .Z(n4967) );
  AND U5226 ( .A(n126), .B(n5256), .Z(n5255) );
  AND U5227 ( .A(n5198), .B(n5179), .Z(n5245) );
  XNOR U5228 ( .A(n5257), .B(n5258), .Z(n5179) );
  AND U5229 ( .A(n118), .B(n5259), .Z(n5258) );
  XNOR U5230 ( .A(n5260), .B(n5257), .Z(n5259) );
  XNOR U5231 ( .A(n5261), .B(n5262), .Z(n118) );
  AND U5232 ( .A(n5263), .B(n5264), .Z(n5262) );
  XOR U5233 ( .A(n5208), .B(n5261), .Z(n5264) );
  AND U5234 ( .A(n5265), .B(n5266), .Z(n5208) );
  XOR U5235 ( .A(n5261), .B(n5205), .Z(n5263) );
  XNOR U5236 ( .A(n5267), .B(n5268), .Z(n5205) );
  AND U5237 ( .A(n122), .B(n5211), .Z(n5268) );
  XOR U5238 ( .A(n5209), .B(n5267), .Z(n5211) );
  XOR U5239 ( .A(n5269), .B(n5270), .Z(n5261) );
  AND U5240 ( .A(n5271), .B(n5272), .Z(n5270) );
  XNOR U5241 ( .A(n5269), .B(n5265), .Z(n5272) );
  IV U5242 ( .A(n5219), .Z(n5265) );
  XOR U5243 ( .A(n5273), .B(n5274), .Z(n5219) );
  XOR U5244 ( .A(n5275), .B(n5266), .Z(n5274) );
  AND U5245 ( .A(n5231), .B(n5276), .Z(n5266) );
  AND U5246 ( .A(n5277), .B(n5278), .Z(n5275) );
  XOR U5247 ( .A(n5279), .B(n5273), .Z(n5277) );
  XNOR U5248 ( .A(n5216), .B(n5269), .Z(n5271) );
  XNOR U5249 ( .A(n5280), .B(n5281), .Z(n5216) );
  AND U5250 ( .A(n122), .B(n5223), .Z(n5281) );
  XOR U5251 ( .A(n5280), .B(n5221), .Z(n5223) );
  XOR U5252 ( .A(n5282), .B(n5283), .Z(n5269) );
  AND U5253 ( .A(n5284), .B(n5285), .Z(n5283) );
  XNOR U5254 ( .A(n5282), .B(n5231), .Z(n5285) );
  XOR U5255 ( .A(n5286), .B(n5278), .Z(n5231) );
  XNOR U5256 ( .A(n5287), .B(n5273), .Z(n5278) );
  XOR U5257 ( .A(n5288), .B(n5289), .Z(n5273) );
  AND U5258 ( .A(n5290), .B(n5291), .Z(n5289) );
  XOR U5259 ( .A(n5292), .B(n5288), .Z(n5290) );
  XNOR U5260 ( .A(n5293), .B(n5294), .Z(n5287) );
  AND U5261 ( .A(n5295), .B(n5296), .Z(n5294) );
  XOR U5262 ( .A(n5293), .B(n5297), .Z(n5295) );
  XNOR U5263 ( .A(n5279), .B(n5276), .Z(n5286) );
  AND U5264 ( .A(n5298), .B(n5299), .Z(n5276) );
  XOR U5265 ( .A(n5300), .B(n5301), .Z(n5279) );
  AND U5266 ( .A(n5302), .B(n5303), .Z(n5301) );
  XOR U5267 ( .A(n5300), .B(n5304), .Z(n5302) );
  XNOR U5268 ( .A(n5228), .B(n5282), .Z(n5284) );
  XNOR U5269 ( .A(n5305), .B(n5306), .Z(n5228) );
  AND U5270 ( .A(n122), .B(n5234), .Z(n5306) );
  XOR U5271 ( .A(n5305), .B(n5232), .Z(n5234) );
  XOR U5272 ( .A(n5307), .B(n5308), .Z(n5282) );
  AND U5273 ( .A(n5309), .B(n5310), .Z(n5308) );
  XNOR U5274 ( .A(n5307), .B(n5298), .Z(n5310) );
  IV U5275 ( .A(n5240), .Z(n5298) );
  XNOR U5276 ( .A(n5311), .B(n5291), .Z(n5240) );
  XNOR U5277 ( .A(n5312), .B(n5297), .Z(n5291) );
  XOR U5278 ( .A(n5313), .B(n5314), .Z(n5297) );
  AND U5279 ( .A(n5315), .B(n5316), .Z(n5314) );
  XOR U5280 ( .A(n5313), .B(n5317), .Z(n5315) );
  XNOR U5281 ( .A(n5296), .B(n5288), .Z(n5312) );
  XOR U5282 ( .A(n5318), .B(n5319), .Z(n5288) );
  AND U5283 ( .A(n5320), .B(n5321), .Z(n5319) );
  XNOR U5284 ( .A(n5322), .B(n5318), .Z(n5320) );
  XNOR U5285 ( .A(n5323), .B(n5293), .Z(n5296) );
  XOR U5286 ( .A(n5324), .B(n5325), .Z(n5293) );
  AND U5287 ( .A(n5326), .B(n5327), .Z(n5325) );
  XOR U5288 ( .A(n5324), .B(n5328), .Z(n5326) );
  XNOR U5289 ( .A(n5329), .B(n5330), .Z(n5323) );
  AND U5290 ( .A(n5331), .B(n5332), .Z(n5330) );
  XNOR U5291 ( .A(n5329), .B(n5333), .Z(n5331) );
  XNOR U5292 ( .A(n5292), .B(n5299), .Z(n5311) );
  AND U5293 ( .A(n5252), .B(n5334), .Z(n5299) );
  XOR U5294 ( .A(n5304), .B(n5303), .Z(n5292) );
  XNOR U5295 ( .A(n5335), .B(n5300), .Z(n5303) );
  XOR U5296 ( .A(n5336), .B(n5337), .Z(n5300) );
  AND U5297 ( .A(n5338), .B(n5339), .Z(n5337) );
  XOR U5298 ( .A(n5336), .B(n5340), .Z(n5338) );
  XNOR U5299 ( .A(n5341), .B(n5342), .Z(n5335) );
  AND U5300 ( .A(n5343), .B(n5344), .Z(n5342) );
  XOR U5301 ( .A(n5341), .B(n5345), .Z(n5343) );
  XOR U5302 ( .A(n5346), .B(n5347), .Z(n5304) );
  AND U5303 ( .A(n5348), .B(n5349), .Z(n5347) );
  XOR U5304 ( .A(n5346), .B(n5350), .Z(n5348) );
  XNOR U5305 ( .A(n5237), .B(n5307), .Z(n5309) );
  XNOR U5306 ( .A(n5351), .B(n5352), .Z(n5237) );
  AND U5307 ( .A(n122), .B(n5244), .Z(n5352) );
  XOR U5308 ( .A(n5351), .B(n5242), .Z(n5244) );
  XOR U5309 ( .A(n5353), .B(n5354), .Z(n5307) );
  AND U5310 ( .A(n5355), .B(n5356), .Z(n5354) );
  XNOR U5311 ( .A(n5353), .B(n5252), .Z(n5356) );
  XOR U5312 ( .A(n5357), .B(n5321), .Z(n5252) );
  XNOR U5313 ( .A(n5358), .B(n5328), .Z(n5321) );
  XOR U5314 ( .A(n5317), .B(n5316), .Z(n5328) );
  XNOR U5315 ( .A(n5359), .B(n5313), .Z(n5316) );
  XOR U5316 ( .A(n5360), .B(n5361), .Z(n5313) );
  AND U5317 ( .A(n5362), .B(n5363), .Z(n5361) );
  XNOR U5318 ( .A(n5364), .B(n5365), .Z(n5362) );
  IV U5319 ( .A(n5360), .Z(n5364) );
  XNOR U5320 ( .A(n5366), .B(n5367), .Z(n5359) );
  NOR U5321 ( .A(n5368), .B(n5369), .Z(n5367) );
  XNOR U5322 ( .A(n5366), .B(n5370), .Z(n5368) );
  XOR U5323 ( .A(n5371), .B(n5372), .Z(n5317) );
  NOR U5324 ( .A(n5373), .B(n5374), .Z(n5372) );
  XNOR U5325 ( .A(n5371), .B(n5375), .Z(n5373) );
  XNOR U5326 ( .A(n5327), .B(n5318), .Z(n5358) );
  XOR U5327 ( .A(n5376), .B(n5377), .Z(n5318) );
  AND U5328 ( .A(n5378), .B(n5379), .Z(n5377) );
  XOR U5329 ( .A(n5376), .B(n5380), .Z(n5378) );
  XOR U5330 ( .A(n5381), .B(n5333), .Z(n5327) );
  XOR U5331 ( .A(n5382), .B(n5383), .Z(n5333) );
  NOR U5332 ( .A(n5384), .B(n5385), .Z(n5383) );
  XOR U5333 ( .A(n5382), .B(n5386), .Z(n5384) );
  XNOR U5334 ( .A(n5332), .B(n5324), .Z(n5381) );
  XOR U5335 ( .A(n5387), .B(n5388), .Z(n5324) );
  AND U5336 ( .A(n5389), .B(n5390), .Z(n5388) );
  XOR U5337 ( .A(n5387), .B(n5391), .Z(n5389) );
  XNOR U5338 ( .A(n5392), .B(n5329), .Z(n5332) );
  XOR U5339 ( .A(n5393), .B(n5394), .Z(n5329) );
  AND U5340 ( .A(n5395), .B(n5396), .Z(n5394) );
  XNOR U5341 ( .A(n5397), .B(n5398), .Z(n5395) );
  IV U5342 ( .A(n5393), .Z(n5397) );
  XNOR U5343 ( .A(n5399), .B(n5400), .Z(n5392) );
  NOR U5344 ( .A(n5401), .B(n5402), .Z(n5400) );
  XNOR U5345 ( .A(n5399), .B(n5403), .Z(n5401) );
  XOR U5346 ( .A(n5322), .B(n5334), .Z(n5357) );
  NOR U5347 ( .A(n5260), .B(n5404), .Z(n5334) );
  XNOR U5348 ( .A(n5340), .B(n5339), .Z(n5322) );
  XNOR U5349 ( .A(n5405), .B(n5345), .Z(n5339) );
  XNOR U5350 ( .A(n5406), .B(n5407), .Z(n5345) );
  NOR U5351 ( .A(n5408), .B(n5409), .Z(n5407) );
  XOR U5352 ( .A(n5406), .B(n5410), .Z(n5408) );
  XNOR U5353 ( .A(n5344), .B(n5336), .Z(n5405) );
  XOR U5354 ( .A(n5411), .B(n5412), .Z(n5336) );
  AND U5355 ( .A(n5413), .B(n5414), .Z(n5412) );
  XOR U5356 ( .A(n5411), .B(n5415), .Z(n5413) );
  XNOR U5357 ( .A(n5416), .B(n5341), .Z(n5344) );
  XOR U5358 ( .A(n5417), .B(n5418), .Z(n5341) );
  AND U5359 ( .A(n5419), .B(n5420), .Z(n5418) );
  XNOR U5360 ( .A(n5421), .B(n5422), .Z(n5419) );
  IV U5361 ( .A(n5417), .Z(n5421) );
  XNOR U5362 ( .A(n5423), .B(n5424), .Z(n5416) );
  NOR U5363 ( .A(n5425), .B(n5426), .Z(n5424) );
  XNOR U5364 ( .A(n5423), .B(n5427), .Z(n5425) );
  XOR U5365 ( .A(n5350), .B(n5349), .Z(n5340) );
  XNOR U5366 ( .A(n5428), .B(n5346), .Z(n5349) );
  XOR U5367 ( .A(n5429), .B(n5430), .Z(n5346) );
  AND U5368 ( .A(n5431), .B(n5432), .Z(n5430) );
  XNOR U5369 ( .A(n5433), .B(n5434), .Z(n5431) );
  IV U5370 ( .A(n5429), .Z(n5433) );
  XNOR U5371 ( .A(n5435), .B(n5436), .Z(n5428) );
  NOR U5372 ( .A(n5437), .B(n5438), .Z(n5436) );
  XNOR U5373 ( .A(n5435), .B(n5439), .Z(n5437) );
  XOR U5374 ( .A(n5440), .B(n5441), .Z(n5350) );
  NOR U5375 ( .A(n5442), .B(n5443), .Z(n5441) );
  XNOR U5376 ( .A(n5440), .B(n5444), .Z(n5442) );
  XNOR U5377 ( .A(n5249), .B(n5353), .Z(n5355) );
  XNOR U5378 ( .A(n5445), .B(n5446), .Z(n5249) );
  AND U5379 ( .A(n122), .B(n5256), .Z(n5446) );
  XOR U5380 ( .A(n5445), .B(n5254), .Z(n5256) );
  AND U5381 ( .A(n5257), .B(n5260), .Z(n5353) );
  XOR U5382 ( .A(n5447), .B(n5404), .Z(n5260) );
  XNOR U5383 ( .A(p_input[160]), .B(p_input[512]), .Z(n5404) );
  XNOR U5384 ( .A(n5380), .B(n5379), .Z(n5447) );
  XNOR U5385 ( .A(n5448), .B(n5391), .Z(n5379) );
  XOR U5386 ( .A(n5365), .B(n5363), .Z(n5391) );
  XNOR U5387 ( .A(n5449), .B(n5370), .Z(n5363) );
  XOR U5388 ( .A(p_input[184]), .B(p_input[536]), .Z(n5370) );
  XOR U5389 ( .A(n5360), .B(n5369), .Z(n5449) );
  XOR U5390 ( .A(n5450), .B(n5366), .Z(n5369) );
  XOR U5391 ( .A(p_input[182]), .B(p_input[534]), .Z(n5366) );
  XOR U5392 ( .A(p_input[183]), .B(n4010), .Z(n5450) );
  XOR U5393 ( .A(p_input[178]), .B(p_input[530]), .Z(n5360) );
  XNOR U5394 ( .A(n5375), .B(n5374), .Z(n5365) );
  XOR U5395 ( .A(n5451), .B(n5371), .Z(n5374) );
  XOR U5396 ( .A(p_input[179]), .B(p_input[531]), .Z(n5371) );
  XOR U5397 ( .A(p_input[180]), .B(n4012), .Z(n5451) );
  XOR U5398 ( .A(p_input[181]), .B(p_input[533]), .Z(n5375) );
  XOR U5399 ( .A(n5390), .B(n5452), .Z(n5448) );
  IV U5400 ( .A(n5376), .Z(n5452) );
  XOR U5401 ( .A(p_input[161]), .B(p_input[513]), .Z(n5376) );
  XNOR U5402 ( .A(n5453), .B(n5398), .Z(n5390) );
  XNOR U5403 ( .A(n5386), .B(n5385), .Z(n5398) );
  XNOR U5404 ( .A(n5454), .B(n5382), .Z(n5385) );
  XNOR U5405 ( .A(p_input[186]), .B(p_input[538]), .Z(n5382) );
  XOR U5406 ( .A(p_input[187]), .B(n4016), .Z(n5454) );
  XOR U5407 ( .A(p_input[188]), .B(p_input[540]), .Z(n5386) );
  XOR U5408 ( .A(n5396), .B(n5455), .Z(n5453) );
  IV U5409 ( .A(n5387), .Z(n5455) );
  XOR U5410 ( .A(p_input[177]), .B(p_input[529]), .Z(n5387) );
  XNOR U5411 ( .A(n5456), .B(n5403), .Z(n5396) );
  XNOR U5412 ( .A(p_input[191]), .B(n4019), .Z(n5403) );
  XOR U5413 ( .A(n5393), .B(n5402), .Z(n5456) );
  XOR U5414 ( .A(n5457), .B(n5399), .Z(n5402) );
  XOR U5415 ( .A(p_input[189]), .B(p_input[541]), .Z(n5399) );
  XOR U5416 ( .A(p_input[190]), .B(n4021), .Z(n5457) );
  XOR U5417 ( .A(p_input[185]), .B(p_input[537]), .Z(n5393) );
  XOR U5418 ( .A(n5415), .B(n5414), .Z(n5380) );
  XNOR U5419 ( .A(n5458), .B(n5422), .Z(n5414) );
  XNOR U5420 ( .A(n5410), .B(n5409), .Z(n5422) );
  XNOR U5421 ( .A(n5459), .B(n5406), .Z(n5409) );
  XNOR U5422 ( .A(p_input[171]), .B(p_input[523]), .Z(n5406) );
  XOR U5423 ( .A(p_input[172]), .B(n4024), .Z(n5459) );
  XOR U5424 ( .A(p_input[173]), .B(p_input[525]), .Z(n5410) );
  XOR U5425 ( .A(n5420), .B(n5460), .Z(n5458) );
  IV U5426 ( .A(n5411), .Z(n5460) );
  XOR U5427 ( .A(p_input[162]), .B(p_input[514]), .Z(n5411) );
  XNOR U5428 ( .A(n5461), .B(n5427), .Z(n5420) );
  XNOR U5429 ( .A(p_input[176]), .B(n4027), .Z(n5427) );
  XOR U5430 ( .A(n5417), .B(n5426), .Z(n5461) );
  XOR U5431 ( .A(n5462), .B(n5423), .Z(n5426) );
  XOR U5432 ( .A(p_input[174]), .B(p_input[526]), .Z(n5423) );
  XOR U5433 ( .A(p_input[175]), .B(n4029), .Z(n5462) );
  XOR U5434 ( .A(p_input[170]), .B(p_input[522]), .Z(n5417) );
  XOR U5435 ( .A(n5434), .B(n5432), .Z(n5415) );
  XNOR U5436 ( .A(n5463), .B(n5439), .Z(n5432) );
  XOR U5437 ( .A(p_input[169]), .B(p_input[521]), .Z(n5439) );
  XOR U5438 ( .A(n5429), .B(n5438), .Z(n5463) );
  XOR U5439 ( .A(n5464), .B(n5435), .Z(n5438) );
  XOR U5440 ( .A(p_input[167]), .B(p_input[519]), .Z(n5435) );
  XOR U5441 ( .A(p_input[168]), .B(n4318), .Z(n5464) );
  XOR U5442 ( .A(p_input[163]), .B(p_input[515]), .Z(n5429) );
  XNOR U5443 ( .A(n5444), .B(n5443), .Z(n5434) );
  XOR U5444 ( .A(n5465), .B(n5440), .Z(n5443) );
  XOR U5445 ( .A(p_input[164]), .B(p_input[516]), .Z(n5440) );
  XOR U5446 ( .A(p_input[165]), .B(n4320), .Z(n5465) );
  XOR U5447 ( .A(p_input[166]), .B(p_input[518]), .Z(n5444) );
  XNOR U5448 ( .A(n5466), .B(n5467), .Z(n5257) );
  AND U5449 ( .A(n122), .B(n5468), .Z(n5467) );
  XNOR U5450 ( .A(n5469), .B(n5470), .Z(n122) );
  AND U5451 ( .A(n5471), .B(n5472), .Z(n5470) );
  XOR U5452 ( .A(n5469), .B(n5267), .Z(n5472) );
  XNOR U5453 ( .A(n5469), .B(n5209), .Z(n5471) );
  XOR U5454 ( .A(n5473), .B(n5474), .Z(n5469) );
  AND U5455 ( .A(n5475), .B(n5476), .Z(n5474) );
  XNOR U5456 ( .A(n5280), .B(n5473), .Z(n5476) );
  XOR U5457 ( .A(n5473), .B(n5221), .Z(n5475) );
  XOR U5458 ( .A(n5477), .B(n5478), .Z(n5473) );
  AND U5459 ( .A(n5479), .B(n5480), .Z(n5478) );
  XNOR U5460 ( .A(n5305), .B(n5477), .Z(n5480) );
  XOR U5461 ( .A(n5477), .B(n5232), .Z(n5479) );
  XOR U5462 ( .A(n5481), .B(n5482), .Z(n5477) );
  AND U5463 ( .A(n5483), .B(n5484), .Z(n5482) );
  XOR U5464 ( .A(n5481), .B(n5242), .Z(n5483) );
  XOR U5465 ( .A(n5485), .B(n5486), .Z(n5198) );
  AND U5466 ( .A(n126), .B(n5468), .Z(n5486) );
  XNOR U5467 ( .A(n5466), .B(n5485), .Z(n5468) );
  XNOR U5468 ( .A(n5487), .B(n5488), .Z(n126) );
  AND U5469 ( .A(n5489), .B(n5490), .Z(n5488) );
  XNOR U5470 ( .A(n5491), .B(n5487), .Z(n5490) );
  IV U5471 ( .A(n5267), .Z(n5491) );
  XNOR U5472 ( .A(n5492), .B(n5493), .Z(n5267) );
  AND U5473 ( .A(n129), .B(n5494), .Z(n5493) );
  XNOR U5474 ( .A(n5492), .B(n5495), .Z(n5494) );
  XNOR U5475 ( .A(n5209), .B(n5487), .Z(n5489) );
  XOR U5476 ( .A(n5496), .B(n5497), .Z(n5209) );
  AND U5477 ( .A(n137), .B(n5498), .Z(n5497) );
  XOR U5478 ( .A(n5499), .B(n5500), .Z(n5487) );
  AND U5479 ( .A(n5501), .B(n5502), .Z(n5500) );
  XNOR U5480 ( .A(n5499), .B(n5280), .Z(n5502) );
  XNOR U5481 ( .A(n5503), .B(n5504), .Z(n5280) );
  AND U5482 ( .A(n129), .B(n5505), .Z(n5504) );
  XOR U5483 ( .A(n5506), .B(n5503), .Z(n5505) );
  XNOR U5484 ( .A(n5507), .B(n5499), .Z(n5501) );
  IV U5485 ( .A(n5221), .Z(n5507) );
  XOR U5486 ( .A(n5508), .B(n5509), .Z(n5221) );
  AND U5487 ( .A(n137), .B(n5510), .Z(n5509) );
  XOR U5488 ( .A(n5511), .B(n5512), .Z(n5499) );
  AND U5489 ( .A(n5513), .B(n5514), .Z(n5512) );
  XNOR U5490 ( .A(n5511), .B(n5305), .Z(n5514) );
  XNOR U5491 ( .A(n5515), .B(n5516), .Z(n5305) );
  AND U5492 ( .A(n129), .B(n5517), .Z(n5516) );
  XNOR U5493 ( .A(n5518), .B(n5515), .Z(n5517) );
  XOR U5494 ( .A(n5232), .B(n5511), .Z(n5513) );
  XOR U5495 ( .A(n5519), .B(n5520), .Z(n5232) );
  AND U5496 ( .A(n137), .B(n5521), .Z(n5520) );
  XOR U5497 ( .A(n5481), .B(n5522), .Z(n5511) );
  AND U5498 ( .A(n5523), .B(n5484), .Z(n5522) );
  XNOR U5499 ( .A(n5351), .B(n5481), .Z(n5484) );
  XNOR U5500 ( .A(n5524), .B(n5525), .Z(n5351) );
  AND U5501 ( .A(n129), .B(n5526), .Z(n5525) );
  XOR U5502 ( .A(n5527), .B(n5524), .Z(n5526) );
  XNOR U5503 ( .A(n5528), .B(n5481), .Z(n5523) );
  IV U5504 ( .A(n5242), .Z(n5528) );
  XOR U5505 ( .A(n5529), .B(n5530), .Z(n5242) );
  AND U5506 ( .A(n137), .B(n5531), .Z(n5530) );
  XOR U5507 ( .A(n5532), .B(n5533), .Z(n5481) );
  AND U5508 ( .A(n5534), .B(n5535), .Z(n5533) );
  XNOR U5509 ( .A(n5532), .B(n5445), .Z(n5535) );
  XNOR U5510 ( .A(n5536), .B(n5537), .Z(n5445) );
  AND U5511 ( .A(n129), .B(n5538), .Z(n5537) );
  XNOR U5512 ( .A(n5539), .B(n5536), .Z(n5538) );
  XNOR U5513 ( .A(n5540), .B(n5532), .Z(n5534) );
  IV U5514 ( .A(n5254), .Z(n5540) );
  XOR U5515 ( .A(n5541), .B(n5542), .Z(n5254) );
  AND U5516 ( .A(n137), .B(n5543), .Z(n5542) );
  AND U5517 ( .A(n5485), .B(n5466), .Z(n5532) );
  XNOR U5518 ( .A(n5544), .B(n5545), .Z(n5466) );
  AND U5519 ( .A(n129), .B(n5546), .Z(n5545) );
  XNOR U5520 ( .A(n5547), .B(n5544), .Z(n5546) );
  XNOR U5521 ( .A(n5548), .B(n5549), .Z(n129) );
  AND U5522 ( .A(n5550), .B(n5551), .Z(n5549) );
  XOR U5523 ( .A(n5495), .B(n5548), .Z(n5551) );
  AND U5524 ( .A(n5552), .B(n5553), .Z(n5495) );
  XOR U5525 ( .A(n5548), .B(n5492), .Z(n5550) );
  XNOR U5526 ( .A(n5554), .B(n5555), .Z(n5492) );
  AND U5527 ( .A(n133), .B(n5498), .Z(n5555) );
  XOR U5528 ( .A(n5496), .B(n5554), .Z(n5498) );
  XOR U5529 ( .A(n5556), .B(n5557), .Z(n5548) );
  AND U5530 ( .A(n5558), .B(n5559), .Z(n5557) );
  XNOR U5531 ( .A(n5556), .B(n5552), .Z(n5559) );
  IV U5532 ( .A(n5506), .Z(n5552) );
  XOR U5533 ( .A(n5560), .B(n5561), .Z(n5506) );
  XOR U5534 ( .A(n5562), .B(n5553), .Z(n5561) );
  AND U5535 ( .A(n5518), .B(n5563), .Z(n5553) );
  AND U5536 ( .A(n5564), .B(n5565), .Z(n5562) );
  XOR U5537 ( .A(n5566), .B(n5560), .Z(n5564) );
  XNOR U5538 ( .A(n5503), .B(n5556), .Z(n5558) );
  XNOR U5539 ( .A(n5567), .B(n5568), .Z(n5503) );
  AND U5540 ( .A(n133), .B(n5510), .Z(n5568) );
  XOR U5541 ( .A(n5567), .B(n5508), .Z(n5510) );
  XOR U5542 ( .A(n5569), .B(n5570), .Z(n5556) );
  AND U5543 ( .A(n5571), .B(n5572), .Z(n5570) );
  XNOR U5544 ( .A(n5569), .B(n5518), .Z(n5572) );
  XOR U5545 ( .A(n5573), .B(n5565), .Z(n5518) );
  XNOR U5546 ( .A(n5574), .B(n5560), .Z(n5565) );
  XOR U5547 ( .A(n5575), .B(n5576), .Z(n5560) );
  AND U5548 ( .A(n5577), .B(n5578), .Z(n5576) );
  XOR U5549 ( .A(n5579), .B(n5575), .Z(n5577) );
  XNOR U5550 ( .A(n5580), .B(n5581), .Z(n5574) );
  AND U5551 ( .A(n5582), .B(n5583), .Z(n5581) );
  XOR U5552 ( .A(n5580), .B(n5584), .Z(n5582) );
  XNOR U5553 ( .A(n5566), .B(n5563), .Z(n5573) );
  AND U5554 ( .A(n5585), .B(n5586), .Z(n5563) );
  XOR U5555 ( .A(n5587), .B(n5588), .Z(n5566) );
  AND U5556 ( .A(n5589), .B(n5590), .Z(n5588) );
  XOR U5557 ( .A(n5587), .B(n5591), .Z(n5589) );
  XNOR U5558 ( .A(n5515), .B(n5569), .Z(n5571) );
  XNOR U5559 ( .A(n5592), .B(n5593), .Z(n5515) );
  AND U5560 ( .A(n133), .B(n5521), .Z(n5593) );
  XOR U5561 ( .A(n5592), .B(n5519), .Z(n5521) );
  XOR U5562 ( .A(n5594), .B(n5595), .Z(n5569) );
  AND U5563 ( .A(n5596), .B(n5597), .Z(n5595) );
  XNOR U5564 ( .A(n5594), .B(n5585), .Z(n5597) );
  IV U5565 ( .A(n5527), .Z(n5585) );
  XNOR U5566 ( .A(n5598), .B(n5578), .Z(n5527) );
  XNOR U5567 ( .A(n5599), .B(n5584), .Z(n5578) );
  XOR U5568 ( .A(n5600), .B(n5601), .Z(n5584) );
  AND U5569 ( .A(n5602), .B(n5603), .Z(n5601) );
  XOR U5570 ( .A(n5600), .B(n5604), .Z(n5602) );
  XNOR U5571 ( .A(n5583), .B(n5575), .Z(n5599) );
  XOR U5572 ( .A(n5605), .B(n5606), .Z(n5575) );
  AND U5573 ( .A(n5607), .B(n5608), .Z(n5606) );
  XNOR U5574 ( .A(n5609), .B(n5605), .Z(n5607) );
  XNOR U5575 ( .A(n5610), .B(n5580), .Z(n5583) );
  XOR U5576 ( .A(n5611), .B(n5612), .Z(n5580) );
  AND U5577 ( .A(n5613), .B(n5614), .Z(n5612) );
  XOR U5578 ( .A(n5611), .B(n5615), .Z(n5613) );
  XNOR U5579 ( .A(n5616), .B(n5617), .Z(n5610) );
  AND U5580 ( .A(n5618), .B(n5619), .Z(n5617) );
  XNOR U5581 ( .A(n5616), .B(n5620), .Z(n5618) );
  XNOR U5582 ( .A(n5579), .B(n5586), .Z(n5598) );
  AND U5583 ( .A(n5539), .B(n5621), .Z(n5586) );
  XOR U5584 ( .A(n5591), .B(n5590), .Z(n5579) );
  XNOR U5585 ( .A(n5622), .B(n5587), .Z(n5590) );
  XOR U5586 ( .A(n5623), .B(n5624), .Z(n5587) );
  AND U5587 ( .A(n5625), .B(n5626), .Z(n5624) );
  XOR U5588 ( .A(n5623), .B(n5627), .Z(n5625) );
  XNOR U5589 ( .A(n5628), .B(n5629), .Z(n5622) );
  AND U5590 ( .A(n5630), .B(n5631), .Z(n5629) );
  XOR U5591 ( .A(n5628), .B(n5632), .Z(n5630) );
  XOR U5592 ( .A(n5633), .B(n5634), .Z(n5591) );
  AND U5593 ( .A(n5635), .B(n5636), .Z(n5634) );
  XOR U5594 ( .A(n5633), .B(n5637), .Z(n5635) );
  XNOR U5595 ( .A(n5524), .B(n5594), .Z(n5596) );
  XNOR U5596 ( .A(n5638), .B(n5639), .Z(n5524) );
  AND U5597 ( .A(n133), .B(n5531), .Z(n5639) );
  XOR U5598 ( .A(n5638), .B(n5529), .Z(n5531) );
  XOR U5599 ( .A(n5640), .B(n5641), .Z(n5594) );
  AND U5600 ( .A(n5642), .B(n5643), .Z(n5641) );
  XNOR U5601 ( .A(n5640), .B(n5539), .Z(n5643) );
  XOR U5602 ( .A(n5644), .B(n5608), .Z(n5539) );
  XNOR U5603 ( .A(n5645), .B(n5615), .Z(n5608) );
  XOR U5604 ( .A(n5604), .B(n5603), .Z(n5615) );
  XNOR U5605 ( .A(n5646), .B(n5600), .Z(n5603) );
  XOR U5606 ( .A(n5647), .B(n5648), .Z(n5600) );
  AND U5607 ( .A(n5649), .B(n5650), .Z(n5648) );
  XNOR U5608 ( .A(n5651), .B(n5652), .Z(n5649) );
  IV U5609 ( .A(n5647), .Z(n5651) );
  XNOR U5610 ( .A(n5653), .B(n5654), .Z(n5646) );
  NOR U5611 ( .A(n5655), .B(n5656), .Z(n5654) );
  XNOR U5612 ( .A(n5653), .B(n5657), .Z(n5655) );
  XOR U5613 ( .A(n5658), .B(n5659), .Z(n5604) );
  NOR U5614 ( .A(n5660), .B(n5661), .Z(n5659) );
  XNOR U5615 ( .A(n5658), .B(n5662), .Z(n5660) );
  XNOR U5616 ( .A(n5614), .B(n5605), .Z(n5645) );
  XOR U5617 ( .A(n5663), .B(n5664), .Z(n5605) );
  AND U5618 ( .A(n5665), .B(n5666), .Z(n5664) );
  XOR U5619 ( .A(n5663), .B(n5667), .Z(n5665) );
  XOR U5620 ( .A(n5668), .B(n5620), .Z(n5614) );
  XOR U5621 ( .A(n5669), .B(n5670), .Z(n5620) );
  NOR U5622 ( .A(n5671), .B(n5672), .Z(n5670) );
  XOR U5623 ( .A(n5669), .B(n5673), .Z(n5671) );
  XNOR U5624 ( .A(n5619), .B(n5611), .Z(n5668) );
  XOR U5625 ( .A(n5674), .B(n5675), .Z(n5611) );
  AND U5626 ( .A(n5676), .B(n5677), .Z(n5675) );
  XOR U5627 ( .A(n5674), .B(n5678), .Z(n5676) );
  XNOR U5628 ( .A(n5679), .B(n5616), .Z(n5619) );
  XOR U5629 ( .A(n5680), .B(n5681), .Z(n5616) );
  AND U5630 ( .A(n5682), .B(n5683), .Z(n5681) );
  XNOR U5631 ( .A(n5684), .B(n5685), .Z(n5682) );
  IV U5632 ( .A(n5680), .Z(n5684) );
  XNOR U5633 ( .A(n5686), .B(n5687), .Z(n5679) );
  NOR U5634 ( .A(n5688), .B(n5689), .Z(n5687) );
  XNOR U5635 ( .A(n5686), .B(n5690), .Z(n5688) );
  XOR U5636 ( .A(n5609), .B(n5621), .Z(n5644) );
  NOR U5637 ( .A(n5547), .B(n5691), .Z(n5621) );
  XNOR U5638 ( .A(n5627), .B(n5626), .Z(n5609) );
  XNOR U5639 ( .A(n5692), .B(n5632), .Z(n5626) );
  XNOR U5640 ( .A(n5693), .B(n5694), .Z(n5632) );
  NOR U5641 ( .A(n5695), .B(n5696), .Z(n5694) );
  XOR U5642 ( .A(n5693), .B(n5697), .Z(n5695) );
  XNOR U5643 ( .A(n5631), .B(n5623), .Z(n5692) );
  XOR U5644 ( .A(n5698), .B(n5699), .Z(n5623) );
  AND U5645 ( .A(n5700), .B(n5701), .Z(n5699) );
  XOR U5646 ( .A(n5698), .B(n5702), .Z(n5700) );
  XNOR U5647 ( .A(n5703), .B(n5628), .Z(n5631) );
  XOR U5648 ( .A(n5704), .B(n5705), .Z(n5628) );
  AND U5649 ( .A(n5706), .B(n5707), .Z(n5705) );
  XNOR U5650 ( .A(n5708), .B(n5709), .Z(n5706) );
  IV U5651 ( .A(n5704), .Z(n5708) );
  XNOR U5652 ( .A(n5710), .B(n5711), .Z(n5703) );
  NOR U5653 ( .A(n5712), .B(n5713), .Z(n5711) );
  XNOR U5654 ( .A(n5710), .B(n5714), .Z(n5712) );
  XOR U5655 ( .A(n5637), .B(n5636), .Z(n5627) );
  XNOR U5656 ( .A(n5715), .B(n5633), .Z(n5636) );
  XOR U5657 ( .A(n5716), .B(n5717), .Z(n5633) );
  AND U5658 ( .A(n5718), .B(n5719), .Z(n5717) );
  XNOR U5659 ( .A(n5720), .B(n5721), .Z(n5718) );
  IV U5660 ( .A(n5716), .Z(n5720) );
  XNOR U5661 ( .A(n5722), .B(n5723), .Z(n5715) );
  NOR U5662 ( .A(n5724), .B(n5725), .Z(n5723) );
  XNOR U5663 ( .A(n5722), .B(n5726), .Z(n5724) );
  XOR U5664 ( .A(n5727), .B(n5728), .Z(n5637) );
  NOR U5665 ( .A(n5729), .B(n5730), .Z(n5728) );
  XNOR U5666 ( .A(n5727), .B(n5731), .Z(n5729) );
  XNOR U5667 ( .A(n5536), .B(n5640), .Z(n5642) );
  XNOR U5668 ( .A(n5732), .B(n5733), .Z(n5536) );
  AND U5669 ( .A(n133), .B(n5543), .Z(n5733) );
  XOR U5670 ( .A(n5732), .B(n5541), .Z(n5543) );
  AND U5671 ( .A(n5544), .B(n5547), .Z(n5640) );
  XOR U5672 ( .A(n5734), .B(n5691), .Z(n5547) );
  XNOR U5673 ( .A(p_input[192]), .B(p_input[512]), .Z(n5691) );
  XNOR U5674 ( .A(n5667), .B(n5666), .Z(n5734) );
  XNOR U5675 ( .A(n5735), .B(n5678), .Z(n5666) );
  XOR U5676 ( .A(n5652), .B(n5650), .Z(n5678) );
  XNOR U5677 ( .A(n5736), .B(n5657), .Z(n5650) );
  XOR U5678 ( .A(p_input[216]), .B(p_input[536]), .Z(n5657) );
  XOR U5679 ( .A(n5647), .B(n5656), .Z(n5736) );
  XOR U5680 ( .A(n5737), .B(n5653), .Z(n5656) );
  XOR U5681 ( .A(p_input[214]), .B(p_input[534]), .Z(n5653) );
  XOR U5682 ( .A(p_input[215]), .B(n4010), .Z(n5737) );
  XOR U5683 ( .A(p_input[210]), .B(p_input[530]), .Z(n5647) );
  XNOR U5684 ( .A(n5662), .B(n5661), .Z(n5652) );
  XOR U5685 ( .A(n5738), .B(n5658), .Z(n5661) );
  XOR U5686 ( .A(p_input[211]), .B(p_input[531]), .Z(n5658) );
  XOR U5687 ( .A(p_input[212]), .B(n4012), .Z(n5738) );
  XOR U5688 ( .A(p_input[213]), .B(p_input[533]), .Z(n5662) );
  XOR U5689 ( .A(n5677), .B(n5739), .Z(n5735) );
  IV U5690 ( .A(n5663), .Z(n5739) );
  XOR U5691 ( .A(p_input[193]), .B(p_input[513]), .Z(n5663) );
  XNOR U5692 ( .A(n5740), .B(n5685), .Z(n5677) );
  XNOR U5693 ( .A(n5673), .B(n5672), .Z(n5685) );
  XNOR U5694 ( .A(n5741), .B(n5669), .Z(n5672) );
  XNOR U5695 ( .A(p_input[218]), .B(p_input[538]), .Z(n5669) );
  XOR U5696 ( .A(p_input[219]), .B(n4016), .Z(n5741) );
  XOR U5697 ( .A(p_input[220]), .B(p_input[540]), .Z(n5673) );
  XOR U5698 ( .A(n5683), .B(n5742), .Z(n5740) );
  IV U5699 ( .A(n5674), .Z(n5742) );
  XOR U5700 ( .A(p_input[209]), .B(p_input[529]), .Z(n5674) );
  XNOR U5701 ( .A(n5743), .B(n5690), .Z(n5683) );
  XNOR U5702 ( .A(p_input[223]), .B(n4019), .Z(n5690) );
  XOR U5703 ( .A(n5680), .B(n5689), .Z(n5743) );
  XOR U5704 ( .A(n5744), .B(n5686), .Z(n5689) );
  XOR U5705 ( .A(p_input[221]), .B(p_input[541]), .Z(n5686) );
  XOR U5706 ( .A(p_input[222]), .B(n4021), .Z(n5744) );
  XOR U5707 ( .A(p_input[217]), .B(p_input[537]), .Z(n5680) );
  XOR U5708 ( .A(n5702), .B(n5701), .Z(n5667) );
  XNOR U5709 ( .A(n5745), .B(n5709), .Z(n5701) );
  XNOR U5710 ( .A(n5697), .B(n5696), .Z(n5709) );
  XNOR U5711 ( .A(n5746), .B(n5693), .Z(n5696) );
  XNOR U5712 ( .A(p_input[203]), .B(p_input[523]), .Z(n5693) );
  XOR U5713 ( .A(p_input[204]), .B(n4024), .Z(n5746) );
  XOR U5714 ( .A(p_input[205]), .B(p_input[525]), .Z(n5697) );
  XOR U5715 ( .A(n5707), .B(n5747), .Z(n5745) );
  IV U5716 ( .A(n5698), .Z(n5747) );
  XOR U5717 ( .A(p_input[194]), .B(p_input[514]), .Z(n5698) );
  XNOR U5718 ( .A(n5748), .B(n5714), .Z(n5707) );
  XNOR U5719 ( .A(p_input[208]), .B(n4027), .Z(n5714) );
  XOR U5720 ( .A(n5704), .B(n5713), .Z(n5748) );
  XOR U5721 ( .A(n5749), .B(n5710), .Z(n5713) );
  XOR U5722 ( .A(p_input[206]), .B(p_input[526]), .Z(n5710) );
  XOR U5723 ( .A(p_input[207]), .B(n4029), .Z(n5749) );
  XOR U5724 ( .A(p_input[202]), .B(p_input[522]), .Z(n5704) );
  XOR U5725 ( .A(n5721), .B(n5719), .Z(n5702) );
  XNOR U5726 ( .A(n5750), .B(n5726), .Z(n5719) );
  XOR U5727 ( .A(p_input[201]), .B(p_input[521]), .Z(n5726) );
  XOR U5728 ( .A(n5716), .B(n5725), .Z(n5750) );
  XOR U5729 ( .A(n5751), .B(n5722), .Z(n5725) );
  XOR U5730 ( .A(p_input[199]), .B(p_input[519]), .Z(n5722) );
  XOR U5731 ( .A(p_input[200]), .B(n4318), .Z(n5751) );
  XOR U5732 ( .A(p_input[195]), .B(p_input[515]), .Z(n5716) );
  XNOR U5733 ( .A(n5731), .B(n5730), .Z(n5721) );
  XOR U5734 ( .A(n5752), .B(n5727), .Z(n5730) );
  XOR U5735 ( .A(p_input[196]), .B(p_input[516]), .Z(n5727) );
  XOR U5736 ( .A(p_input[197]), .B(n4320), .Z(n5752) );
  XOR U5737 ( .A(p_input[198]), .B(p_input[518]), .Z(n5731) );
  XNOR U5738 ( .A(n5753), .B(n5754), .Z(n5544) );
  AND U5739 ( .A(n133), .B(n5755), .Z(n5754) );
  XNOR U5740 ( .A(n5756), .B(n5757), .Z(n133) );
  AND U5741 ( .A(n5758), .B(n5759), .Z(n5757) );
  XOR U5742 ( .A(n5756), .B(n5554), .Z(n5759) );
  XNOR U5743 ( .A(n5756), .B(n5496), .Z(n5758) );
  XOR U5744 ( .A(n5760), .B(n5761), .Z(n5756) );
  AND U5745 ( .A(n5762), .B(n5763), .Z(n5761) );
  XNOR U5746 ( .A(n5567), .B(n5760), .Z(n5763) );
  XOR U5747 ( .A(n5760), .B(n5508), .Z(n5762) );
  XOR U5748 ( .A(n5764), .B(n5765), .Z(n5760) );
  AND U5749 ( .A(n5766), .B(n5767), .Z(n5765) );
  XNOR U5750 ( .A(n5592), .B(n5764), .Z(n5767) );
  XOR U5751 ( .A(n5764), .B(n5519), .Z(n5766) );
  XOR U5752 ( .A(n5768), .B(n5769), .Z(n5764) );
  AND U5753 ( .A(n5770), .B(n5771), .Z(n5769) );
  XOR U5754 ( .A(n5768), .B(n5529), .Z(n5770) );
  XOR U5755 ( .A(n5772), .B(n5773), .Z(n5485) );
  AND U5756 ( .A(n137), .B(n5755), .Z(n5773) );
  XNOR U5757 ( .A(n5753), .B(n5772), .Z(n5755) );
  XNOR U5758 ( .A(n5774), .B(n5775), .Z(n137) );
  AND U5759 ( .A(n5776), .B(n5777), .Z(n5775) );
  XNOR U5760 ( .A(n5778), .B(n5774), .Z(n5777) );
  IV U5761 ( .A(n5554), .Z(n5778) );
  XNOR U5762 ( .A(n5779), .B(n5780), .Z(n5554) );
  AND U5763 ( .A(n140), .B(n5781), .Z(n5780) );
  XNOR U5764 ( .A(n5779), .B(n5782), .Z(n5781) );
  XNOR U5765 ( .A(n5496), .B(n5774), .Z(n5776) );
  XOR U5766 ( .A(n5783), .B(n5784), .Z(n5496) );
  AND U5767 ( .A(n148), .B(n5785), .Z(n5784) );
  XOR U5768 ( .A(n5786), .B(n5787), .Z(n5774) );
  AND U5769 ( .A(n5788), .B(n5789), .Z(n5787) );
  XNOR U5770 ( .A(n5786), .B(n5567), .Z(n5789) );
  XNOR U5771 ( .A(n5790), .B(n5791), .Z(n5567) );
  AND U5772 ( .A(n140), .B(n5792), .Z(n5791) );
  XOR U5773 ( .A(n5793), .B(n5790), .Z(n5792) );
  XNOR U5774 ( .A(n5794), .B(n5786), .Z(n5788) );
  IV U5775 ( .A(n5508), .Z(n5794) );
  XOR U5776 ( .A(n5795), .B(n5796), .Z(n5508) );
  AND U5777 ( .A(n148), .B(n5797), .Z(n5796) );
  XOR U5778 ( .A(n5798), .B(n5799), .Z(n5786) );
  AND U5779 ( .A(n5800), .B(n5801), .Z(n5799) );
  XNOR U5780 ( .A(n5798), .B(n5592), .Z(n5801) );
  XNOR U5781 ( .A(n5802), .B(n5803), .Z(n5592) );
  AND U5782 ( .A(n140), .B(n5804), .Z(n5803) );
  XNOR U5783 ( .A(n5805), .B(n5802), .Z(n5804) );
  XOR U5784 ( .A(n5519), .B(n5798), .Z(n5800) );
  XOR U5785 ( .A(n5806), .B(n5807), .Z(n5519) );
  AND U5786 ( .A(n148), .B(n5808), .Z(n5807) );
  XOR U5787 ( .A(n5768), .B(n5809), .Z(n5798) );
  AND U5788 ( .A(n5810), .B(n5771), .Z(n5809) );
  XNOR U5789 ( .A(n5638), .B(n5768), .Z(n5771) );
  XNOR U5790 ( .A(n5811), .B(n5812), .Z(n5638) );
  AND U5791 ( .A(n140), .B(n5813), .Z(n5812) );
  XOR U5792 ( .A(n5814), .B(n5811), .Z(n5813) );
  XNOR U5793 ( .A(n5815), .B(n5768), .Z(n5810) );
  IV U5794 ( .A(n5529), .Z(n5815) );
  XOR U5795 ( .A(n5816), .B(n5817), .Z(n5529) );
  AND U5796 ( .A(n148), .B(n5818), .Z(n5817) );
  XOR U5797 ( .A(n5819), .B(n5820), .Z(n5768) );
  AND U5798 ( .A(n5821), .B(n5822), .Z(n5820) );
  XNOR U5799 ( .A(n5819), .B(n5732), .Z(n5822) );
  XNOR U5800 ( .A(n5823), .B(n5824), .Z(n5732) );
  AND U5801 ( .A(n140), .B(n5825), .Z(n5824) );
  XNOR U5802 ( .A(n5826), .B(n5823), .Z(n5825) );
  XNOR U5803 ( .A(n5827), .B(n5819), .Z(n5821) );
  IV U5804 ( .A(n5541), .Z(n5827) );
  XOR U5805 ( .A(n5828), .B(n5829), .Z(n5541) );
  AND U5806 ( .A(n148), .B(n5830), .Z(n5829) );
  AND U5807 ( .A(n5772), .B(n5753), .Z(n5819) );
  XNOR U5808 ( .A(n5831), .B(n5832), .Z(n5753) );
  AND U5809 ( .A(n140), .B(n5833), .Z(n5832) );
  XNOR U5810 ( .A(n5834), .B(n5831), .Z(n5833) );
  XNOR U5811 ( .A(n5835), .B(n5836), .Z(n140) );
  AND U5812 ( .A(n5837), .B(n5838), .Z(n5836) );
  XOR U5813 ( .A(n5782), .B(n5835), .Z(n5838) );
  AND U5814 ( .A(n5839), .B(n5840), .Z(n5782) );
  XOR U5815 ( .A(n5835), .B(n5779), .Z(n5837) );
  XNOR U5816 ( .A(n5841), .B(n5842), .Z(n5779) );
  AND U5817 ( .A(n144), .B(n5785), .Z(n5842) );
  XOR U5818 ( .A(n5783), .B(n5841), .Z(n5785) );
  XOR U5819 ( .A(n5843), .B(n5844), .Z(n5835) );
  AND U5820 ( .A(n5845), .B(n5846), .Z(n5844) );
  XNOR U5821 ( .A(n5843), .B(n5839), .Z(n5846) );
  IV U5822 ( .A(n5793), .Z(n5839) );
  XOR U5823 ( .A(n5847), .B(n5848), .Z(n5793) );
  XOR U5824 ( .A(n5849), .B(n5840), .Z(n5848) );
  AND U5825 ( .A(n5805), .B(n5850), .Z(n5840) );
  AND U5826 ( .A(n5851), .B(n5852), .Z(n5849) );
  XOR U5827 ( .A(n5853), .B(n5847), .Z(n5851) );
  XNOR U5828 ( .A(n5790), .B(n5843), .Z(n5845) );
  XNOR U5829 ( .A(n5854), .B(n5855), .Z(n5790) );
  AND U5830 ( .A(n144), .B(n5797), .Z(n5855) );
  XOR U5831 ( .A(n5854), .B(n5795), .Z(n5797) );
  XOR U5832 ( .A(n5856), .B(n5857), .Z(n5843) );
  AND U5833 ( .A(n5858), .B(n5859), .Z(n5857) );
  XNOR U5834 ( .A(n5856), .B(n5805), .Z(n5859) );
  XOR U5835 ( .A(n5860), .B(n5852), .Z(n5805) );
  XNOR U5836 ( .A(n5861), .B(n5847), .Z(n5852) );
  XOR U5837 ( .A(n5862), .B(n5863), .Z(n5847) );
  AND U5838 ( .A(n5864), .B(n5865), .Z(n5863) );
  XOR U5839 ( .A(n5866), .B(n5862), .Z(n5864) );
  XNOR U5840 ( .A(n5867), .B(n5868), .Z(n5861) );
  AND U5841 ( .A(n5869), .B(n5870), .Z(n5868) );
  XOR U5842 ( .A(n5867), .B(n5871), .Z(n5869) );
  XNOR U5843 ( .A(n5853), .B(n5850), .Z(n5860) );
  AND U5844 ( .A(n5872), .B(n5873), .Z(n5850) );
  XOR U5845 ( .A(n5874), .B(n5875), .Z(n5853) );
  AND U5846 ( .A(n5876), .B(n5877), .Z(n5875) );
  XOR U5847 ( .A(n5874), .B(n5878), .Z(n5876) );
  XNOR U5848 ( .A(n5802), .B(n5856), .Z(n5858) );
  XNOR U5849 ( .A(n5879), .B(n5880), .Z(n5802) );
  AND U5850 ( .A(n144), .B(n5808), .Z(n5880) );
  XOR U5851 ( .A(n5879), .B(n5806), .Z(n5808) );
  XOR U5852 ( .A(n5881), .B(n5882), .Z(n5856) );
  AND U5853 ( .A(n5883), .B(n5884), .Z(n5882) );
  XNOR U5854 ( .A(n5881), .B(n5872), .Z(n5884) );
  IV U5855 ( .A(n5814), .Z(n5872) );
  XNOR U5856 ( .A(n5885), .B(n5865), .Z(n5814) );
  XNOR U5857 ( .A(n5886), .B(n5871), .Z(n5865) );
  XOR U5858 ( .A(n5887), .B(n5888), .Z(n5871) );
  AND U5859 ( .A(n5889), .B(n5890), .Z(n5888) );
  XOR U5860 ( .A(n5887), .B(n5891), .Z(n5889) );
  XNOR U5861 ( .A(n5870), .B(n5862), .Z(n5886) );
  XOR U5862 ( .A(n5892), .B(n5893), .Z(n5862) );
  AND U5863 ( .A(n5894), .B(n5895), .Z(n5893) );
  XNOR U5864 ( .A(n5896), .B(n5892), .Z(n5894) );
  XNOR U5865 ( .A(n5897), .B(n5867), .Z(n5870) );
  XOR U5866 ( .A(n5898), .B(n5899), .Z(n5867) );
  AND U5867 ( .A(n5900), .B(n5901), .Z(n5899) );
  XOR U5868 ( .A(n5898), .B(n5902), .Z(n5900) );
  XNOR U5869 ( .A(n5903), .B(n5904), .Z(n5897) );
  AND U5870 ( .A(n5905), .B(n5906), .Z(n5904) );
  XNOR U5871 ( .A(n5903), .B(n5907), .Z(n5905) );
  XNOR U5872 ( .A(n5866), .B(n5873), .Z(n5885) );
  AND U5873 ( .A(n5826), .B(n5908), .Z(n5873) );
  XOR U5874 ( .A(n5878), .B(n5877), .Z(n5866) );
  XNOR U5875 ( .A(n5909), .B(n5874), .Z(n5877) );
  XOR U5876 ( .A(n5910), .B(n5911), .Z(n5874) );
  AND U5877 ( .A(n5912), .B(n5913), .Z(n5911) );
  XOR U5878 ( .A(n5910), .B(n5914), .Z(n5912) );
  XNOR U5879 ( .A(n5915), .B(n5916), .Z(n5909) );
  AND U5880 ( .A(n5917), .B(n5918), .Z(n5916) );
  XOR U5881 ( .A(n5915), .B(n5919), .Z(n5917) );
  XOR U5882 ( .A(n5920), .B(n5921), .Z(n5878) );
  AND U5883 ( .A(n5922), .B(n5923), .Z(n5921) );
  XOR U5884 ( .A(n5920), .B(n5924), .Z(n5922) );
  XNOR U5885 ( .A(n5811), .B(n5881), .Z(n5883) );
  XNOR U5886 ( .A(n5925), .B(n5926), .Z(n5811) );
  AND U5887 ( .A(n144), .B(n5818), .Z(n5926) );
  XOR U5888 ( .A(n5925), .B(n5816), .Z(n5818) );
  XOR U5889 ( .A(n5927), .B(n5928), .Z(n5881) );
  AND U5890 ( .A(n5929), .B(n5930), .Z(n5928) );
  XNOR U5891 ( .A(n5927), .B(n5826), .Z(n5930) );
  XOR U5892 ( .A(n5931), .B(n5895), .Z(n5826) );
  XNOR U5893 ( .A(n5932), .B(n5902), .Z(n5895) );
  XOR U5894 ( .A(n5891), .B(n5890), .Z(n5902) );
  XNOR U5895 ( .A(n5933), .B(n5887), .Z(n5890) );
  XOR U5896 ( .A(n5934), .B(n5935), .Z(n5887) );
  AND U5897 ( .A(n5936), .B(n5937), .Z(n5935) );
  XNOR U5898 ( .A(n5938), .B(n5939), .Z(n5936) );
  IV U5899 ( .A(n5934), .Z(n5938) );
  XNOR U5900 ( .A(n5940), .B(n5941), .Z(n5933) );
  NOR U5901 ( .A(n5942), .B(n5943), .Z(n5941) );
  XNOR U5902 ( .A(n5940), .B(n5944), .Z(n5942) );
  XOR U5903 ( .A(n5945), .B(n5946), .Z(n5891) );
  NOR U5904 ( .A(n5947), .B(n5948), .Z(n5946) );
  XNOR U5905 ( .A(n5945), .B(n5949), .Z(n5947) );
  XNOR U5906 ( .A(n5901), .B(n5892), .Z(n5932) );
  XOR U5907 ( .A(n5950), .B(n5951), .Z(n5892) );
  AND U5908 ( .A(n5952), .B(n5953), .Z(n5951) );
  XOR U5909 ( .A(n5950), .B(n5954), .Z(n5952) );
  XOR U5910 ( .A(n5955), .B(n5907), .Z(n5901) );
  XOR U5911 ( .A(n5956), .B(n5957), .Z(n5907) );
  NOR U5912 ( .A(n5958), .B(n5959), .Z(n5957) );
  XOR U5913 ( .A(n5956), .B(n5960), .Z(n5958) );
  XNOR U5914 ( .A(n5906), .B(n5898), .Z(n5955) );
  XOR U5915 ( .A(n5961), .B(n5962), .Z(n5898) );
  AND U5916 ( .A(n5963), .B(n5964), .Z(n5962) );
  XOR U5917 ( .A(n5961), .B(n5965), .Z(n5963) );
  XNOR U5918 ( .A(n5966), .B(n5903), .Z(n5906) );
  XOR U5919 ( .A(n5967), .B(n5968), .Z(n5903) );
  AND U5920 ( .A(n5969), .B(n5970), .Z(n5968) );
  XNOR U5921 ( .A(n5971), .B(n5972), .Z(n5969) );
  IV U5922 ( .A(n5967), .Z(n5971) );
  XNOR U5923 ( .A(n5973), .B(n5974), .Z(n5966) );
  NOR U5924 ( .A(n5975), .B(n5976), .Z(n5974) );
  XNOR U5925 ( .A(n5973), .B(n5977), .Z(n5975) );
  XOR U5926 ( .A(n5896), .B(n5908), .Z(n5931) );
  NOR U5927 ( .A(n5834), .B(n5978), .Z(n5908) );
  XNOR U5928 ( .A(n5914), .B(n5913), .Z(n5896) );
  XNOR U5929 ( .A(n5979), .B(n5919), .Z(n5913) );
  XNOR U5930 ( .A(n5980), .B(n5981), .Z(n5919) );
  NOR U5931 ( .A(n5982), .B(n5983), .Z(n5981) );
  XOR U5932 ( .A(n5980), .B(n5984), .Z(n5982) );
  XNOR U5933 ( .A(n5918), .B(n5910), .Z(n5979) );
  XOR U5934 ( .A(n5985), .B(n5986), .Z(n5910) );
  AND U5935 ( .A(n5987), .B(n5988), .Z(n5986) );
  XOR U5936 ( .A(n5985), .B(n5989), .Z(n5987) );
  XNOR U5937 ( .A(n5990), .B(n5915), .Z(n5918) );
  XOR U5938 ( .A(n5991), .B(n5992), .Z(n5915) );
  AND U5939 ( .A(n5993), .B(n5994), .Z(n5992) );
  XNOR U5940 ( .A(n5995), .B(n5996), .Z(n5993) );
  IV U5941 ( .A(n5991), .Z(n5995) );
  XNOR U5942 ( .A(n5997), .B(n5998), .Z(n5990) );
  NOR U5943 ( .A(n5999), .B(n6000), .Z(n5998) );
  XNOR U5944 ( .A(n5997), .B(n6001), .Z(n5999) );
  XOR U5945 ( .A(n5924), .B(n5923), .Z(n5914) );
  XNOR U5946 ( .A(n6002), .B(n5920), .Z(n5923) );
  XOR U5947 ( .A(n6003), .B(n6004), .Z(n5920) );
  AND U5948 ( .A(n6005), .B(n6006), .Z(n6004) );
  XNOR U5949 ( .A(n6007), .B(n6008), .Z(n6005) );
  IV U5950 ( .A(n6003), .Z(n6007) );
  XNOR U5951 ( .A(n6009), .B(n6010), .Z(n6002) );
  NOR U5952 ( .A(n6011), .B(n6012), .Z(n6010) );
  XNOR U5953 ( .A(n6009), .B(n6013), .Z(n6011) );
  XOR U5954 ( .A(n6014), .B(n6015), .Z(n5924) );
  NOR U5955 ( .A(n6016), .B(n6017), .Z(n6015) );
  XNOR U5956 ( .A(n6014), .B(n6018), .Z(n6016) );
  XNOR U5957 ( .A(n5823), .B(n5927), .Z(n5929) );
  XNOR U5958 ( .A(n6019), .B(n6020), .Z(n5823) );
  AND U5959 ( .A(n144), .B(n5830), .Z(n6020) );
  XOR U5960 ( .A(n6019), .B(n5828), .Z(n5830) );
  AND U5961 ( .A(n5831), .B(n5834), .Z(n5927) );
  XOR U5962 ( .A(n6021), .B(n5978), .Z(n5834) );
  XNOR U5963 ( .A(p_input[224]), .B(p_input[512]), .Z(n5978) );
  XNOR U5964 ( .A(n5954), .B(n5953), .Z(n6021) );
  XNOR U5965 ( .A(n6022), .B(n5965), .Z(n5953) );
  XOR U5966 ( .A(n5939), .B(n5937), .Z(n5965) );
  XNOR U5967 ( .A(n6023), .B(n5944), .Z(n5937) );
  XOR U5968 ( .A(p_input[248]), .B(p_input[536]), .Z(n5944) );
  XOR U5969 ( .A(n5934), .B(n5943), .Z(n6023) );
  XOR U5970 ( .A(n6024), .B(n5940), .Z(n5943) );
  XOR U5971 ( .A(p_input[246]), .B(p_input[534]), .Z(n5940) );
  XOR U5972 ( .A(p_input[247]), .B(n4010), .Z(n6024) );
  XOR U5973 ( .A(p_input[242]), .B(p_input[530]), .Z(n5934) );
  XNOR U5974 ( .A(n5949), .B(n5948), .Z(n5939) );
  XOR U5975 ( .A(n6025), .B(n5945), .Z(n5948) );
  XOR U5976 ( .A(p_input[243]), .B(p_input[531]), .Z(n5945) );
  XOR U5977 ( .A(p_input[244]), .B(n4012), .Z(n6025) );
  XOR U5978 ( .A(p_input[245]), .B(p_input[533]), .Z(n5949) );
  XOR U5979 ( .A(n5964), .B(n6026), .Z(n6022) );
  IV U5980 ( .A(n5950), .Z(n6026) );
  XOR U5981 ( .A(p_input[225]), .B(p_input[513]), .Z(n5950) );
  XNOR U5982 ( .A(n6027), .B(n5972), .Z(n5964) );
  XNOR U5983 ( .A(n5960), .B(n5959), .Z(n5972) );
  XNOR U5984 ( .A(n6028), .B(n5956), .Z(n5959) );
  XNOR U5985 ( .A(p_input[250]), .B(p_input[538]), .Z(n5956) );
  XOR U5986 ( .A(p_input[251]), .B(n4016), .Z(n6028) );
  XOR U5987 ( .A(p_input[252]), .B(p_input[540]), .Z(n5960) );
  XOR U5988 ( .A(n5970), .B(n6029), .Z(n6027) );
  IV U5989 ( .A(n5961), .Z(n6029) );
  XOR U5990 ( .A(p_input[241]), .B(p_input[529]), .Z(n5961) );
  XNOR U5991 ( .A(n6030), .B(n5977), .Z(n5970) );
  XNOR U5992 ( .A(p_input[255]), .B(n4019), .Z(n5977) );
  XOR U5993 ( .A(n5967), .B(n5976), .Z(n6030) );
  XOR U5994 ( .A(n6031), .B(n5973), .Z(n5976) );
  XOR U5995 ( .A(p_input[253]), .B(p_input[541]), .Z(n5973) );
  XOR U5996 ( .A(p_input[254]), .B(n4021), .Z(n6031) );
  XOR U5997 ( .A(p_input[249]), .B(p_input[537]), .Z(n5967) );
  XOR U5998 ( .A(n5989), .B(n5988), .Z(n5954) );
  XNOR U5999 ( .A(n6032), .B(n5996), .Z(n5988) );
  XNOR U6000 ( .A(n5984), .B(n5983), .Z(n5996) );
  XNOR U6001 ( .A(n6033), .B(n5980), .Z(n5983) );
  XNOR U6002 ( .A(p_input[235]), .B(p_input[523]), .Z(n5980) );
  XOR U6003 ( .A(p_input[236]), .B(n4024), .Z(n6033) );
  XOR U6004 ( .A(p_input[237]), .B(p_input[525]), .Z(n5984) );
  XOR U6005 ( .A(n5994), .B(n6034), .Z(n6032) );
  IV U6006 ( .A(n5985), .Z(n6034) );
  XOR U6007 ( .A(p_input[226]), .B(p_input[514]), .Z(n5985) );
  XNOR U6008 ( .A(n6035), .B(n6001), .Z(n5994) );
  XNOR U6009 ( .A(p_input[240]), .B(n4027), .Z(n6001) );
  XOR U6010 ( .A(n5991), .B(n6000), .Z(n6035) );
  XOR U6011 ( .A(n6036), .B(n5997), .Z(n6000) );
  XOR U6012 ( .A(p_input[238]), .B(p_input[526]), .Z(n5997) );
  XOR U6013 ( .A(p_input[239]), .B(n4029), .Z(n6036) );
  XOR U6014 ( .A(p_input[234]), .B(p_input[522]), .Z(n5991) );
  XOR U6015 ( .A(n6008), .B(n6006), .Z(n5989) );
  XNOR U6016 ( .A(n6037), .B(n6013), .Z(n6006) );
  XOR U6017 ( .A(p_input[233]), .B(p_input[521]), .Z(n6013) );
  XOR U6018 ( .A(n6003), .B(n6012), .Z(n6037) );
  XOR U6019 ( .A(n6038), .B(n6009), .Z(n6012) );
  XOR U6020 ( .A(p_input[231]), .B(p_input[519]), .Z(n6009) );
  XOR U6021 ( .A(p_input[232]), .B(n4318), .Z(n6038) );
  XOR U6022 ( .A(p_input[227]), .B(p_input[515]), .Z(n6003) );
  XNOR U6023 ( .A(n6018), .B(n6017), .Z(n6008) );
  XOR U6024 ( .A(n6039), .B(n6014), .Z(n6017) );
  XOR U6025 ( .A(p_input[228]), .B(p_input[516]), .Z(n6014) );
  XOR U6026 ( .A(p_input[229]), .B(n4320), .Z(n6039) );
  XOR U6027 ( .A(p_input[230]), .B(p_input[518]), .Z(n6018) );
  XNOR U6028 ( .A(n6040), .B(n6041), .Z(n5831) );
  AND U6029 ( .A(n144), .B(n6042), .Z(n6041) );
  XNOR U6030 ( .A(n6043), .B(n6044), .Z(n144) );
  AND U6031 ( .A(n6045), .B(n6046), .Z(n6044) );
  XOR U6032 ( .A(n6043), .B(n5841), .Z(n6046) );
  XNOR U6033 ( .A(n6043), .B(n5783), .Z(n6045) );
  XOR U6034 ( .A(n6047), .B(n6048), .Z(n6043) );
  AND U6035 ( .A(n6049), .B(n6050), .Z(n6048) );
  XNOR U6036 ( .A(n5854), .B(n6047), .Z(n6050) );
  XOR U6037 ( .A(n6047), .B(n5795), .Z(n6049) );
  XOR U6038 ( .A(n6051), .B(n6052), .Z(n6047) );
  AND U6039 ( .A(n6053), .B(n6054), .Z(n6052) );
  XNOR U6040 ( .A(n5879), .B(n6051), .Z(n6054) );
  XOR U6041 ( .A(n6051), .B(n5806), .Z(n6053) );
  XOR U6042 ( .A(n6055), .B(n6056), .Z(n6051) );
  AND U6043 ( .A(n6057), .B(n6058), .Z(n6056) );
  XOR U6044 ( .A(n6055), .B(n5816), .Z(n6057) );
  XOR U6045 ( .A(n6059), .B(n6060), .Z(n5772) );
  AND U6046 ( .A(n148), .B(n6042), .Z(n6060) );
  XNOR U6047 ( .A(n6040), .B(n6059), .Z(n6042) );
  XNOR U6048 ( .A(n6061), .B(n6062), .Z(n148) );
  AND U6049 ( .A(n6063), .B(n6064), .Z(n6062) );
  XNOR U6050 ( .A(n6065), .B(n6061), .Z(n6064) );
  IV U6051 ( .A(n5841), .Z(n6065) );
  XNOR U6052 ( .A(n6066), .B(n6067), .Z(n5841) );
  AND U6053 ( .A(n151), .B(n6068), .Z(n6067) );
  XNOR U6054 ( .A(n6066), .B(n6069), .Z(n6068) );
  XNOR U6055 ( .A(n5783), .B(n6061), .Z(n6063) );
  XOR U6056 ( .A(n6070), .B(n6071), .Z(n5783) );
  AND U6057 ( .A(n159), .B(n6072), .Z(n6071) );
  XOR U6058 ( .A(n6073), .B(n6074), .Z(n6061) );
  AND U6059 ( .A(n6075), .B(n6076), .Z(n6074) );
  XNOR U6060 ( .A(n6073), .B(n5854), .Z(n6076) );
  XNOR U6061 ( .A(n6077), .B(n6078), .Z(n5854) );
  AND U6062 ( .A(n151), .B(n6079), .Z(n6078) );
  XOR U6063 ( .A(n6080), .B(n6077), .Z(n6079) );
  XNOR U6064 ( .A(n6081), .B(n6073), .Z(n6075) );
  IV U6065 ( .A(n5795), .Z(n6081) );
  XOR U6066 ( .A(n6082), .B(n6083), .Z(n5795) );
  AND U6067 ( .A(n159), .B(n6084), .Z(n6083) );
  XOR U6068 ( .A(n6085), .B(n6086), .Z(n6073) );
  AND U6069 ( .A(n6087), .B(n6088), .Z(n6086) );
  XNOR U6070 ( .A(n6085), .B(n5879), .Z(n6088) );
  XNOR U6071 ( .A(n6089), .B(n6090), .Z(n5879) );
  AND U6072 ( .A(n151), .B(n6091), .Z(n6090) );
  XNOR U6073 ( .A(n6092), .B(n6089), .Z(n6091) );
  XOR U6074 ( .A(n5806), .B(n6085), .Z(n6087) );
  XOR U6075 ( .A(n6093), .B(n6094), .Z(n5806) );
  AND U6076 ( .A(n159), .B(n6095), .Z(n6094) );
  XOR U6077 ( .A(n6055), .B(n6096), .Z(n6085) );
  AND U6078 ( .A(n6097), .B(n6058), .Z(n6096) );
  XNOR U6079 ( .A(n5925), .B(n6055), .Z(n6058) );
  XNOR U6080 ( .A(n6098), .B(n6099), .Z(n5925) );
  AND U6081 ( .A(n151), .B(n6100), .Z(n6099) );
  XOR U6082 ( .A(n6101), .B(n6098), .Z(n6100) );
  XNOR U6083 ( .A(n6102), .B(n6055), .Z(n6097) );
  IV U6084 ( .A(n5816), .Z(n6102) );
  XOR U6085 ( .A(n6103), .B(n6104), .Z(n5816) );
  AND U6086 ( .A(n159), .B(n6105), .Z(n6104) );
  XOR U6087 ( .A(n6106), .B(n6107), .Z(n6055) );
  AND U6088 ( .A(n6108), .B(n6109), .Z(n6107) );
  XNOR U6089 ( .A(n6106), .B(n6019), .Z(n6109) );
  XNOR U6090 ( .A(n6110), .B(n6111), .Z(n6019) );
  AND U6091 ( .A(n151), .B(n6112), .Z(n6111) );
  XNOR U6092 ( .A(n6113), .B(n6110), .Z(n6112) );
  XNOR U6093 ( .A(n6114), .B(n6106), .Z(n6108) );
  IV U6094 ( .A(n5828), .Z(n6114) );
  XOR U6095 ( .A(n6115), .B(n6116), .Z(n5828) );
  AND U6096 ( .A(n159), .B(n6117), .Z(n6116) );
  AND U6097 ( .A(n6059), .B(n6040), .Z(n6106) );
  XNOR U6098 ( .A(n6118), .B(n6119), .Z(n6040) );
  AND U6099 ( .A(n151), .B(n6120), .Z(n6119) );
  XNOR U6100 ( .A(n6121), .B(n6118), .Z(n6120) );
  XNOR U6101 ( .A(n6122), .B(n6123), .Z(n151) );
  AND U6102 ( .A(n6124), .B(n6125), .Z(n6123) );
  XOR U6103 ( .A(n6069), .B(n6122), .Z(n6125) );
  AND U6104 ( .A(n6126), .B(n6127), .Z(n6069) );
  XOR U6105 ( .A(n6122), .B(n6066), .Z(n6124) );
  XNOR U6106 ( .A(n6128), .B(n6129), .Z(n6066) );
  AND U6107 ( .A(n155), .B(n6072), .Z(n6129) );
  XOR U6108 ( .A(n6070), .B(n6128), .Z(n6072) );
  XOR U6109 ( .A(n6130), .B(n6131), .Z(n6122) );
  AND U6110 ( .A(n6132), .B(n6133), .Z(n6131) );
  XNOR U6111 ( .A(n6130), .B(n6126), .Z(n6133) );
  IV U6112 ( .A(n6080), .Z(n6126) );
  XOR U6113 ( .A(n6134), .B(n6135), .Z(n6080) );
  XOR U6114 ( .A(n6136), .B(n6127), .Z(n6135) );
  AND U6115 ( .A(n6092), .B(n6137), .Z(n6127) );
  AND U6116 ( .A(n6138), .B(n6139), .Z(n6136) );
  XOR U6117 ( .A(n6140), .B(n6134), .Z(n6138) );
  XNOR U6118 ( .A(n6077), .B(n6130), .Z(n6132) );
  XNOR U6119 ( .A(n6141), .B(n6142), .Z(n6077) );
  AND U6120 ( .A(n155), .B(n6084), .Z(n6142) );
  XOR U6121 ( .A(n6141), .B(n6082), .Z(n6084) );
  XOR U6122 ( .A(n6143), .B(n6144), .Z(n6130) );
  AND U6123 ( .A(n6145), .B(n6146), .Z(n6144) );
  XNOR U6124 ( .A(n6143), .B(n6092), .Z(n6146) );
  XOR U6125 ( .A(n6147), .B(n6139), .Z(n6092) );
  XNOR U6126 ( .A(n6148), .B(n6134), .Z(n6139) );
  XOR U6127 ( .A(n6149), .B(n6150), .Z(n6134) );
  AND U6128 ( .A(n6151), .B(n6152), .Z(n6150) );
  XOR U6129 ( .A(n6153), .B(n6149), .Z(n6151) );
  XNOR U6130 ( .A(n6154), .B(n6155), .Z(n6148) );
  AND U6131 ( .A(n6156), .B(n6157), .Z(n6155) );
  XOR U6132 ( .A(n6154), .B(n6158), .Z(n6156) );
  XNOR U6133 ( .A(n6140), .B(n6137), .Z(n6147) );
  AND U6134 ( .A(n6159), .B(n6160), .Z(n6137) );
  XOR U6135 ( .A(n6161), .B(n6162), .Z(n6140) );
  AND U6136 ( .A(n6163), .B(n6164), .Z(n6162) );
  XOR U6137 ( .A(n6161), .B(n6165), .Z(n6163) );
  XNOR U6138 ( .A(n6089), .B(n6143), .Z(n6145) );
  XNOR U6139 ( .A(n6166), .B(n6167), .Z(n6089) );
  AND U6140 ( .A(n155), .B(n6095), .Z(n6167) );
  XOR U6141 ( .A(n6166), .B(n6093), .Z(n6095) );
  XOR U6142 ( .A(n6168), .B(n6169), .Z(n6143) );
  AND U6143 ( .A(n6170), .B(n6171), .Z(n6169) );
  XNOR U6144 ( .A(n6168), .B(n6159), .Z(n6171) );
  IV U6145 ( .A(n6101), .Z(n6159) );
  XNOR U6146 ( .A(n6172), .B(n6152), .Z(n6101) );
  XNOR U6147 ( .A(n6173), .B(n6158), .Z(n6152) );
  XOR U6148 ( .A(n6174), .B(n6175), .Z(n6158) );
  AND U6149 ( .A(n6176), .B(n6177), .Z(n6175) );
  XOR U6150 ( .A(n6174), .B(n6178), .Z(n6176) );
  XNOR U6151 ( .A(n6157), .B(n6149), .Z(n6173) );
  XOR U6152 ( .A(n6179), .B(n6180), .Z(n6149) );
  AND U6153 ( .A(n6181), .B(n6182), .Z(n6180) );
  XNOR U6154 ( .A(n6183), .B(n6179), .Z(n6181) );
  XNOR U6155 ( .A(n6184), .B(n6154), .Z(n6157) );
  XOR U6156 ( .A(n6185), .B(n6186), .Z(n6154) );
  AND U6157 ( .A(n6187), .B(n6188), .Z(n6186) );
  XOR U6158 ( .A(n6185), .B(n6189), .Z(n6187) );
  XNOR U6159 ( .A(n6190), .B(n6191), .Z(n6184) );
  AND U6160 ( .A(n6192), .B(n6193), .Z(n6191) );
  XNOR U6161 ( .A(n6190), .B(n6194), .Z(n6192) );
  XNOR U6162 ( .A(n6153), .B(n6160), .Z(n6172) );
  AND U6163 ( .A(n6113), .B(n6195), .Z(n6160) );
  XOR U6164 ( .A(n6165), .B(n6164), .Z(n6153) );
  XNOR U6165 ( .A(n6196), .B(n6161), .Z(n6164) );
  XOR U6166 ( .A(n6197), .B(n6198), .Z(n6161) );
  AND U6167 ( .A(n6199), .B(n6200), .Z(n6198) );
  XOR U6168 ( .A(n6197), .B(n6201), .Z(n6199) );
  XNOR U6169 ( .A(n6202), .B(n6203), .Z(n6196) );
  AND U6170 ( .A(n6204), .B(n6205), .Z(n6203) );
  XOR U6171 ( .A(n6202), .B(n6206), .Z(n6204) );
  XOR U6172 ( .A(n6207), .B(n6208), .Z(n6165) );
  AND U6173 ( .A(n6209), .B(n6210), .Z(n6208) );
  XOR U6174 ( .A(n6207), .B(n6211), .Z(n6209) );
  XNOR U6175 ( .A(n6098), .B(n6168), .Z(n6170) );
  XNOR U6176 ( .A(n6212), .B(n6213), .Z(n6098) );
  AND U6177 ( .A(n155), .B(n6105), .Z(n6213) );
  XOR U6178 ( .A(n6212), .B(n6103), .Z(n6105) );
  XOR U6179 ( .A(n6214), .B(n6215), .Z(n6168) );
  AND U6180 ( .A(n6216), .B(n6217), .Z(n6215) );
  XNOR U6181 ( .A(n6214), .B(n6113), .Z(n6217) );
  XOR U6182 ( .A(n6218), .B(n6182), .Z(n6113) );
  XNOR U6183 ( .A(n6219), .B(n6189), .Z(n6182) );
  XOR U6184 ( .A(n6178), .B(n6177), .Z(n6189) );
  XNOR U6185 ( .A(n6220), .B(n6174), .Z(n6177) );
  XOR U6186 ( .A(n6221), .B(n6222), .Z(n6174) );
  AND U6187 ( .A(n6223), .B(n6224), .Z(n6222) );
  XNOR U6188 ( .A(n6225), .B(n6226), .Z(n6223) );
  IV U6189 ( .A(n6221), .Z(n6225) );
  XNOR U6190 ( .A(n6227), .B(n6228), .Z(n6220) );
  NOR U6191 ( .A(n6229), .B(n6230), .Z(n6228) );
  XNOR U6192 ( .A(n6227), .B(n6231), .Z(n6229) );
  XOR U6193 ( .A(n6232), .B(n6233), .Z(n6178) );
  NOR U6194 ( .A(n6234), .B(n6235), .Z(n6233) );
  XNOR U6195 ( .A(n6232), .B(n6236), .Z(n6234) );
  XNOR U6196 ( .A(n6188), .B(n6179), .Z(n6219) );
  XOR U6197 ( .A(n6237), .B(n6238), .Z(n6179) );
  AND U6198 ( .A(n6239), .B(n6240), .Z(n6238) );
  XOR U6199 ( .A(n6237), .B(n6241), .Z(n6239) );
  XOR U6200 ( .A(n6242), .B(n6194), .Z(n6188) );
  XOR U6201 ( .A(n6243), .B(n6244), .Z(n6194) );
  NOR U6202 ( .A(n6245), .B(n6246), .Z(n6244) );
  XOR U6203 ( .A(n6243), .B(n6247), .Z(n6245) );
  XNOR U6204 ( .A(n6193), .B(n6185), .Z(n6242) );
  XOR U6205 ( .A(n6248), .B(n6249), .Z(n6185) );
  AND U6206 ( .A(n6250), .B(n6251), .Z(n6249) );
  XOR U6207 ( .A(n6248), .B(n6252), .Z(n6250) );
  XNOR U6208 ( .A(n6253), .B(n6190), .Z(n6193) );
  XOR U6209 ( .A(n6254), .B(n6255), .Z(n6190) );
  AND U6210 ( .A(n6256), .B(n6257), .Z(n6255) );
  XNOR U6211 ( .A(n6258), .B(n6259), .Z(n6256) );
  IV U6212 ( .A(n6254), .Z(n6258) );
  XNOR U6213 ( .A(n6260), .B(n6261), .Z(n6253) );
  NOR U6214 ( .A(n6262), .B(n6263), .Z(n6261) );
  XNOR U6215 ( .A(n6260), .B(n6264), .Z(n6262) );
  XOR U6216 ( .A(n6183), .B(n6195), .Z(n6218) );
  NOR U6217 ( .A(n6121), .B(n6265), .Z(n6195) );
  XNOR U6218 ( .A(n6201), .B(n6200), .Z(n6183) );
  XNOR U6219 ( .A(n6266), .B(n6206), .Z(n6200) );
  XNOR U6220 ( .A(n6267), .B(n6268), .Z(n6206) );
  NOR U6221 ( .A(n6269), .B(n6270), .Z(n6268) );
  XOR U6222 ( .A(n6267), .B(n6271), .Z(n6269) );
  XNOR U6223 ( .A(n6205), .B(n6197), .Z(n6266) );
  XOR U6224 ( .A(n6272), .B(n6273), .Z(n6197) );
  AND U6225 ( .A(n6274), .B(n6275), .Z(n6273) );
  XOR U6226 ( .A(n6272), .B(n6276), .Z(n6274) );
  XNOR U6227 ( .A(n6277), .B(n6202), .Z(n6205) );
  XOR U6228 ( .A(n6278), .B(n6279), .Z(n6202) );
  AND U6229 ( .A(n6280), .B(n6281), .Z(n6279) );
  XNOR U6230 ( .A(n6282), .B(n6283), .Z(n6280) );
  IV U6231 ( .A(n6278), .Z(n6282) );
  XNOR U6232 ( .A(n6284), .B(n6285), .Z(n6277) );
  NOR U6233 ( .A(n6286), .B(n6287), .Z(n6285) );
  XNOR U6234 ( .A(n6284), .B(n6288), .Z(n6286) );
  XOR U6235 ( .A(n6211), .B(n6210), .Z(n6201) );
  XNOR U6236 ( .A(n6289), .B(n6207), .Z(n6210) );
  XOR U6237 ( .A(n6290), .B(n6291), .Z(n6207) );
  AND U6238 ( .A(n6292), .B(n6293), .Z(n6291) );
  XNOR U6239 ( .A(n6294), .B(n6295), .Z(n6292) );
  IV U6240 ( .A(n6290), .Z(n6294) );
  XNOR U6241 ( .A(n6296), .B(n6297), .Z(n6289) );
  NOR U6242 ( .A(n6298), .B(n6299), .Z(n6297) );
  XNOR U6243 ( .A(n6296), .B(n6300), .Z(n6298) );
  XOR U6244 ( .A(n6301), .B(n6302), .Z(n6211) );
  NOR U6245 ( .A(n6303), .B(n6304), .Z(n6302) );
  XNOR U6246 ( .A(n6301), .B(n6305), .Z(n6303) );
  XNOR U6247 ( .A(n6110), .B(n6214), .Z(n6216) );
  XNOR U6248 ( .A(n6306), .B(n6307), .Z(n6110) );
  AND U6249 ( .A(n155), .B(n6117), .Z(n6307) );
  XOR U6250 ( .A(n6306), .B(n6115), .Z(n6117) );
  AND U6251 ( .A(n6118), .B(n6121), .Z(n6214) );
  XOR U6252 ( .A(n6308), .B(n6265), .Z(n6121) );
  XNOR U6253 ( .A(p_input[256]), .B(p_input[512]), .Z(n6265) );
  XNOR U6254 ( .A(n6241), .B(n6240), .Z(n6308) );
  XNOR U6255 ( .A(n6309), .B(n6252), .Z(n6240) );
  XOR U6256 ( .A(n6226), .B(n6224), .Z(n6252) );
  XNOR U6257 ( .A(n6310), .B(n6231), .Z(n6224) );
  XOR U6258 ( .A(p_input[280]), .B(p_input[536]), .Z(n6231) );
  XOR U6259 ( .A(n6221), .B(n6230), .Z(n6310) );
  XOR U6260 ( .A(n6311), .B(n6227), .Z(n6230) );
  XOR U6261 ( .A(p_input[278]), .B(p_input[534]), .Z(n6227) );
  XOR U6262 ( .A(p_input[279]), .B(n4010), .Z(n6311) );
  XOR U6263 ( .A(p_input[274]), .B(p_input[530]), .Z(n6221) );
  XNOR U6264 ( .A(n6236), .B(n6235), .Z(n6226) );
  XOR U6265 ( .A(n6312), .B(n6232), .Z(n6235) );
  XOR U6266 ( .A(p_input[275]), .B(p_input[531]), .Z(n6232) );
  XOR U6267 ( .A(p_input[276]), .B(n4012), .Z(n6312) );
  XOR U6268 ( .A(p_input[277]), .B(p_input[533]), .Z(n6236) );
  XOR U6269 ( .A(n6251), .B(n6313), .Z(n6309) );
  IV U6270 ( .A(n6237), .Z(n6313) );
  XOR U6271 ( .A(p_input[257]), .B(p_input[513]), .Z(n6237) );
  XNOR U6272 ( .A(n6314), .B(n6259), .Z(n6251) );
  XNOR U6273 ( .A(n6247), .B(n6246), .Z(n6259) );
  XNOR U6274 ( .A(n6315), .B(n6243), .Z(n6246) );
  XNOR U6275 ( .A(p_input[282]), .B(p_input[538]), .Z(n6243) );
  XOR U6276 ( .A(p_input[283]), .B(n4016), .Z(n6315) );
  XOR U6277 ( .A(p_input[284]), .B(p_input[540]), .Z(n6247) );
  XOR U6278 ( .A(n6257), .B(n6316), .Z(n6314) );
  IV U6279 ( .A(n6248), .Z(n6316) );
  XOR U6280 ( .A(p_input[273]), .B(p_input[529]), .Z(n6248) );
  XNOR U6281 ( .A(n6317), .B(n6264), .Z(n6257) );
  XNOR U6282 ( .A(p_input[287]), .B(n4019), .Z(n6264) );
  XOR U6283 ( .A(n6254), .B(n6263), .Z(n6317) );
  XOR U6284 ( .A(n6318), .B(n6260), .Z(n6263) );
  XOR U6285 ( .A(p_input[285]), .B(p_input[541]), .Z(n6260) );
  XOR U6286 ( .A(p_input[286]), .B(n4021), .Z(n6318) );
  XOR U6287 ( .A(p_input[281]), .B(p_input[537]), .Z(n6254) );
  XOR U6288 ( .A(n6276), .B(n6275), .Z(n6241) );
  XNOR U6289 ( .A(n6319), .B(n6283), .Z(n6275) );
  XNOR U6290 ( .A(n6271), .B(n6270), .Z(n6283) );
  XNOR U6291 ( .A(n6320), .B(n6267), .Z(n6270) );
  XNOR U6292 ( .A(p_input[267]), .B(p_input[523]), .Z(n6267) );
  XOR U6293 ( .A(p_input[268]), .B(n4024), .Z(n6320) );
  XOR U6294 ( .A(p_input[269]), .B(p_input[525]), .Z(n6271) );
  XOR U6295 ( .A(n6281), .B(n6321), .Z(n6319) );
  IV U6296 ( .A(n6272), .Z(n6321) );
  XOR U6297 ( .A(p_input[258]), .B(p_input[514]), .Z(n6272) );
  XNOR U6298 ( .A(n6322), .B(n6288), .Z(n6281) );
  XNOR U6299 ( .A(p_input[272]), .B(n4027), .Z(n6288) );
  XOR U6300 ( .A(n6278), .B(n6287), .Z(n6322) );
  XOR U6301 ( .A(n6323), .B(n6284), .Z(n6287) );
  XOR U6302 ( .A(p_input[270]), .B(p_input[526]), .Z(n6284) );
  XOR U6303 ( .A(p_input[271]), .B(n4029), .Z(n6323) );
  XOR U6304 ( .A(p_input[266]), .B(p_input[522]), .Z(n6278) );
  XOR U6305 ( .A(n6295), .B(n6293), .Z(n6276) );
  XNOR U6306 ( .A(n6324), .B(n6300), .Z(n6293) );
  XOR U6307 ( .A(p_input[265]), .B(p_input[521]), .Z(n6300) );
  XOR U6308 ( .A(n6290), .B(n6299), .Z(n6324) );
  XOR U6309 ( .A(n6325), .B(n6296), .Z(n6299) );
  XOR U6310 ( .A(p_input[263]), .B(p_input[519]), .Z(n6296) );
  XOR U6311 ( .A(p_input[264]), .B(n4318), .Z(n6325) );
  XOR U6312 ( .A(p_input[259]), .B(p_input[515]), .Z(n6290) );
  XNOR U6313 ( .A(n6305), .B(n6304), .Z(n6295) );
  XOR U6314 ( .A(n6326), .B(n6301), .Z(n6304) );
  XOR U6315 ( .A(p_input[260]), .B(p_input[516]), .Z(n6301) );
  XOR U6316 ( .A(p_input[261]), .B(n4320), .Z(n6326) );
  XOR U6317 ( .A(p_input[262]), .B(p_input[518]), .Z(n6305) );
  XNOR U6318 ( .A(n6327), .B(n6328), .Z(n6118) );
  AND U6319 ( .A(n155), .B(n6329), .Z(n6328) );
  XNOR U6320 ( .A(n6330), .B(n6331), .Z(n155) );
  AND U6321 ( .A(n6332), .B(n6333), .Z(n6331) );
  XOR U6322 ( .A(n6330), .B(n6128), .Z(n6333) );
  XNOR U6323 ( .A(n6330), .B(n6070), .Z(n6332) );
  XOR U6324 ( .A(n6334), .B(n6335), .Z(n6330) );
  AND U6325 ( .A(n6336), .B(n6337), .Z(n6335) );
  XNOR U6326 ( .A(n6141), .B(n6334), .Z(n6337) );
  XOR U6327 ( .A(n6334), .B(n6082), .Z(n6336) );
  XOR U6328 ( .A(n6338), .B(n6339), .Z(n6334) );
  AND U6329 ( .A(n6340), .B(n6341), .Z(n6339) );
  XNOR U6330 ( .A(n6166), .B(n6338), .Z(n6341) );
  XOR U6331 ( .A(n6338), .B(n6093), .Z(n6340) );
  XOR U6332 ( .A(n6342), .B(n6343), .Z(n6338) );
  AND U6333 ( .A(n6344), .B(n6345), .Z(n6343) );
  XOR U6334 ( .A(n6342), .B(n6103), .Z(n6344) );
  XOR U6335 ( .A(n6346), .B(n6347), .Z(n6059) );
  AND U6336 ( .A(n159), .B(n6329), .Z(n6347) );
  XNOR U6337 ( .A(n6327), .B(n6346), .Z(n6329) );
  XNOR U6338 ( .A(n6348), .B(n6349), .Z(n159) );
  AND U6339 ( .A(n6350), .B(n6351), .Z(n6349) );
  XNOR U6340 ( .A(n6352), .B(n6348), .Z(n6351) );
  IV U6341 ( .A(n6128), .Z(n6352) );
  XNOR U6342 ( .A(n6353), .B(n6354), .Z(n6128) );
  AND U6343 ( .A(n162), .B(n6355), .Z(n6354) );
  XNOR U6344 ( .A(n6353), .B(n6356), .Z(n6355) );
  XNOR U6345 ( .A(n6070), .B(n6348), .Z(n6350) );
  XNOR U6346 ( .A(n6357), .B(n6358), .Z(n6070) );
  AND U6347 ( .A(n170), .B(n6359), .Z(n6358) );
  XNOR U6348 ( .A(n6360), .B(n6361), .Z(n6359) );
  XOR U6349 ( .A(n6362), .B(n6363), .Z(n6348) );
  AND U6350 ( .A(n6364), .B(n6365), .Z(n6363) );
  XNOR U6351 ( .A(n6362), .B(n6141), .Z(n6365) );
  XNOR U6352 ( .A(n6366), .B(n6367), .Z(n6141) );
  AND U6353 ( .A(n162), .B(n6368), .Z(n6367) );
  XOR U6354 ( .A(n6369), .B(n6366), .Z(n6368) );
  XNOR U6355 ( .A(n6370), .B(n6362), .Z(n6364) );
  IV U6356 ( .A(n6082), .Z(n6370) );
  XOR U6357 ( .A(n6371), .B(n6372), .Z(n6082) );
  AND U6358 ( .A(n170), .B(n6373), .Z(n6372) );
  XOR U6359 ( .A(n6374), .B(n6375), .Z(n6362) );
  AND U6360 ( .A(n6376), .B(n6377), .Z(n6375) );
  XNOR U6361 ( .A(n6374), .B(n6166), .Z(n6377) );
  XNOR U6362 ( .A(n6378), .B(n6379), .Z(n6166) );
  AND U6363 ( .A(n162), .B(n6380), .Z(n6379) );
  XNOR U6364 ( .A(n6381), .B(n6378), .Z(n6380) );
  XOR U6365 ( .A(n6093), .B(n6374), .Z(n6376) );
  XOR U6366 ( .A(n6382), .B(n6383), .Z(n6093) );
  AND U6367 ( .A(n170), .B(n6384), .Z(n6383) );
  XOR U6368 ( .A(n6342), .B(n6385), .Z(n6374) );
  AND U6369 ( .A(n6386), .B(n6345), .Z(n6385) );
  XNOR U6370 ( .A(n6212), .B(n6342), .Z(n6345) );
  XNOR U6371 ( .A(n6387), .B(n6388), .Z(n6212) );
  AND U6372 ( .A(n162), .B(n6389), .Z(n6388) );
  XOR U6373 ( .A(n6390), .B(n6387), .Z(n6389) );
  XNOR U6374 ( .A(n6391), .B(n6342), .Z(n6386) );
  IV U6375 ( .A(n6103), .Z(n6391) );
  XOR U6376 ( .A(n6392), .B(n6393), .Z(n6103) );
  AND U6377 ( .A(n170), .B(n6394), .Z(n6393) );
  XOR U6378 ( .A(n6395), .B(n6396), .Z(n6342) );
  AND U6379 ( .A(n6397), .B(n6398), .Z(n6396) );
  XNOR U6380 ( .A(n6395), .B(n6306), .Z(n6398) );
  XNOR U6381 ( .A(n6399), .B(n6400), .Z(n6306) );
  AND U6382 ( .A(n162), .B(n6401), .Z(n6400) );
  XNOR U6383 ( .A(n6402), .B(n6399), .Z(n6401) );
  XNOR U6384 ( .A(n6403), .B(n6395), .Z(n6397) );
  IV U6385 ( .A(n6115), .Z(n6403) );
  XOR U6386 ( .A(n6404), .B(n6405), .Z(n6115) );
  AND U6387 ( .A(n170), .B(n6406), .Z(n6405) );
  AND U6388 ( .A(n6346), .B(n6327), .Z(n6395) );
  XNOR U6389 ( .A(n6407), .B(n6408), .Z(n6327) );
  AND U6390 ( .A(n162), .B(n6409), .Z(n6408) );
  XNOR U6391 ( .A(n6410), .B(n6407), .Z(n6409) );
  XNOR U6392 ( .A(n6411), .B(n6412), .Z(n162) );
  AND U6393 ( .A(n6413), .B(n6414), .Z(n6412) );
  XOR U6394 ( .A(n6356), .B(n6411), .Z(n6414) );
  AND U6395 ( .A(n6415), .B(n6416), .Z(n6356) );
  XOR U6396 ( .A(n6411), .B(n6353), .Z(n6413) );
  XOR U6397 ( .A(n6360), .B(n6417), .Z(n6353) );
  AND U6398 ( .A(n166), .B(n6418), .Z(n6417) );
  XOR U6399 ( .A(n6360), .B(n6357), .Z(n6418) );
  XOR U6400 ( .A(n6419), .B(n6420), .Z(n6411) );
  AND U6401 ( .A(n6421), .B(n6422), .Z(n6420) );
  XNOR U6402 ( .A(n6419), .B(n6415), .Z(n6422) );
  IV U6403 ( .A(n6369), .Z(n6415) );
  XOR U6404 ( .A(n6423), .B(n6424), .Z(n6369) );
  XOR U6405 ( .A(n6425), .B(n6416), .Z(n6424) );
  AND U6406 ( .A(n6381), .B(n6426), .Z(n6416) );
  AND U6407 ( .A(n6427), .B(n6428), .Z(n6425) );
  XOR U6408 ( .A(n6429), .B(n6423), .Z(n6427) );
  XNOR U6409 ( .A(n6366), .B(n6419), .Z(n6421) );
  XNOR U6410 ( .A(n6430), .B(n6431), .Z(n6366) );
  AND U6411 ( .A(n166), .B(n6373), .Z(n6431) );
  XOR U6412 ( .A(n6430), .B(n6371), .Z(n6373) );
  XOR U6413 ( .A(n6432), .B(n6433), .Z(n6419) );
  AND U6414 ( .A(n6434), .B(n6435), .Z(n6433) );
  XNOR U6415 ( .A(n6432), .B(n6381), .Z(n6435) );
  XOR U6416 ( .A(n6436), .B(n6428), .Z(n6381) );
  XNOR U6417 ( .A(n6437), .B(n6423), .Z(n6428) );
  XOR U6418 ( .A(n6438), .B(n6439), .Z(n6423) );
  AND U6419 ( .A(n6440), .B(n6441), .Z(n6439) );
  XOR U6420 ( .A(n6442), .B(n6438), .Z(n6440) );
  XNOR U6421 ( .A(n6443), .B(n6444), .Z(n6437) );
  AND U6422 ( .A(n6445), .B(n6446), .Z(n6444) );
  XOR U6423 ( .A(n6443), .B(n6447), .Z(n6445) );
  XNOR U6424 ( .A(n6429), .B(n6426), .Z(n6436) );
  AND U6425 ( .A(n6448), .B(n6449), .Z(n6426) );
  XOR U6426 ( .A(n6450), .B(n6451), .Z(n6429) );
  AND U6427 ( .A(n6452), .B(n6453), .Z(n6451) );
  XOR U6428 ( .A(n6450), .B(n6454), .Z(n6452) );
  XNOR U6429 ( .A(n6378), .B(n6432), .Z(n6434) );
  XNOR U6430 ( .A(n6455), .B(n6456), .Z(n6378) );
  AND U6431 ( .A(n166), .B(n6384), .Z(n6456) );
  XOR U6432 ( .A(n6455), .B(n6382), .Z(n6384) );
  XOR U6433 ( .A(n6457), .B(n6458), .Z(n6432) );
  AND U6434 ( .A(n6459), .B(n6460), .Z(n6458) );
  XNOR U6435 ( .A(n6457), .B(n6448), .Z(n6460) );
  IV U6436 ( .A(n6390), .Z(n6448) );
  XNOR U6437 ( .A(n6461), .B(n6441), .Z(n6390) );
  XNOR U6438 ( .A(n6462), .B(n6447), .Z(n6441) );
  XOR U6439 ( .A(n6463), .B(n6464), .Z(n6447) );
  AND U6440 ( .A(n6465), .B(n6466), .Z(n6464) );
  XOR U6441 ( .A(n6463), .B(n6467), .Z(n6465) );
  XNOR U6442 ( .A(n6446), .B(n6438), .Z(n6462) );
  XOR U6443 ( .A(n6468), .B(n6469), .Z(n6438) );
  AND U6444 ( .A(n6470), .B(n6471), .Z(n6469) );
  XNOR U6445 ( .A(n6472), .B(n6468), .Z(n6470) );
  XNOR U6446 ( .A(n6473), .B(n6443), .Z(n6446) );
  XOR U6447 ( .A(n6474), .B(n6475), .Z(n6443) );
  AND U6448 ( .A(n6476), .B(n6477), .Z(n6475) );
  XOR U6449 ( .A(n6474), .B(n6478), .Z(n6476) );
  XNOR U6450 ( .A(n6479), .B(n6480), .Z(n6473) );
  AND U6451 ( .A(n6481), .B(n6482), .Z(n6480) );
  XNOR U6452 ( .A(n6479), .B(n6483), .Z(n6481) );
  XNOR U6453 ( .A(n6442), .B(n6449), .Z(n6461) );
  AND U6454 ( .A(n6402), .B(n6484), .Z(n6449) );
  XOR U6455 ( .A(n6454), .B(n6453), .Z(n6442) );
  XNOR U6456 ( .A(n6485), .B(n6450), .Z(n6453) );
  XOR U6457 ( .A(n6486), .B(n6487), .Z(n6450) );
  AND U6458 ( .A(n6488), .B(n6489), .Z(n6487) );
  XOR U6459 ( .A(n6486), .B(n6490), .Z(n6488) );
  XNOR U6460 ( .A(n6491), .B(n6492), .Z(n6485) );
  AND U6461 ( .A(n6493), .B(n6494), .Z(n6492) );
  XOR U6462 ( .A(n6491), .B(n6495), .Z(n6493) );
  XOR U6463 ( .A(n6496), .B(n6497), .Z(n6454) );
  AND U6464 ( .A(n6498), .B(n6499), .Z(n6497) );
  XOR U6465 ( .A(n6496), .B(n6500), .Z(n6498) );
  XNOR U6466 ( .A(n6387), .B(n6457), .Z(n6459) );
  XNOR U6467 ( .A(n6501), .B(n6502), .Z(n6387) );
  AND U6468 ( .A(n166), .B(n6394), .Z(n6502) );
  XOR U6469 ( .A(n6501), .B(n6392), .Z(n6394) );
  XOR U6470 ( .A(n6503), .B(n6504), .Z(n6457) );
  AND U6471 ( .A(n6505), .B(n6506), .Z(n6504) );
  XNOR U6472 ( .A(n6503), .B(n6402), .Z(n6506) );
  XOR U6473 ( .A(n6507), .B(n6471), .Z(n6402) );
  XNOR U6474 ( .A(n6508), .B(n6478), .Z(n6471) );
  XOR U6475 ( .A(n6467), .B(n6466), .Z(n6478) );
  XNOR U6476 ( .A(n6509), .B(n6463), .Z(n6466) );
  XOR U6477 ( .A(n6510), .B(n6511), .Z(n6463) );
  AND U6478 ( .A(n6512), .B(n6513), .Z(n6511) );
  XNOR U6479 ( .A(n6514), .B(n6515), .Z(n6512) );
  IV U6480 ( .A(n6510), .Z(n6514) );
  XNOR U6481 ( .A(n6516), .B(n6517), .Z(n6509) );
  NOR U6482 ( .A(n6518), .B(n6519), .Z(n6517) );
  XNOR U6483 ( .A(n6516), .B(n6520), .Z(n6518) );
  XOR U6484 ( .A(n6521), .B(n6522), .Z(n6467) );
  NOR U6485 ( .A(n6523), .B(n6524), .Z(n6522) );
  XNOR U6486 ( .A(n6521), .B(n6525), .Z(n6523) );
  XNOR U6487 ( .A(n6477), .B(n6468), .Z(n6508) );
  XOR U6488 ( .A(n6526), .B(n6527), .Z(n6468) );
  AND U6489 ( .A(n6528), .B(n6529), .Z(n6527) );
  XOR U6490 ( .A(n6526), .B(n6530), .Z(n6528) );
  XOR U6491 ( .A(n6531), .B(n6483), .Z(n6477) );
  XOR U6492 ( .A(n6532), .B(n6533), .Z(n6483) );
  NOR U6493 ( .A(n6534), .B(n6535), .Z(n6533) );
  XOR U6494 ( .A(n6532), .B(n6536), .Z(n6534) );
  XNOR U6495 ( .A(n6482), .B(n6474), .Z(n6531) );
  XOR U6496 ( .A(n6537), .B(n6538), .Z(n6474) );
  AND U6497 ( .A(n6539), .B(n6540), .Z(n6538) );
  XOR U6498 ( .A(n6537), .B(n6541), .Z(n6539) );
  XNOR U6499 ( .A(n6542), .B(n6479), .Z(n6482) );
  XOR U6500 ( .A(n6543), .B(n6544), .Z(n6479) );
  AND U6501 ( .A(n6545), .B(n6546), .Z(n6544) );
  XNOR U6502 ( .A(n6547), .B(n6548), .Z(n6545) );
  IV U6503 ( .A(n6543), .Z(n6547) );
  XNOR U6504 ( .A(n6549), .B(n6550), .Z(n6542) );
  NOR U6505 ( .A(n6551), .B(n6552), .Z(n6550) );
  XNOR U6506 ( .A(n6549), .B(n6553), .Z(n6551) );
  XOR U6507 ( .A(n6472), .B(n6484), .Z(n6507) );
  NOR U6508 ( .A(n6410), .B(n6554), .Z(n6484) );
  XNOR U6509 ( .A(n6490), .B(n6489), .Z(n6472) );
  XNOR U6510 ( .A(n6555), .B(n6495), .Z(n6489) );
  XNOR U6511 ( .A(n6556), .B(n6557), .Z(n6495) );
  NOR U6512 ( .A(n6558), .B(n6559), .Z(n6557) );
  XOR U6513 ( .A(n6556), .B(n6560), .Z(n6558) );
  XNOR U6514 ( .A(n6494), .B(n6486), .Z(n6555) );
  XOR U6515 ( .A(n6561), .B(n6562), .Z(n6486) );
  AND U6516 ( .A(n6563), .B(n6564), .Z(n6562) );
  XOR U6517 ( .A(n6561), .B(n6565), .Z(n6563) );
  XNOR U6518 ( .A(n6566), .B(n6491), .Z(n6494) );
  XOR U6519 ( .A(n6567), .B(n6568), .Z(n6491) );
  AND U6520 ( .A(n6569), .B(n6570), .Z(n6568) );
  XNOR U6521 ( .A(n6571), .B(n6572), .Z(n6569) );
  IV U6522 ( .A(n6567), .Z(n6571) );
  XNOR U6523 ( .A(n6573), .B(n6574), .Z(n6566) );
  NOR U6524 ( .A(n6575), .B(n6576), .Z(n6574) );
  XNOR U6525 ( .A(n6573), .B(n6577), .Z(n6575) );
  XOR U6526 ( .A(n6500), .B(n6499), .Z(n6490) );
  XNOR U6527 ( .A(n6578), .B(n6496), .Z(n6499) );
  XOR U6528 ( .A(n6579), .B(n6580), .Z(n6496) );
  AND U6529 ( .A(n6581), .B(n6582), .Z(n6580) );
  XNOR U6530 ( .A(n6583), .B(n6584), .Z(n6581) );
  IV U6531 ( .A(n6579), .Z(n6583) );
  XNOR U6532 ( .A(n6585), .B(n6586), .Z(n6578) );
  NOR U6533 ( .A(n6587), .B(n6588), .Z(n6586) );
  XNOR U6534 ( .A(n6585), .B(n6589), .Z(n6587) );
  XOR U6535 ( .A(n6590), .B(n6591), .Z(n6500) );
  NOR U6536 ( .A(n6592), .B(n6593), .Z(n6591) );
  XNOR U6537 ( .A(n6590), .B(n6594), .Z(n6592) );
  XNOR U6538 ( .A(n6399), .B(n6503), .Z(n6505) );
  XNOR U6539 ( .A(n6595), .B(n6596), .Z(n6399) );
  AND U6540 ( .A(n166), .B(n6406), .Z(n6596) );
  XOR U6541 ( .A(n6595), .B(n6404), .Z(n6406) );
  AND U6542 ( .A(n6407), .B(n6410), .Z(n6503) );
  XOR U6543 ( .A(n6597), .B(n6554), .Z(n6410) );
  XNOR U6544 ( .A(p_input[288]), .B(p_input[512]), .Z(n6554) );
  XNOR U6545 ( .A(n6530), .B(n6529), .Z(n6597) );
  XNOR U6546 ( .A(n6598), .B(n6541), .Z(n6529) );
  XOR U6547 ( .A(n6515), .B(n6513), .Z(n6541) );
  XNOR U6548 ( .A(n6599), .B(n6520), .Z(n6513) );
  XOR U6549 ( .A(p_input[312]), .B(p_input[536]), .Z(n6520) );
  XOR U6550 ( .A(n6510), .B(n6519), .Z(n6599) );
  XOR U6551 ( .A(n6600), .B(n6516), .Z(n6519) );
  XOR U6552 ( .A(p_input[310]), .B(p_input[534]), .Z(n6516) );
  XOR U6553 ( .A(p_input[311]), .B(n4010), .Z(n6600) );
  XOR U6554 ( .A(p_input[306]), .B(p_input[530]), .Z(n6510) );
  XNOR U6555 ( .A(n6525), .B(n6524), .Z(n6515) );
  XOR U6556 ( .A(n6601), .B(n6521), .Z(n6524) );
  XOR U6557 ( .A(p_input[307]), .B(p_input[531]), .Z(n6521) );
  XOR U6558 ( .A(p_input[308]), .B(n4012), .Z(n6601) );
  XOR U6559 ( .A(p_input[309]), .B(p_input[533]), .Z(n6525) );
  XOR U6560 ( .A(n6540), .B(n6602), .Z(n6598) );
  IV U6561 ( .A(n6526), .Z(n6602) );
  XOR U6562 ( .A(p_input[289]), .B(p_input[513]), .Z(n6526) );
  XNOR U6563 ( .A(n6603), .B(n6548), .Z(n6540) );
  XNOR U6564 ( .A(n6536), .B(n6535), .Z(n6548) );
  XNOR U6565 ( .A(n6604), .B(n6532), .Z(n6535) );
  XNOR U6566 ( .A(p_input[314]), .B(p_input[538]), .Z(n6532) );
  XOR U6567 ( .A(p_input[315]), .B(n4016), .Z(n6604) );
  XOR U6568 ( .A(p_input[316]), .B(p_input[540]), .Z(n6536) );
  XOR U6569 ( .A(n6546), .B(n6605), .Z(n6603) );
  IV U6570 ( .A(n6537), .Z(n6605) );
  XOR U6571 ( .A(p_input[305]), .B(p_input[529]), .Z(n6537) );
  XNOR U6572 ( .A(n6606), .B(n6553), .Z(n6546) );
  XNOR U6573 ( .A(p_input[319]), .B(n4019), .Z(n6553) );
  XOR U6574 ( .A(n6543), .B(n6552), .Z(n6606) );
  XOR U6575 ( .A(n6607), .B(n6549), .Z(n6552) );
  XOR U6576 ( .A(p_input[317]), .B(p_input[541]), .Z(n6549) );
  XOR U6577 ( .A(p_input[318]), .B(n4021), .Z(n6607) );
  XOR U6578 ( .A(p_input[313]), .B(p_input[537]), .Z(n6543) );
  XOR U6579 ( .A(n6565), .B(n6564), .Z(n6530) );
  XNOR U6580 ( .A(n6608), .B(n6572), .Z(n6564) );
  XNOR U6581 ( .A(n6560), .B(n6559), .Z(n6572) );
  XNOR U6582 ( .A(n6609), .B(n6556), .Z(n6559) );
  XNOR U6583 ( .A(p_input[299]), .B(p_input[523]), .Z(n6556) );
  XOR U6584 ( .A(p_input[300]), .B(n4024), .Z(n6609) );
  XOR U6585 ( .A(p_input[301]), .B(p_input[525]), .Z(n6560) );
  XOR U6586 ( .A(n6570), .B(n6610), .Z(n6608) );
  IV U6587 ( .A(n6561), .Z(n6610) );
  XOR U6588 ( .A(p_input[290]), .B(p_input[514]), .Z(n6561) );
  XNOR U6589 ( .A(n6611), .B(n6577), .Z(n6570) );
  XNOR U6590 ( .A(p_input[304]), .B(n4027), .Z(n6577) );
  XOR U6591 ( .A(n6567), .B(n6576), .Z(n6611) );
  XOR U6592 ( .A(n6612), .B(n6573), .Z(n6576) );
  XOR U6593 ( .A(p_input[302]), .B(p_input[526]), .Z(n6573) );
  XOR U6594 ( .A(p_input[303]), .B(n4029), .Z(n6612) );
  XOR U6595 ( .A(p_input[298]), .B(p_input[522]), .Z(n6567) );
  XOR U6596 ( .A(n6584), .B(n6582), .Z(n6565) );
  XNOR U6597 ( .A(n6613), .B(n6589), .Z(n6582) );
  XOR U6598 ( .A(p_input[297]), .B(p_input[521]), .Z(n6589) );
  XOR U6599 ( .A(n6579), .B(n6588), .Z(n6613) );
  XOR U6600 ( .A(n6614), .B(n6585), .Z(n6588) );
  XOR U6601 ( .A(p_input[295]), .B(p_input[519]), .Z(n6585) );
  XOR U6602 ( .A(p_input[296]), .B(n4318), .Z(n6614) );
  XOR U6603 ( .A(p_input[291]), .B(p_input[515]), .Z(n6579) );
  XNOR U6604 ( .A(n6594), .B(n6593), .Z(n6584) );
  XOR U6605 ( .A(n6615), .B(n6590), .Z(n6593) );
  XOR U6606 ( .A(p_input[292]), .B(p_input[516]), .Z(n6590) );
  XOR U6607 ( .A(p_input[293]), .B(n4320), .Z(n6615) );
  XOR U6608 ( .A(p_input[294]), .B(p_input[518]), .Z(n6594) );
  XNOR U6609 ( .A(n6616), .B(n6617), .Z(n6407) );
  AND U6610 ( .A(n166), .B(n6618), .Z(n6617) );
  XNOR U6611 ( .A(n6619), .B(n6620), .Z(n166) );
  AND U6612 ( .A(n6621), .B(n6622), .Z(n6620) );
  XNOR U6613 ( .A(n6619), .B(n6360), .Z(n6622) );
  XOR U6614 ( .A(n6619), .B(n6357), .Z(n6621) );
  XOR U6615 ( .A(n6623), .B(n6624), .Z(n6619) );
  AND U6616 ( .A(n6625), .B(n6626), .Z(n6624) );
  XNOR U6617 ( .A(n6430), .B(n6623), .Z(n6626) );
  XOR U6618 ( .A(n6623), .B(n6371), .Z(n6625) );
  XOR U6619 ( .A(n6627), .B(n6628), .Z(n6623) );
  AND U6620 ( .A(n6629), .B(n6630), .Z(n6628) );
  XNOR U6621 ( .A(n6455), .B(n6627), .Z(n6630) );
  XOR U6622 ( .A(n6627), .B(n6382), .Z(n6629) );
  XOR U6623 ( .A(n6631), .B(n6632), .Z(n6627) );
  AND U6624 ( .A(n6633), .B(n6634), .Z(n6632) );
  XOR U6625 ( .A(n6631), .B(n6392), .Z(n6633) );
  XOR U6626 ( .A(n6635), .B(n6636), .Z(n6346) );
  AND U6627 ( .A(n170), .B(n6618), .Z(n6636) );
  XNOR U6628 ( .A(n6616), .B(n6635), .Z(n6618) );
  XNOR U6629 ( .A(n6637), .B(n6638), .Z(n170) );
  AND U6630 ( .A(n6639), .B(n6640), .Z(n6638) );
  XNOR U6631 ( .A(n6360), .B(n6637), .Z(n6640) );
  XOR U6632 ( .A(n6641), .B(n6642), .Z(n6360) );
  AND U6633 ( .A(n6643), .B(n173), .Z(n6642) );
  NOR U6634 ( .A(n6644), .B(n6641), .Z(n6643) );
  XOR U6635 ( .A(n6637), .B(n6357), .Z(n6639) );
  IV U6636 ( .A(n6361), .Z(n6357) );
  AND U6637 ( .A(n6645), .B(n6646), .Z(n6361) );
  XOR U6638 ( .A(n6647), .B(n6648), .Z(n6637) );
  AND U6639 ( .A(n6649), .B(n6650), .Z(n6648) );
  XNOR U6640 ( .A(n6647), .B(n6430), .Z(n6650) );
  XNOR U6641 ( .A(n6651), .B(n6652), .Z(n6430) );
  AND U6642 ( .A(n173), .B(n6653), .Z(n6652) );
  XOR U6643 ( .A(n6654), .B(n6651), .Z(n6653) );
  XNOR U6644 ( .A(n6655), .B(n6647), .Z(n6649) );
  IV U6645 ( .A(n6371), .Z(n6655) );
  XOR U6646 ( .A(n6656), .B(n6657), .Z(n6371) );
  AND U6647 ( .A(n181), .B(n6658), .Z(n6657) );
  XOR U6648 ( .A(n6659), .B(n6660), .Z(n6647) );
  AND U6649 ( .A(n6661), .B(n6662), .Z(n6660) );
  XNOR U6650 ( .A(n6659), .B(n6455), .Z(n6662) );
  XNOR U6651 ( .A(n6663), .B(n6664), .Z(n6455) );
  AND U6652 ( .A(n173), .B(n6665), .Z(n6664) );
  XNOR U6653 ( .A(n6666), .B(n6663), .Z(n6665) );
  XOR U6654 ( .A(n6382), .B(n6659), .Z(n6661) );
  XOR U6655 ( .A(n6667), .B(n6668), .Z(n6382) );
  AND U6656 ( .A(n181), .B(n6669), .Z(n6668) );
  XOR U6657 ( .A(n6631), .B(n6670), .Z(n6659) );
  AND U6658 ( .A(n6671), .B(n6634), .Z(n6670) );
  XNOR U6659 ( .A(n6501), .B(n6631), .Z(n6634) );
  XNOR U6660 ( .A(n6672), .B(n6673), .Z(n6501) );
  AND U6661 ( .A(n173), .B(n6674), .Z(n6673) );
  XOR U6662 ( .A(n6675), .B(n6672), .Z(n6674) );
  XNOR U6663 ( .A(n6676), .B(n6631), .Z(n6671) );
  IV U6664 ( .A(n6392), .Z(n6676) );
  XOR U6665 ( .A(n6677), .B(n6678), .Z(n6392) );
  AND U6666 ( .A(n181), .B(n6679), .Z(n6678) );
  XOR U6667 ( .A(n6680), .B(n6681), .Z(n6631) );
  AND U6668 ( .A(n6682), .B(n6683), .Z(n6681) );
  XNOR U6669 ( .A(n6680), .B(n6595), .Z(n6683) );
  XNOR U6670 ( .A(n6684), .B(n6685), .Z(n6595) );
  AND U6671 ( .A(n173), .B(n6686), .Z(n6685) );
  XNOR U6672 ( .A(n6687), .B(n6684), .Z(n6686) );
  XNOR U6673 ( .A(n6688), .B(n6680), .Z(n6682) );
  IV U6674 ( .A(n6404), .Z(n6688) );
  XOR U6675 ( .A(n6689), .B(n6690), .Z(n6404) );
  AND U6676 ( .A(n181), .B(n6691), .Z(n6690) );
  AND U6677 ( .A(n6635), .B(n6616), .Z(n6680) );
  XNOR U6678 ( .A(n6692), .B(n6693), .Z(n6616) );
  AND U6679 ( .A(n173), .B(n6694), .Z(n6693) );
  XNOR U6680 ( .A(n6695), .B(n6692), .Z(n6694) );
  XNOR U6681 ( .A(n6696), .B(n6697), .Z(n173) );
  NOR U6682 ( .A(n6698), .B(n6699), .Z(n6697) );
  XNOR U6683 ( .A(n6696), .B(n6641), .Z(n6699) );
  NOR U6684 ( .A(n6645), .B(n6646), .Z(n6641) );
  NOR U6685 ( .A(n6696), .B(n6644), .Z(n6698) );
  AND U6686 ( .A(n6700), .B(n6701), .Z(n6644) );
  XOR U6687 ( .A(n6702), .B(n6703), .Z(n6696) );
  AND U6688 ( .A(n6704), .B(n6705), .Z(n6703) );
  XNOR U6689 ( .A(n6702), .B(n6700), .Z(n6705) );
  IV U6690 ( .A(n6654), .Z(n6700) );
  XOR U6691 ( .A(n6706), .B(n6707), .Z(n6654) );
  XOR U6692 ( .A(n6708), .B(n6701), .Z(n6707) );
  AND U6693 ( .A(n6666), .B(n6709), .Z(n6701) );
  AND U6694 ( .A(n6710), .B(n6711), .Z(n6708) );
  XOR U6695 ( .A(n6712), .B(n6706), .Z(n6710) );
  XNOR U6696 ( .A(n6651), .B(n6702), .Z(n6704) );
  XNOR U6697 ( .A(n6713), .B(n6714), .Z(n6651) );
  AND U6698 ( .A(n177), .B(n6658), .Z(n6714) );
  XOR U6699 ( .A(n6713), .B(n6656), .Z(n6658) );
  XOR U6700 ( .A(n6715), .B(n6716), .Z(n6702) );
  AND U6701 ( .A(n6717), .B(n6718), .Z(n6716) );
  XNOR U6702 ( .A(n6715), .B(n6666), .Z(n6718) );
  XOR U6703 ( .A(n6719), .B(n6711), .Z(n6666) );
  XNOR U6704 ( .A(n6720), .B(n6706), .Z(n6711) );
  XOR U6705 ( .A(n6721), .B(n6722), .Z(n6706) );
  AND U6706 ( .A(n6723), .B(n6724), .Z(n6722) );
  XOR U6707 ( .A(n6725), .B(n6721), .Z(n6723) );
  XNOR U6708 ( .A(n6726), .B(n6727), .Z(n6720) );
  AND U6709 ( .A(n6728), .B(n6729), .Z(n6727) );
  XOR U6710 ( .A(n6726), .B(n6730), .Z(n6728) );
  XNOR U6711 ( .A(n6712), .B(n6709), .Z(n6719) );
  AND U6712 ( .A(n6731), .B(n6732), .Z(n6709) );
  XOR U6713 ( .A(n6733), .B(n6734), .Z(n6712) );
  AND U6714 ( .A(n6735), .B(n6736), .Z(n6734) );
  XOR U6715 ( .A(n6733), .B(n6737), .Z(n6735) );
  XNOR U6716 ( .A(n6663), .B(n6715), .Z(n6717) );
  XNOR U6717 ( .A(n6738), .B(n6739), .Z(n6663) );
  AND U6718 ( .A(n177), .B(n6669), .Z(n6739) );
  XOR U6719 ( .A(n6738), .B(n6667), .Z(n6669) );
  XOR U6720 ( .A(n6740), .B(n6741), .Z(n6715) );
  AND U6721 ( .A(n6742), .B(n6743), .Z(n6741) );
  XNOR U6722 ( .A(n6740), .B(n6731), .Z(n6743) );
  IV U6723 ( .A(n6675), .Z(n6731) );
  XNOR U6724 ( .A(n6744), .B(n6724), .Z(n6675) );
  XNOR U6725 ( .A(n6745), .B(n6730), .Z(n6724) );
  XOR U6726 ( .A(n6746), .B(n6747), .Z(n6730) );
  AND U6727 ( .A(n6748), .B(n6749), .Z(n6747) );
  XOR U6728 ( .A(n6746), .B(n6750), .Z(n6748) );
  XNOR U6729 ( .A(n6729), .B(n6721), .Z(n6745) );
  XOR U6730 ( .A(n6751), .B(n6752), .Z(n6721) );
  AND U6731 ( .A(n6753), .B(n6754), .Z(n6752) );
  XNOR U6732 ( .A(n6755), .B(n6751), .Z(n6753) );
  XNOR U6733 ( .A(n6756), .B(n6726), .Z(n6729) );
  XOR U6734 ( .A(n6757), .B(n6758), .Z(n6726) );
  AND U6735 ( .A(n6759), .B(n6760), .Z(n6758) );
  XOR U6736 ( .A(n6757), .B(n6761), .Z(n6759) );
  XNOR U6737 ( .A(n6762), .B(n6763), .Z(n6756) );
  AND U6738 ( .A(n6764), .B(n6765), .Z(n6763) );
  XNOR U6739 ( .A(n6762), .B(n6766), .Z(n6764) );
  XNOR U6740 ( .A(n6725), .B(n6732), .Z(n6744) );
  AND U6741 ( .A(n6687), .B(n6767), .Z(n6732) );
  XOR U6742 ( .A(n6737), .B(n6736), .Z(n6725) );
  XNOR U6743 ( .A(n6768), .B(n6733), .Z(n6736) );
  XOR U6744 ( .A(n6769), .B(n6770), .Z(n6733) );
  AND U6745 ( .A(n6771), .B(n6772), .Z(n6770) );
  XOR U6746 ( .A(n6769), .B(n6773), .Z(n6771) );
  XNOR U6747 ( .A(n6774), .B(n6775), .Z(n6768) );
  AND U6748 ( .A(n6776), .B(n6777), .Z(n6775) );
  XOR U6749 ( .A(n6774), .B(n6778), .Z(n6776) );
  XOR U6750 ( .A(n6779), .B(n6780), .Z(n6737) );
  AND U6751 ( .A(n6781), .B(n6782), .Z(n6780) );
  XOR U6752 ( .A(n6779), .B(n6783), .Z(n6781) );
  XNOR U6753 ( .A(n6672), .B(n6740), .Z(n6742) );
  XNOR U6754 ( .A(n6784), .B(n6785), .Z(n6672) );
  AND U6755 ( .A(n177), .B(n6679), .Z(n6785) );
  XOR U6756 ( .A(n6784), .B(n6677), .Z(n6679) );
  XOR U6757 ( .A(n6786), .B(n6787), .Z(n6740) );
  AND U6758 ( .A(n6788), .B(n6789), .Z(n6787) );
  XNOR U6759 ( .A(n6786), .B(n6687), .Z(n6789) );
  XOR U6760 ( .A(n6790), .B(n6754), .Z(n6687) );
  XNOR U6761 ( .A(n6791), .B(n6761), .Z(n6754) );
  XOR U6762 ( .A(n6750), .B(n6749), .Z(n6761) );
  XNOR U6763 ( .A(n6792), .B(n6746), .Z(n6749) );
  XOR U6764 ( .A(n6793), .B(n6794), .Z(n6746) );
  AND U6765 ( .A(n6795), .B(n6796), .Z(n6794) );
  XNOR U6766 ( .A(n6797), .B(n6798), .Z(n6795) );
  IV U6767 ( .A(n6793), .Z(n6797) );
  XNOR U6768 ( .A(n6799), .B(n6800), .Z(n6792) );
  NOR U6769 ( .A(n6801), .B(n6802), .Z(n6800) );
  XNOR U6770 ( .A(n6799), .B(n6803), .Z(n6801) );
  XOR U6771 ( .A(n6804), .B(n6805), .Z(n6750) );
  NOR U6772 ( .A(n6806), .B(n6807), .Z(n6805) );
  XNOR U6773 ( .A(n6804), .B(n6808), .Z(n6806) );
  XNOR U6774 ( .A(n6760), .B(n6751), .Z(n6791) );
  XOR U6775 ( .A(n6809), .B(n6810), .Z(n6751) );
  AND U6776 ( .A(n6811), .B(n6812), .Z(n6810) );
  XOR U6777 ( .A(n6809), .B(n6813), .Z(n6811) );
  XOR U6778 ( .A(n6814), .B(n6766), .Z(n6760) );
  XOR U6779 ( .A(n6815), .B(n6816), .Z(n6766) );
  NOR U6780 ( .A(n6817), .B(n6818), .Z(n6816) );
  XOR U6781 ( .A(n6815), .B(n6819), .Z(n6817) );
  XNOR U6782 ( .A(n6765), .B(n6757), .Z(n6814) );
  XOR U6783 ( .A(n6820), .B(n6821), .Z(n6757) );
  AND U6784 ( .A(n6822), .B(n6823), .Z(n6821) );
  XOR U6785 ( .A(n6820), .B(n6824), .Z(n6822) );
  XNOR U6786 ( .A(n6825), .B(n6762), .Z(n6765) );
  XOR U6787 ( .A(n6826), .B(n6827), .Z(n6762) );
  AND U6788 ( .A(n6828), .B(n6829), .Z(n6827) );
  XNOR U6789 ( .A(n6830), .B(n6831), .Z(n6828) );
  IV U6790 ( .A(n6826), .Z(n6830) );
  XNOR U6791 ( .A(n6832), .B(n6833), .Z(n6825) );
  NOR U6792 ( .A(n6834), .B(n6835), .Z(n6833) );
  XNOR U6793 ( .A(n6832), .B(n6836), .Z(n6834) );
  XOR U6794 ( .A(n6755), .B(n6767), .Z(n6790) );
  NOR U6795 ( .A(n6695), .B(n6837), .Z(n6767) );
  XNOR U6796 ( .A(n6773), .B(n6772), .Z(n6755) );
  XNOR U6797 ( .A(n6838), .B(n6778), .Z(n6772) );
  XNOR U6798 ( .A(n6839), .B(n6840), .Z(n6778) );
  NOR U6799 ( .A(n6841), .B(n6842), .Z(n6840) );
  XOR U6800 ( .A(n6839), .B(n6843), .Z(n6841) );
  XNOR U6801 ( .A(n6777), .B(n6769), .Z(n6838) );
  XOR U6802 ( .A(n6844), .B(n6845), .Z(n6769) );
  AND U6803 ( .A(n6846), .B(n6847), .Z(n6845) );
  XOR U6804 ( .A(n6844), .B(n6848), .Z(n6846) );
  XNOR U6805 ( .A(n6849), .B(n6774), .Z(n6777) );
  XOR U6806 ( .A(n6850), .B(n6851), .Z(n6774) );
  AND U6807 ( .A(n6852), .B(n6853), .Z(n6851) );
  XNOR U6808 ( .A(n6854), .B(n6855), .Z(n6852) );
  IV U6809 ( .A(n6850), .Z(n6854) );
  XNOR U6810 ( .A(n6856), .B(n6857), .Z(n6849) );
  NOR U6811 ( .A(n6858), .B(n6859), .Z(n6857) );
  XNOR U6812 ( .A(n6856), .B(n6860), .Z(n6858) );
  XOR U6813 ( .A(n6783), .B(n6782), .Z(n6773) );
  XNOR U6814 ( .A(n6861), .B(n6779), .Z(n6782) );
  XOR U6815 ( .A(n6862), .B(n6863), .Z(n6779) );
  AND U6816 ( .A(n6864), .B(n6865), .Z(n6863) );
  XNOR U6817 ( .A(n6866), .B(n6867), .Z(n6864) );
  IV U6818 ( .A(n6862), .Z(n6866) );
  XNOR U6819 ( .A(n6868), .B(n6869), .Z(n6861) );
  NOR U6820 ( .A(n6870), .B(n6871), .Z(n6869) );
  XNOR U6821 ( .A(n6868), .B(n6872), .Z(n6870) );
  XOR U6822 ( .A(n6873), .B(n6874), .Z(n6783) );
  NOR U6823 ( .A(n6875), .B(n6876), .Z(n6874) );
  XNOR U6824 ( .A(n6873), .B(n6877), .Z(n6875) );
  XNOR U6825 ( .A(n6684), .B(n6786), .Z(n6788) );
  XNOR U6826 ( .A(n6878), .B(n6879), .Z(n6684) );
  AND U6827 ( .A(n177), .B(n6691), .Z(n6879) );
  XOR U6828 ( .A(n6878), .B(n6689), .Z(n6691) );
  AND U6829 ( .A(n6692), .B(n6695), .Z(n6786) );
  XOR U6830 ( .A(n6880), .B(n6837), .Z(n6695) );
  XNOR U6831 ( .A(p_input[320]), .B(p_input[512]), .Z(n6837) );
  XNOR U6832 ( .A(n6813), .B(n6812), .Z(n6880) );
  XNOR U6833 ( .A(n6881), .B(n6824), .Z(n6812) );
  XOR U6834 ( .A(n6798), .B(n6796), .Z(n6824) );
  XNOR U6835 ( .A(n6882), .B(n6803), .Z(n6796) );
  XOR U6836 ( .A(p_input[344]), .B(p_input[536]), .Z(n6803) );
  XOR U6837 ( .A(n6793), .B(n6802), .Z(n6882) );
  XOR U6838 ( .A(n6883), .B(n6799), .Z(n6802) );
  XOR U6839 ( .A(p_input[342]), .B(p_input[534]), .Z(n6799) );
  XOR U6840 ( .A(p_input[343]), .B(n4010), .Z(n6883) );
  XOR U6841 ( .A(p_input[338]), .B(p_input[530]), .Z(n6793) );
  XNOR U6842 ( .A(n6808), .B(n6807), .Z(n6798) );
  XOR U6843 ( .A(n6884), .B(n6804), .Z(n6807) );
  XOR U6844 ( .A(p_input[339]), .B(p_input[531]), .Z(n6804) );
  XOR U6845 ( .A(p_input[340]), .B(n4012), .Z(n6884) );
  XOR U6846 ( .A(p_input[341]), .B(p_input[533]), .Z(n6808) );
  XOR U6847 ( .A(n6823), .B(n6885), .Z(n6881) );
  IV U6848 ( .A(n6809), .Z(n6885) );
  XOR U6849 ( .A(p_input[321]), .B(p_input[513]), .Z(n6809) );
  XNOR U6850 ( .A(n6886), .B(n6831), .Z(n6823) );
  XNOR U6851 ( .A(n6819), .B(n6818), .Z(n6831) );
  XNOR U6852 ( .A(n6887), .B(n6815), .Z(n6818) );
  XNOR U6853 ( .A(p_input[346]), .B(p_input[538]), .Z(n6815) );
  XOR U6854 ( .A(p_input[347]), .B(n4016), .Z(n6887) );
  XOR U6855 ( .A(p_input[348]), .B(p_input[540]), .Z(n6819) );
  XOR U6856 ( .A(n6829), .B(n6888), .Z(n6886) );
  IV U6857 ( .A(n6820), .Z(n6888) );
  XOR U6858 ( .A(p_input[337]), .B(p_input[529]), .Z(n6820) );
  XNOR U6859 ( .A(n6889), .B(n6836), .Z(n6829) );
  XNOR U6860 ( .A(p_input[351]), .B(n4019), .Z(n6836) );
  XOR U6861 ( .A(n6826), .B(n6835), .Z(n6889) );
  XOR U6862 ( .A(n6890), .B(n6832), .Z(n6835) );
  XOR U6863 ( .A(p_input[349]), .B(p_input[541]), .Z(n6832) );
  XOR U6864 ( .A(p_input[350]), .B(n4021), .Z(n6890) );
  XOR U6865 ( .A(p_input[345]), .B(p_input[537]), .Z(n6826) );
  XOR U6866 ( .A(n6848), .B(n6847), .Z(n6813) );
  XNOR U6867 ( .A(n6891), .B(n6855), .Z(n6847) );
  XNOR U6868 ( .A(n6843), .B(n6842), .Z(n6855) );
  XNOR U6869 ( .A(n6892), .B(n6839), .Z(n6842) );
  XNOR U6870 ( .A(p_input[331]), .B(p_input[523]), .Z(n6839) );
  XOR U6871 ( .A(p_input[332]), .B(n4024), .Z(n6892) );
  XOR U6872 ( .A(p_input[333]), .B(p_input[525]), .Z(n6843) );
  XOR U6873 ( .A(n6853), .B(n6893), .Z(n6891) );
  IV U6874 ( .A(n6844), .Z(n6893) );
  XOR U6875 ( .A(p_input[322]), .B(p_input[514]), .Z(n6844) );
  XNOR U6876 ( .A(n6894), .B(n6860), .Z(n6853) );
  XNOR U6877 ( .A(p_input[336]), .B(n4027), .Z(n6860) );
  XOR U6878 ( .A(n6850), .B(n6859), .Z(n6894) );
  XOR U6879 ( .A(n6895), .B(n6856), .Z(n6859) );
  XOR U6880 ( .A(p_input[334]), .B(p_input[526]), .Z(n6856) );
  XOR U6881 ( .A(p_input[335]), .B(n4029), .Z(n6895) );
  XOR U6882 ( .A(p_input[330]), .B(p_input[522]), .Z(n6850) );
  XOR U6883 ( .A(n6867), .B(n6865), .Z(n6848) );
  XNOR U6884 ( .A(n6896), .B(n6872), .Z(n6865) );
  XOR U6885 ( .A(p_input[329]), .B(p_input[521]), .Z(n6872) );
  XOR U6886 ( .A(n6862), .B(n6871), .Z(n6896) );
  XOR U6887 ( .A(n6897), .B(n6868), .Z(n6871) );
  XOR U6888 ( .A(p_input[327]), .B(p_input[519]), .Z(n6868) );
  XOR U6889 ( .A(p_input[328]), .B(n4318), .Z(n6897) );
  XOR U6890 ( .A(p_input[323]), .B(p_input[515]), .Z(n6862) );
  XNOR U6891 ( .A(n6877), .B(n6876), .Z(n6867) );
  XOR U6892 ( .A(n6898), .B(n6873), .Z(n6876) );
  XOR U6893 ( .A(p_input[324]), .B(p_input[516]), .Z(n6873) );
  XOR U6894 ( .A(p_input[325]), .B(n4320), .Z(n6898) );
  XOR U6895 ( .A(p_input[326]), .B(p_input[518]), .Z(n6877) );
  XNOR U6896 ( .A(n6899), .B(n6900), .Z(n6692) );
  AND U6897 ( .A(n177), .B(n6901), .Z(n6900) );
  XNOR U6898 ( .A(n6902), .B(n6903), .Z(n177) );
  NOR U6899 ( .A(n6904), .B(n6905), .Z(n6903) );
  XOR U6900 ( .A(n6646), .B(n6902), .Z(n6905) );
  NOR U6901 ( .A(n6902), .B(n6645), .Z(n6904) );
  XOR U6902 ( .A(n6906), .B(n6907), .Z(n6902) );
  AND U6903 ( .A(n6908), .B(n6909), .Z(n6907) );
  XNOR U6904 ( .A(n6713), .B(n6906), .Z(n6909) );
  XOR U6905 ( .A(n6906), .B(n6656), .Z(n6908) );
  XOR U6906 ( .A(n6910), .B(n6911), .Z(n6906) );
  AND U6907 ( .A(n6912), .B(n6913), .Z(n6911) );
  XNOR U6908 ( .A(n6738), .B(n6910), .Z(n6913) );
  XOR U6909 ( .A(n6910), .B(n6667), .Z(n6912) );
  XOR U6910 ( .A(n6914), .B(n6915), .Z(n6910) );
  AND U6911 ( .A(n6916), .B(n6917), .Z(n6915) );
  XOR U6912 ( .A(n6914), .B(n6677), .Z(n6916) );
  XOR U6913 ( .A(n6918), .B(n6919), .Z(n6635) );
  AND U6914 ( .A(n181), .B(n6901), .Z(n6919) );
  XNOR U6915 ( .A(n6899), .B(n6918), .Z(n6901) );
  XNOR U6916 ( .A(n6920), .B(n6921), .Z(n181) );
  NOR U6917 ( .A(n6922), .B(n6923), .Z(n6921) );
  XNOR U6918 ( .A(n6646), .B(n6924), .Z(n6923) );
  IV U6919 ( .A(n6920), .Z(n6924) );
  AND U6920 ( .A(n6925), .B(n6926), .Z(n6646) );
  NOR U6921 ( .A(n6920), .B(n6645), .Z(n6922) );
  AND U6922 ( .A(n6927), .B(n6928), .Z(n6645) );
  IV U6923 ( .A(n6929), .Z(n6927) );
  XOR U6924 ( .A(n6930), .B(n6931), .Z(n6920) );
  AND U6925 ( .A(n6932), .B(n6933), .Z(n6931) );
  XNOR U6926 ( .A(n6930), .B(n6713), .Z(n6933) );
  XNOR U6927 ( .A(n6934), .B(n6935), .Z(n6713) );
  AND U6928 ( .A(n184), .B(n6936), .Z(n6935) );
  XOR U6929 ( .A(n6937), .B(n6934), .Z(n6936) );
  XNOR U6930 ( .A(n6938), .B(n6930), .Z(n6932) );
  IV U6931 ( .A(n6656), .Z(n6938) );
  XOR U6932 ( .A(n6939), .B(n6940), .Z(n6656) );
  AND U6933 ( .A(n192), .B(n6941), .Z(n6940) );
  XOR U6934 ( .A(n6942), .B(n6943), .Z(n6930) );
  AND U6935 ( .A(n6944), .B(n6945), .Z(n6943) );
  XNOR U6936 ( .A(n6942), .B(n6738), .Z(n6945) );
  XNOR U6937 ( .A(n6946), .B(n6947), .Z(n6738) );
  AND U6938 ( .A(n184), .B(n6948), .Z(n6947) );
  XNOR U6939 ( .A(n6949), .B(n6946), .Z(n6948) );
  XOR U6940 ( .A(n6667), .B(n6942), .Z(n6944) );
  XOR U6941 ( .A(n6950), .B(n6951), .Z(n6667) );
  AND U6942 ( .A(n192), .B(n6952), .Z(n6951) );
  XOR U6943 ( .A(n6914), .B(n6953), .Z(n6942) );
  AND U6944 ( .A(n6954), .B(n6917), .Z(n6953) );
  XNOR U6945 ( .A(n6784), .B(n6914), .Z(n6917) );
  XNOR U6946 ( .A(n6955), .B(n6956), .Z(n6784) );
  AND U6947 ( .A(n184), .B(n6957), .Z(n6956) );
  XOR U6948 ( .A(n6958), .B(n6955), .Z(n6957) );
  XNOR U6949 ( .A(n6959), .B(n6914), .Z(n6954) );
  IV U6950 ( .A(n6677), .Z(n6959) );
  XOR U6951 ( .A(n6960), .B(n6961), .Z(n6677) );
  AND U6952 ( .A(n192), .B(n6962), .Z(n6961) );
  XOR U6953 ( .A(n6963), .B(n6964), .Z(n6914) );
  AND U6954 ( .A(n6965), .B(n6966), .Z(n6964) );
  XNOR U6955 ( .A(n6963), .B(n6878), .Z(n6966) );
  XNOR U6956 ( .A(n6967), .B(n6968), .Z(n6878) );
  AND U6957 ( .A(n184), .B(n6969), .Z(n6968) );
  XNOR U6958 ( .A(n6970), .B(n6967), .Z(n6969) );
  XNOR U6959 ( .A(n6971), .B(n6963), .Z(n6965) );
  IV U6960 ( .A(n6689), .Z(n6971) );
  XOR U6961 ( .A(n6972), .B(n6973), .Z(n6689) );
  AND U6962 ( .A(n192), .B(n6974), .Z(n6973) );
  AND U6963 ( .A(n6918), .B(n6899), .Z(n6963) );
  XNOR U6964 ( .A(n6975), .B(n6976), .Z(n6899) );
  AND U6965 ( .A(n184), .B(n6977), .Z(n6976) );
  XNOR U6966 ( .A(n6978), .B(n6975), .Z(n6977) );
  XNOR U6967 ( .A(n6979), .B(n6980), .Z(n184) );
  NOR U6968 ( .A(n6981), .B(n6982), .Z(n6980) );
  XNOR U6969 ( .A(n6979), .B(n6929), .Z(n6982) );
  NOR U6970 ( .A(n6925), .B(n6926), .Z(n6929) );
  NOR U6971 ( .A(n6979), .B(n6928), .Z(n6981) );
  AND U6972 ( .A(n6983), .B(n6984), .Z(n6928) );
  XOR U6973 ( .A(n6985), .B(n6986), .Z(n6979) );
  AND U6974 ( .A(n6987), .B(n6988), .Z(n6986) );
  XNOR U6975 ( .A(n6985), .B(n6983), .Z(n6988) );
  IV U6976 ( .A(n6937), .Z(n6983) );
  XOR U6977 ( .A(n6989), .B(n6990), .Z(n6937) );
  XOR U6978 ( .A(n6991), .B(n6984), .Z(n6990) );
  AND U6979 ( .A(n6949), .B(n6992), .Z(n6984) );
  AND U6980 ( .A(n6993), .B(n6994), .Z(n6991) );
  XOR U6981 ( .A(n6995), .B(n6989), .Z(n6993) );
  XNOR U6982 ( .A(n6934), .B(n6985), .Z(n6987) );
  XNOR U6983 ( .A(n6996), .B(n6997), .Z(n6934) );
  AND U6984 ( .A(n188), .B(n6941), .Z(n6997) );
  XOR U6985 ( .A(n6996), .B(n6939), .Z(n6941) );
  XOR U6986 ( .A(n6998), .B(n6999), .Z(n6985) );
  AND U6987 ( .A(n7000), .B(n7001), .Z(n6999) );
  XNOR U6988 ( .A(n6998), .B(n6949), .Z(n7001) );
  XOR U6989 ( .A(n7002), .B(n6994), .Z(n6949) );
  XNOR U6990 ( .A(n7003), .B(n6989), .Z(n6994) );
  XOR U6991 ( .A(n7004), .B(n7005), .Z(n6989) );
  AND U6992 ( .A(n7006), .B(n7007), .Z(n7005) );
  XOR U6993 ( .A(n7008), .B(n7004), .Z(n7006) );
  XNOR U6994 ( .A(n7009), .B(n7010), .Z(n7003) );
  AND U6995 ( .A(n7011), .B(n7012), .Z(n7010) );
  XOR U6996 ( .A(n7009), .B(n7013), .Z(n7011) );
  XNOR U6997 ( .A(n6995), .B(n6992), .Z(n7002) );
  AND U6998 ( .A(n7014), .B(n7015), .Z(n6992) );
  XOR U6999 ( .A(n7016), .B(n7017), .Z(n6995) );
  AND U7000 ( .A(n7018), .B(n7019), .Z(n7017) );
  XOR U7001 ( .A(n7016), .B(n7020), .Z(n7018) );
  XNOR U7002 ( .A(n6946), .B(n6998), .Z(n7000) );
  XNOR U7003 ( .A(n7021), .B(n7022), .Z(n6946) );
  AND U7004 ( .A(n188), .B(n6952), .Z(n7022) );
  XOR U7005 ( .A(n7021), .B(n6950), .Z(n6952) );
  XOR U7006 ( .A(n7023), .B(n7024), .Z(n6998) );
  AND U7007 ( .A(n7025), .B(n7026), .Z(n7024) );
  XNOR U7008 ( .A(n7023), .B(n7014), .Z(n7026) );
  IV U7009 ( .A(n6958), .Z(n7014) );
  XNOR U7010 ( .A(n7027), .B(n7007), .Z(n6958) );
  XNOR U7011 ( .A(n7028), .B(n7013), .Z(n7007) );
  XOR U7012 ( .A(n7029), .B(n7030), .Z(n7013) );
  AND U7013 ( .A(n7031), .B(n7032), .Z(n7030) );
  XOR U7014 ( .A(n7029), .B(n7033), .Z(n7031) );
  XNOR U7015 ( .A(n7012), .B(n7004), .Z(n7028) );
  XOR U7016 ( .A(n7034), .B(n7035), .Z(n7004) );
  AND U7017 ( .A(n7036), .B(n7037), .Z(n7035) );
  XNOR U7018 ( .A(n7038), .B(n7034), .Z(n7036) );
  XNOR U7019 ( .A(n7039), .B(n7009), .Z(n7012) );
  XOR U7020 ( .A(n7040), .B(n7041), .Z(n7009) );
  AND U7021 ( .A(n7042), .B(n7043), .Z(n7041) );
  XOR U7022 ( .A(n7040), .B(n7044), .Z(n7042) );
  XNOR U7023 ( .A(n7045), .B(n7046), .Z(n7039) );
  AND U7024 ( .A(n7047), .B(n7048), .Z(n7046) );
  XNOR U7025 ( .A(n7045), .B(n7049), .Z(n7047) );
  XNOR U7026 ( .A(n7008), .B(n7015), .Z(n7027) );
  AND U7027 ( .A(n6970), .B(n7050), .Z(n7015) );
  XOR U7028 ( .A(n7020), .B(n7019), .Z(n7008) );
  XNOR U7029 ( .A(n7051), .B(n7016), .Z(n7019) );
  XOR U7030 ( .A(n7052), .B(n7053), .Z(n7016) );
  AND U7031 ( .A(n7054), .B(n7055), .Z(n7053) );
  XOR U7032 ( .A(n7052), .B(n7056), .Z(n7054) );
  XNOR U7033 ( .A(n7057), .B(n7058), .Z(n7051) );
  AND U7034 ( .A(n7059), .B(n7060), .Z(n7058) );
  XOR U7035 ( .A(n7057), .B(n7061), .Z(n7059) );
  XOR U7036 ( .A(n7062), .B(n7063), .Z(n7020) );
  AND U7037 ( .A(n7064), .B(n7065), .Z(n7063) );
  XOR U7038 ( .A(n7062), .B(n7066), .Z(n7064) );
  XNOR U7039 ( .A(n6955), .B(n7023), .Z(n7025) );
  XNOR U7040 ( .A(n7067), .B(n7068), .Z(n6955) );
  AND U7041 ( .A(n188), .B(n6962), .Z(n7068) );
  XOR U7042 ( .A(n7067), .B(n6960), .Z(n6962) );
  XOR U7043 ( .A(n7069), .B(n7070), .Z(n7023) );
  AND U7044 ( .A(n7071), .B(n7072), .Z(n7070) );
  XNOR U7045 ( .A(n7069), .B(n6970), .Z(n7072) );
  XOR U7046 ( .A(n7073), .B(n7037), .Z(n6970) );
  XNOR U7047 ( .A(n7074), .B(n7044), .Z(n7037) );
  XOR U7048 ( .A(n7033), .B(n7032), .Z(n7044) );
  XNOR U7049 ( .A(n7075), .B(n7029), .Z(n7032) );
  XOR U7050 ( .A(n7076), .B(n7077), .Z(n7029) );
  AND U7051 ( .A(n7078), .B(n7079), .Z(n7077) );
  XNOR U7052 ( .A(n7080), .B(n7081), .Z(n7078) );
  IV U7053 ( .A(n7076), .Z(n7080) );
  XNOR U7054 ( .A(n7082), .B(n7083), .Z(n7075) );
  NOR U7055 ( .A(n7084), .B(n7085), .Z(n7083) );
  XNOR U7056 ( .A(n7082), .B(n7086), .Z(n7084) );
  XOR U7057 ( .A(n7087), .B(n7088), .Z(n7033) );
  NOR U7058 ( .A(n7089), .B(n7090), .Z(n7088) );
  XNOR U7059 ( .A(n7087), .B(n7091), .Z(n7089) );
  XNOR U7060 ( .A(n7043), .B(n7034), .Z(n7074) );
  XOR U7061 ( .A(n7092), .B(n7093), .Z(n7034) );
  AND U7062 ( .A(n7094), .B(n7095), .Z(n7093) );
  XOR U7063 ( .A(n7092), .B(n7096), .Z(n7094) );
  XOR U7064 ( .A(n7097), .B(n7049), .Z(n7043) );
  XOR U7065 ( .A(n7098), .B(n7099), .Z(n7049) );
  NOR U7066 ( .A(n7100), .B(n7101), .Z(n7099) );
  XOR U7067 ( .A(n7098), .B(n7102), .Z(n7100) );
  XNOR U7068 ( .A(n7048), .B(n7040), .Z(n7097) );
  XOR U7069 ( .A(n7103), .B(n7104), .Z(n7040) );
  AND U7070 ( .A(n7105), .B(n7106), .Z(n7104) );
  XOR U7071 ( .A(n7103), .B(n7107), .Z(n7105) );
  XNOR U7072 ( .A(n7108), .B(n7045), .Z(n7048) );
  XOR U7073 ( .A(n7109), .B(n7110), .Z(n7045) );
  AND U7074 ( .A(n7111), .B(n7112), .Z(n7110) );
  XNOR U7075 ( .A(n7113), .B(n7114), .Z(n7111) );
  IV U7076 ( .A(n7109), .Z(n7113) );
  XNOR U7077 ( .A(n7115), .B(n7116), .Z(n7108) );
  NOR U7078 ( .A(n7117), .B(n7118), .Z(n7116) );
  XNOR U7079 ( .A(n7115), .B(n7119), .Z(n7117) );
  XOR U7080 ( .A(n7038), .B(n7050), .Z(n7073) );
  NOR U7081 ( .A(n6978), .B(n7120), .Z(n7050) );
  XNOR U7082 ( .A(n7056), .B(n7055), .Z(n7038) );
  XNOR U7083 ( .A(n7121), .B(n7061), .Z(n7055) );
  XNOR U7084 ( .A(n7122), .B(n7123), .Z(n7061) );
  NOR U7085 ( .A(n7124), .B(n7125), .Z(n7123) );
  XOR U7086 ( .A(n7122), .B(n7126), .Z(n7124) );
  XNOR U7087 ( .A(n7060), .B(n7052), .Z(n7121) );
  XOR U7088 ( .A(n7127), .B(n7128), .Z(n7052) );
  AND U7089 ( .A(n7129), .B(n7130), .Z(n7128) );
  XOR U7090 ( .A(n7127), .B(n7131), .Z(n7129) );
  XNOR U7091 ( .A(n7132), .B(n7057), .Z(n7060) );
  XOR U7092 ( .A(n7133), .B(n7134), .Z(n7057) );
  AND U7093 ( .A(n7135), .B(n7136), .Z(n7134) );
  XNOR U7094 ( .A(n7137), .B(n7138), .Z(n7135) );
  IV U7095 ( .A(n7133), .Z(n7137) );
  XNOR U7096 ( .A(n7139), .B(n7140), .Z(n7132) );
  NOR U7097 ( .A(n7141), .B(n7142), .Z(n7140) );
  XNOR U7098 ( .A(n7139), .B(n7143), .Z(n7141) );
  XOR U7099 ( .A(n7066), .B(n7065), .Z(n7056) );
  XNOR U7100 ( .A(n7144), .B(n7062), .Z(n7065) );
  XOR U7101 ( .A(n7145), .B(n7146), .Z(n7062) );
  AND U7102 ( .A(n7147), .B(n7148), .Z(n7146) );
  XNOR U7103 ( .A(n7149), .B(n7150), .Z(n7147) );
  IV U7104 ( .A(n7145), .Z(n7149) );
  XNOR U7105 ( .A(n7151), .B(n7152), .Z(n7144) );
  NOR U7106 ( .A(n7153), .B(n7154), .Z(n7152) );
  XNOR U7107 ( .A(n7151), .B(n7155), .Z(n7153) );
  XOR U7108 ( .A(n7156), .B(n7157), .Z(n7066) );
  NOR U7109 ( .A(n7158), .B(n7159), .Z(n7157) );
  XNOR U7110 ( .A(n7156), .B(n7160), .Z(n7158) );
  XNOR U7111 ( .A(n6967), .B(n7069), .Z(n7071) );
  XNOR U7112 ( .A(n7161), .B(n7162), .Z(n6967) );
  AND U7113 ( .A(n188), .B(n6974), .Z(n7162) );
  XOR U7114 ( .A(n7161), .B(n6972), .Z(n6974) );
  AND U7115 ( .A(n6975), .B(n6978), .Z(n7069) );
  XOR U7116 ( .A(n7163), .B(n7120), .Z(n6978) );
  XNOR U7117 ( .A(p_input[352]), .B(p_input[512]), .Z(n7120) );
  XNOR U7118 ( .A(n7096), .B(n7095), .Z(n7163) );
  XNOR U7119 ( .A(n7164), .B(n7107), .Z(n7095) );
  XOR U7120 ( .A(n7081), .B(n7079), .Z(n7107) );
  XNOR U7121 ( .A(n7165), .B(n7086), .Z(n7079) );
  XOR U7122 ( .A(p_input[376]), .B(p_input[536]), .Z(n7086) );
  XOR U7123 ( .A(n7076), .B(n7085), .Z(n7165) );
  XOR U7124 ( .A(n7166), .B(n7082), .Z(n7085) );
  XOR U7125 ( .A(p_input[374]), .B(p_input[534]), .Z(n7082) );
  XOR U7126 ( .A(p_input[375]), .B(n4010), .Z(n7166) );
  XOR U7127 ( .A(p_input[370]), .B(p_input[530]), .Z(n7076) );
  XNOR U7128 ( .A(n7091), .B(n7090), .Z(n7081) );
  XOR U7129 ( .A(n7167), .B(n7087), .Z(n7090) );
  XOR U7130 ( .A(p_input[371]), .B(p_input[531]), .Z(n7087) );
  XOR U7131 ( .A(p_input[372]), .B(n4012), .Z(n7167) );
  XOR U7132 ( .A(p_input[373]), .B(p_input[533]), .Z(n7091) );
  XOR U7133 ( .A(n7106), .B(n7168), .Z(n7164) );
  IV U7134 ( .A(n7092), .Z(n7168) );
  XOR U7135 ( .A(p_input[353]), .B(p_input[513]), .Z(n7092) );
  XNOR U7136 ( .A(n7169), .B(n7114), .Z(n7106) );
  XNOR U7137 ( .A(n7102), .B(n7101), .Z(n7114) );
  XNOR U7138 ( .A(n7170), .B(n7098), .Z(n7101) );
  XNOR U7139 ( .A(p_input[378]), .B(p_input[538]), .Z(n7098) );
  XOR U7140 ( .A(p_input[379]), .B(n4016), .Z(n7170) );
  XOR U7141 ( .A(p_input[380]), .B(p_input[540]), .Z(n7102) );
  XOR U7142 ( .A(n7112), .B(n7171), .Z(n7169) );
  IV U7143 ( .A(n7103), .Z(n7171) );
  XOR U7144 ( .A(p_input[369]), .B(p_input[529]), .Z(n7103) );
  XNOR U7145 ( .A(n7172), .B(n7119), .Z(n7112) );
  XNOR U7146 ( .A(p_input[383]), .B(n4019), .Z(n7119) );
  XOR U7147 ( .A(n7109), .B(n7118), .Z(n7172) );
  XOR U7148 ( .A(n7173), .B(n7115), .Z(n7118) );
  XOR U7149 ( .A(p_input[381]), .B(p_input[541]), .Z(n7115) );
  XOR U7150 ( .A(p_input[382]), .B(n4021), .Z(n7173) );
  XOR U7151 ( .A(p_input[377]), .B(p_input[537]), .Z(n7109) );
  XOR U7152 ( .A(n7131), .B(n7130), .Z(n7096) );
  XNOR U7153 ( .A(n7174), .B(n7138), .Z(n7130) );
  XNOR U7154 ( .A(n7126), .B(n7125), .Z(n7138) );
  XNOR U7155 ( .A(n7175), .B(n7122), .Z(n7125) );
  XNOR U7156 ( .A(p_input[363]), .B(p_input[523]), .Z(n7122) );
  XOR U7157 ( .A(p_input[364]), .B(n4024), .Z(n7175) );
  XOR U7158 ( .A(p_input[365]), .B(p_input[525]), .Z(n7126) );
  XOR U7159 ( .A(n7136), .B(n7176), .Z(n7174) );
  IV U7160 ( .A(n7127), .Z(n7176) );
  XOR U7161 ( .A(p_input[354]), .B(p_input[514]), .Z(n7127) );
  XNOR U7162 ( .A(n7177), .B(n7143), .Z(n7136) );
  XNOR U7163 ( .A(p_input[368]), .B(n4027), .Z(n7143) );
  XOR U7164 ( .A(n7133), .B(n7142), .Z(n7177) );
  XOR U7165 ( .A(n7178), .B(n7139), .Z(n7142) );
  XOR U7166 ( .A(p_input[366]), .B(p_input[526]), .Z(n7139) );
  XOR U7167 ( .A(p_input[367]), .B(n4029), .Z(n7178) );
  XOR U7168 ( .A(p_input[362]), .B(p_input[522]), .Z(n7133) );
  XOR U7169 ( .A(n7150), .B(n7148), .Z(n7131) );
  XNOR U7170 ( .A(n7179), .B(n7155), .Z(n7148) );
  XOR U7171 ( .A(p_input[361]), .B(p_input[521]), .Z(n7155) );
  XOR U7172 ( .A(n7145), .B(n7154), .Z(n7179) );
  XOR U7173 ( .A(n7180), .B(n7151), .Z(n7154) );
  XOR U7174 ( .A(p_input[359]), .B(p_input[519]), .Z(n7151) );
  XOR U7175 ( .A(p_input[360]), .B(n4318), .Z(n7180) );
  XOR U7176 ( .A(p_input[355]), .B(p_input[515]), .Z(n7145) );
  XNOR U7177 ( .A(n7160), .B(n7159), .Z(n7150) );
  XOR U7178 ( .A(n7181), .B(n7156), .Z(n7159) );
  XOR U7179 ( .A(p_input[356]), .B(p_input[516]), .Z(n7156) );
  XOR U7180 ( .A(p_input[357]), .B(n4320), .Z(n7181) );
  XOR U7181 ( .A(p_input[358]), .B(p_input[518]), .Z(n7160) );
  XNOR U7182 ( .A(n7182), .B(n7183), .Z(n6975) );
  AND U7183 ( .A(n188), .B(n7184), .Z(n7183) );
  XNOR U7184 ( .A(n7185), .B(n7186), .Z(n188) );
  NOR U7185 ( .A(n7187), .B(n7188), .Z(n7186) );
  XOR U7186 ( .A(n6926), .B(n7185), .Z(n7188) );
  NOR U7187 ( .A(n7185), .B(n6925), .Z(n7187) );
  XOR U7188 ( .A(n7189), .B(n7190), .Z(n7185) );
  AND U7189 ( .A(n7191), .B(n7192), .Z(n7190) );
  XNOR U7190 ( .A(n6996), .B(n7189), .Z(n7192) );
  XOR U7191 ( .A(n7189), .B(n6939), .Z(n7191) );
  XOR U7192 ( .A(n7193), .B(n7194), .Z(n7189) );
  AND U7193 ( .A(n7195), .B(n7196), .Z(n7194) );
  XNOR U7194 ( .A(n7021), .B(n7193), .Z(n7196) );
  XOR U7195 ( .A(n7193), .B(n6950), .Z(n7195) );
  XOR U7196 ( .A(n7197), .B(n7198), .Z(n7193) );
  AND U7197 ( .A(n7199), .B(n7200), .Z(n7198) );
  XOR U7198 ( .A(n7197), .B(n6960), .Z(n7199) );
  XOR U7199 ( .A(n7201), .B(n7202), .Z(n6918) );
  AND U7200 ( .A(n192), .B(n7184), .Z(n7202) );
  XNOR U7201 ( .A(n7182), .B(n7201), .Z(n7184) );
  XNOR U7202 ( .A(n7203), .B(n7204), .Z(n192) );
  NOR U7203 ( .A(n7205), .B(n7206), .Z(n7204) );
  XNOR U7204 ( .A(n6926), .B(n7207), .Z(n7206) );
  IV U7205 ( .A(n7203), .Z(n7207) );
  AND U7206 ( .A(n7208), .B(n7209), .Z(n6926) );
  NOR U7207 ( .A(n7203), .B(n6925), .Z(n7205) );
  AND U7208 ( .A(n7210), .B(n7211), .Z(n6925) );
  IV U7209 ( .A(n7212), .Z(n7210) );
  XOR U7210 ( .A(n7213), .B(n7214), .Z(n7203) );
  AND U7211 ( .A(n7215), .B(n7216), .Z(n7214) );
  XNOR U7212 ( .A(n7213), .B(n6996), .Z(n7216) );
  XNOR U7213 ( .A(n7217), .B(n7218), .Z(n6996) );
  AND U7214 ( .A(n195), .B(n7219), .Z(n7218) );
  XOR U7215 ( .A(n7220), .B(n7217), .Z(n7219) );
  XNOR U7216 ( .A(n7221), .B(n7213), .Z(n7215) );
  IV U7217 ( .A(n6939), .Z(n7221) );
  XOR U7218 ( .A(n7222), .B(n7223), .Z(n6939) );
  AND U7219 ( .A(n203), .B(n7224), .Z(n7223) );
  XOR U7220 ( .A(n7225), .B(n7226), .Z(n7213) );
  AND U7221 ( .A(n7227), .B(n7228), .Z(n7226) );
  XNOR U7222 ( .A(n7225), .B(n7021), .Z(n7228) );
  XNOR U7223 ( .A(n7229), .B(n7230), .Z(n7021) );
  AND U7224 ( .A(n195), .B(n7231), .Z(n7230) );
  XNOR U7225 ( .A(n7232), .B(n7229), .Z(n7231) );
  XOR U7226 ( .A(n6950), .B(n7225), .Z(n7227) );
  XOR U7227 ( .A(n7233), .B(n7234), .Z(n6950) );
  AND U7228 ( .A(n203), .B(n7235), .Z(n7234) );
  XOR U7229 ( .A(n7197), .B(n7236), .Z(n7225) );
  AND U7230 ( .A(n7237), .B(n7200), .Z(n7236) );
  XNOR U7231 ( .A(n7067), .B(n7197), .Z(n7200) );
  XNOR U7232 ( .A(n7238), .B(n7239), .Z(n7067) );
  AND U7233 ( .A(n195), .B(n7240), .Z(n7239) );
  XOR U7234 ( .A(n7241), .B(n7238), .Z(n7240) );
  XNOR U7235 ( .A(n7242), .B(n7197), .Z(n7237) );
  IV U7236 ( .A(n6960), .Z(n7242) );
  XOR U7237 ( .A(n7243), .B(n7244), .Z(n6960) );
  AND U7238 ( .A(n203), .B(n7245), .Z(n7244) );
  XOR U7239 ( .A(n7246), .B(n7247), .Z(n7197) );
  AND U7240 ( .A(n7248), .B(n7249), .Z(n7247) );
  XNOR U7241 ( .A(n7246), .B(n7161), .Z(n7249) );
  XNOR U7242 ( .A(n7250), .B(n7251), .Z(n7161) );
  AND U7243 ( .A(n195), .B(n7252), .Z(n7251) );
  XNOR U7244 ( .A(n7253), .B(n7250), .Z(n7252) );
  XNOR U7245 ( .A(n7254), .B(n7246), .Z(n7248) );
  IV U7246 ( .A(n6972), .Z(n7254) );
  XOR U7247 ( .A(n7255), .B(n7256), .Z(n6972) );
  AND U7248 ( .A(n203), .B(n7257), .Z(n7256) );
  AND U7249 ( .A(n7201), .B(n7182), .Z(n7246) );
  XNOR U7250 ( .A(n7258), .B(n7259), .Z(n7182) );
  AND U7251 ( .A(n195), .B(n7260), .Z(n7259) );
  XNOR U7252 ( .A(n7261), .B(n7258), .Z(n7260) );
  XNOR U7253 ( .A(n7262), .B(n7263), .Z(n195) );
  NOR U7254 ( .A(n7264), .B(n7265), .Z(n7263) );
  XNOR U7255 ( .A(n7262), .B(n7212), .Z(n7265) );
  NOR U7256 ( .A(n7208), .B(n7209), .Z(n7212) );
  NOR U7257 ( .A(n7262), .B(n7211), .Z(n7264) );
  AND U7258 ( .A(n7266), .B(n7267), .Z(n7211) );
  XOR U7259 ( .A(n7268), .B(n7269), .Z(n7262) );
  AND U7260 ( .A(n7270), .B(n7271), .Z(n7269) );
  XNOR U7261 ( .A(n7268), .B(n7266), .Z(n7271) );
  IV U7262 ( .A(n7220), .Z(n7266) );
  XOR U7263 ( .A(n7272), .B(n7273), .Z(n7220) );
  XOR U7264 ( .A(n7274), .B(n7267), .Z(n7273) );
  AND U7265 ( .A(n7232), .B(n7275), .Z(n7267) );
  AND U7266 ( .A(n7276), .B(n7277), .Z(n7274) );
  XOR U7267 ( .A(n7278), .B(n7272), .Z(n7276) );
  XNOR U7268 ( .A(n7217), .B(n7268), .Z(n7270) );
  XNOR U7269 ( .A(n7279), .B(n7280), .Z(n7217) );
  AND U7270 ( .A(n199), .B(n7224), .Z(n7280) );
  XOR U7271 ( .A(n7279), .B(n7222), .Z(n7224) );
  XOR U7272 ( .A(n7281), .B(n7282), .Z(n7268) );
  AND U7273 ( .A(n7283), .B(n7284), .Z(n7282) );
  XNOR U7274 ( .A(n7281), .B(n7232), .Z(n7284) );
  XOR U7275 ( .A(n7285), .B(n7277), .Z(n7232) );
  XNOR U7276 ( .A(n7286), .B(n7272), .Z(n7277) );
  XOR U7277 ( .A(n7287), .B(n7288), .Z(n7272) );
  AND U7278 ( .A(n7289), .B(n7290), .Z(n7288) );
  XOR U7279 ( .A(n7291), .B(n7287), .Z(n7289) );
  XNOR U7280 ( .A(n7292), .B(n7293), .Z(n7286) );
  AND U7281 ( .A(n7294), .B(n7295), .Z(n7293) );
  XOR U7282 ( .A(n7292), .B(n7296), .Z(n7294) );
  XNOR U7283 ( .A(n7278), .B(n7275), .Z(n7285) );
  AND U7284 ( .A(n7297), .B(n7298), .Z(n7275) );
  XOR U7285 ( .A(n7299), .B(n7300), .Z(n7278) );
  AND U7286 ( .A(n7301), .B(n7302), .Z(n7300) );
  XOR U7287 ( .A(n7299), .B(n7303), .Z(n7301) );
  XNOR U7288 ( .A(n7229), .B(n7281), .Z(n7283) );
  XNOR U7289 ( .A(n7304), .B(n7305), .Z(n7229) );
  AND U7290 ( .A(n199), .B(n7235), .Z(n7305) );
  XOR U7291 ( .A(n7304), .B(n7233), .Z(n7235) );
  XOR U7292 ( .A(n7306), .B(n7307), .Z(n7281) );
  AND U7293 ( .A(n7308), .B(n7309), .Z(n7307) );
  XNOR U7294 ( .A(n7306), .B(n7297), .Z(n7309) );
  IV U7295 ( .A(n7241), .Z(n7297) );
  XNOR U7296 ( .A(n7310), .B(n7290), .Z(n7241) );
  XNOR U7297 ( .A(n7311), .B(n7296), .Z(n7290) );
  XOR U7298 ( .A(n7312), .B(n7313), .Z(n7296) );
  AND U7299 ( .A(n7314), .B(n7315), .Z(n7313) );
  XOR U7300 ( .A(n7312), .B(n7316), .Z(n7314) );
  XNOR U7301 ( .A(n7295), .B(n7287), .Z(n7311) );
  XOR U7302 ( .A(n7317), .B(n7318), .Z(n7287) );
  AND U7303 ( .A(n7319), .B(n7320), .Z(n7318) );
  XNOR U7304 ( .A(n7321), .B(n7317), .Z(n7319) );
  XNOR U7305 ( .A(n7322), .B(n7292), .Z(n7295) );
  XOR U7306 ( .A(n7323), .B(n7324), .Z(n7292) );
  AND U7307 ( .A(n7325), .B(n7326), .Z(n7324) );
  XOR U7308 ( .A(n7323), .B(n7327), .Z(n7325) );
  XNOR U7309 ( .A(n7328), .B(n7329), .Z(n7322) );
  AND U7310 ( .A(n7330), .B(n7331), .Z(n7329) );
  XNOR U7311 ( .A(n7328), .B(n7332), .Z(n7330) );
  XNOR U7312 ( .A(n7291), .B(n7298), .Z(n7310) );
  AND U7313 ( .A(n7253), .B(n7333), .Z(n7298) );
  XOR U7314 ( .A(n7303), .B(n7302), .Z(n7291) );
  XNOR U7315 ( .A(n7334), .B(n7299), .Z(n7302) );
  XOR U7316 ( .A(n7335), .B(n7336), .Z(n7299) );
  AND U7317 ( .A(n7337), .B(n7338), .Z(n7336) );
  XOR U7318 ( .A(n7335), .B(n7339), .Z(n7337) );
  XNOR U7319 ( .A(n7340), .B(n7341), .Z(n7334) );
  AND U7320 ( .A(n7342), .B(n7343), .Z(n7341) );
  XOR U7321 ( .A(n7340), .B(n7344), .Z(n7342) );
  XOR U7322 ( .A(n7345), .B(n7346), .Z(n7303) );
  AND U7323 ( .A(n7347), .B(n7348), .Z(n7346) );
  XOR U7324 ( .A(n7345), .B(n7349), .Z(n7347) );
  XNOR U7325 ( .A(n7238), .B(n7306), .Z(n7308) );
  XNOR U7326 ( .A(n7350), .B(n7351), .Z(n7238) );
  AND U7327 ( .A(n199), .B(n7245), .Z(n7351) );
  XOR U7328 ( .A(n7350), .B(n7243), .Z(n7245) );
  XOR U7329 ( .A(n7352), .B(n7353), .Z(n7306) );
  AND U7330 ( .A(n7354), .B(n7355), .Z(n7353) );
  XNOR U7331 ( .A(n7352), .B(n7253), .Z(n7355) );
  XOR U7332 ( .A(n7356), .B(n7320), .Z(n7253) );
  XNOR U7333 ( .A(n7357), .B(n7327), .Z(n7320) );
  XOR U7334 ( .A(n7316), .B(n7315), .Z(n7327) );
  XNOR U7335 ( .A(n7358), .B(n7312), .Z(n7315) );
  XOR U7336 ( .A(n7359), .B(n7360), .Z(n7312) );
  AND U7337 ( .A(n7361), .B(n7362), .Z(n7360) );
  XNOR U7338 ( .A(n7363), .B(n7364), .Z(n7361) );
  IV U7339 ( .A(n7359), .Z(n7363) );
  XNOR U7340 ( .A(n7365), .B(n7366), .Z(n7358) );
  NOR U7341 ( .A(n7367), .B(n7368), .Z(n7366) );
  XNOR U7342 ( .A(n7365), .B(n7369), .Z(n7367) );
  XOR U7343 ( .A(n7370), .B(n7371), .Z(n7316) );
  NOR U7344 ( .A(n7372), .B(n7373), .Z(n7371) );
  XNOR U7345 ( .A(n7370), .B(n7374), .Z(n7372) );
  XNOR U7346 ( .A(n7326), .B(n7317), .Z(n7357) );
  XOR U7347 ( .A(n7375), .B(n7376), .Z(n7317) );
  AND U7348 ( .A(n7377), .B(n7378), .Z(n7376) );
  XOR U7349 ( .A(n7375), .B(n7379), .Z(n7377) );
  XOR U7350 ( .A(n7380), .B(n7332), .Z(n7326) );
  XOR U7351 ( .A(n7381), .B(n7382), .Z(n7332) );
  NOR U7352 ( .A(n7383), .B(n7384), .Z(n7382) );
  XOR U7353 ( .A(n7381), .B(n7385), .Z(n7383) );
  XNOR U7354 ( .A(n7331), .B(n7323), .Z(n7380) );
  XOR U7355 ( .A(n7386), .B(n7387), .Z(n7323) );
  AND U7356 ( .A(n7388), .B(n7389), .Z(n7387) );
  XOR U7357 ( .A(n7386), .B(n7390), .Z(n7388) );
  XNOR U7358 ( .A(n7391), .B(n7328), .Z(n7331) );
  XOR U7359 ( .A(n7392), .B(n7393), .Z(n7328) );
  AND U7360 ( .A(n7394), .B(n7395), .Z(n7393) );
  XNOR U7361 ( .A(n7396), .B(n7397), .Z(n7394) );
  IV U7362 ( .A(n7392), .Z(n7396) );
  XNOR U7363 ( .A(n7398), .B(n7399), .Z(n7391) );
  NOR U7364 ( .A(n7400), .B(n7401), .Z(n7399) );
  XNOR U7365 ( .A(n7398), .B(n7402), .Z(n7400) );
  XOR U7366 ( .A(n7321), .B(n7333), .Z(n7356) );
  NOR U7367 ( .A(n7261), .B(n7403), .Z(n7333) );
  XNOR U7368 ( .A(n7339), .B(n7338), .Z(n7321) );
  XNOR U7369 ( .A(n7404), .B(n7344), .Z(n7338) );
  XNOR U7370 ( .A(n7405), .B(n7406), .Z(n7344) );
  NOR U7371 ( .A(n7407), .B(n7408), .Z(n7406) );
  XOR U7372 ( .A(n7405), .B(n7409), .Z(n7407) );
  XNOR U7373 ( .A(n7343), .B(n7335), .Z(n7404) );
  XOR U7374 ( .A(n7410), .B(n7411), .Z(n7335) );
  AND U7375 ( .A(n7412), .B(n7413), .Z(n7411) );
  XOR U7376 ( .A(n7410), .B(n7414), .Z(n7412) );
  XNOR U7377 ( .A(n7415), .B(n7340), .Z(n7343) );
  XOR U7378 ( .A(n7416), .B(n7417), .Z(n7340) );
  AND U7379 ( .A(n7418), .B(n7419), .Z(n7417) );
  XNOR U7380 ( .A(n7420), .B(n7421), .Z(n7418) );
  IV U7381 ( .A(n7416), .Z(n7420) );
  XNOR U7382 ( .A(n7422), .B(n7423), .Z(n7415) );
  NOR U7383 ( .A(n7424), .B(n7425), .Z(n7423) );
  XNOR U7384 ( .A(n7422), .B(n7426), .Z(n7424) );
  XOR U7385 ( .A(n7349), .B(n7348), .Z(n7339) );
  XNOR U7386 ( .A(n7427), .B(n7345), .Z(n7348) );
  XOR U7387 ( .A(n7428), .B(n7429), .Z(n7345) );
  AND U7388 ( .A(n7430), .B(n7431), .Z(n7429) );
  XNOR U7389 ( .A(n7432), .B(n7433), .Z(n7430) );
  IV U7390 ( .A(n7428), .Z(n7432) );
  XNOR U7391 ( .A(n7434), .B(n7435), .Z(n7427) );
  NOR U7392 ( .A(n7436), .B(n7437), .Z(n7435) );
  XNOR U7393 ( .A(n7434), .B(n7438), .Z(n7436) );
  XOR U7394 ( .A(n7439), .B(n7440), .Z(n7349) );
  NOR U7395 ( .A(n7441), .B(n7442), .Z(n7440) );
  XNOR U7396 ( .A(n7439), .B(n7443), .Z(n7441) );
  XNOR U7397 ( .A(n7250), .B(n7352), .Z(n7354) );
  XNOR U7398 ( .A(n7444), .B(n7445), .Z(n7250) );
  AND U7399 ( .A(n199), .B(n7257), .Z(n7445) );
  XOR U7400 ( .A(n7444), .B(n7255), .Z(n7257) );
  AND U7401 ( .A(n7258), .B(n7261), .Z(n7352) );
  XOR U7402 ( .A(n7446), .B(n7403), .Z(n7261) );
  XNOR U7403 ( .A(p_input[384]), .B(p_input[512]), .Z(n7403) );
  XNOR U7404 ( .A(n7379), .B(n7378), .Z(n7446) );
  XNOR U7405 ( .A(n7447), .B(n7390), .Z(n7378) );
  XOR U7406 ( .A(n7364), .B(n7362), .Z(n7390) );
  XNOR U7407 ( .A(n7448), .B(n7369), .Z(n7362) );
  XOR U7408 ( .A(p_input[408]), .B(p_input[536]), .Z(n7369) );
  XOR U7409 ( .A(n7359), .B(n7368), .Z(n7448) );
  XOR U7410 ( .A(n7449), .B(n7365), .Z(n7368) );
  XOR U7411 ( .A(p_input[406]), .B(p_input[534]), .Z(n7365) );
  XOR U7412 ( .A(p_input[407]), .B(n4010), .Z(n7449) );
  XOR U7413 ( .A(p_input[402]), .B(p_input[530]), .Z(n7359) );
  XNOR U7414 ( .A(n7374), .B(n7373), .Z(n7364) );
  XOR U7415 ( .A(n7450), .B(n7370), .Z(n7373) );
  XOR U7416 ( .A(p_input[403]), .B(p_input[531]), .Z(n7370) );
  XOR U7417 ( .A(p_input[404]), .B(n4012), .Z(n7450) );
  XOR U7418 ( .A(p_input[405]), .B(p_input[533]), .Z(n7374) );
  XOR U7419 ( .A(n7389), .B(n7451), .Z(n7447) );
  IV U7420 ( .A(n7375), .Z(n7451) );
  XOR U7421 ( .A(p_input[385]), .B(p_input[513]), .Z(n7375) );
  XNOR U7422 ( .A(n7452), .B(n7397), .Z(n7389) );
  XNOR U7423 ( .A(n7385), .B(n7384), .Z(n7397) );
  XNOR U7424 ( .A(n7453), .B(n7381), .Z(n7384) );
  XNOR U7425 ( .A(p_input[410]), .B(p_input[538]), .Z(n7381) );
  XOR U7426 ( .A(p_input[411]), .B(n4016), .Z(n7453) );
  XOR U7427 ( .A(p_input[412]), .B(p_input[540]), .Z(n7385) );
  XOR U7428 ( .A(n7395), .B(n7454), .Z(n7452) );
  IV U7429 ( .A(n7386), .Z(n7454) );
  XOR U7430 ( .A(p_input[401]), .B(p_input[529]), .Z(n7386) );
  XNOR U7431 ( .A(n7455), .B(n7402), .Z(n7395) );
  XNOR U7432 ( .A(p_input[415]), .B(n4019), .Z(n7402) );
  XOR U7433 ( .A(n7392), .B(n7401), .Z(n7455) );
  XOR U7434 ( .A(n7456), .B(n7398), .Z(n7401) );
  XOR U7435 ( .A(p_input[413]), .B(p_input[541]), .Z(n7398) );
  XOR U7436 ( .A(p_input[414]), .B(n4021), .Z(n7456) );
  XOR U7437 ( .A(p_input[409]), .B(p_input[537]), .Z(n7392) );
  XOR U7438 ( .A(n7414), .B(n7413), .Z(n7379) );
  XNOR U7439 ( .A(n7457), .B(n7421), .Z(n7413) );
  XNOR U7440 ( .A(n7409), .B(n7408), .Z(n7421) );
  XNOR U7441 ( .A(n7458), .B(n7405), .Z(n7408) );
  XNOR U7442 ( .A(p_input[395]), .B(p_input[523]), .Z(n7405) );
  XOR U7443 ( .A(p_input[396]), .B(n4024), .Z(n7458) );
  XOR U7444 ( .A(p_input[397]), .B(p_input[525]), .Z(n7409) );
  XOR U7445 ( .A(n7419), .B(n7459), .Z(n7457) );
  IV U7446 ( .A(n7410), .Z(n7459) );
  XOR U7447 ( .A(p_input[386]), .B(p_input[514]), .Z(n7410) );
  XNOR U7448 ( .A(n7460), .B(n7426), .Z(n7419) );
  XNOR U7449 ( .A(p_input[400]), .B(n4027), .Z(n7426) );
  XOR U7450 ( .A(n7416), .B(n7425), .Z(n7460) );
  XOR U7451 ( .A(n7461), .B(n7422), .Z(n7425) );
  XOR U7452 ( .A(p_input[398]), .B(p_input[526]), .Z(n7422) );
  XOR U7453 ( .A(p_input[399]), .B(n4029), .Z(n7461) );
  XOR U7454 ( .A(p_input[394]), .B(p_input[522]), .Z(n7416) );
  XOR U7455 ( .A(n7433), .B(n7431), .Z(n7414) );
  XNOR U7456 ( .A(n7462), .B(n7438), .Z(n7431) );
  XOR U7457 ( .A(p_input[393]), .B(p_input[521]), .Z(n7438) );
  XOR U7458 ( .A(n7428), .B(n7437), .Z(n7462) );
  XOR U7459 ( .A(n7463), .B(n7434), .Z(n7437) );
  XOR U7460 ( .A(p_input[391]), .B(p_input[519]), .Z(n7434) );
  XOR U7461 ( .A(p_input[392]), .B(n4318), .Z(n7463) );
  XOR U7462 ( .A(p_input[387]), .B(p_input[515]), .Z(n7428) );
  XNOR U7463 ( .A(n7443), .B(n7442), .Z(n7433) );
  XOR U7464 ( .A(n7464), .B(n7439), .Z(n7442) );
  XOR U7465 ( .A(p_input[388]), .B(p_input[516]), .Z(n7439) );
  XOR U7466 ( .A(p_input[389]), .B(n4320), .Z(n7464) );
  XOR U7467 ( .A(p_input[390]), .B(p_input[518]), .Z(n7443) );
  XNOR U7468 ( .A(n7465), .B(n7466), .Z(n7258) );
  AND U7469 ( .A(n199), .B(n7467), .Z(n7466) );
  XNOR U7470 ( .A(n7468), .B(n7469), .Z(n199) );
  NOR U7471 ( .A(n7470), .B(n7471), .Z(n7469) );
  XOR U7472 ( .A(n7209), .B(n7468), .Z(n7471) );
  NOR U7473 ( .A(n7468), .B(n7208), .Z(n7470) );
  XOR U7474 ( .A(n7472), .B(n7473), .Z(n7468) );
  AND U7475 ( .A(n7474), .B(n7475), .Z(n7473) );
  XNOR U7476 ( .A(n7279), .B(n7472), .Z(n7475) );
  XOR U7477 ( .A(n7472), .B(n7222), .Z(n7474) );
  XOR U7478 ( .A(n7476), .B(n7477), .Z(n7472) );
  AND U7479 ( .A(n7478), .B(n7479), .Z(n7477) );
  XNOR U7480 ( .A(n7304), .B(n7476), .Z(n7479) );
  XOR U7481 ( .A(n7476), .B(n7233), .Z(n7478) );
  XOR U7482 ( .A(n7480), .B(n7481), .Z(n7476) );
  AND U7483 ( .A(n7482), .B(n7483), .Z(n7481) );
  XOR U7484 ( .A(n7480), .B(n7243), .Z(n7482) );
  XOR U7485 ( .A(n7484), .B(n7485), .Z(n7201) );
  AND U7486 ( .A(n203), .B(n7467), .Z(n7485) );
  XNOR U7487 ( .A(n7465), .B(n7484), .Z(n7467) );
  XNOR U7488 ( .A(n7486), .B(n7487), .Z(n203) );
  NOR U7489 ( .A(n7488), .B(n7489), .Z(n7487) );
  XNOR U7490 ( .A(n7209), .B(n7490), .Z(n7489) );
  IV U7491 ( .A(n7486), .Z(n7490) );
  AND U7492 ( .A(n7491), .B(n7492), .Z(n7209) );
  NOR U7493 ( .A(n7486), .B(n7208), .Z(n7488) );
  AND U7494 ( .A(n7493), .B(n7494), .Z(n7208) );
  IV U7495 ( .A(n7495), .Z(n7493) );
  XOR U7496 ( .A(n7496), .B(n7497), .Z(n7486) );
  AND U7497 ( .A(n7498), .B(n7499), .Z(n7497) );
  XNOR U7498 ( .A(n7496), .B(n7279), .Z(n7499) );
  XNOR U7499 ( .A(n7500), .B(n7501), .Z(n7279) );
  AND U7500 ( .A(n206), .B(n7502), .Z(n7501) );
  XOR U7501 ( .A(n7503), .B(n7500), .Z(n7502) );
  XNOR U7502 ( .A(n7504), .B(n7496), .Z(n7498) );
  IV U7503 ( .A(n7222), .Z(n7504) );
  XOR U7504 ( .A(n7505), .B(n7506), .Z(n7222) );
  AND U7505 ( .A(n213), .B(n7507), .Z(n7506) );
  XOR U7506 ( .A(n7508), .B(n7509), .Z(n7496) );
  AND U7507 ( .A(n7510), .B(n7511), .Z(n7509) );
  XNOR U7508 ( .A(n7508), .B(n7304), .Z(n7511) );
  XNOR U7509 ( .A(n7512), .B(n7513), .Z(n7304) );
  AND U7510 ( .A(n206), .B(n7514), .Z(n7513) );
  XNOR U7511 ( .A(n7515), .B(n7512), .Z(n7514) );
  XOR U7512 ( .A(n7233), .B(n7508), .Z(n7510) );
  XOR U7513 ( .A(n7516), .B(n7517), .Z(n7233) );
  AND U7514 ( .A(n213), .B(n7518), .Z(n7517) );
  XOR U7515 ( .A(n7480), .B(n7519), .Z(n7508) );
  AND U7516 ( .A(n7520), .B(n7483), .Z(n7519) );
  XNOR U7517 ( .A(n7350), .B(n7480), .Z(n7483) );
  XNOR U7518 ( .A(n7521), .B(n7522), .Z(n7350) );
  AND U7519 ( .A(n206), .B(n7523), .Z(n7522) );
  XOR U7520 ( .A(n7524), .B(n7521), .Z(n7523) );
  XNOR U7521 ( .A(n7525), .B(n7480), .Z(n7520) );
  IV U7522 ( .A(n7243), .Z(n7525) );
  XOR U7523 ( .A(n7526), .B(n7527), .Z(n7243) );
  AND U7524 ( .A(n213), .B(n7528), .Z(n7527) );
  XOR U7525 ( .A(n7529), .B(n7530), .Z(n7480) );
  AND U7526 ( .A(n7531), .B(n7532), .Z(n7530) );
  XNOR U7527 ( .A(n7529), .B(n7444), .Z(n7532) );
  XNOR U7528 ( .A(n7533), .B(n7534), .Z(n7444) );
  AND U7529 ( .A(n206), .B(n7535), .Z(n7534) );
  XNOR U7530 ( .A(n7536), .B(n7533), .Z(n7535) );
  XNOR U7531 ( .A(n7537), .B(n7529), .Z(n7531) );
  IV U7532 ( .A(n7255), .Z(n7537) );
  XOR U7533 ( .A(n7538), .B(n7539), .Z(n7255) );
  AND U7534 ( .A(n213), .B(n7540), .Z(n7539) );
  AND U7535 ( .A(n7484), .B(n7465), .Z(n7529) );
  XNOR U7536 ( .A(n7541), .B(n7542), .Z(n7465) );
  AND U7537 ( .A(n206), .B(n7543), .Z(n7542) );
  XNOR U7538 ( .A(n7544), .B(n7541), .Z(n7543) );
  XNOR U7539 ( .A(n7545), .B(n7546), .Z(n206) );
  NOR U7540 ( .A(n7547), .B(n7548), .Z(n7546) );
  XNOR U7541 ( .A(n7545), .B(n7495), .Z(n7548) );
  NOR U7542 ( .A(n7491), .B(n7492), .Z(n7495) );
  NOR U7543 ( .A(n7545), .B(n7494), .Z(n7547) );
  AND U7544 ( .A(n7549), .B(n7550), .Z(n7494) );
  XOR U7545 ( .A(n7551), .B(n7552), .Z(n7545) );
  AND U7546 ( .A(n7553), .B(n7554), .Z(n7552) );
  XNOR U7547 ( .A(n7551), .B(n7549), .Z(n7554) );
  IV U7548 ( .A(n7503), .Z(n7549) );
  XOR U7549 ( .A(n7555), .B(n7556), .Z(n7503) );
  XOR U7550 ( .A(n7557), .B(n7550), .Z(n7556) );
  AND U7551 ( .A(n7515), .B(n7558), .Z(n7550) );
  AND U7552 ( .A(n7559), .B(n7560), .Z(n7557) );
  XOR U7553 ( .A(n7561), .B(n7555), .Z(n7559) );
  XNOR U7554 ( .A(n7500), .B(n7551), .Z(n7553) );
  XNOR U7555 ( .A(n7562), .B(n7563), .Z(n7500) );
  AND U7556 ( .A(n210), .B(n7507), .Z(n7563) );
  XOR U7557 ( .A(n7562), .B(n7505), .Z(n7507) );
  XOR U7558 ( .A(n7564), .B(n7565), .Z(n7551) );
  AND U7559 ( .A(n7566), .B(n7567), .Z(n7565) );
  XNOR U7560 ( .A(n7564), .B(n7515), .Z(n7567) );
  XOR U7561 ( .A(n7568), .B(n7560), .Z(n7515) );
  XNOR U7562 ( .A(n7569), .B(n7555), .Z(n7560) );
  XOR U7563 ( .A(n7570), .B(n7571), .Z(n7555) );
  AND U7564 ( .A(n7572), .B(n7573), .Z(n7571) );
  XOR U7565 ( .A(n7574), .B(n7570), .Z(n7572) );
  XNOR U7566 ( .A(n7575), .B(n7576), .Z(n7569) );
  AND U7567 ( .A(n7577), .B(n7578), .Z(n7576) );
  XOR U7568 ( .A(n7575), .B(n7579), .Z(n7577) );
  XNOR U7569 ( .A(n7561), .B(n7558), .Z(n7568) );
  AND U7570 ( .A(n7580), .B(n7581), .Z(n7558) );
  XOR U7571 ( .A(n7582), .B(n7583), .Z(n7561) );
  AND U7572 ( .A(n7584), .B(n7585), .Z(n7583) );
  XOR U7573 ( .A(n7582), .B(n7586), .Z(n7584) );
  XNOR U7574 ( .A(n7512), .B(n7564), .Z(n7566) );
  XNOR U7575 ( .A(n7587), .B(n7588), .Z(n7512) );
  AND U7576 ( .A(n210), .B(n7518), .Z(n7588) );
  XOR U7577 ( .A(n7587), .B(n7516), .Z(n7518) );
  XOR U7578 ( .A(n7589), .B(n7590), .Z(n7564) );
  AND U7579 ( .A(n7591), .B(n7592), .Z(n7590) );
  XNOR U7580 ( .A(n7589), .B(n7580), .Z(n7592) );
  IV U7581 ( .A(n7524), .Z(n7580) );
  XNOR U7582 ( .A(n7593), .B(n7573), .Z(n7524) );
  XNOR U7583 ( .A(n7594), .B(n7579), .Z(n7573) );
  XOR U7584 ( .A(n7595), .B(n7596), .Z(n7579) );
  AND U7585 ( .A(n7597), .B(n7598), .Z(n7596) );
  XOR U7586 ( .A(n7595), .B(n7599), .Z(n7597) );
  XNOR U7587 ( .A(n7578), .B(n7570), .Z(n7594) );
  XOR U7588 ( .A(n7600), .B(n7601), .Z(n7570) );
  AND U7589 ( .A(n7602), .B(n7603), .Z(n7601) );
  XNOR U7590 ( .A(n7604), .B(n7600), .Z(n7602) );
  XNOR U7591 ( .A(n7605), .B(n7575), .Z(n7578) );
  XOR U7592 ( .A(n7606), .B(n7607), .Z(n7575) );
  AND U7593 ( .A(n7608), .B(n7609), .Z(n7607) );
  XOR U7594 ( .A(n7606), .B(n7610), .Z(n7608) );
  XNOR U7595 ( .A(n7611), .B(n7612), .Z(n7605) );
  AND U7596 ( .A(n7613), .B(n7614), .Z(n7612) );
  XNOR U7597 ( .A(n7611), .B(n7615), .Z(n7613) );
  XNOR U7598 ( .A(n7574), .B(n7581), .Z(n7593) );
  AND U7599 ( .A(n7536), .B(n7616), .Z(n7581) );
  XOR U7600 ( .A(n7586), .B(n7585), .Z(n7574) );
  XNOR U7601 ( .A(n7617), .B(n7582), .Z(n7585) );
  XOR U7602 ( .A(n7618), .B(n7619), .Z(n7582) );
  AND U7603 ( .A(n7620), .B(n7621), .Z(n7619) );
  XOR U7604 ( .A(n7618), .B(n7622), .Z(n7620) );
  XNOR U7605 ( .A(n7623), .B(n7624), .Z(n7617) );
  AND U7606 ( .A(n7625), .B(n7626), .Z(n7624) );
  XOR U7607 ( .A(n7623), .B(n7627), .Z(n7625) );
  XOR U7608 ( .A(n7628), .B(n7629), .Z(n7586) );
  AND U7609 ( .A(n7630), .B(n7631), .Z(n7629) );
  XOR U7610 ( .A(n7628), .B(n7632), .Z(n7630) );
  XNOR U7611 ( .A(n7521), .B(n7589), .Z(n7591) );
  XNOR U7612 ( .A(n7633), .B(n7634), .Z(n7521) );
  AND U7613 ( .A(n210), .B(n7528), .Z(n7634) );
  XOR U7614 ( .A(n7633), .B(n7526), .Z(n7528) );
  XOR U7615 ( .A(n7635), .B(n7636), .Z(n7589) );
  AND U7616 ( .A(n7637), .B(n7638), .Z(n7636) );
  XNOR U7617 ( .A(n7635), .B(n7536), .Z(n7638) );
  XOR U7618 ( .A(n7639), .B(n7603), .Z(n7536) );
  XNOR U7619 ( .A(n7640), .B(n7610), .Z(n7603) );
  XOR U7620 ( .A(n7599), .B(n7598), .Z(n7610) );
  XNOR U7621 ( .A(n7641), .B(n7595), .Z(n7598) );
  XOR U7622 ( .A(n7642), .B(n7643), .Z(n7595) );
  AND U7623 ( .A(n7644), .B(n7645), .Z(n7643) );
  XNOR U7624 ( .A(n7646), .B(n7647), .Z(n7644) );
  IV U7625 ( .A(n7642), .Z(n7646) );
  XNOR U7626 ( .A(n7648), .B(n7649), .Z(n7641) );
  NOR U7627 ( .A(n7650), .B(n7651), .Z(n7649) );
  XNOR U7628 ( .A(n7648), .B(n7652), .Z(n7650) );
  XOR U7629 ( .A(n7653), .B(n7654), .Z(n7599) );
  NOR U7630 ( .A(n7655), .B(n7656), .Z(n7654) );
  XNOR U7631 ( .A(n7653), .B(n7657), .Z(n7655) );
  XNOR U7632 ( .A(n7609), .B(n7600), .Z(n7640) );
  XOR U7633 ( .A(n7658), .B(n7659), .Z(n7600) );
  AND U7634 ( .A(n7660), .B(n7661), .Z(n7659) );
  XOR U7635 ( .A(n7658), .B(n7662), .Z(n7660) );
  XOR U7636 ( .A(n7663), .B(n7615), .Z(n7609) );
  XOR U7637 ( .A(n7664), .B(n7665), .Z(n7615) );
  NOR U7638 ( .A(n7666), .B(n7667), .Z(n7665) );
  XOR U7639 ( .A(n7664), .B(n7668), .Z(n7666) );
  XNOR U7640 ( .A(n7614), .B(n7606), .Z(n7663) );
  XOR U7641 ( .A(n7669), .B(n7670), .Z(n7606) );
  AND U7642 ( .A(n7671), .B(n7672), .Z(n7670) );
  XOR U7643 ( .A(n7669), .B(n7673), .Z(n7671) );
  XNOR U7644 ( .A(n7674), .B(n7611), .Z(n7614) );
  XOR U7645 ( .A(n7675), .B(n7676), .Z(n7611) );
  AND U7646 ( .A(n7677), .B(n7678), .Z(n7676) );
  XNOR U7647 ( .A(n7679), .B(n7680), .Z(n7677) );
  IV U7648 ( .A(n7675), .Z(n7679) );
  XNOR U7649 ( .A(n7681), .B(n7682), .Z(n7674) );
  NOR U7650 ( .A(n7683), .B(n7684), .Z(n7682) );
  XNOR U7651 ( .A(n7681), .B(n7685), .Z(n7683) );
  XOR U7652 ( .A(n7604), .B(n7616), .Z(n7639) );
  NOR U7653 ( .A(n7544), .B(n7686), .Z(n7616) );
  XNOR U7654 ( .A(n7622), .B(n7621), .Z(n7604) );
  XNOR U7655 ( .A(n7687), .B(n7627), .Z(n7621) );
  XNOR U7656 ( .A(n7688), .B(n7689), .Z(n7627) );
  NOR U7657 ( .A(n7690), .B(n7691), .Z(n7689) );
  XOR U7658 ( .A(n7688), .B(n7692), .Z(n7690) );
  XNOR U7659 ( .A(n7626), .B(n7618), .Z(n7687) );
  XOR U7660 ( .A(n7693), .B(n7694), .Z(n7618) );
  AND U7661 ( .A(n7695), .B(n7696), .Z(n7694) );
  XOR U7662 ( .A(n7693), .B(n7697), .Z(n7695) );
  XNOR U7663 ( .A(n7698), .B(n7623), .Z(n7626) );
  XOR U7664 ( .A(n7699), .B(n7700), .Z(n7623) );
  AND U7665 ( .A(n7701), .B(n7702), .Z(n7700) );
  XNOR U7666 ( .A(n7703), .B(n7704), .Z(n7701) );
  IV U7667 ( .A(n7699), .Z(n7703) );
  XNOR U7668 ( .A(n7705), .B(n7706), .Z(n7698) );
  NOR U7669 ( .A(n7707), .B(n7708), .Z(n7706) );
  XNOR U7670 ( .A(n7705), .B(n7709), .Z(n7707) );
  XOR U7671 ( .A(n7632), .B(n7631), .Z(n7622) );
  XNOR U7672 ( .A(n7710), .B(n7628), .Z(n7631) );
  XOR U7673 ( .A(n7711), .B(n7712), .Z(n7628) );
  AND U7674 ( .A(n7713), .B(n7714), .Z(n7712) );
  XNOR U7675 ( .A(n7715), .B(n7716), .Z(n7713) );
  IV U7676 ( .A(n7711), .Z(n7715) );
  XNOR U7677 ( .A(n7717), .B(n7718), .Z(n7710) );
  NOR U7678 ( .A(n7719), .B(n7720), .Z(n7718) );
  XNOR U7679 ( .A(n7717), .B(n7721), .Z(n7719) );
  XOR U7680 ( .A(n7722), .B(n7723), .Z(n7632) );
  NOR U7681 ( .A(n7724), .B(n7725), .Z(n7723) );
  XNOR U7682 ( .A(n7722), .B(n7726), .Z(n7724) );
  XNOR U7683 ( .A(n7533), .B(n7635), .Z(n7637) );
  XNOR U7684 ( .A(n7727), .B(n7728), .Z(n7533) );
  AND U7685 ( .A(n210), .B(n7540), .Z(n7728) );
  XOR U7686 ( .A(n7727), .B(n7538), .Z(n7540) );
  AND U7687 ( .A(n7541), .B(n7544), .Z(n7635) );
  XOR U7688 ( .A(n7729), .B(n7686), .Z(n7544) );
  XNOR U7689 ( .A(p_input[416]), .B(p_input[512]), .Z(n7686) );
  XNOR U7690 ( .A(n7662), .B(n7661), .Z(n7729) );
  XNOR U7691 ( .A(n7730), .B(n7673), .Z(n7661) );
  XOR U7692 ( .A(n7647), .B(n7645), .Z(n7673) );
  XNOR U7693 ( .A(n7731), .B(n7652), .Z(n7645) );
  XOR U7694 ( .A(p_input[440]), .B(p_input[536]), .Z(n7652) );
  XOR U7695 ( .A(n7642), .B(n7651), .Z(n7731) );
  XOR U7696 ( .A(n7732), .B(n7648), .Z(n7651) );
  XOR U7697 ( .A(p_input[438]), .B(p_input[534]), .Z(n7648) );
  XOR U7698 ( .A(p_input[439]), .B(n4010), .Z(n7732) );
  XOR U7699 ( .A(p_input[434]), .B(p_input[530]), .Z(n7642) );
  XNOR U7700 ( .A(n7657), .B(n7656), .Z(n7647) );
  XOR U7701 ( .A(n7733), .B(n7653), .Z(n7656) );
  XOR U7702 ( .A(p_input[435]), .B(p_input[531]), .Z(n7653) );
  XOR U7703 ( .A(p_input[436]), .B(n4012), .Z(n7733) );
  XOR U7704 ( .A(p_input[437]), .B(p_input[533]), .Z(n7657) );
  XOR U7705 ( .A(n7672), .B(n7734), .Z(n7730) );
  IV U7706 ( .A(n7658), .Z(n7734) );
  XOR U7707 ( .A(p_input[417]), .B(p_input[513]), .Z(n7658) );
  XNOR U7708 ( .A(n7735), .B(n7680), .Z(n7672) );
  XNOR U7709 ( .A(n7668), .B(n7667), .Z(n7680) );
  XNOR U7710 ( .A(n7736), .B(n7664), .Z(n7667) );
  XNOR U7711 ( .A(p_input[442]), .B(p_input[538]), .Z(n7664) );
  XOR U7712 ( .A(p_input[443]), .B(n4016), .Z(n7736) );
  XOR U7713 ( .A(p_input[444]), .B(p_input[540]), .Z(n7668) );
  XOR U7714 ( .A(n7678), .B(n7737), .Z(n7735) );
  IV U7715 ( .A(n7669), .Z(n7737) );
  XOR U7716 ( .A(p_input[433]), .B(p_input[529]), .Z(n7669) );
  XNOR U7717 ( .A(n7738), .B(n7685), .Z(n7678) );
  XNOR U7718 ( .A(p_input[447]), .B(n4019), .Z(n7685) );
  IV U7719 ( .A(p_input[543]), .Z(n4019) );
  XOR U7720 ( .A(n7675), .B(n7684), .Z(n7738) );
  XOR U7721 ( .A(n7739), .B(n7681), .Z(n7684) );
  XOR U7722 ( .A(p_input[445]), .B(p_input[541]), .Z(n7681) );
  XOR U7723 ( .A(p_input[446]), .B(n4021), .Z(n7739) );
  XOR U7724 ( .A(p_input[441]), .B(p_input[537]), .Z(n7675) );
  XOR U7725 ( .A(n7697), .B(n7696), .Z(n7662) );
  XNOR U7726 ( .A(n7740), .B(n7704), .Z(n7696) );
  XNOR U7727 ( .A(n7692), .B(n7691), .Z(n7704) );
  XNOR U7728 ( .A(n7741), .B(n7688), .Z(n7691) );
  XNOR U7729 ( .A(p_input[427]), .B(p_input[523]), .Z(n7688) );
  XOR U7730 ( .A(p_input[428]), .B(n4024), .Z(n7741) );
  XOR U7731 ( .A(p_input[429]), .B(p_input[525]), .Z(n7692) );
  XOR U7732 ( .A(n7702), .B(n7742), .Z(n7740) );
  IV U7733 ( .A(n7693), .Z(n7742) );
  XOR U7734 ( .A(p_input[418]), .B(p_input[514]), .Z(n7693) );
  XNOR U7735 ( .A(n7743), .B(n7709), .Z(n7702) );
  XNOR U7736 ( .A(p_input[432]), .B(n4027), .Z(n7709) );
  IV U7737 ( .A(p_input[528]), .Z(n4027) );
  XOR U7738 ( .A(n7699), .B(n7708), .Z(n7743) );
  XOR U7739 ( .A(n7744), .B(n7705), .Z(n7708) );
  XOR U7740 ( .A(p_input[430]), .B(p_input[526]), .Z(n7705) );
  XOR U7741 ( .A(p_input[431]), .B(n4029), .Z(n7744) );
  XOR U7742 ( .A(p_input[426]), .B(p_input[522]), .Z(n7699) );
  XOR U7743 ( .A(n7716), .B(n7714), .Z(n7697) );
  XNOR U7744 ( .A(n7745), .B(n7721), .Z(n7714) );
  XOR U7745 ( .A(p_input[425]), .B(p_input[521]), .Z(n7721) );
  XOR U7746 ( .A(n7711), .B(n7720), .Z(n7745) );
  XOR U7747 ( .A(n7746), .B(n7717), .Z(n7720) );
  XOR U7748 ( .A(p_input[423]), .B(p_input[519]), .Z(n7717) );
  XOR U7749 ( .A(p_input[424]), .B(n4318), .Z(n7746) );
  XOR U7750 ( .A(p_input[419]), .B(p_input[515]), .Z(n7711) );
  XNOR U7751 ( .A(n7726), .B(n7725), .Z(n7716) );
  XOR U7752 ( .A(n7747), .B(n7722), .Z(n7725) );
  XOR U7753 ( .A(p_input[420]), .B(p_input[516]), .Z(n7722) );
  XOR U7754 ( .A(p_input[421]), .B(n4320), .Z(n7747) );
  XOR U7755 ( .A(p_input[422]), .B(p_input[518]), .Z(n7726) );
  XNOR U7756 ( .A(n7748), .B(n7749), .Z(n7541) );
  AND U7757 ( .A(n210), .B(n7750), .Z(n7749) );
  XNOR U7758 ( .A(n7751), .B(n7752), .Z(n210) );
  NOR U7759 ( .A(n7753), .B(n7754), .Z(n7752) );
  XOR U7760 ( .A(n7492), .B(n7751), .Z(n7754) );
  NOR U7761 ( .A(n7751), .B(n7491), .Z(n7753) );
  XOR U7762 ( .A(n7755), .B(n7756), .Z(n7751) );
  AND U7763 ( .A(n7757), .B(n7758), .Z(n7756) );
  XNOR U7764 ( .A(n7562), .B(n7755), .Z(n7758) );
  XOR U7765 ( .A(n7755), .B(n7505), .Z(n7757) );
  XOR U7766 ( .A(n7759), .B(n7760), .Z(n7755) );
  AND U7767 ( .A(n7761), .B(n7762), .Z(n7760) );
  XNOR U7768 ( .A(n7587), .B(n7759), .Z(n7762) );
  XOR U7769 ( .A(n7759), .B(n7516), .Z(n7761) );
  XOR U7770 ( .A(n7763), .B(n7764), .Z(n7759) );
  AND U7771 ( .A(n7765), .B(n7766), .Z(n7764) );
  XOR U7772 ( .A(n7763), .B(n7526), .Z(n7765) );
  XOR U7773 ( .A(n7767), .B(n7768), .Z(n7484) );
  AND U7774 ( .A(n213), .B(n7750), .Z(n7768) );
  XOR U7775 ( .A(n7769), .B(n7767), .Z(n7750) );
  XNOR U7776 ( .A(n7770), .B(n7771), .Z(n213) );
  NOR U7777 ( .A(n7772), .B(n7773), .Z(n7771) );
  XNOR U7778 ( .A(n7492), .B(n7774), .Z(n7773) );
  IV U7779 ( .A(n7770), .Z(n7774) );
  AND U7780 ( .A(n7505), .B(n7775), .Z(n7492) );
  NOR U7781 ( .A(n7770), .B(n7491), .Z(n7772) );
  AND U7782 ( .A(n7562), .B(n7776), .Z(n7491) );
  XOR U7783 ( .A(n7777), .B(n7778), .Z(n7770) );
  AND U7784 ( .A(n7779), .B(n7780), .Z(n7778) );
  XNOR U7785 ( .A(n7777), .B(n7562), .Z(n7780) );
  XNOR U7786 ( .A(n7781), .B(n7782), .Z(n7562) );
  XOR U7787 ( .A(n7783), .B(n7776), .Z(n7782) );
  AND U7788 ( .A(n7587), .B(n7784), .Z(n7776) );
  AND U7789 ( .A(n7785), .B(n7786), .Z(n7783) );
  XOR U7790 ( .A(n7787), .B(n7781), .Z(n7785) );
  XNOR U7791 ( .A(n7788), .B(n7777), .Z(n7779) );
  IV U7792 ( .A(n7505), .Z(n7788) );
  XNOR U7793 ( .A(n7789), .B(n7790), .Z(n7505) );
  XOR U7794 ( .A(n7791), .B(n7775), .Z(n7790) );
  AND U7795 ( .A(n7516), .B(n7792), .Z(n7775) );
  AND U7796 ( .A(n7793), .B(n7794), .Z(n7791) );
  XNOR U7797 ( .A(n7789), .B(n7795), .Z(n7793) );
  XOR U7798 ( .A(n7796), .B(n7797), .Z(n7777) );
  AND U7799 ( .A(n7798), .B(n7799), .Z(n7797) );
  XNOR U7800 ( .A(n7796), .B(n7587), .Z(n7799) );
  XOR U7801 ( .A(n7800), .B(n7786), .Z(n7587) );
  XNOR U7802 ( .A(n7801), .B(n7781), .Z(n7786) );
  XOR U7803 ( .A(n7802), .B(n7803), .Z(n7781) );
  AND U7804 ( .A(n7804), .B(n7805), .Z(n7803) );
  XOR U7805 ( .A(n7806), .B(n7802), .Z(n7804) );
  XNOR U7806 ( .A(n7807), .B(n7808), .Z(n7801) );
  AND U7807 ( .A(n7809), .B(n7810), .Z(n7808) );
  XOR U7808 ( .A(n7807), .B(n7811), .Z(n7809) );
  XNOR U7809 ( .A(n7787), .B(n7784), .Z(n7800) );
  AND U7810 ( .A(n7633), .B(n7812), .Z(n7784) );
  XOR U7811 ( .A(n7813), .B(n7814), .Z(n7787) );
  AND U7812 ( .A(n7815), .B(n7816), .Z(n7814) );
  XOR U7813 ( .A(n7813), .B(n7817), .Z(n7815) );
  XOR U7814 ( .A(n7516), .B(n7796), .Z(n7798) );
  XNOR U7815 ( .A(n7818), .B(n7795), .Z(n7516) );
  XNOR U7816 ( .A(n7819), .B(n7820), .Z(n7795) );
  AND U7817 ( .A(n7821), .B(n7822), .Z(n7820) );
  XOR U7818 ( .A(n7819), .B(n7823), .Z(n7821) );
  XNOR U7819 ( .A(n7794), .B(n7792), .Z(n7818) );
  AND U7820 ( .A(n7526), .B(n7824), .Z(n7792) );
  XNOR U7821 ( .A(n7825), .B(n7789), .Z(n7794) );
  XOR U7822 ( .A(n7826), .B(n7827), .Z(n7789) );
  AND U7823 ( .A(n7828), .B(n7829), .Z(n7827) );
  XOR U7824 ( .A(n7826), .B(n7830), .Z(n7828) );
  XNOR U7825 ( .A(n7831), .B(n7832), .Z(n7825) );
  AND U7826 ( .A(n7833), .B(n7834), .Z(n7832) );
  XNOR U7827 ( .A(n7831), .B(n7835), .Z(n7833) );
  XOR U7828 ( .A(n7763), .B(n7836), .Z(n7796) );
  AND U7829 ( .A(n7837), .B(n7766), .Z(n7836) );
  XNOR U7830 ( .A(n7633), .B(n7763), .Z(n7766) );
  XOR U7831 ( .A(n7838), .B(n7805), .Z(n7633) );
  XNOR U7832 ( .A(n7839), .B(n7811), .Z(n7805) );
  XOR U7833 ( .A(n7840), .B(n7841), .Z(n7811) );
  AND U7834 ( .A(n7842), .B(n7843), .Z(n7841) );
  XOR U7835 ( .A(n7840), .B(n7844), .Z(n7842) );
  XNOR U7836 ( .A(n7810), .B(n7802), .Z(n7839) );
  XOR U7837 ( .A(n7845), .B(n7846), .Z(n7802) );
  AND U7838 ( .A(n7847), .B(n7848), .Z(n7846) );
  XNOR U7839 ( .A(n7849), .B(n7845), .Z(n7847) );
  XNOR U7840 ( .A(n7850), .B(n7807), .Z(n7810) );
  XOR U7841 ( .A(n7851), .B(n7852), .Z(n7807) );
  AND U7842 ( .A(n7853), .B(n7854), .Z(n7852) );
  XOR U7843 ( .A(n7851), .B(n7855), .Z(n7853) );
  XNOR U7844 ( .A(n7856), .B(n7857), .Z(n7850) );
  AND U7845 ( .A(n7858), .B(n7859), .Z(n7857) );
  XNOR U7846 ( .A(n7856), .B(n7860), .Z(n7858) );
  XNOR U7847 ( .A(n7806), .B(n7812), .Z(n7838) );
  AND U7848 ( .A(n7727), .B(n7861), .Z(n7812) );
  XOR U7849 ( .A(n7817), .B(n7816), .Z(n7806) );
  XNOR U7850 ( .A(n7862), .B(n7813), .Z(n7816) );
  XOR U7851 ( .A(n7863), .B(n7864), .Z(n7813) );
  AND U7852 ( .A(n7865), .B(n7866), .Z(n7864) );
  XOR U7853 ( .A(n7863), .B(n7867), .Z(n7865) );
  XNOR U7854 ( .A(n7868), .B(n7869), .Z(n7862) );
  AND U7855 ( .A(n7870), .B(n7871), .Z(n7869) );
  XOR U7856 ( .A(n7868), .B(n7872), .Z(n7870) );
  XOR U7857 ( .A(n7873), .B(n7874), .Z(n7817) );
  AND U7858 ( .A(n7875), .B(n7876), .Z(n7874) );
  XOR U7859 ( .A(n7873), .B(n7877), .Z(n7875) );
  XNOR U7860 ( .A(n7878), .B(n7763), .Z(n7837) );
  IV U7861 ( .A(n7526), .Z(n7878) );
  XOR U7862 ( .A(n7879), .B(n7830), .Z(n7526) );
  XOR U7863 ( .A(n7823), .B(n7822), .Z(n7830) );
  XNOR U7864 ( .A(n7880), .B(n7819), .Z(n7822) );
  XOR U7865 ( .A(n7881), .B(n7882), .Z(n7819) );
  AND U7866 ( .A(n7883), .B(n7884), .Z(n7882) );
  XOR U7867 ( .A(n7881), .B(n7885), .Z(n7883) );
  XNOR U7868 ( .A(n7886), .B(n7887), .Z(n7880) );
  AND U7869 ( .A(n7888), .B(n7889), .Z(n7887) );
  XOR U7870 ( .A(n7886), .B(n7890), .Z(n7888) );
  XOR U7871 ( .A(n7891), .B(n7892), .Z(n7823) );
  AND U7872 ( .A(n7893), .B(n7894), .Z(n7892) );
  XOR U7873 ( .A(n7891), .B(n7895), .Z(n7893) );
  XNOR U7874 ( .A(n7829), .B(n7824), .Z(n7879) );
  AND U7875 ( .A(n7538), .B(n7896), .Z(n7824) );
  XOR U7876 ( .A(n7897), .B(n7835), .Z(n7829) );
  XNOR U7877 ( .A(n7898), .B(n7899), .Z(n7835) );
  AND U7878 ( .A(n7900), .B(n7901), .Z(n7899) );
  XOR U7879 ( .A(n7898), .B(n7902), .Z(n7900) );
  XNOR U7880 ( .A(n7834), .B(n7826), .Z(n7897) );
  XOR U7881 ( .A(n7903), .B(n7904), .Z(n7826) );
  AND U7882 ( .A(n7905), .B(n7906), .Z(n7904) );
  XOR U7883 ( .A(n7903), .B(n7907), .Z(n7905) );
  XNOR U7884 ( .A(n7908), .B(n7831), .Z(n7834) );
  XOR U7885 ( .A(n7909), .B(n7910), .Z(n7831) );
  AND U7886 ( .A(n7911), .B(n7912), .Z(n7910) );
  XOR U7887 ( .A(n7909), .B(n7913), .Z(n7911) );
  XNOR U7888 ( .A(n7914), .B(n7915), .Z(n7908) );
  AND U7889 ( .A(n7916), .B(n7917), .Z(n7915) );
  XNOR U7890 ( .A(n7914), .B(n7918), .Z(n7916) );
  XOR U7891 ( .A(n7919), .B(n7920), .Z(n7763) );
  AND U7892 ( .A(n7921), .B(n7922), .Z(n7920) );
  XNOR U7893 ( .A(n7919), .B(n7727), .Z(n7922) );
  XOR U7894 ( .A(n7923), .B(n7848), .Z(n7727) );
  XNOR U7895 ( .A(n7924), .B(n7855), .Z(n7848) );
  XOR U7896 ( .A(n7844), .B(n7843), .Z(n7855) );
  XNOR U7897 ( .A(n7925), .B(n7840), .Z(n7843) );
  XOR U7898 ( .A(n7926), .B(n7927), .Z(n7840) );
  AND U7899 ( .A(n7928), .B(n7929), .Z(n7927) );
  XOR U7900 ( .A(n7926), .B(n7930), .Z(n7928) );
  XNOR U7901 ( .A(n7931), .B(n7932), .Z(n7925) );
  NOR U7902 ( .A(n7933), .B(n7934), .Z(n7932) );
  XNOR U7903 ( .A(n7931), .B(n7935), .Z(n7933) );
  XOR U7904 ( .A(n7936), .B(n7937), .Z(n7844) );
  NOR U7905 ( .A(n7938), .B(n7939), .Z(n7937) );
  XNOR U7906 ( .A(n7936), .B(n7940), .Z(n7938) );
  XNOR U7907 ( .A(n7854), .B(n7845), .Z(n7924) );
  XOR U7908 ( .A(n7941), .B(n7942), .Z(n7845) );
  NOR U7909 ( .A(n7943), .B(n7944), .Z(n7942) );
  XNOR U7910 ( .A(n7941), .B(n7945), .Z(n7943) );
  XOR U7911 ( .A(n7946), .B(n7860), .Z(n7854) );
  XNOR U7912 ( .A(n7947), .B(n7948), .Z(n7860) );
  NOR U7913 ( .A(n7949), .B(n7950), .Z(n7948) );
  XNOR U7914 ( .A(n7947), .B(n7951), .Z(n7949) );
  XNOR U7915 ( .A(n7859), .B(n7851), .Z(n7946) );
  XOR U7916 ( .A(n7952), .B(n7953), .Z(n7851) );
  AND U7917 ( .A(n7954), .B(n7955), .Z(n7953) );
  XOR U7918 ( .A(n7952), .B(n7956), .Z(n7954) );
  XNOR U7919 ( .A(n7957), .B(n7856), .Z(n7859) );
  XOR U7920 ( .A(n7958), .B(n7959), .Z(n7856) );
  AND U7921 ( .A(n7960), .B(n7961), .Z(n7959) );
  XOR U7922 ( .A(n7958), .B(n7962), .Z(n7960) );
  XNOR U7923 ( .A(n7963), .B(n7964), .Z(n7957) );
  NOR U7924 ( .A(n7965), .B(n7966), .Z(n7964) );
  XOR U7925 ( .A(n7963), .B(n7967), .Z(n7965) );
  XOR U7926 ( .A(n7849), .B(n7861), .Z(n7923) );
  AND U7927 ( .A(n7769), .B(n7968), .Z(n7861) );
  IV U7928 ( .A(n7748), .Z(n7769) );
  XNOR U7929 ( .A(n7867), .B(n7866), .Z(n7849) );
  XNOR U7930 ( .A(n7969), .B(n7872), .Z(n7866) );
  XOR U7931 ( .A(n7970), .B(n7971), .Z(n7872) );
  NOR U7932 ( .A(n7972), .B(n7973), .Z(n7971) );
  XNOR U7933 ( .A(n7970), .B(n7974), .Z(n7972) );
  XNOR U7934 ( .A(n7871), .B(n7863), .Z(n7969) );
  XOR U7935 ( .A(n7975), .B(n7976), .Z(n7863) );
  AND U7936 ( .A(n7977), .B(n7978), .Z(n7976) );
  XNOR U7937 ( .A(n7975), .B(n7979), .Z(n7977) );
  XNOR U7938 ( .A(n7980), .B(n7868), .Z(n7871) );
  XOR U7939 ( .A(n7981), .B(n7982), .Z(n7868) );
  AND U7940 ( .A(n7983), .B(n7984), .Z(n7982) );
  XOR U7941 ( .A(n7981), .B(n7985), .Z(n7983) );
  XNOR U7942 ( .A(n7986), .B(n7987), .Z(n7980) );
  NOR U7943 ( .A(n7988), .B(n7989), .Z(n7987) );
  XOR U7944 ( .A(n7986), .B(n7990), .Z(n7988) );
  XOR U7945 ( .A(n7877), .B(n7876), .Z(n7867) );
  XNOR U7946 ( .A(n7991), .B(n7873), .Z(n7876) );
  XOR U7947 ( .A(n7992), .B(n7993), .Z(n7873) );
  AND U7948 ( .A(n7994), .B(n7995), .Z(n7993) );
  XOR U7949 ( .A(n7992), .B(n7996), .Z(n7994) );
  XNOR U7950 ( .A(n7997), .B(n7998), .Z(n7991) );
  NOR U7951 ( .A(n7999), .B(n8000), .Z(n7998) );
  XNOR U7952 ( .A(n7997), .B(n8001), .Z(n7999) );
  XOR U7953 ( .A(n8002), .B(n8003), .Z(n7877) );
  NOR U7954 ( .A(n8004), .B(n8005), .Z(n8003) );
  XNOR U7955 ( .A(n8002), .B(n8006), .Z(n8004) );
  XNOR U7956 ( .A(n8007), .B(n7919), .Z(n7921) );
  IV U7957 ( .A(n7538), .Z(n8007) );
  XOR U7958 ( .A(n8008), .B(n7907), .Z(n7538) );
  XOR U7959 ( .A(n7885), .B(n7884), .Z(n7907) );
  XNOR U7960 ( .A(n8009), .B(n7890), .Z(n7884) );
  XOR U7961 ( .A(n8010), .B(n8011), .Z(n7890) );
  NOR U7962 ( .A(n8012), .B(n8013), .Z(n8011) );
  XNOR U7963 ( .A(n8010), .B(n8014), .Z(n8012) );
  XNOR U7964 ( .A(n7889), .B(n7881), .Z(n8009) );
  XOR U7965 ( .A(n8015), .B(n8016), .Z(n7881) );
  AND U7966 ( .A(n8017), .B(n8018), .Z(n8016) );
  XNOR U7967 ( .A(n8015), .B(n8019), .Z(n8017) );
  XNOR U7968 ( .A(n8020), .B(n7886), .Z(n7889) );
  XOR U7969 ( .A(n8021), .B(n8022), .Z(n7886) );
  AND U7970 ( .A(n8023), .B(n8024), .Z(n8022) );
  XOR U7971 ( .A(n8021), .B(n8025), .Z(n8023) );
  XNOR U7972 ( .A(n8026), .B(n8027), .Z(n8020) );
  NOR U7973 ( .A(n8028), .B(n8029), .Z(n8027) );
  XOR U7974 ( .A(n8026), .B(n8030), .Z(n8028) );
  XOR U7975 ( .A(n7895), .B(n7894), .Z(n7885) );
  XNOR U7976 ( .A(n8031), .B(n7891), .Z(n7894) );
  XOR U7977 ( .A(n8032), .B(n8033), .Z(n7891) );
  AND U7978 ( .A(n8034), .B(n8035), .Z(n8033) );
  XOR U7979 ( .A(n8032), .B(n8036), .Z(n8034) );
  XNOR U7980 ( .A(n8037), .B(n8038), .Z(n8031) );
  NOR U7981 ( .A(n8039), .B(n8040), .Z(n8038) );
  XNOR U7982 ( .A(n8037), .B(n8041), .Z(n8039) );
  XOR U7983 ( .A(n8042), .B(n8043), .Z(n7895) );
  NOR U7984 ( .A(n8044), .B(n8045), .Z(n8043) );
  XNOR U7985 ( .A(n8042), .B(n8046), .Z(n8044) );
  XNOR U7986 ( .A(n7906), .B(n7896), .Z(n8008) );
  AND U7987 ( .A(n7767), .B(n8047), .Z(n7896) );
  XNOR U7988 ( .A(n8048), .B(n7913), .Z(n7906) );
  XOR U7989 ( .A(n7902), .B(n7901), .Z(n7913) );
  XNOR U7990 ( .A(n8049), .B(n7898), .Z(n7901) );
  XOR U7991 ( .A(n8050), .B(n8051), .Z(n7898) );
  AND U7992 ( .A(n8052), .B(n8053), .Z(n8051) );
  XOR U7993 ( .A(n8050), .B(n8054), .Z(n8052) );
  XNOR U7994 ( .A(n8055), .B(n8056), .Z(n8049) );
  NOR U7995 ( .A(n8057), .B(n8058), .Z(n8056) );
  XNOR U7996 ( .A(n8055), .B(n8059), .Z(n8057) );
  XOR U7997 ( .A(n8060), .B(n8061), .Z(n7902) );
  NOR U7998 ( .A(n8062), .B(n8063), .Z(n8061) );
  XNOR U7999 ( .A(n8060), .B(n8064), .Z(n8062) );
  XNOR U8000 ( .A(n7912), .B(n7903), .Z(n8048) );
  XOR U8001 ( .A(n8065), .B(n8066), .Z(n7903) );
  NOR U8002 ( .A(n8067), .B(n8068), .Z(n8066) );
  XNOR U8003 ( .A(n8065), .B(n8069), .Z(n8067) );
  XOR U8004 ( .A(n8070), .B(n7918), .Z(n7912) );
  XNOR U8005 ( .A(n8071), .B(n8072), .Z(n7918) );
  NOR U8006 ( .A(n8073), .B(n8074), .Z(n8072) );
  XNOR U8007 ( .A(n8071), .B(n8075), .Z(n8073) );
  XNOR U8008 ( .A(n7917), .B(n7909), .Z(n8070) );
  XOR U8009 ( .A(n8076), .B(n8077), .Z(n7909) );
  AND U8010 ( .A(n8078), .B(n8079), .Z(n8077) );
  XOR U8011 ( .A(n8076), .B(n8080), .Z(n8078) );
  XNOR U8012 ( .A(n8081), .B(n7914), .Z(n7917) );
  XOR U8013 ( .A(n8082), .B(n8083), .Z(n7914) );
  AND U8014 ( .A(n8084), .B(n8085), .Z(n8083) );
  XOR U8015 ( .A(n8082), .B(n8086), .Z(n8084) );
  XNOR U8016 ( .A(n8087), .B(n8088), .Z(n8081) );
  NOR U8017 ( .A(n8089), .B(n8090), .Z(n8088) );
  XOR U8018 ( .A(n8087), .B(n8091), .Z(n8089) );
  AND U8019 ( .A(n7767), .B(n7748), .Z(n7919) );
  XNOR U8020 ( .A(n8092), .B(n7968), .Z(n7748) );
  XOR U8021 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(
        p_input[512]), .Z(n7968) );
  XOR U8022 ( .A(n7945), .B(n7944), .Z(n8092) );
  XOR U8023 ( .A(n8093), .B(n7956), .Z(n7944) );
  XOR U8024 ( .A(n7930), .B(n7929), .Z(n7956) );
  XNOR U8025 ( .A(n8094), .B(n7935), .Z(n7929) );
  XNOR U8026 ( .A(n1931), .B(p_input[536]), .Z(n7935) );
  IV U8027 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .Z(n1931) );
  XOR U8028 ( .A(n7926), .B(n7934), .Z(n8094) );
  XOR U8029 ( .A(n8095), .B(n7931), .Z(n7934) );
  XNOR U8030 ( .A(n2158), .B(p_input[534]), .Z(n7931) );
  IV U8031 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .Z(n2158) );
  XOR U8032 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .B(n4010), 
        .Z(n8095) );
  XNOR U8033 ( .A(n2724), .B(p_input[530]), .Z(n7926) );
  IV U8034 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .Z(n2724) );
  XNOR U8035 ( .A(n7940), .B(n7939), .Z(n7930) );
  XOR U8036 ( .A(n8096), .B(n7936), .Z(n7939) );
  XNOR U8037 ( .A(n2611), .B(p_input[531]), .Z(n7936) );
  IV U8038 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .Z(n2611) );
  XOR U8039 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .B(n4012), 
        .Z(n8096) );
  XNOR U8040 ( .A(n2271), .B(p_input[533]), .Z(n7940) );
  IV U8041 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .Z(n2271) );
  XNOR U8042 ( .A(n7955), .B(n7941), .Z(n8093) );
  XNOR U8043 ( .A(n2498), .B(p_input[513]), .Z(n7941) );
  IV U8044 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n2498) );
  XNOR U8045 ( .A(n8097), .B(n7962), .Z(n7955) );
  XNOR U8046 ( .A(n7951), .B(n7950), .Z(n7962) );
  XOR U8047 ( .A(n8098), .B(n7947), .Z(n7950) );
  XNOR U8048 ( .A(n1705), .B(p_input[538]), .Z(n7947) );
  IV U8049 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .Z(n1705) );
  XOR U8050 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .B(n4016), 
        .Z(n8098) );
  XNOR U8051 ( .A(n1478), .B(p_input[540]), .Z(n7951) );
  IV U8052 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .Z(n1478) );
  XNOR U8053 ( .A(n7961), .B(n7952), .Z(n8097) );
  XNOR U8054 ( .A(n2837), .B(p_input[529]), .Z(n7952) );
  IV U8055 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .Z(n2837) );
  XOR U8056 ( .A(n8099), .B(n7967), .Z(n7961) );
  XNOR U8057 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .B(
        p_input[543]), .Z(n7967) );
  XOR U8058 ( .A(n7958), .B(n7966), .Z(n8099) );
  XOR U8059 ( .A(n8100), .B(n7963), .Z(n7966) );
  XNOR U8060 ( .A(n1365), .B(p_input[541]), .Z(n7963) );
  IV U8061 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .Z(n1365) );
  XOR U8062 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .B(n4021), 
        .Z(n8100) );
  XNOR U8063 ( .A(n1818), .B(p_input[537]), .Z(n7958) );
  IV U8064 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .Z(n1818) );
  XNOR U8065 ( .A(n7979), .B(n7978), .Z(n7945) );
  XNOR U8066 ( .A(n8101), .B(n7985), .Z(n7978) );
  XNOR U8067 ( .A(n7974), .B(n7973), .Z(n7985) );
  XOR U8068 ( .A(n8102), .B(n7970), .Z(n7973) );
  XNOR U8069 ( .A(n3518), .B(p_input[523]), .Z(n7970) );
  IV U8070 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n3518) );
  XOR U8071 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(n4024), 
        .Z(n8102) );
  XNOR U8072 ( .A(n3291), .B(p_input[525]), .Z(n7974) );
  IV U8073 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n3291) );
  XNOR U8074 ( .A(n7984), .B(n7975), .Z(n8101) );
  XNOR U8075 ( .A(n1252), .B(p_input[514]), .Z(n7975) );
  IV U8076 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n1252) );
  XOR U8077 ( .A(n8103), .B(n7990), .Z(n7984) );
  XNOR U8078 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .B(
        p_input[528]), .Z(n7990) );
  XOR U8079 ( .A(n7981), .B(n7989), .Z(n8103) );
  XOR U8080 ( .A(n8104), .B(n7986), .Z(n7989) );
  XNOR U8081 ( .A(n3178), .B(p_input[526]), .Z(n7986) );
  IV U8082 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n3178) );
  XOR U8083 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(n4029), 
        .Z(n8104) );
  XNOR U8084 ( .A(n3631), .B(p_input[522]), .Z(n7981) );
  IV U8085 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n3631) );
  XNOR U8086 ( .A(n7996), .B(n7995), .Z(n7979) );
  XNOR U8087 ( .A(n8105), .B(n8001), .Z(n7995) );
  XNOR U8088 ( .A(n208), .B(p_input[521]), .Z(n8001) );
  IV U8089 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .Z(n208) );
  XOR U8090 ( .A(n7992), .B(n8000), .Z(n8105) );
  XOR U8091 ( .A(n8106), .B(n7997), .Z(n8000) );
  XNOR U8092 ( .A(n442), .B(p_input[519]), .Z(n7997) );
  IV U8093 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .Z(n442) );
  XOR U8094 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(n4318), 
        .Z(n8106) );
  XNOR U8095 ( .A(n902), .B(p_input[515]), .Z(n7992) );
  IV U8096 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .Z(n902) );
  XNOR U8097 ( .A(n8006), .B(n8005), .Z(n7996) );
  XOR U8098 ( .A(n8107), .B(n8002), .Z(n8005) );
  XNOR U8099 ( .A(n787), .B(p_input[516]), .Z(n8002) );
  IV U8100 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .Z(n787) );
  XOR U8101 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(n4320), 
        .Z(n8107) );
  XNOR U8102 ( .A(n557), .B(p_input[518]), .Z(n8006) );
  IV U8103 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .Z(n557) );
  XOR U8104 ( .A(n8108), .B(n8069), .Z(n7767) );
  XNOR U8105 ( .A(n8019), .B(n8018), .Z(n8069) );
  XNOR U8106 ( .A(n8109), .B(n8025), .Z(n8018) );
  XNOR U8107 ( .A(n8014), .B(n8013), .Z(n8025) );
  XOR U8108 ( .A(n8110), .B(n8010), .Z(n8013) );
  XNOR U8109 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n4599), .Z(n8010) );
  IV U8110 ( .A(p_input[523]), .Z(n4599) );
  XOR U8111 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n4024), .Z(n8110) );
  IV U8112 ( .A(p_input[524]), .Z(n4024) );
  XOR U8113 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[525]), .Z(n8014)
         );
  XNOR U8114 ( .A(n8024), .B(n8015), .Z(n8109) );
  XNOR U8115 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n4600), .Z(n8015) );
  IV U8116 ( .A(p_input[514]), .Z(n4600) );
  XOR U8117 ( .A(n8111), .B(n8030), .Z(n8024) );
  XNOR U8118 ( .A(\knn_comb_/min_val_out[0][16] ), .B(p_input[528]), .Z(n8030)
         );
  XOR U8119 ( .A(n8021), .B(n8029), .Z(n8111) );
  XOR U8120 ( .A(n8112), .B(n8026), .Z(n8029) );
  XOR U8121 ( .A(\knn_comb_/min_val_out[0][14] ), .B(p_input[526]), .Z(n8026)
         );
  XOR U8122 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n4029), .Z(n8112) );
  IV U8123 ( .A(p_input[527]), .Z(n4029) );
  XNOR U8124 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n4603), .Z(n8021) );
  IV U8125 ( .A(p_input[522]), .Z(n4603) );
  XNOR U8126 ( .A(n8036), .B(n8035), .Z(n8019) );
  XNOR U8127 ( .A(n8113), .B(n8041), .Z(n8035) );
  XNOR U8128 ( .A(n214), .B(p_input[521]), .Z(n8041) );
  IV U8129 ( .A(\knn_comb_/min_val_out[0][9] ), .Z(n214) );
  XOR U8130 ( .A(n8032), .B(n8040), .Z(n8113) );
  XOR U8131 ( .A(n8114), .B(n8037), .Z(n8040) );
  XNOR U8132 ( .A(n446), .B(p_input[519]), .Z(n8037) );
  IV U8133 ( .A(\knn_comb_/min_val_out[0][7] ), .Z(n446) );
  XOR U8134 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n4318), .Z(n8114) );
  IV U8135 ( .A(p_input[520]), .Z(n4318) );
  XNOR U8136 ( .A(n906), .B(p_input[515]), .Z(n8032) );
  IV U8137 ( .A(\knn_comb_/min_val_out[0][3] ), .Z(n906) );
  XNOR U8138 ( .A(n8046), .B(n8045), .Z(n8036) );
  XOR U8139 ( .A(n8115), .B(n8042), .Z(n8045) );
  XNOR U8140 ( .A(n791), .B(p_input[516]), .Z(n8042) );
  IV U8141 ( .A(\knn_comb_/min_val_out[0][4] ), .Z(n791) );
  XOR U8142 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n4320), .Z(n8115) );
  IV U8143 ( .A(p_input[517]), .Z(n4320) );
  XNOR U8144 ( .A(n561), .B(p_input[518]), .Z(n8046) );
  IV U8145 ( .A(\knn_comb_/min_val_out[0][6] ), .Z(n561) );
  XOR U8146 ( .A(n8068), .B(n8047), .Z(n8108) );
  XOR U8147 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[512]), .Z(n8047)
         );
  XOR U8148 ( .A(n8116), .B(n8080), .Z(n8068) );
  XOR U8149 ( .A(n8054), .B(n8053), .Z(n8080) );
  XNOR U8150 ( .A(n8117), .B(n8059), .Z(n8053) );
  XOR U8151 ( .A(\knn_comb_/min_val_out[0][24] ), .B(p_input[536]), .Z(n8059)
         );
  XOR U8152 ( .A(n8050), .B(n8058), .Z(n8117) );
  XOR U8153 ( .A(n8118), .B(n8055), .Z(n8058) );
  XOR U8154 ( .A(\knn_comb_/min_val_out[0][22] ), .B(p_input[534]), .Z(n8055)
         );
  XOR U8155 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n4010), .Z(n8118) );
  IV U8156 ( .A(p_input[535]), .Z(n4010) );
  XNOR U8157 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n4589), .Z(n8050) );
  IV U8158 ( .A(p_input[530]), .Z(n4589) );
  XNOR U8159 ( .A(n8064), .B(n8063), .Z(n8054) );
  XOR U8160 ( .A(n8119), .B(n8060), .Z(n8063) );
  XOR U8161 ( .A(\knn_comb_/min_val_out[0][19] ), .B(p_input[531]), .Z(n8060)
         );
  XOR U8162 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n4012), .Z(n8119) );
  IV U8163 ( .A(p_input[532]), .Z(n4012) );
  XOR U8164 ( .A(\knn_comb_/min_val_out[0][21] ), .B(p_input[533]), .Z(n8064)
         );
  XNOR U8165 ( .A(n8079), .B(n8065), .Z(n8116) );
  XNOR U8166 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n4591), .Z(n8065) );
  IV U8167 ( .A(p_input[513]), .Z(n4591) );
  XNOR U8168 ( .A(n8120), .B(n8086), .Z(n8079) );
  XNOR U8169 ( .A(n8075), .B(n8074), .Z(n8086) );
  XOR U8170 ( .A(n8121), .B(n8071), .Z(n8074) );
  XNOR U8171 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n4306), .Z(n8071) );
  IV U8172 ( .A(p_input[538]), .Z(n4306) );
  XOR U8173 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n4016), .Z(n8121) );
  IV U8174 ( .A(p_input[539]), .Z(n4016) );
  XOR U8175 ( .A(\knn_comb_/min_val_out[0][28] ), .B(p_input[540]), .Z(n8075)
         );
  XNOR U8176 ( .A(n8085), .B(n8076), .Z(n8120) );
  XNOR U8177 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n4594), .Z(n8076) );
  IV U8178 ( .A(p_input[529]), .Z(n4594) );
  XOR U8179 ( .A(n8122), .B(n8091), .Z(n8085) );
  XNOR U8180 ( .A(\knn_comb_/min_val_out[0][31] ), .B(p_input[543]), .Z(n8091)
         );
  XOR U8181 ( .A(n8082), .B(n8090), .Z(n8122) );
  XOR U8182 ( .A(n8123), .B(n8087), .Z(n8090) );
  XOR U8183 ( .A(\knn_comb_/min_val_out[0][29] ), .B(p_input[541]), .Z(n8087)
         );
  XOR U8184 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n4021), .Z(n8123) );
  IV U8185 ( .A(p_input[542]), .Z(n4021) );
  XNOR U8186 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n4310), .Z(n8082) );
  IV U8187 ( .A(p_input[537]), .Z(n4310) );
endmodule

