
module auction_BMR_N3_W16 ( p_input, o );
  input [127:0] p_input;
  output [18:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789;

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(o[2]), .B(n3), .Z(n1) );
  XOR U3 ( .A(n2), .B(n4), .Z(n3) );
  XOR U4 ( .A(n5), .B(n6), .Z(o[8]) );
  AND U5 ( .A(o[2]), .B(n7), .Z(n5) );
  XOR U6 ( .A(n8), .B(n9), .Z(n7) );
  XOR U7 ( .A(n10), .B(n11), .Z(o[7]) );
  AND U8 ( .A(o[2]), .B(n12), .Z(n10) );
  XOR U9 ( .A(n13), .B(n14), .Z(n12) );
  XOR U10 ( .A(n15), .B(n16), .Z(o[6]) );
  AND U11 ( .A(o[2]), .B(n17), .Z(n15) );
  XOR U12 ( .A(n18), .B(n19), .Z(n17) );
  XOR U13 ( .A(n20), .B(n21), .Z(o[5]) );
  AND U14 ( .A(o[2]), .B(n22), .Z(n20) );
  XOR U15 ( .A(n23), .B(n24), .Z(n22) );
  XOR U16 ( .A(n25), .B(n26), .Z(o[4]) );
  AND U17 ( .A(o[2]), .B(n27), .Z(n25) );
  XOR U18 ( .A(n28), .B(n29), .Z(n27) );
  XNOR U19 ( .A(n30), .B(n31), .Z(o[3]) );
  AND U20 ( .A(o[2]), .B(n32), .Z(n30) );
  XNOR U21 ( .A(n33), .B(n31), .Z(n32) );
  AND U22 ( .A(n34), .B(n35), .Z(o[18]) );
  XOR U23 ( .A(n36), .B(n37), .Z(o[17]) );
  AND U24 ( .A(o[2]), .B(n38), .Z(n36) );
  XOR U25 ( .A(n39), .B(n40), .Z(n38) );
  XOR U26 ( .A(n41), .B(n42), .Z(o[16]) );
  AND U27 ( .A(o[2]), .B(n43), .Z(n41) );
  XOR U28 ( .A(n44), .B(n45), .Z(n43) );
  XOR U29 ( .A(n46), .B(n47), .Z(o[15]) );
  AND U30 ( .A(o[2]), .B(n48), .Z(n46) );
  XOR U31 ( .A(n49), .B(n50), .Z(n48) );
  XOR U32 ( .A(n51), .B(n52), .Z(o[14]) );
  AND U33 ( .A(o[2]), .B(n53), .Z(n51) );
  XOR U34 ( .A(n54), .B(n55), .Z(n53) );
  XOR U35 ( .A(n56), .B(n57), .Z(o[13]) );
  AND U36 ( .A(o[2]), .B(n58), .Z(n56) );
  XOR U37 ( .A(n59), .B(n60), .Z(n58) );
  XOR U38 ( .A(n61), .B(n62), .Z(o[12]) );
  AND U39 ( .A(o[2]), .B(n63), .Z(n61) );
  XOR U40 ( .A(n64), .B(n65), .Z(n63) );
  XOR U41 ( .A(n66), .B(n67), .Z(o[11]) );
  AND U42 ( .A(o[2]), .B(n68), .Z(n66) );
  XOR U43 ( .A(n69), .B(n70), .Z(n68) );
  XOR U44 ( .A(n71), .B(n72), .Z(o[10]) );
  AND U45 ( .A(o[2]), .B(n73), .Z(n71) );
  XOR U46 ( .A(n74), .B(n75), .Z(n73) );
  XOR U47 ( .A(n76), .B(n77), .Z(o[0]) );
  AND U48 ( .A(o[1]), .B(n78), .Z(n77) );
  XNOR U49 ( .A(n76), .B(n79), .Z(n78) );
  XNOR U50 ( .A(n80), .B(n81), .Z(n79) );
  AND U51 ( .A(o[2]), .B(n82), .Z(n80) );
  XOR U52 ( .A(n81), .B(n83), .Z(n82) );
  XOR U53 ( .A(n84), .B(n85), .Z(o[1]) );
  AND U54 ( .A(o[2]), .B(n86), .Z(n85) );
  XOR U55 ( .A(n84), .B(n87), .Z(n86) );
  XOR U56 ( .A(n88), .B(n89), .Z(n76) );
  AND U57 ( .A(o[2]), .B(n90), .Z(n89) );
  XOR U58 ( .A(n88), .B(n91), .Z(n90) );
  XOR U59 ( .A(n92), .B(n93), .Z(o[2]) );
  AND U60 ( .A(n94), .B(n95), .Z(n93) );
  XNOR U61 ( .A(n35), .B(n92), .Z(n95) );
  AND U62 ( .A(n96), .B(n97), .Z(n35) );
  XOR U63 ( .A(n92), .B(n34), .Z(n94) );
  AND U64 ( .A(n98), .B(n99), .Z(n34) );
  XOR U65 ( .A(n100), .B(n101), .Z(n92) );
  AND U66 ( .A(n102), .B(n103), .Z(n101) );
  XOR U67 ( .A(n100), .B(n39), .Z(n103) );
  XOR U68 ( .A(n104), .B(n105), .Z(n39) );
  AND U69 ( .A(n87), .B(n106), .Z(n105) );
  XOR U70 ( .A(n107), .B(n104), .Z(n106) );
  XNOR U71 ( .A(n40), .B(n100), .Z(n102) );
  IV U72 ( .A(n37), .Z(n40) );
  XNOR U73 ( .A(n108), .B(n109), .Z(n37) );
  AND U74 ( .A(n84), .B(n110), .Z(n109) );
  XOR U75 ( .A(n111), .B(n108), .Z(n110) );
  XOR U76 ( .A(n112), .B(n113), .Z(n100) );
  AND U77 ( .A(n114), .B(n115), .Z(n113) );
  XOR U78 ( .A(n112), .B(n44), .Z(n115) );
  XOR U79 ( .A(n116), .B(n117), .Z(n44) );
  AND U80 ( .A(n87), .B(n118), .Z(n117) );
  XOR U81 ( .A(n119), .B(n116), .Z(n118) );
  XNOR U82 ( .A(n45), .B(n112), .Z(n114) );
  IV U83 ( .A(n42), .Z(n45) );
  XNOR U84 ( .A(n120), .B(n121), .Z(n42) );
  AND U85 ( .A(n84), .B(n122), .Z(n121) );
  XOR U86 ( .A(n123), .B(n120), .Z(n122) );
  XOR U87 ( .A(n124), .B(n125), .Z(n112) );
  AND U88 ( .A(n126), .B(n127), .Z(n125) );
  XOR U89 ( .A(n124), .B(n49), .Z(n127) );
  XOR U90 ( .A(n128), .B(n129), .Z(n49) );
  AND U91 ( .A(n87), .B(n130), .Z(n129) );
  XOR U92 ( .A(n131), .B(n128), .Z(n130) );
  XNOR U93 ( .A(n50), .B(n124), .Z(n126) );
  IV U94 ( .A(n47), .Z(n50) );
  XNOR U95 ( .A(n132), .B(n133), .Z(n47) );
  AND U96 ( .A(n84), .B(n134), .Z(n133) );
  XOR U97 ( .A(n135), .B(n132), .Z(n134) );
  XOR U98 ( .A(n136), .B(n137), .Z(n124) );
  AND U99 ( .A(n138), .B(n139), .Z(n137) );
  XOR U100 ( .A(n136), .B(n54), .Z(n139) );
  XOR U101 ( .A(n140), .B(n141), .Z(n54) );
  AND U102 ( .A(n87), .B(n142), .Z(n141) );
  XOR U103 ( .A(n143), .B(n140), .Z(n142) );
  XNOR U104 ( .A(n55), .B(n136), .Z(n138) );
  IV U105 ( .A(n52), .Z(n55) );
  XNOR U106 ( .A(n144), .B(n145), .Z(n52) );
  AND U107 ( .A(n84), .B(n146), .Z(n145) );
  XOR U108 ( .A(n147), .B(n144), .Z(n146) );
  XOR U109 ( .A(n148), .B(n149), .Z(n136) );
  AND U110 ( .A(n150), .B(n151), .Z(n149) );
  XOR U111 ( .A(n148), .B(n59), .Z(n151) );
  XOR U112 ( .A(n152), .B(n153), .Z(n59) );
  AND U113 ( .A(n87), .B(n154), .Z(n153) );
  XOR U114 ( .A(n155), .B(n152), .Z(n154) );
  XNOR U115 ( .A(n60), .B(n148), .Z(n150) );
  IV U116 ( .A(n57), .Z(n60) );
  XNOR U117 ( .A(n156), .B(n157), .Z(n57) );
  AND U118 ( .A(n84), .B(n158), .Z(n157) );
  XOR U119 ( .A(n159), .B(n156), .Z(n158) );
  XOR U120 ( .A(n160), .B(n161), .Z(n148) );
  AND U121 ( .A(n162), .B(n163), .Z(n161) );
  XOR U122 ( .A(n160), .B(n64), .Z(n163) );
  XOR U123 ( .A(n164), .B(n165), .Z(n64) );
  AND U124 ( .A(n87), .B(n166), .Z(n165) );
  XOR U125 ( .A(n167), .B(n164), .Z(n166) );
  XNOR U126 ( .A(n65), .B(n160), .Z(n162) );
  IV U127 ( .A(n62), .Z(n65) );
  XNOR U128 ( .A(n168), .B(n169), .Z(n62) );
  AND U129 ( .A(n84), .B(n170), .Z(n169) );
  XOR U130 ( .A(n171), .B(n168), .Z(n170) );
  XOR U131 ( .A(n172), .B(n173), .Z(n160) );
  AND U132 ( .A(n174), .B(n175), .Z(n173) );
  XOR U133 ( .A(n172), .B(n69), .Z(n175) );
  XOR U134 ( .A(n176), .B(n177), .Z(n69) );
  AND U135 ( .A(n87), .B(n178), .Z(n177) );
  XOR U136 ( .A(n179), .B(n176), .Z(n178) );
  XNOR U137 ( .A(n70), .B(n172), .Z(n174) );
  IV U138 ( .A(n67), .Z(n70) );
  XNOR U139 ( .A(n180), .B(n181), .Z(n67) );
  AND U140 ( .A(n84), .B(n182), .Z(n181) );
  XOR U141 ( .A(n183), .B(n180), .Z(n182) );
  XOR U142 ( .A(n184), .B(n185), .Z(n172) );
  AND U143 ( .A(n186), .B(n187), .Z(n185) );
  XOR U144 ( .A(n184), .B(n74), .Z(n187) );
  XOR U145 ( .A(n188), .B(n189), .Z(n74) );
  AND U146 ( .A(n87), .B(n190), .Z(n189) );
  XOR U147 ( .A(n191), .B(n188), .Z(n190) );
  XNOR U148 ( .A(n75), .B(n184), .Z(n186) );
  IV U149 ( .A(n72), .Z(n75) );
  XNOR U150 ( .A(n192), .B(n193), .Z(n72) );
  AND U151 ( .A(n84), .B(n194), .Z(n193) );
  XOR U152 ( .A(n195), .B(n192), .Z(n194) );
  XOR U153 ( .A(n196), .B(n197), .Z(n184) );
  AND U154 ( .A(n198), .B(n199), .Z(n197) );
  XOR U155 ( .A(n4), .B(n196), .Z(n199) );
  XOR U156 ( .A(n200), .B(n201), .Z(n4) );
  AND U157 ( .A(n87), .B(n202), .Z(n201) );
  XOR U158 ( .A(n200), .B(n203), .Z(n202) );
  XNOR U159 ( .A(n196), .B(n2), .Z(n198) );
  XOR U160 ( .A(n204), .B(n205), .Z(n2) );
  AND U161 ( .A(n84), .B(n206), .Z(n205) );
  XOR U162 ( .A(n204), .B(n207), .Z(n206) );
  XOR U163 ( .A(n208), .B(n209), .Z(n196) );
  AND U164 ( .A(n210), .B(n211), .Z(n209) );
  XOR U165 ( .A(n208), .B(n8), .Z(n211) );
  XOR U166 ( .A(n212), .B(n213), .Z(n8) );
  AND U167 ( .A(n87), .B(n214), .Z(n213) );
  XOR U168 ( .A(n215), .B(n212), .Z(n214) );
  XNOR U169 ( .A(n9), .B(n208), .Z(n210) );
  IV U170 ( .A(n6), .Z(n9) );
  XNOR U171 ( .A(n216), .B(n217), .Z(n6) );
  AND U172 ( .A(n84), .B(n218), .Z(n217) );
  XOR U173 ( .A(n219), .B(n216), .Z(n218) );
  XOR U174 ( .A(n220), .B(n221), .Z(n208) );
  AND U175 ( .A(n222), .B(n223), .Z(n221) );
  XOR U176 ( .A(n220), .B(n13), .Z(n223) );
  XOR U177 ( .A(n224), .B(n225), .Z(n13) );
  AND U178 ( .A(n87), .B(n226), .Z(n225) );
  XOR U179 ( .A(n227), .B(n224), .Z(n226) );
  XNOR U180 ( .A(n14), .B(n220), .Z(n222) );
  IV U181 ( .A(n11), .Z(n14) );
  XNOR U182 ( .A(n228), .B(n229), .Z(n11) );
  AND U183 ( .A(n84), .B(n230), .Z(n229) );
  XOR U184 ( .A(n231), .B(n228), .Z(n230) );
  XOR U185 ( .A(n232), .B(n233), .Z(n220) );
  AND U186 ( .A(n234), .B(n235), .Z(n233) );
  XOR U187 ( .A(n232), .B(n18), .Z(n235) );
  XOR U188 ( .A(n236), .B(n237), .Z(n18) );
  AND U189 ( .A(n87), .B(n238), .Z(n237) );
  XOR U190 ( .A(n239), .B(n236), .Z(n238) );
  XNOR U191 ( .A(n19), .B(n232), .Z(n234) );
  IV U192 ( .A(n16), .Z(n19) );
  XNOR U193 ( .A(n240), .B(n241), .Z(n16) );
  AND U194 ( .A(n84), .B(n242), .Z(n241) );
  XOR U195 ( .A(n243), .B(n240), .Z(n242) );
  XOR U196 ( .A(n244), .B(n245), .Z(n232) );
  AND U197 ( .A(n246), .B(n247), .Z(n245) );
  XOR U198 ( .A(n244), .B(n23), .Z(n247) );
  XOR U199 ( .A(n248), .B(n249), .Z(n23) );
  AND U200 ( .A(n87), .B(n250), .Z(n249) );
  XOR U201 ( .A(n251), .B(n248), .Z(n250) );
  XNOR U202 ( .A(n24), .B(n244), .Z(n246) );
  IV U203 ( .A(n21), .Z(n24) );
  XNOR U204 ( .A(n252), .B(n253), .Z(n21) );
  AND U205 ( .A(n84), .B(n254), .Z(n253) );
  XOR U206 ( .A(n255), .B(n252), .Z(n254) );
  XNOR U207 ( .A(n256), .B(n257), .Z(n244) );
  AND U208 ( .A(n258), .B(n259), .Z(n257) );
  XNOR U209 ( .A(n256), .B(n28), .Z(n259) );
  XOR U210 ( .A(n260), .B(n261), .Z(n28) );
  AND U211 ( .A(n87), .B(n262), .Z(n261) );
  XOR U212 ( .A(n263), .B(n260), .Z(n262) );
  XOR U213 ( .A(n29), .B(n256), .Z(n258) );
  IV U214 ( .A(n26), .Z(n29) );
  XNOR U215 ( .A(n264), .B(n265), .Z(n26) );
  AND U216 ( .A(n84), .B(n266), .Z(n265) );
  XOR U217 ( .A(n267), .B(n264), .Z(n266) );
  AND U218 ( .A(n31), .B(n33), .Z(n256) );
  XNOR U219 ( .A(n268), .B(n269), .Z(n33) );
  AND U220 ( .A(n87), .B(n270), .Z(n269) );
  XNOR U221 ( .A(n271), .B(n268), .Z(n270) );
  XOR U222 ( .A(n272), .B(n273), .Z(n87) );
  AND U223 ( .A(n274), .B(n275), .Z(n273) );
  XNOR U224 ( .A(n96), .B(n272), .Z(n275) );
  AND U225 ( .A(p_input[127]), .B(p_input[111]), .Z(n96) );
  XOR U226 ( .A(n272), .B(n97), .Z(n274) );
  AND U227 ( .A(p_input[95]), .B(p_input[79]), .Z(n97) );
  XOR U228 ( .A(n276), .B(n277), .Z(n272) );
  AND U229 ( .A(n278), .B(n279), .Z(n277) );
  XOR U230 ( .A(n276), .B(n107), .Z(n279) );
  XNOR U231 ( .A(p_input[110]), .B(n280), .Z(n107) );
  AND U232 ( .A(n83), .B(n281), .Z(n280) );
  XOR U233 ( .A(p_input[126]), .B(p_input[110]), .Z(n281) );
  XNOR U234 ( .A(n104), .B(n276), .Z(n278) );
  XOR U235 ( .A(n282), .B(n283), .Z(n104) );
  AND U236 ( .A(n81), .B(n284), .Z(n283) );
  XOR U237 ( .A(p_input[94]), .B(p_input[78]), .Z(n284) );
  XOR U238 ( .A(n285), .B(n286), .Z(n276) );
  AND U239 ( .A(n287), .B(n288), .Z(n286) );
  XOR U240 ( .A(n285), .B(n119), .Z(n288) );
  XNOR U241 ( .A(p_input[109]), .B(n289), .Z(n119) );
  AND U242 ( .A(n83), .B(n290), .Z(n289) );
  XOR U243 ( .A(p_input[125]), .B(p_input[109]), .Z(n290) );
  XNOR U244 ( .A(n116), .B(n285), .Z(n287) );
  XOR U245 ( .A(n291), .B(n292), .Z(n116) );
  AND U246 ( .A(n81), .B(n293), .Z(n292) );
  XOR U247 ( .A(p_input[93]), .B(p_input[77]), .Z(n293) );
  XOR U248 ( .A(n294), .B(n295), .Z(n285) );
  AND U249 ( .A(n296), .B(n297), .Z(n295) );
  XOR U250 ( .A(n294), .B(n131), .Z(n297) );
  XNOR U251 ( .A(p_input[108]), .B(n298), .Z(n131) );
  AND U252 ( .A(n83), .B(n299), .Z(n298) );
  XOR U253 ( .A(p_input[124]), .B(p_input[108]), .Z(n299) );
  XNOR U254 ( .A(n128), .B(n294), .Z(n296) );
  XOR U255 ( .A(n300), .B(n301), .Z(n128) );
  AND U256 ( .A(n81), .B(n302), .Z(n301) );
  XOR U257 ( .A(p_input[92]), .B(p_input[76]), .Z(n302) );
  XOR U258 ( .A(n303), .B(n304), .Z(n294) );
  AND U259 ( .A(n305), .B(n306), .Z(n304) );
  XOR U260 ( .A(n303), .B(n143), .Z(n306) );
  XNOR U261 ( .A(p_input[107]), .B(n307), .Z(n143) );
  AND U262 ( .A(n83), .B(n308), .Z(n307) );
  XOR U263 ( .A(p_input[123]), .B(p_input[107]), .Z(n308) );
  XNOR U264 ( .A(n140), .B(n303), .Z(n305) );
  XOR U265 ( .A(n309), .B(n310), .Z(n140) );
  AND U266 ( .A(n81), .B(n311), .Z(n310) );
  XOR U267 ( .A(p_input[91]), .B(p_input[75]), .Z(n311) );
  XOR U268 ( .A(n312), .B(n313), .Z(n303) );
  AND U269 ( .A(n314), .B(n315), .Z(n313) );
  XOR U270 ( .A(n312), .B(n155), .Z(n315) );
  XNOR U271 ( .A(p_input[106]), .B(n316), .Z(n155) );
  AND U272 ( .A(n83), .B(n317), .Z(n316) );
  XOR U273 ( .A(p_input[122]), .B(p_input[106]), .Z(n317) );
  XNOR U274 ( .A(n152), .B(n312), .Z(n314) );
  XOR U275 ( .A(n318), .B(n319), .Z(n152) );
  AND U276 ( .A(n81), .B(n320), .Z(n319) );
  XOR U277 ( .A(p_input[90]), .B(p_input[74]), .Z(n320) );
  XOR U278 ( .A(n321), .B(n322), .Z(n312) );
  AND U279 ( .A(n323), .B(n324), .Z(n322) );
  XOR U280 ( .A(n321), .B(n167), .Z(n324) );
  XNOR U281 ( .A(p_input[105]), .B(n325), .Z(n167) );
  AND U282 ( .A(n83), .B(n326), .Z(n325) );
  XOR U283 ( .A(p_input[121]), .B(p_input[105]), .Z(n326) );
  XNOR U284 ( .A(n164), .B(n321), .Z(n323) );
  XOR U285 ( .A(n327), .B(n328), .Z(n164) );
  AND U286 ( .A(n81), .B(n329), .Z(n328) );
  XOR U287 ( .A(p_input[89]), .B(p_input[73]), .Z(n329) );
  XOR U288 ( .A(n330), .B(n331), .Z(n321) );
  AND U289 ( .A(n332), .B(n333), .Z(n331) );
  XOR U290 ( .A(n330), .B(n179), .Z(n333) );
  XNOR U291 ( .A(p_input[104]), .B(n334), .Z(n179) );
  AND U292 ( .A(n83), .B(n335), .Z(n334) );
  XOR U293 ( .A(p_input[120]), .B(p_input[104]), .Z(n335) );
  XNOR U294 ( .A(n176), .B(n330), .Z(n332) );
  XOR U295 ( .A(n336), .B(n337), .Z(n176) );
  AND U296 ( .A(n81), .B(n338), .Z(n337) );
  XOR U297 ( .A(p_input[88]), .B(p_input[72]), .Z(n338) );
  XOR U298 ( .A(n339), .B(n340), .Z(n330) );
  AND U299 ( .A(n341), .B(n342), .Z(n340) );
  XOR U300 ( .A(n339), .B(n191), .Z(n342) );
  XNOR U301 ( .A(p_input[103]), .B(n343), .Z(n191) );
  AND U302 ( .A(n83), .B(n344), .Z(n343) );
  XOR U303 ( .A(p_input[119]), .B(p_input[103]), .Z(n344) );
  XNOR U304 ( .A(n188), .B(n339), .Z(n341) );
  XOR U305 ( .A(n345), .B(n346), .Z(n188) );
  AND U306 ( .A(n81), .B(n347), .Z(n346) );
  XOR U307 ( .A(p_input[87]), .B(p_input[71]), .Z(n347) );
  XOR U308 ( .A(n348), .B(n349), .Z(n339) );
  AND U309 ( .A(n350), .B(n351), .Z(n349) );
  XOR U310 ( .A(n203), .B(n348), .Z(n351) );
  XNOR U311 ( .A(p_input[102]), .B(n352), .Z(n203) );
  AND U312 ( .A(n83), .B(n353), .Z(n352) );
  XOR U313 ( .A(p_input[118]), .B(p_input[102]), .Z(n353) );
  XNOR U314 ( .A(n348), .B(n200), .Z(n350) );
  XOR U315 ( .A(n354), .B(n355), .Z(n200) );
  AND U316 ( .A(n81), .B(n356), .Z(n355) );
  XOR U317 ( .A(p_input[86]), .B(p_input[70]), .Z(n356) );
  XOR U318 ( .A(n357), .B(n358), .Z(n348) );
  AND U319 ( .A(n359), .B(n360), .Z(n358) );
  XOR U320 ( .A(n357), .B(n215), .Z(n360) );
  XNOR U321 ( .A(p_input[101]), .B(n361), .Z(n215) );
  AND U322 ( .A(n83), .B(n362), .Z(n361) );
  XOR U323 ( .A(p_input[117]), .B(p_input[101]), .Z(n362) );
  XNOR U324 ( .A(n212), .B(n357), .Z(n359) );
  XOR U325 ( .A(n363), .B(n364), .Z(n212) );
  AND U326 ( .A(n81), .B(n365), .Z(n364) );
  XOR U327 ( .A(p_input[85]), .B(p_input[69]), .Z(n365) );
  XOR U328 ( .A(n366), .B(n367), .Z(n357) );
  AND U329 ( .A(n368), .B(n369), .Z(n367) );
  XOR U330 ( .A(n366), .B(n227), .Z(n369) );
  XNOR U331 ( .A(p_input[100]), .B(n370), .Z(n227) );
  AND U332 ( .A(n83), .B(n371), .Z(n370) );
  XOR U333 ( .A(p_input[116]), .B(p_input[100]), .Z(n371) );
  XNOR U334 ( .A(n224), .B(n366), .Z(n368) );
  XOR U335 ( .A(n372), .B(n373), .Z(n224) );
  AND U336 ( .A(n81), .B(n374), .Z(n373) );
  XOR U337 ( .A(p_input[84]), .B(p_input[68]), .Z(n374) );
  XOR U338 ( .A(n375), .B(n376), .Z(n366) );
  AND U339 ( .A(n377), .B(n378), .Z(n376) );
  XOR U340 ( .A(n375), .B(n239), .Z(n378) );
  XNOR U341 ( .A(p_input[99]), .B(n379), .Z(n239) );
  AND U342 ( .A(n83), .B(n380), .Z(n379) );
  XOR U343 ( .A(p_input[99]), .B(p_input[115]), .Z(n380) );
  XNOR U344 ( .A(n236), .B(n375), .Z(n377) );
  XOR U345 ( .A(n381), .B(n382), .Z(n236) );
  AND U346 ( .A(n81), .B(n383), .Z(n382) );
  XOR U347 ( .A(p_input[83]), .B(p_input[67]), .Z(n383) );
  XOR U348 ( .A(n384), .B(n385), .Z(n375) );
  AND U349 ( .A(n386), .B(n387), .Z(n385) );
  XOR U350 ( .A(n384), .B(n251), .Z(n387) );
  XNOR U351 ( .A(p_input[98]), .B(n388), .Z(n251) );
  AND U352 ( .A(n83), .B(n389), .Z(n388) );
  XOR U353 ( .A(p_input[98]), .B(p_input[114]), .Z(n389) );
  XNOR U354 ( .A(n248), .B(n384), .Z(n386) );
  XOR U355 ( .A(n390), .B(n391), .Z(n248) );
  AND U356 ( .A(n81), .B(n392), .Z(n391) );
  XOR U357 ( .A(p_input[82]), .B(p_input[66]), .Z(n392) );
  XOR U358 ( .A(n393), .B(n394), .Z(n384) );
  AND U359 ( .A(n395), .B(n396), .Z(n394) );
  XNOR U360 ( .A(n397), .B(n263), .Z(n396) );
  XNOR U361 ( .A(p_input[97]), .B(n398), .Z(n263) );
  AND U362 ( .A(n83), .B(n399), .Z(n398) );
  XNOR U363 ( .A(n400), .B(p_input[113]), .Z(n399) );
  IV U364 ( .A(p_input[97]), .Z(n400) );
  XNOR U365 ( .A(n260), .B(n393), .Z(n395) );
  XNOR U366 ( .A(p_input[65]), .B(n401), .Z(n260) );
  AND U367 ( .A(n81), .B(n402), .Z(n401) );
  XOR U368 ( .A(p_input[81]), .B(p_input[65]), .Z(n402) );
  IV U369 ( .A(n397), .Z(n393) );
  AND U370 ( .A(n268), .B(n271), .Z(n397) );
  XOR U371 ( .A(p_input[96]), .B(n403), .Z(n271) );
  AND U372 ( .A(n83), .B(n404), .Z(n403) );
  XOR U373 ( .A(p_input[96]), .B(p_input[112]), .Z(n404) );
  XOR U374 ( .A(n405), .B(n406), .Z(n83) );
  AND U375 ( .A(n407), .B(n408), .Z(n406) );
  XNOR U376 ( .A(p_input[127]), .B(n405), .Z(n408) );
  XOR U377 ( .A(n405), .B(p_input[111]), .Z(n407) );
  XOR U378 ( .A(n409), .B(n410), .Z(n405) );
  AND U379 ( .A(n411), .B(n412), .Z(n410) );
  XNOR U380 ( .A(p_input[126]), .B(n409), .Z(n412) );
  XOR U381 ( .A(n409), .B(p_input[110]), .Z(n411) );
  XOR U382 ( .A(n413), .B(n414), .Z(n409) );
  AND U383 ( .A(n415), .B(n416), .Z(n414) );
  XNOR U384 ( .A(p_input[125]), .B(n413), .Z(n416) );
  XOR U385 ( .A(n413), .B(p_input[109]), .Z(n415) );
  XOR U386 ( .A(n417), .B(n418), .Z(n413) );
  AND U387 ( .A(n419), .B(n420), .Z(n418) );
  XNOR U388 ( .A(p_input[124]), .B(n417), .Z(n420) );
  XOR U389 ( .A(n417), .B(p_input[108]), .Z(n419) );
  XOR U390 ( .A(n421), .B(n422), .Z(n417) );
  AND U391 ( .A(n423), .B(n424), .Z(n422) );
  XNOR U392 ( .A(p_input[123]), .B(n421), .Z(n424) );
  XOR U393 ( .A(n421), .B(p_input[107]), .Z(n423) );
  XOR U394 ( .A(n425), .B(n426), .Z(n421) );
  AND U395 ( .A(n427), .B(n428), .Z(n426) );
  XNOR U396 ( .A(p_input[122]), .B(n425), .Z(n428) );
  XOR U397 ( .A(n425), .B(p_input[106]), .Z(n427) );
  XOR U398 ( .A(n429), .B(n430), .Z(n425) );
  AND U399 ( .A(n431), .B(n432), .Z(n430) );
  XNOR U400 ( .A(p_input[121]), .B(n429), .Z(n432) );
  XOR U401 ( .A(n429), .B(p_input[105]), .Z(n431) );
  XOR U402 ( .A(n433), .B(n434), .Z(n429) );
  AND U403 ( .A(n435), .B(n436), .Z(n434) );
  XNOR U404 ( .A(p_input[120]), .B(n433), .Z(n436) );
  XOR U405 ( .A(n433), .B(p_input[104]), .Z(n435) );
  XOR U406 ( .A(n437), .B(n438), .Z(n433) );
  AND U407 ( .A(n439), .B(n440), .Z(n438) );
  XNOR U408 ( .A(p_input[119]), .B(n437), .Z(n440) );
  XOR U409 ( .A(n437), .B(p_input[103]), .Z(n439) );
  XOR U410 ( .A(n441), .B(n442), .Z(n437) );
  AND U411 ( .A(n443), .B(n444), .Z(n442) );
  XNOR U412 ( .A(p_input[118]), .B(n441), .Z(n444) );
  XOR U413 ( .A(n441), .B(p_input[102]), .Z(n443) );
  XOR U414 ( .A(n445), .B(n446), .Z(n441) );
  AND U415 ( .A(n447), .B(n448), .Z(n446) );
  XNOR U416 ( .A(p_input[117]), .B(n445), .Z(n448) );
  XOR U417 ( .A(n445), .B(p_input[101]), .Z(n447) );
  XOR U418 ( .A(n449), .B(n450), .Z(n445) );
  AND U419 ( .A(n451), .B(n452), .Z(n450) );
  XNOR U420 ( .A(p_input[116]), .B(n449), .Z(n452) );
  XOR U421 ( .A(n449), .B(p_input[100]), .Z(n451) );
  XOR U422 ( .A(n453), .B(n454), .Z(n449) );
  AND U423 ( .A(n455), .B(n456), .Z(n454) );
  XNOR U424 ( .A(p_input[115]), .B(n453), .Z(n456) );
  XOR U425 ( .A(n453), .B(p_input[99]), .Z(n455) );
  XOR U426 ( .A(n457), .B(n458), .Z(n453) );
  AND U427 ( .A(n459), .B(n460), .Z(n458) );
  XNOR U428 ( .A(p_input[114]), .B(n457), .Z(n460) );
  XOR U429 ( .A(n457), .B(p_input[98]), .Z(n459) );
  XNOR U430 ( .A(n461), .B(n462), .Z(n457) );
  AND U431 ( .A(n463), .B(n464), .Z(n462) );
  XOR U432 ( .A(p_input[113]), .B(n461), .Z(n464) );
  XNOR U433 ( .A(p_input[97]), .B(n461), .Z(n463) );
  AND U434 ( .A(p_input[112]), .B(n465), .Z(n461) );
  IV U435 ( .A(p_input[96]), .Z(n465) );
  XNOR U436 ( .A(p_input[64]), .B(n466), .Z(n268) );
  AND U437 ( .A(n81), .B(n467), .Z(n466) );
  XOR U438 ( .A(p_input[80]), .B(p_input[64]), .Z(n467) );
  XOR U439 ( .A(n468), .B(n469), .Z(n81) );
  AND U440 ( .A(n470), .B(n471), .Z(n469) );
  XNOR U441 ( .A(p_input[95]), .B(n468), .Z(n471) );
  XOR U442 ( .A(n468), .B(p_input[79]), .Z(n470) );
  XOR U443 ( .A(n472), .B(n473), .Z(n468) );
  AND U444 ( .A(n474), .B(n475), .Z(n473) );
  XNOR U445 ( .A(p_input[94]), .B(n472), .Z(n475) );
  XNOR U446 ( .A(n472), .B(n282), .Z(n474) );
  IV U447 ( .A(p_input[78]), .Z(n282) );
  XOR U448 ( .A(n476), .B(n477), .Z(n472) );
  AND U449 ( .A(n478), .B(n479), .Z(n477) );
  XNOR U450 ( .A(p_input[93]), .B(n476), .Z(n479) );
  XNOR U451 ( .A(n476), .B(n291), .Z(n478) );
  IV U452 ( .A(p_input[77]), .Z(n291) );
  XOR U453 ( .A(n480), .B(n481), .Z(n476) );
  AND U454 ( .A(n482), .B(n483), .Z(n481) );
  XNOR U455 ( .A(p_input[92]), .B(n480), .Z(n483) );
  XNOR U456 ( .A(n480), .B(n300), .Z(n482) );
  IV U457 ( .A(p_input[76]), .Z(n300) );
  XOR U458 ( .A(n484), .B(n485), .Z(n480) );
  AND U459 ( .A(n486), .B(n487), .Z(n485) );
  XNOR U460 ( .A(p_input[91]), .B(n484), .Z(n487) );
  XNOR U461 ( .A(n484), .B(n309), .Z(n486) );
  IV U462 ( .A(p_input[75]), .Z(n309) );
  XOR U463 ( .A(n488), .B(n489), .Z(n484) );
  AND U464 ( .A(n490), .B(n491), .Z(n489) );
  XNOR U465 ( .A(p_input[90]), .B(n488), .Z(n491) );
  XNOR U466 ( .A(n488), .B(n318), .Z(n490) );
  IV U467 ( .A(p_input[74]), .Z(n318) );
  XOR U468 ( .A(n492), .B(n493), .Z(n488) );
  AND U469 ( .A(n494), .B(n495), .Z(n493) );
  XNOR U470 ( .A(p_input[89]), .B(n492), .Z(n495) );
  XNOR U471 ( .A(n492), .B(n327), .Z(n494) );
  IV U472 ( .A(p_input[73]), .Z(n327) );
  XOR U473 ( .A(n496), .B(n497), .Z(n492) );
  AND U474 ( .A(n498), .B(n499), .Z(n497) );
  XNOR U475 ( .A(p_input[88]), .B(n496), .Z(n499) );
  XNOR U476 ( .A(n496), .B(n336), .Z(n498) );
  IV U477 ( .A(p_input[72]), .Z(n336) );
  XOR U478 ( .A(n500), .B(n501), .Z(n496) );
  AND U479 ( .A(n502), .B(n503), .Z(n501) );
  XNOR U480 ( .A(p_input[87]), .B(n500), .Z(n503) );
  XNOR U481 ( .A(n500), .B(n345), .Z(n502) );
  IV U482 ( .A(p_input[71]), .Z(n345) );
  XOR U483 ( .A(n504), .B(n505), .Z(n500) );
  AND U484 ( .A(n506), .B(n507), .Z(n505) );
  XNOR U485 ( .A(p_input[86]), .B(n504), .Z(n507) );
  XNOR U486 ( .A(n504), .B(n354), .Z(n506) );
  IV U487 ( .A(p_input[70]), .Z(n354) );
  XOR U488 ( .A(n508), .B(n509), .Z(n504) );
  AND U489 ( .A(n510), .B(n511), .Z(n509) );
  XNOR U490 ( .A(p_input[85]), .B(n508), .Z(n511) );
  XNOR U491 ( .A(n508), .B(n363), .Z(n510) );
  IV U492 ( .A(p_input[69]), .Z(n363) );
  XOR U493 ( .A(n512), .B(n513), .Z(n508) );
  AND U494 ( .A(n514), .B(n515), .Z(n513) );
  XNOR U495 ( .A(p_input[84]), .B(n512), .Z(n515) );
  XNOR U496 ( .A(n512), .B(n372), .Z(n514) );
  IV U497 ( .A(p_input[68]), .Z(n372) );
  XOR U498 ( .A(n516), .B(n517), .Z(n512) );
  AND U499 ( .A(n518), .B(n519), .Z(n517) );
  XNOR U500 ( .A(p_input[83]), .B(n516), .Z(n519) );
  XNOR U501 ( .A(n516), .B(n381), .Z(n518) );
  IV U502 ( .A(p_input[67]), .Z(n381) );
  XOR U503 ( .A(n520), .B(n521), .Z(n516) );
  AND U504 ( .A(n522), .B(n523), .Z(n521) );
  XNOR U505 ( .A(p_input[82]), .B(n520), .Z(n523) );
  XNOR U506 ( .A(n520), .B(n390), .Z(n522) );
  IV U507 ( .A(p_input[66]), .Z(n390) );
  XNOR U508 ( .A(n524), .B(n525), .Z(n520) );
  AND U509 ( .A(n526), .B(n527), .Z(n525) );
  XOR U510 ( .A(p_input[81]), .B(n524), .Z(n527) );
  XNOR U511 ( .A(p_input[65]), .B(n524), .Z(n526) );
  AND U512 ( .A(p_input[80]), .B(n528), .Z(n524) );
  IV U513 ( .A(p_input[64]), .Z(n528) );
  XOR U514 ( .A(n529), .B(n530), .Z(n31) );
  AND U515 ( .A(n84), .B(n531), .Z(n530) );
  XNOR U516 ( .A(n532), .B(n529), .Z(n531) );
  XOR U517 ( .A(n533), .B(n534), .Z(n84) );
  AND U518 ( .A(n535), .B(n536), .Z(n534) );
  XNOR U519 ( .A(n99), .B(n533), .Z(n536) );
  AND U520 ( .A(p_input[63]), .B(p_input[47]), .Z(n99) );
  XOR U521 ( .A(n533), .B(n98), .Z(n535) );
  AND U522 ( .A(p_input[15]), .B(p_input[31]), .Z(n98) );
  XOR U523 ( .A(n537), .B(n538), .Z(n533) );
  AND U524 ( .A(n539), .B(n540), .Z(n538) );
  XOR U525 ( .A(n537), .B(n111), .Z(n540) );
  XNOR U526 ( .A(p_input[46]), .B(n541), .Z(n111) );
  AND U527 ( .A(n91), .B(n542), .Z(n541) );
  XOR U528 ( .A(p_input[62]), .B(p_input[46]), .Z(n542) );
  XNOR U529 ( .A(n108), .B(n537), .Z(n539) );
  XOR U530 ( .A(n543), .B(n544), .Z(n108) );
  AND U531 ( .A(n88), .B(n545), .Z(n544) );
  XOR U532 ( .A(p_input[30]), .B(p_input[14]), .Z(n545) );
  XOR U533 ( .A(n546), .B(n547), .Z(n537) );
  AND U534 ( .A(n548), .B(n549), .Z(n547) );
  XOR U535 ( .A(n546), .B(n123), .Z(n549) );
  XNOR U536 ( .A(p_input[45]), .B(n550), .Z(n123) );
  AND U537 ( .A(n91), .B(n551), .Z(n550) );
  XOR U538 ( .A(p_input[61]), .B(p_input[45]), .Z(n551) );
  XNOR U539 ( .A(n120), .B(n546), .Z(n548) );
  XOR U540 ( .A(n552), .B(n553), .Z(n120) );
  AND U541 ( .A(n88), .B(n554), .Z(n553) );
  XOR U542 ( .A(p_input[29]), .B(p_input[13]), .Z(n554) );
  XOR U543 ( .A(n555), .B(n556), .Z(n546) );
  AND U544 ( .A(n557), .B(n558), .Z(n556) );
  XOR U545 ( .A(n555), .B(n135), .Z(n558) );
  XNOR U546 ( .A(p_input[44]), .B(n559), .Z(n135) );
  AND U547 ( .A(n91), .B(n560), .Z(n559) );
  XOR U548 ( .A(p_input[60]), .B(p_input[44]), .Z(n560) );
  XNOR U549 ( .A(n132), .B(n555), .Z(n557) );
  XOR U550 ( .A(n561), .B(n562), .Z(n132) );
  AND U551 ( .A(n88), .B(n563), .Z(n562) );
  XOR U552 ( .A(p_input[28]), .B(p_input[12]), .Z(n563) );
  XOR U553 ( .A(n564), .B(n565), .Z(n555) );
  AND U554 ( .A(n566), .B(n567), .Z(n565) );
  XOR U555 ( .A(n564), .B(n147), .Z(n567) );
  XNOR U556 ( .A(p_input[43]), .B(n568), .Z(n147) );
  AND U557 ( .A(n91), .B(n569), .Z(n568) );
  XOR U558 ( .A(p_input[59]), .B(p_input[43]), .Z(n569) );
  XNOR U559 ( .A(n144), .B(n564), .Z(n566) );
  XOR U560 ( .A(n570), .B(n571), .Z(n144) );
  AND U561 ( .A(n88), .B(n572), .Z(n571) );
  XOR U562 ( .A(p_input[27]), .B(p_input[11]), .Z(n572) );
  XOR U563 ( .A(n573), .B(n574), .Z(n564) );
  AND U564 ( .A(n575), .B(n576), .Z(n574) );
  XOR U565 ( .A(n573), .B(n159), .Z(n576) );
  XNOR U566 ( .A(p_input[42]), .B(n577), .Z(n159) );
  AND U567 ( .A(n91), .B(n578), .Z(n577) );
  XOR U568 ( .A(p_input[58]), .B(p_input[42]), .Z(n578) );
  XNOR U569 ( .A(n156), .B(n573), .Z(n575) );
  XOR U570 ( .A(n579), .B(n580), .Z(n156) );
  AND U571 ( .A(n88), .B(n581), .Z(n580) );
  XOR U572 ( .A(p_input[26]), .B(p_input[10]), .Z(n581) );
  XOR U573 ( .A(n582), .B(n583), .Z(n573) );
  AND U574 ( .A(n584), .B(n585), .Z(n583) );
  XOR U575 ( .A(n582), .B(n171), .Z(n585) );
  XNOR U576 ( .A(p_input[41]), .B(n586), .Z(n171) );
  AND U577 ( .A(n91), .B(n587), .Z(n586) );
  XOR U578 ( .A(p_input[57]), .B(p_input[41]), .Z(n587) );
  XNOR U579 ( .A(n168), .B(n582), .Z(n584) );
  XOR U580 ( .A(n588), .B(n589), .Z(n168) );
  AND U581 ( .A(n88), .B(n590), .Z(n589) );
  XOR U582 ( .A(p_input[9]), .B(p_input[25]), .Z(n590) );
  XOR U583 ( .A(n591), .B(n592), .Z(n582) );
  AND U584 ( .A(n593), .B(n594), .Z(n592) );
  XOR U585 ( .A(n591), .B(n183), .Z(n594) );
  XNOR U586 ( .A(p_input[40]), .B(n595), .Z(n183) );
  AND U587 ( .A(n91), .B(n596), .Z(n595) );
  XOR U588 ( .A(p_input[56]), .B(p_input[40]), .Z(n596) );
  XNOR U589 ( .A(n180), .B(n591), .Z(n593) );
  XOR U590 ( .A(n597), .B(n598), .Z(n180) );
  AND U591 ( .A(n88), .B(n599), .Z(n598) );
  XOR U592 ( .A(p_input[8]), .B(p_input[24]), .Z(n599) );
  XOR U593 ( .A(n600), .B(n601), .Z(n591) );
  AND U594 ( .A(n602), .B(n603), .Z(n601) );
  XOR U595 ( .A(n600), .B(n195), .Z(n603) );
  XNOR U596 ( .A(p_input[39]), .B(n604), .Z(n195) );
  AND U597 ( .A(n91), .B(n605), .Z(n604) );
  XOR U598 ( .A(p_input[55]), .B(p_input[39]), .Z(n605) );
  XNOR U599 ( .A(n192), .B(n600), .Z(n602) );
  XOR U600 ( .A(n606), .B(n607), .Z(n192) );
  AND U601 ( .A(n88), .B(n608), .Z(n607) );
  XOR U602 ( .A(p_input[7]), .B(p_input[23]), .Z(n608) );
  XOR U603 ( .A(n609), .B(n610), .Z(n600) );
  AND U604 ( .A(n611), .B(n612), .Z(n610) );
  XOR U605 ( .A(n207), .B(n609), .Z(n612) );
  XNOR U606 ( .A(p_input[38]), .B(n613), .Z(n207) );
  AND U607 ( .A(n91), .B(n614), .Z(n613) );
  XOR U608 ( .A(p_input[54]), .B(p_input[38]), .Z(n614) );
  XNOR U609 ( .A(n609), .B(n204), .Z(n611) );
  XOR U610 ( .A(n615), .B(n616), .Z(n204) );
  AND U611 ( .A(n88), .B(n617), .Z(n616) );
  XOR U612 ( .A(p_input[6]), .B(p_input[22]), .Z(n617) );
  XOR U613 ( .A(n618), .B(n619), .Z(n609) );
  AND U614 ( .A(n620), .B(n621), .Z(n619) );
  XOR U615 ( .A(n618), .B(n219), .Z(n621) );
  XNOR U616 ( .A(p_input[37]), .B(n622), .Z(n219) );
  AND U617 ( .A(n91), .B(n623), .Z(n622) );
  XOR U618 ( .A(p_input[53]), .B(p_input[37]), .Z(n623) );
  XNOR U619 ( .A(n216), .B(n618), .Z(n620) );
  XOR U620 ( .A(n624), .B(n625), .Z(n216) );
  AND U621 ( .A(n88), .B(n626), .Z(n625) );
  XOR U622 ( .A(p_input[5]), .B(p_input[21]), .Z(n626) );
  XOR U623 ( .A(n627), .B(n628), .Z(n618) );
  AND U624 ( .A(n629), .B(n630), .Z(n628) );
  XOR U625 ( .A(n627), .B(n231), .Z(n630) );
  XNOR U626 ( .A(p_input[36]), .B(n631), .Z(n231) );
  AND U627 ( .A(n91), .B(n632), .Z(n631) );
  XOR U628 ( .A(p_input[52]), .B(p_input[36]), .Z(n632) );
  XNOR U629 ( .A(n228), .B(n627), .Z(n629) );
  XOR U630 ( .A(n633), .B(n634), .Z(n228) );
  AND U631 ( .A(n88), .B(n635), .Z(n634) );
  XOR U632 ( .A(p_input[4]), .B(p_input[20]), .Z(n635) );
  XOR U633 ( .A(n636), .B(n637), .Z(n627) );
  AND U634 ( .A(n638), .B(n639), .Z(n637) );
  XOR U635 ( .A(n636), .B(n243), .Z(n639) );
  XNOR U636 ( .A(p_input[35]), .B(n640), .Z(n243) );
  AND U637 ( .A(n91), .B(n641), .Z(n640) );
  XOR U638 ( .A(p_input[51]), .B(p_input[35]), .Z(n641) );
  XNOR U639 ( .A(n240), .B(n636), .Z(n638) );
  XOR U640 ( .A(n642), .B(n643), .Z(n240) );
  AND U641 ( .A(n88), .B(n644), .Z(n643) );
  XOR U642 ( .A(p_input[3]), .B(p_input[19]), .Z(n644) );
  XOR U643 ( .A(n645), .B(n646), .Z(n636) );
  AND U644 ( .A(n647), .B(n648), .Z(n646) );
  XOR U645 ( .A(n645), .B(n255), .Z(n648) );
  XNOR U646 ( .A(p_input[34]), .B(n649), .Z(n255) );
  AND U647 ( .A(n91), .B(n650), .Z(n649) );
  XOR U648 ( .A(p_input[50]), .B(p_input[34]), .Z(n650) );
  XNOR U649 ( .A(n252), .B(n645), .Z(n647) );
  XOR U650 ( .A(n651), .B(n652), .Z(n252) );
  AND U651 ( .A(n88), .B(n653), .Z(n652) );
  XOR U652 ( .A(p_input[2]), .B(p_input[18]), .Z(n653) );
  XOR U653 ( .A(n654), .B(n655), .Z(n645) );
  AND U654 ( .A(n656), .B(n657), .Z(n655) );
  XNOR U655 ( .A(n658), .B(n267), .Z(n657) );
  XNOR U656 ( .A(p_input[33]), .B(n659), .Z(n267) );
  AND U657 ( .A(n91), .B(n660), .Z(n659) );
  XNOR U658 ( .A(p_input[49]), .B(n661), .Z(n660) );
  IV U659 ( .A(p_input[33]), .Z(n661) );
  XNOR U660 ( .A(n264), .B(n654), .Z(n656) );
  XNOR U661 ( .A(p_input[1]), .B(n662), .Z(n264) );
  AND U662 ( .A(n88), .B(n663), .Z(n662) );
  XOR U663 ( .A(p_input[1]), .B(p_input[17]), .Z(n663) );
  IV U664 ( .A(n658), .Z(n654) );
  AND U665 ( .A(n529), .B(n532), .Z(n658) );
  XOR U666 ( .A(p_input[32]), .B(n664), .Z(n532) );
  AND U667 ( .A(n91), .B(n665), .Z(n664) );
  XOR U668 ( .A(p_input[48]), .B(p_input[32]), .Z(n665) );
  XOR U669 ( .A(n666), .B(n667), .Z(n91) );
  AND U670 ( .A(n668), .B(n669), .Z(n667) );
  XNOR U671 ( .A(p_input[63]), .B(n666), .Z(n669) );
  XOR U672 ( .A(n666), .B(p_input[47]), .Z(n668) );
  XOR U673 ( .A(n670), .B(n671), .Z(n666) );
  AND U674 ( .A(n672), .B(n673), .Z(n671) );
  XNOR U675 ( .A(p_input[62]), .B(n670), .Z(n673) );
  XOR U676 ( .A(n670), .B(p_input[46]), .Z(n672) );
  XOR U677 ( .A(n674), .B(n675), .Z(n670) );
  AND U678 ( .A(n676), .B(n677), .Z(n675) );
  XNOR U679 ( .A(p_input[61]), .B(n674), .Z(n677) );
  XOR U680 ( .A(n674), .B(p_input[45]), .Z(n676) );
  XOR U681 ( .A(n678), .B(n679), .Z(n674) );
  AND U682 ( .A(n680), .B(n681), .Z(n679) );
  XNOR U683 ( .A(p_input[60]), .B(n678), .Z(n681) );
  XOR U684 ( .A(n678), .B(p_input[44]), .Z(n680) );
  XOR U685 ( .A(n682), .B(n683), .Z(n678) );
  AND U686 ( .A(n684), .B(n685), .Z(n683) );
  XNOR U687 ( .A(p_input[59]), .B(n682), .Z(n685) );
  XOR U688 ( .A(n682), .B(p_input[43]), .Z(n684) );
  XOR U689 ( .A(n686), .B(n687), .Z(n682) );
  AND U690 ( .A(n688), .B(n689), .Z(n687) );
  XNOR U691 ( .A(p_input[58]), .B(n686), .Z(n689) );
  XOR U692 ( .A(n686), .B(p_input[42]), .Z(n688) );
  XOR U693 ( .A(n690), .B(n691), .Z(n686) );
  AND U694 ( .A(n692), .B(n693), .Z(n691) );
  XNOR U695 ( .A(p_input[57]), .B(n690), .Z(n693) );
  XOR U696 ( .A(n690), .B(p_input[41]), .Z(n692) );
  XOR U697 ( .A(n694), .B(n695), .Z(n690) );
  AND U698 ( .A(n696), .B(n697), .Z(n695) );
  XNOR U699 ( .A(p_input[56]), .B(n694), .Z(n697) );
  XOR U700 ( .A(n694), .B(p_input[40]), .Z(n696) );
  XOR U701 ( .A(n698), .B(n699), .Z(n694) );
  AND U702 ( .A(n700), .B(n701), .Z(n699) );
  XNOR U703 ( .A(p_input[55]), .B(n698), .Z(n701) );
  XOR U704 ( .A(n698), .B(p_input[39]), .Z(n700) );
  XOR U705 ( .A(n702), .B(n703), .Z(n698) );
  AND U706 ( .A(n704), .B(n705), .Z(n703) );
  XNOR U707 ( .A(p_input[54]), .B(n702), .Z(n705) );
  XOR U708 ( .A(n702), .B(p_input[38]), .Z(n704) );
  XOR U709 ( .A(n706), .B(n707), .Z(n702) );
  AND U710 ( .A(n708), .B(n709), .Z(n707) );
  XNOR U711 ( .A(p_input[53]), .B(n706), .Z(n709) );
  XOR U712 ( .A(n706), .B(p_input[37]), .Z(n708) );
  XOR U713 ( .A(n710), .B(n711), .Z(n706) );
  AND U714 ( .A(n712), .B(n713), .Z(n711) );
  XNOR U715 ( .A(p_input[52]), .B(n710), .Z(n713) );
  XOR U716 ( .A(n710), .B(p_input[36]), .Z(n712) );
  XOR U717 ( .A(n714), .B(n715), .Z(n710) );
  AND U718 ( .A(n716), .B(n717), .Z(n715) );
  XNOR U719 ( .A(p_input[51]), .B(n714), .Z(n717) );
  XOR U720 ( .A(n714), .B(p_input[35]), .Z(n716) );
  XOR U721 ( .A(n718), .B(n719), .Z(n714) );
  AND U722 ( .A(n720), .B(n721), .Z(n719) );
  XNOR U723 ( .A(p_input[50]), .B(n718), .Z(n721) );
  XOR U724 ( .A(n718), .B(p_input[34]), .Z(n720) );
  XNOR U725 ( .A(n722), .B(n723), .Z(n718) );
  AND U726 ( .A(n724), .B(n725), .Z(n723) );
  XOR U727 ( .A(p_input[49]), .B(n722), .Z(n725) );
  XNOR U728 ( .A(p_input[33]), .B(n722), .Z(n724) );
  AND U729 ( .A(p_input[48]), .B(n726), .Z(n722) );
  IV U730 ( .A(p_input[32]), .Z(n726) );
  XNOR U731 ( .A(p_input[0]), .B(n727), .Z(n529) );
  AND U732 ( .A(n88), .B(n728), .Z(n727) );
  XOR U733 ( .A(p_input[16]), .B(p_input[0]), .Z(n728) );
  XOR U734 ( .A(n729), .B(n730), .Z(n88) );
  AND U735 ( .A(n731), .B(n732), .Z(n730) );
  XNOR U736 ( .A(p_input[31]), .B(n729), .Z(n732) );
  XOR U737 ( .A(n729), .B(p_input[15]), .Z(n731) );
  XOR U738 ( .A(n733), .B(n734), .Z(n729) );
  AND U739 ( .A(n735), .B(n736), .Z(n734) );
  XNOR U740 ( .A(p_input[30]), .B(n733), .Z(n736) );
  XNOR U741 ( .A(n733), .B(n543), .Z(n735) );
  IV U742 ( .A(p_input[14]), .Z(n543) );
  XOR U743 ( .A(n737), .B(n738), .Z(n733) );
  AND U744 ( .A(n739), .B(n740), .Z(n738) );
  XNOR U745 ( .A(p_input[29]), .B(n737), .Z(n740) );
  XNOR U746 ( .A(n737), .B(n552), .Z(n739) );
  IV U747 ( .A(p_input[13]), .Z(n552) );
  XOR U748 ( .A(n741), .B(n742), .Z(n737) );
  AND U749 ( .A(n743), .B(n744), .Z(n742) );
  XNOR U750 ( .A(p_input[28]), .B(n741), .Z(n744) );
  XNOR U751 ( .A(n741), .B(n561), .Z(n743) );
  IV U752 ( .A(p_input[12]), .Z(n561) );
  XOR U753 ( .A(n745), .B(n746), .Z(n741) );
  AND U754 ( .A(n747), .B(n748), .Z(n746) );
  XNOR U755 ( .A(p_input[27]), .B(n745), .Z(n748) );
  XNOR U756 ( .A(n745), .B(n570), .Z(n747) );
  IV U757 ( .A(p_input[11]), .Z(n570) );
  XOR U758 ( .A(n749), .B(n750), .Z(n745) );
  AND U759 ( .A(n751), .B(n752), .Z(n750) );
  XNOR U760 ( .A(p_input[26]), .B(n749), .Z(n752) );
  XNOR U761 ( .A(n749), .B(n579), .Z(n751) );
  IV U762 ( .A(p_input[10]), .Z(n579) );
  XOR U763 ( .A(n753), .B(n754), .Z(n749) );
  AND U764 ( .A(n755), .B(n756), .Z(n754) );
  XNOR U765 ( .A(p_input[25]), .B(n753), .Z(n756) );
  XNOR U766 ( .A(n753), .B(n588), .Z(n755) );
  IV U767 ( .A(p_input[9]), .Z(n588) );
  XOR U768 ( .A(n757), .B(n758), .Z(n753) );
  AND U769 ( .A(n759), .B(n760), .Z(n758) );
  XNOR U770 ( .A(p_input[24]), .B(n757), .Z(n760) );
  XNOR U771 ( .A(n757), .B(n597), .Z(n759) );
  IV U772 ( .A(p_input[8]), .Z(n597) );
  XOR U773 ( .A(n761), .B(n762), .Z(n757) );
  AND U774 ( .A(n763), .B(n764), .Z(n762) );
  XNOR U775 ( .A(p_input[23]), .B(n761), .Z(n764) );
  XNOR U776 ( .A(n761), .B(n606), .Z(n763) );
  IV U777 ( .A(p_input[7]), .Z(n606) );
  XOR U778 ( .A(n765), .B(n766), .Z(n761) );
  AND U779 ( .A(n767), .B(n768), .Z(n766) );
  XNOR U780 ( .A(p_input[22]), .B(n765), .Z(n768) );
  XNOR U781 ( .A(n765), .B(n615), .Z(n767) );
  IV U782 ( .A(p_input[6]), .Z(n615) );
  XOR U783 ( .A(n769), .B(n770), .Z(n765) );
  AND U784 ( .A(n771), .B(n772), .Z(n770) );
  XNOR U785 ( .A(p_input[21]), .B(n769), .Z(n772) );
  XNOR U786 ( .A(n769), .B(n624), .Z(n771) );
  IV U787 ( .A(p_input[5]), .Z(n624) );
  XOR U788 ( .A(n773), .B(n774), .Z(n769) );
  AND U789 ( .A(n775), .B(n776), .Z(n774) );
  XNOR U790 ( .A(p_input[20]), .B(n773), .Z(n776) );
  XNOR U791 ( .A(n773), .B(n633), .Z(n775) );
  IV U792 ( .A(p_input[4]), .Z(n633) );
  XOR U793 ( .A(n777), .B(n778), .Z(n773) );
  AND U794 ( .A(n779), .B(n780), .Z(n778) );
  XNOR U795 ( .A(p_input[19]), .B(n777), .Z(n780) );
  XNOR U796 ( .A(n777), .B(n642), .Z(n779) );
  IV U797 ( .A(p_input[3]), .Z(n642) );
  XOR U798 ( .A(n781), .B(n782), .Z(n777) );
  AND U799 ( .A(n783), .B(n784), .Z(n782) );
  XNOR U800 ( .A(p_input[18]), .B(n781), .Z(n784) );
  XNOR U801 ( .A(n781), .B(n651), .Z(n783) );
  IV U802 ( .A(p_input[2]), .Z(n651) );
  XNOR U803 ( .A(n785), .B(n786), .Z(n781) );
  AND U804 ( .A(n787), .B(n788), .Z(n786) );
  XOR U805 ( .A(p_input[17]), .B(n785), .Z(n788) );
  XNOR U806 ( .A(p_input[1]), .B(n785), .Z(n787) );
  AND U807 ( .A(p_input[16]), .B(n789), .Z(n785) );
  IV U808 ( .A(p_input[0]), .Z(n789) );
endmodule

