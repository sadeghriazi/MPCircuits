
module voting_N2_M4 ( p_input, o );
  input [31:0] p_input;
  output [1:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513;

  XOR U2 ( .A(n1), .B(n2), .Z(o[0]) );
  AND U3 ( .A(o[1]), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(n5), .Z(n3) );
  IV U5 ( .A(n1), .Z(n5) );
  NOR U6 ( .A(n6), .B(n7), .Z(o[1]) );
  XOR U7 ( .A(n8), .B(n9), .Z(n7) );
  AND U8 ( .A(n10), .B(n11), .Z(n8) );
  XOR U9 ( .A(n12), .B(n9), .Z(n11) );
  XNOR U10 ( .A(n9), .B(n13), .Z(n10) );
  AND U11 ( .A(n14), .B(n15), .Z(n13) );
  XOR U12 ( .A(n16), .B(n17), .Z(n9) );
  AND U13 ( .A(n18), .B(n19), .Z(n17) );
  XOR U14 ( .A(n16), .B(n20), .Z(n19) );
  XNOR U15 ( .A(n21), .B(n22), .Z(n20) );
  AND U16 ( .A(n4), .B(n23), .Z(n21) );
  XOR U17 ( .A(n24), .B(n22), .Z(n23) );
  XOR U18 ( .A(n25), .B(n16), .Z(n18) );
  XOR U19 ( .A(n26), .B(n27), .Z(n25) );
  AND U20 ( .A(n1), .B(n28), .Z(n27) );
  XOR U21 ( .A(n29), .B(n26), .Z(n28) );
  XOR U22 ( .A(n30), .B(n31), .Z(n16) );
  AND U23 ( .A(n32), .B(n33), .Z(n31) );
  XNOR U24 ( .A(n34), .B(n35), .Z(n33) );
  XOR U25 ( .A(n30), .B(n36), .Z(n35) );
  AND U26 ( .A(n4), .B(n37), .Z(n36) );
  XOR U27 ( .A(n38), .B(n34), .Z(n37) );
  XOR U28 ( .A(n39), .B(n40), .Z(n32) );
  XOR U29 ( .A(n30), .B(n41), .Z(n40) );
  AND U30 ( .A(n1), .B(n42), .Z(n41) );
  XOR U31 ( .A(n43), .B(n39), .Z(n42) );
  AND U32 ( .A(n44), .B(n45), .Z(n30) );
  XOR U33 ( .A(n46), .B(n47), .Z(n45) );
  AND U34 ( .A(n4), .B(n48), .Z(n46) );
  XNOR U35 ( .A(n49), .B(n47), .Z(n48) );
  XNOR U36 ( .A(n50), .B(n51), .Z(n4) );
  AND U37 ( .A(n52), .B(n53), .Z(n51) );
  XOR U38 ( .A(n54), .B(n50), .Z(n53) );
  XNOR U39 ( .A(n50), .B(n55), .Z(n52) );
  XOR U40 ( .A(n56), .B(n57), .Z(n50) );
  AND U41 ( .A(n58), .B(n59), .Z(n57) );
  XNOR U42 ( .A(n24), .B(n56), .Z(n59) );
  XOR U43 ( .A(n56), .B(n22), .Z(n58) );
  XOR U44 ( .A(n60), .B(n61), .Z(n56) );
  AND U45 ( .A(n62), .B(n63), .Z(n61) );
  XNOR U46 ( .A(n38), .B(n60), .Z(n63) );
  XOR U47 ( .A(n60), .B(n34), .Z(n62) );
  NOR U48 ( .A(n47), .B(n49), .Z(n60) );
  XNOR U49 ( .A(n64), .B(n65), .Z(n49) );
  XOR U50 ( .A(n66), .B(n67), .Z(n47) );
  XNOR U51 ( .A(n68), .B(n69), .Z(n44) );
  AND U52 ( .A(n1), .B(n70), .Z(n69) );
  XNOR U53 ( .A(n68), .B(n71), .Z(n70) );
  NOR U54 ( .A(n72), .B(n73), .Z(n6) );
  AND U55 ( .A(n74), .B(n75), .Z(n73) );
  IV U56 ( .A(n12), .Z(n72) );
  AND U57 ( .A(n55), .B(n54), .Z(n12) );
  XNOR U58 ( .A(n76), .B(n77), .Z(n54) );
  AND U59 ( .A(n24), .B(n78), .Z(n77) );
  XOR U60 ( .A(n79), .B(n78), .Z(n24) );
  AND U61 ( .A(n38), .B(n80), .Z(n78) );
  XOR U62 ( .A(n81), .B(n80), .Z(n38) );
  AND U63 ( .A(n65), .B(n64), .Z(n80) );
  XOR U64 ( .A(n82), .B(n83), .Z(n64) );
  AND U65 ( .A(p_input[31]), .B(p_input[30]), .Z(n65) );
  XNOR U66 ( .A(n84), .B(n85), .Z(n76) );
  AND U67 ( .A(n86), .B(n87), .Z(n85) );
  NOR U68 ( .A(n88), .B(n89), .Z(n87) );
  NOR U69 ( .A(n90), .B(n91), .Z(n86) );
  AND U70 ( .A(n79), .B(n92), .Z(n91) );
  XNOR U71 ( .A(n93), .B(n92), .Z(n79) );
  AND U72 ( .A(n81), .B(n94), .Z(n92) );
  XOR U73 ( .A(n95), .B(n94), .Z(n81) );
  AND U74 ( .A(n83), .B(n82), .Z(n94) );
  XOR U75 ( .A(n96), .B(n97), .Z(n82) );
  AND U76 ( .A(p_input[29]), .B(p_input[28]), .Z(n83) );
  AND U77 ( .A(n98), .B(n99), .Z(n84) );
  NOR U78 ( .A(n100), .B(n101), .Z(n99) );
  AND U79 ( .A(n90), .B(n102), .Z(n101) );
  AND U80 ( .A(n88), .B(n93), .Z(n100) );
  XOR U81 ( .A(n102), .B(n88), .Z(n93) );
  XOR U82 ( .A(n103), .B(n90), .Z(n102) );
  AND U83 ( .A(n104), .B(n105), .Z(n90) );
  AND U84 ( .A(n95), .B(n106), .Z(n88) );
  XOR U85 ( .A(n104), .B(n106), .Z(n95) );
  AND U86 ( .A(n97), .B(n96), .Z(n106) );
  XOR U87 ( .A(n107), .B(n108), .Z(n96) );
  AND U88 ( .A(p_input[27]), .B(p_input[26]), .Z(n97) );
  XOR U89 ( .A(n109), .B(n105), .Z(n104) );
  AND U90 ( .A(n108), .B(n107), .Z(n105) );
  XOR U91 ( .A(n110), .B(n111), .Z(n107) );
  AND U92 ( .A(p_input[25]), .B(p_input[24]), .Z(n108) );
  NOR U93 ( .A(n112), .B(n113), .Z(n98) );
  AND U94 ( .A(n114), .B(n115), .Z(n113) );
  AND U95 ( .A(n116), .B(n117), .Z(n115) );
  IV U96 ( .A(n118), .Z(n117) );
  NOR U97 ( .A(n119), .B(n120), .Z(n116) );
  NOR U98 ( .A(n121), .B(n122), .Z(n114) );
  AND U99 ( .A(n89), .B(n103), .Z(n112) );
  XNOR U100 ( .A(n123), .B(n124), .Z(n103) );
  XOR U101 ( .A(n121), .B(n125), .Z(n124) );
  XOR U102 ( .A(n119), .B(n118), .Z(n125) );
  AND U103 ( .A(n126), .B(n127), .Z(n118) );
  AND U104 ( .A(n128), .B(n129), .Z(n119) );
  AND U105 ( .A(n130), .B(n131), .Z(n121) );
  XNOR U106 ( .A(n132), .B(n120), .Z(n123) );
  XOR U107 ( .A(n133), .B(n134), .Z(n120) );
  XOR U108 ( .A(n135), .B(n136), .Z(n134) );
  AND U109 ( .A(n137), .B(n138), .Z(n136) );
  XNOR U110 ( .A(n139), .B(n140), .Z(n133) );
  NOR U111 ( .A(n141), .B(n142), .Z(n140) );
  AND U112 ( .A(n143), .B(n144), .Z(n142) );
  IV U113 ( .A(n145), .Z(n141) );
  NOR U114 ( .A(n135), .B(n146), .Z(n145) );
  AND U115 ( .A(n147), .B(n148), .Z(n146) );
  NOR U116 ( .A(n137), .B(n147), .Z(n139) );
  XNOR U117 ( .A(n122), .B(n89), .Z(n132) );
  AND U118 ( .A(n149), .B(n150), .Z(n122) );
  AND U119 ( .A(n109), .B(n151), .Z(n89) );
  XOR U120 ( .A(n149), .B(n151), .Z(n109) );
  AND U121 ( .A(n111), .B(n110), .Z(n151) );
  XOR U122 ( .A(n152), .B(n153), .Z(n110) );
  AND U123 ( .A(p_input[23]), .B(p_input[22]), .Z(n111) );
  XOR U124 ( .A(n130), .B(n150), .Z(n149) );
  AND U125 ( .A(n153), .B(n152), .Z(n150) );
  XOR U126 ( .A(n154), .B(n155), .Z(n152) );
  AND U127 ( .A(p_input[21]), .B(p_input[20]), .Z(n153) );
  XOR U128 ( .A(n126), .B(n131), .Z(n130) );
  AND U129 ( .A(n155), .B(n154), .Z(n131) );
  XOR U130 ( .A(n156), .B(n157), .Z(n154) );
  AND U131 ( .A(p_input[19]), .B(p_input[18]), .Z(n155) );
  XOR U132 ( .A(n128), .B(n127), .Z(n126) );
  AND U133 ( .A(n157), .B(n156), .Z(n127) );
  XOR U134 ( .A(n158), .B(n159), .Z(n156) );
  AND U135 ( .A(p_input[17]), .B(p_input[16]), .Z(n157) );
  XNOR U136 ( .A(n138), .B(n129), .Z(n128) );
  AND U137 ( .A(n159), .B(n158), .Z(n129) );
  XOR U138 ( .A(n160), .B(n161), .Z(n158) );
  AND U139 ( .A(p_input[15]), .B(p_input[14]), .Z(n159) );
  XOR U140 ( .A(n148), .B(n137), .Z(n138) );
  AND U141 ( .A(n161), .B(n160), .Z(n137) );
  XOR U142 ( .A(n162), .B(n163), .Z(n160) );
  AND U143 ( .A(p_input[13]), .B(p_input[12]), .Z(n161) );
  XNOR U144 ( .A(n164), .B(n143), .Z(n148) );
  XOR U145 ( .A(n144), .B(n165), .Z(n143) );
  AND U146 ( .A(n166), .B(n167), .Z(n165) );
  XOR U147 ( .A(n168), .B(n169), .Z(n144) );
  NOR U148 ( .A(n170), .B(n171), .Z(n169) );
  AND U149 ( .A(n172), .B(n173), .Z(n171) );
  AND U150 ( .A(n174), .B(n175), .Z(n170) );
  XNOR U151 ( .A(n172), .B(n173), .Z(n168) );
  XNOR U152 ( .A(n135), .B(n147), .Z(n164) );
  AND U153 ( .A(n163), .B(n162), .Z(n147) );
  XOR U154 ( .A(n176), .B(n177), .Z(n162) );
  AND U155 ( .A(p_input[11]), .B(p_input[10]), .Z(n163) );
  AND U156 ( .A(n177), .B(n176), .Z(n135) );
  XOR U157 ( .A(n167), .B(n166), .Z(n176) );
  AND U158 ( .A(p_input[7]), .B(p_input[6]), .Z(n166) );
  XOR U159 ( .A(n174), .B(n175), .Z(n167) );
  XOR U160 ( .A(n172), .B(n173), .Z(n175) );
  AND U161 ( .A(p_input[3]), .B(p_input[2]), .Z(n173) );
  AND U162 ( .A(p_input[1]), .B(p_input[0]), .Z(n172) );
  AND U163 ( .A(p_input[5]), .B(p_input[4]), .Z(n174) );
  AND U164 ( .A(p_input[9]), .B(p_input[8]), .Z(n177) );
  XNOR U165 ( .A(n178), .B(n179), .Z(n55) );
  XOR U166 ( .A(n180), .B(n181), .Z(n179) );
  XOR U167 ( .A(n182), .B(n183), .Z(n181) );
  NOR U168 ( .A(n184), .B(n185), .Z(n183) );
  NOR U169 ( .A(n186), .B(n187), .Z(n182) );
  AND U170 ( .A(n188), .B(n189), .Z(n187) );
  IV U171 ( .A(n190), .Z(n186) );
  NOR U172 ( .A(n191), .B(n192), .Z(n190) );
  AND U173 ( .A(n184), .B(n193), .Z(n192) );
  AND U174 ( .A(n185), .B(n194), .Z(n191) );
  AND U175 ( .A(n195), .B(n196), .Z(n180) );
  AND U176 ( .A(n197), .B(n198), .Z(n196) );
  IV U177 ( .A(n199), .Z(n198) );
  NOR U178 ( .A(n200), .B(n201), .Z(n197) );
  NOR U179 ( .A(n202), .B(n203), .Z(n195) );
  XNOR U180 ( .A(n204), .B(n205), .Z(n178) );
  AND U181 ( .A(n22), .B(n206), .Z(n205) );
  XOR U182 ( .A(n207), .B(n206), .Z(n22) );
  AND U183 ( .A(n34), .B(n208), .Z(n206) );
  XOR U184 ( .A(n209), .B(n208), .Z(n34) );
  AND U185 ( .A(n67), .B(n66), .Z(n208) );
  XOR U186 ( .A(n210), .B(n211), .Z(n66) );
  AND U187 ( .A(p_input[31]), .B(n212), .Z(n67) );
  AND U188 ( .A(n207), .B(n213), .Z(n204) );
  XNOR U189 ( .A(n194), .B(n213), .Z(n207) );
  AND U190 ( .A(n209), .B(n214), .Z(n213) );
  XOR U191 ( .A(n215), .B(n214), .Z(n209) );
  AND U192 ( .A(n211), .B(n210), .Z(n214) );
  XOR U193 ( .A(n216), .B(n217), .Z(n210) );
  AND U194 ( .A(p_input[29]), .B(n218), .Z(n211) );
  XOR U195 ( .A(n193), .B(n185), .Z(n194) );
  AND U196 ( .A(n215), .B(n219), .Z(n185) );
  XOR U197 ( .A(n220), .B(n219), .Z(n215) );
  AND U198 ( .A(n217), .B(n216), .Z(n219) );
  XOR U199 ( .A(n221), .B(n222), .Z(n216) );
  AND U200 ( .A(p_input[27]), .B(n223), .Z(n217) );
  XNOR U201 ( .A(n188), .B(n184), .Z(n193) );
  AND U202 ( .A(n220), .B(n224), .Z(n184) );
  XOR U203 ( .A(n225), .B(n224), .Z(n220) );
  AND U204 ( .A(n222), .B(n221), .Z(n224) );
  XOR U205 ( .A(n226), .B(n227), .Z(n221) );
  AND U206 ( .A(p_input[25]), .B(n228), .Z(n222) );
  XOR U207 ( .A(n229), .B(n230), .Z(n188) );
  XOR U208 ( .A(n202), .B(n231), .Z(n230) );
  XOR U209 ( .A(n200), .B(n199), .Z(n231) );
  AND U210 ( .A(n232), .B(n233), .Z(n199) );
  AND U211 ( .A(n234), .B(n235), .Z(n200) );
  AND U212 ( .A(n236), .B(n237), .Z(n202) );
  XNOR U213 ( .A(n238), .B(n201), .Z(n229) );
  XOR U214 ( .A(n239), .B(n240), .Z(n201) );
  XOR U215 ( .A(n241), .B(n242), .Z(n240) );
  AND U216 ( .A(n243), .B(n244), .Z(n242) );
  XNOR U217 ( .A(n245), .B(n246), .Z(n239) );
  NOR U218 ( .A(n247), .B(n248), .Z(n246) );
  AND U219 ( .A(n249), .B(n250), .Z(n248) );
  IV U220 ( .A(n251), .Z(n247) );
  NOR U221 ( .A(n241), .B(n252), .Z(n251) );
  AND U222 ( .A(n253), .B(n254), .Z(n252) );
  NOR U223 ( .A(n243), .B(n253), .Z(n245) );
  XNOR U224 ( .A(n203), .B(n189), .Z(n238) );
  AND U225 ( .A(n225), .B(n255), .Z(n189) );
  XOR U226 ( .A(n256), .B(n255), .Z(n225) );
  AND U227 ( .A(n227), .B(n226), .Z(n255) );
  XOR U228 ( .A(n257), .B(n258), .Z(n226) );
  AND U229 ( .A(p_input[23]), .B(n259), .Z(n227) );
  AND U230 ( .A(n256), .B(n260), .Z(n203) );
  XOR U231 ( .A(n236), .B(n260), .Z(n256) );
  AND U232 ( .A(n258), .B(n257), .Z(n260) );
  XOR U233 ( .A(n261), .B(n262), .Z(n257) );
  AND U234 ( .A(p_input[21]), .B(n263), .Z(n258) );
  XOR U235 ( .A(n232), .B(n237), .Z(n236) );
  AND U236 ( .A(n262), .B(n261), .Z(n237) );
  XOR U237 ( .A(n264), .B(n265), .Z(n261) );
  AND U238 ( .A(p_input[19]), .B(n266), .Z(n262) );
  XOR U239 ( .A(n234), .B(n233), .Z(n232) );
  AND U240 ( .A(n265), .B(n264), .Z(n233) );
  XOR U241 ( .A(n267), .B(n268), .Z(n264) );
  AND U242 ( .A(p_input[17]), .B(n269), .Z(n265) );
  XNOR U243 ( .A(n244), .B(n235), .Z(n234) );
  AND U244 ( .A(n268), .B(n267), .Z(n235) );
  XOR U245 ( .A(n270), .B(n271), .Z(n267) );
  AND U246 ( .A(p_input[15]), .B(n272), .Z(n268) );
  XOR U247 ( .A(n254), .B(n243), .Z(n244) );
  AND U248 ( .A(n271), .B(n270), .Z(n243) );
  XOR U249 ( .A(n273), .B(n274), .Z(n270) );
  AND U250 ( .A(p_input[13]), .B(n275), .Z(n271) );
  XNOR U251 ( .A(n276), .B(n249), .Z(n254) );
  XOR U252 ( .A(n250), .B(n277), .Z(n249) );
  AND U253 ( .A(n278), .B(n279), .Z(n277) );
  XOR U254 ( .A(n280), .B(n281), .Z(n250) );
  NOR U255 ( .A(n282), .B(n283), .Z(n281) );
  AND U256 ( .A(n284), .B(n285), .Z(n283) );
  AND U257 ( .A(n286), .B(n287), .Z(n282) );
  XNOR U258 ( .A(n284), .B(n285), .Z(n280) );
  XNOR U259 ( .A(n241), .B(n253), .Z(n276) );
  AND U260 ( .A(n274), .B(n273), .Z(n253) );
  XOR U261 ( .A(n288), .B(n289), .Z(n273) );
  AND U262 ( .A(p_input[11]), .B(n290), .Z(n274) );
  AND U263 ( .A(n289), .B(n288), .Z(n241) );
  XOR U264 ( .A(n279), .B(n278), .Z(n288) );
  AND U265 ( .A(p_input[7]), .B(n291), .Z(n278) );
  XOR U266 ( .A(n286), .B(n287), .Z(n279) );
  XOR U267 ( .A(n284), .B(n285), .Z(n287) );
  AND U268 ( .A(p_input[3]), .B(n292), .Z(n285) );
  AND U269 ( .A(p_input[1]), .B(n293), .Z(n284) );
  AND U270 ( .A(p_input[5]), .B(n294), .Z(n286) );
  AND U271 ( .A(p_input[9]), .B(n295), .Z(n289) );
  XNOR U272 ( .A(n296), .B(n297), .Z(n1) );
  AND U273 ( .A(n298), .B(n299), .Z(n297) );
  XOR U274 ( .A(n296), .B(n15), .Z(n299) );
  XOR U275 ( .A(n75), .B(n300), .Z(n15) );
  AND U276 ( .A(n29), .B(n301), .Z(n300) );
  XOR U277 ( .A(n302), .B(n303), .Z(n75) );
  AND U278 ( .A(n304), .B(n305), .Z(n303) );
  NOR U279 ( .A(n306), .B(n307), .Z(n305) );
  NOR U280 ( .A(n308), .B(n309), .Z(n304) );
  AND U281 ( .A(n310), .B(n311), .Z(n309) );
  AND U282 ( .A(n312), .B(n313), .Z(n302) );
  NOR U283 ( .A(n314), .B(n315), .Z(n313) );
  AND U284 ( .A(n308), .B(n316), .Z(n315) );
  AND U285 ( .A(n306), .B(n317), .Z(n314) );
  NOR U286 ( .A(n318), .B(n319), .Z(n312) );
  AND U287 ( .A(n320), .B(n321), .Z(n319) );
  AND U288 ( .A(n322), .B(n323), .Z(n321) );
  IV U289 ( .A(n324), .Z(n323) );
  NOR U290 ( .A(n325), .B(n326), .Z(n322) );
  NOR U291 ( .A(n327), .B(n328), .Z(n320) );
  AND U292 ( .A(n307), .B(n329), .Z(n318) );
  XNOR U293 ( .A(n14), .B(n296), .Z(n298) );
  XOR U294 ( .A(n74), .B(n330), .Z(n14) );
  AND U295 ( .A(n26), .B(n331), .Z(n330) );
  XNOR U296 ( .A(n332), .B(n333), .Z(n74) );
  XOR U297 ( .A(n334), .B(n335), .Z(n333) );
  NOR U298 ( .A(n336), .B(n337), .Z(n335) );
  NOR U299 ( .A(n338), .B(n339), .Z(n334) );
  AND U300 ( .A(n340), .B(n341), .Z(n339) );
  IV U301 ( .A(n342), .Z(n338) );
  NOR U302 ( .A(n343), .B(n344), .Z(n342) );
  AND U303 ( .A(n336), .B(n345), .Z(n344) );
  AND U304 ( .A(n337), .B(n346), .Z(n343) );
  XNOR U305 ( .A(n347), .B(n348), .Z(n332) );
  AND U306 ( .A(n349), .B(n350), .Z(n348) );
  AND U307 ( .A(n351), .B(n352), .Z(n347) );
  NOR U308 ( .A(n353), .B(n354), .Z(n352) );
  IV U309 ( .A(n355), .Z(n353) );
  NOR U310 ( .A(n356), .B(n357), .Z(n355) );
  NOR U311 ( .A(n358), .B(n359), .Z(n351) );
  XOR U312 ( .A(n360), .B(n361), .Z(n296) );
  AND U313 ( .A(n362), .B(n363), .Z(n361) );
  XNOR U314 ( .A(n360), .B(n29), .Z(n363) );
  XOR U315 ( .A(n310), .B(n301), .Z(n29) );
  AND U316 ( .A(n43), .B(n364), .Z(n301) );
  XNOR U317 ( .A(n317), .B(n311), .Z(n310) );
  AND U318 ( .A(n365), .B(n366), .Z(n311) );
  XOR U319 ( .A(n316), .B(n306), .Z(n317) );
  AND U320 ( .A(n367), .B(n368), .Z(n306) );
  XOR U321 ( .A(n329), .B(n308), .Z(n316) );
  AND U322 ( .A(n369), .B(n370), .Z(n308) );
  XNOR U323 ( .A(n371), .B(n372), .Z(n329) );
  XOR U324 ( .A(n327), .B(n373), .Z(n372) );
  XOR U325 ( .A(n325), .B(n324), .Z(n373) );
  AND U326 ( .A(n374), .B(n375), .Z(n324) );
  AND U327 ( .A(n376), .B(n377), .Z(n325) );
  AND U328 ( .A(n378), .B(n379), .Z(n327) );
  XNOR U329 ( .A(n380), .B(n326), .Z(n371) );
  XOR U330 ( .A(n381), .B(n382), .Z(n326) );
  XOR U331 ( .A(n383), .B(n384), .Z(n382) );
  AND U332 ( .A(n385), .B(n386), .Z(n384) );
  XNOR U333 ( .A(n387), .B(n388), .Z(n381) );
  NOR U334 ( .A(n389), .B(n390), .Z(n388) );
  AND U335 ( .A(n391), .B(n392), .Z(n390) );
  IV U336 ( .A(n393), .Z(n389) );
  NOR U337 ( .A(n383), .B(n394), .Z(n393) );
  AND U338 ( .A(n395), .B(n396), .Z(n394) );
  NOR U339 ( .A(n385), .B(n395), .Z(n387) );
  XNOR U340 ( .A(n328), .B(n307), .Z(n380) );
  AND U341 ( .A(n397), .B(n398), .Z(n307) );
  AND U342 ( .A(n399), .B(n400), .Z(n328) );
  XOR U343 ( .A(n26), .B(n360), .Z(n362) );
  XOR U344 ( .A(n349), .B(n331), .Z(n26) );
  AND U345 ( .A(n39), .B(n401), .Z(n331) );
  XNOR U346 ( .A(n346), .B(n350), .Z(n349) );
  AND U347 ( .A(n402), .B(n403), .Z(n350) );
  XOR U348 ( .A(n345), .B(n337), .Z(n346) );
  AND U349 ( .A(n404), .B(n405), .Z(n337) );
  XNOR U350 ( .A(n340), .B(n336), .Z(n345) );
  AND U351 ( .A(n406), .B(n407), .Z(n336) );
  XOR U352 ( .A(n408), .B(n409), .Z(n340) );
  XOR U353 ( .A(n358), .B(n410), .Z(n409) );
  XOR U354 ( .A(n356), .B(n354), .Z(n410) );
  AND U355 ( .A(n411), .B(n412), .Z(n354) );
  AND U356 ( .A(n413), .B(n414), .Z(n356) );
  AND U357 ( .A(n415), .B(n416), .Z(n358) );
  XNOR U358 ( .A(n417), .B(n357), .Z(n408) );
  XOR U359 ( .A(n418), .B(n419), .Z(n357) );
  XOR U360 ( .A(n420), .B(n421), .Z(n419) );
  AND U361 ( .A(n422), .B(n423), .Z(n421) );
  XNOR U362 ( .A(n424), .B(n425), .Z(n418) );
  NOR U363 ( .A(n426), .B(n427), .Z(n425) );
  AND U364 ( .A(n428), .B(n429), .Z(n427) );
  IV U365 ( .A(n430), .Z(n426) );
  NOR U366 ( .A(n420), .B(n431), .Z(n430) );
  AND U367 ( .A(n432), .B(n433), .Z(n431) );
  NOR U368 ( .A(n422), .B(n432), .Z(n424) );
  XNOR U369 ( .A(n359), .B(n341), .Z(n417) );
  AND U370 ( .A(n434), .B(n435), .Z(n341) );
  AND U371 ( .A(n436), .B(n437), .Z(n359) );
  XOR U372 ( .A(n438), .B(n439), .Z(n360) );
  AND U373 ( .A(n440), .B(n441), .Z(n439) );
  XNOR U374 ( .A(n43), .B(n438), .Z(n441) );
  XOR U375 ( .A(n365), .B(n364), .Z(n43) );
  AND U376 ( .A(n442), .B(n443), .Z(n364) );
  XOR U377 ( .A(n367), .B(n366), .Z(n365) );
  AND U378 ( .A(n444), .B(n445), .Z(n366) );
  XOR U379 ( .A(n369), .B(n368), .Z(n367) );
  AND U380 ( .A(n446), .B(n447), .Z(n368) );
  XOR U381 ( .A(n397), .B(n370), .Z(n369) );
  AND U382 ( .A(n448), .B(n449), .Z(n370) );
  XOR U383 ( .A(n399), .B(n398), .Z(n397) );
  AND U384 ( .A(n450), .B(n451), .Z(n398) );
  XOR U385 ( .A(n378), .B(n400), .Z(n399) );
  AND U386 ( .A(n452), .B(n453), .Z(n400) );
  XOR U387 ( .A(n374), .B(n379), .Z(n378) );
  AND U388 ( .A(n454), .B(n455), .Z(n379) );
  XOR U389 ( .A(n376), .B(n375), .Z(n374) );
  AND U390 ( .A(n456), .B(n457), .Z(n375) );
  XNOR U391 ( .A(n386), .B(n377), .Z(n376) );
  AND U392 ( .A(n458), .B(n459), .Z(n377) );
  XOR U393 ( .A(n396), .B(n385), .Z(n386) );
  AND U394 ( .A(n460), .B(n461), .Z(n385) );
  XNOR U395 ( .A(n462), .B(n391), .Z(n396) );
  XOR U396 ( .A(n392), .B(n463), .Z(n391) );
  AND U397 ( .A(n464), .B(n465), .Z(n463) );
  XOR U398 ( .A(n466), .B(n467), .Z(n392) );
  NOR U399 ( .A(n468), .B(n469), .Z(n467) );
  AND U400 ( .A(n470), .B(n471), .Z(n469) );
  AND U401 ( .A(n472), .B(n473), .Z(n468) );
  XNOR U402 ( .A(n470), .B(n471), .Z(n466) );
  XNOR U403 ( .A(n383), .B(n395), .Z(n462) );
  AND U404 ( .A(n474), .B(n475), .Z(n395) );
  AND U405 ( .A(n476), .B(n477), .Z(n383) );
  XOR U406 ( .A(n438), .B(n39), .Z(n440) );
  XOR U407 ( .A(n402), .B(n401), .Z(n39) );
  AND U408 ( .A(n478), .B(n479), .Z(n401) );
  XOR U409 ( .A(n404), .B(n403), .Z(n402) );
  AND U410 ( .A(n480), .B(n481), .Z(n403) );
  XOR U411 ( .A(n406), .B(n405), .Z(n404) );
  AND U412 ( .A(n482), .B(n483), .Z(n405) );
  XOR U413 ( .A(n434), .B(n407), .Z(n406) );
  AND U414 ( .A(n484), .B(n485), .Z(n407) );
  XOR U415 ( .A(n436), .B(n435), .Z(n434) );
  AND U416 ( .A(n486), .B(n487), .Z(n435) );
  XOR U417 ( .A(n415), .B(n437), .Z(n436) );
  AND U418 ( .A(n488), .B(n489), .Z(n437) );
  XOR U419 ( .A(n411), .B(n416), .Z(n415) );
  AND U420 ( .A(n490), .B(n491), .Z(n416) );
  XOR U421 ( .A(n413), .B(n412), .Z(n411) );
  AND U422 ( .A(n492), .B(n493), .Z(n412) );
  XNOR U423 ( .A(n423), .B(n414), .Z(n413) );
  AND U424 ( .A(n494), .B(n495), .Z(n414) );
  XOR U425 ( .A(n433), .B(n422), .Z(n423) );
  AND U426 ( .A(n496), .B(n497), .Z(n422) );
  XNOR U427 ( .A(n498), .B(n428), .Z(n433) );
  XOR U428 ( .A(n429), .B(n499), .Z(n428) );
  AND U429 ( .A(n500), .B(n501), .Z(n499) );
  XOR U430 ( .A(n502), .B(n503), .Z(n429) );
  NOR U431 ( .A(n504), .B(n505), .Z(n503) );
  AND U432 ( .A(n506), .B(n507), .Z(n505) );
  AND U433 ( .A(n508), .B(n509), .Z(n504) );
  XNOR U434 ( .A(n506), .B(n507), .Z(n502) );
  XNOR U435 ( .A(n420), .B(n432), .Z(n498) );
  AND U436 ( .A(n510), .B(n511), .Z(n432) );
  AND U437 ( .A(n512), .B(n513), .Z(n420) );
  NOR U438 ( .A(n68), .B(n71), .Z(n438) );
  XNOR U439 ( .A(n443), .B(n442), .Z(n71) );
  NOR U440 ( .A(n212), .B(p_input[31]), .Z(n442) );
  IV U441 ( .A(p_input[30]), .Z(n212) );
  XOR U442 ( .A(n445), .B(n444), .Z(n443) );
  NOR U443 ( .A(n218), .B(p_input[29]), .Z(n444) );
  IV U444 ( .A(p_input[28]), .Z(n218) );
  XOR U445 ( .A(n447), .B(n446), .Z(n445) );
  NOR U446 ( .A(n223), .B(p_input[27]), .Z(n446) );
  IV U447 ( .A(p_input[26]), .Z(n223) );
  XOR U448 ( .A(n449), .B(n448), .Z(n447) );
  NOR U449 ( .A(n228), .B(p_input[25]), .Z(n448) );
  IV U450 ( .A(p_input[24]), .Z(n228) );
  XOR U451 ( .A(n451), .B(n450), .Z(n449) );
  NOR U452 ( .A(n259), .B(p_input[23]), .Z(n450) );
  IV U453 ( .A(p_input[22]), .Z(n259) );
  XOR U454 ( .A(n453), .B(n452), .Z(n451) );
  NOR U455 ( .A(n263), .B(p_input[21]), .Z(n452) );
  IV U456 ( .A(p_input[20]), .Z(n263) );
  XOR U457 ( .A(n455), .B(n454), .Z(n453) );
  NOR U458 ( .A(n266), .B(p_input[19]), .Z(n454) );
  IV U459 ( .A(p_input[18]), .Z(n266) );
  XOR U460 ( .A(n457), .B(n456), .Z(n455) );
  NOR U461 ( .A(n269), .B(p_input[17]), .Z(n456) );
  IV U462 ( .A(p_input[16]), .Z(n269) );
  XOR U463 ( .A(n459), .B(n458), .Z(n457) );
  NOR U464 ( .A(n272), .B(p_input[15]), .Z(n458) );
  IV U465 ( .A(p_input[14]), .Z(n272) );
  XOR U466 ( .A(n461), .B(n460), .Z(n459) );
  NOR U467 ( .A(n275), .B(p_input[13]), .Z(n460) );
  IV U468 ( .A(p_input[12]), .Z(n275) );
  XOR U469 ( .A(n475), .B(n474), .Z(n461) );
  NOR U470 ( .A(n290), .B(p_input[11]), .Z(n474) );
  IV U471 ( .A(p_input[10]), .Z(n290) );
  XOR U472 ( .A(n477), .B(n476), .Z(n475) );
  NOR U473 ( .A(n295), .B(p_input[9]), .Z(n476) );
  IV U474 ( .A(p_input[8]), .Z(n295) );
  XOR U475 ( .A(n465), .B(n464), .Z(n477) );
  NOR U476 ( .A(n291), .B(p_input[7]), .Z(n464) );
  IV U477 ( .A(p_input[6]), .Z(n291) );
  XOR U478 ( .A(n472), .B(n473), .Z(n465) );
  XOR U479 ( .A(n470), .B(n471), .Z(n473) );
  NOR U480 ( .A(n292), .B(p_input[3]), .Z(n471) );
  IV U481 ( .A(p_input[2]), .Z(n292) );
  NOR U482 ( .A(n293), .B(p_input[1]), .Z(n470) );
  IV U483 ( .A(p_input[0]), .Z(n293) );
  NOR U484 ( .A(n294), .B(p_input[5]), .Z(n472) );
  IV U485 ( .A(p_input[4]), .Z(n294) );
  XOR U486 ( .A(n479), .B(n478), .Z(n68) );
  NOR U487 ( .A(p_input[31]), .B(p_input[30]), .Z(n478) );
  XOR U488 ( .A(n481), .B(n480), .Z(n479) );
  NOR U489 ( .A(p_input[29]), .B(p_input[28]), .Z(n480) );
  XOR U490 ( .A(n483), .B(n482), .Z(n481) );
  NOR U491 ( .A(p_input[27]), .B(p_input[26]), .Z(n482) );
  XOR U492 ( .A(n485), .B(n484), .Z(n483) );
  NOR U493 ( .A(p_input[25]), .B(p_input[24]), .Z(n484) );
  XOR U494 ( .A(n487), .B(n486), .Z(n485) );
  NOR U495 ( .A(p_input[23]), .B(p_input[22]), .Z(n486) );
  XOR U496 ( .A(n489), .B(n488), .Z(n487) );
  NOR U497 ( .A(p_input[21]), .B(p_input[20]), .Z(n488) );
  XOR U498 ( .A(n491), .B(n490), .Z(n489) );
  NOR U499 ( .A(p_input[19]), .B(p_input[18]), .Z(n490) );
  XOR U500 ( .A(n493), .B(n492), .Z(n491) );
  NOR U501 ( .A(p_input[17]), .B(p_input[16]), .Z(n492) );
  XOR U502 ( .A(n495), .B(n494), .Z(n493) );
  NOR U503 ( .A(p_input[15]), .B(p_input[14]), .Z(n494) );
  XOR U504 ( .A(n497), .B(n496), .Z(n495) );
  NOR U505 ( .A(p_input[13]), .B(p_input[12]), .Z(n496) );
  XOR U506 ( .A(n511), .B(n510), .Z(n497) );
  NOR U507 ( .A(p_input[11]), .B(p_input[10]), .Z(n510) );
  XOR U508 ( .A(n513), .B(n512), .Z(n511) );
  NOR U509 ( .A(p_input[9]), .B(p_input[8]), .Z(n512) );
  XOR U510 ( .A(n501), .B(n500), .Z(n513) );
  NOR U511 ( .A(p_input[7]), .B(p_input[6]), .Z(n500) );
  XOR U512 ( .A(n508), .B(n509), .Z(n501) );
  XOR U513 ( .A(n506), .B(n507), .Z(n509) );
  NOR U514 ( .A(p_input[3]), .B(p_input[2]), .Z(n507) );
  NOR U515 ( .A(p_input[1]), .B(p_input[0]), .Z(n506) );
  NOR U516 ( .A(p_input[5]), .B(p_input[4]), .Z(n508) );
endmodule

