
module auction_BMR_N2_W16 ( p_input, o );
  input [63:0] p_input;
  output [17:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323;

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(o[1]), .B(n3), .Z(n1) );
  XOR U3 ( .A(n2), .B(n4), .Z(n3) );
  XNOR U4 ( .A(n5), .B(n6), .Z(o[8]) );
  AND U5 ( .A(o[1]), .B(n7), .Z(n5) );
  XOR U6 ( .A(n8), .B(n6), .Z(n7) );
  XNOR U7 ( .A(n9), .B(n10), .Z(o[7]) );
  AND U8 ( .A(o[1]), .B(n11), .Z(n9) );
  XOR U9 ( .A(n12), .B(n10), .Z(n11) );
  XNOR U10 ( .A(n13), .B(n14), .Z(o[6]) );
  AND U11 ( .A(o[1]), .B(n15), .Z(n13) );
  XOR U12 ( .A(n16), .B(n14), .Z(n15) );
  XNOR U13 ( .A(n17), .B(n18), .Z(o[5]) );
  AND U14 ( .A(o[1]), .B(n19), .Z(n17) );
  XOR U15 ( .A(n20), .B(n18), .Z(n19) );
  XNOR U16 ( .A(n21), .B(n22), .Z(o[4]) );
  AND U17 ( .A(o[1]), .B(n23), .Z(n21) );
  XOR U18 ( .A(n24), .B(n22), .Z(n23) );
  XOR U19 ( .A(n25), .B(n26), .Z(o[3]) );
  AND U20 ( .A(o[1]), .B(n27), .Z(n25) );
  XOR U21 ( .A(n28), .B(n29), .Z(n27) );
  XNOR U22 ( .A(n30), .B(n31), .Z(o[2]) );
  AND U23 ( .A(o[1]), .B(n32), .Z(n30) );
  XNOR U24 ( .A(n33), .B(n31), .Z(n32) );
  AND U25 ( .A(n34), .B(n35), .Z(o[17]) );
  XNOR U26 ( .A(n36), .B(n37), .Z(o[16]) );
  AND U27 ( .A(o[1]), .B(n38), .Z(n36) );
  XOR U28 ( .A(n39), .B(n37), .Z(n38) );
  XNOR U29 ( .A(n40), .B(n41), .Z(o[15]) );
  AND U30 ( .A(o[1]), .B(n42), .Z(n40) );
  XOR U31 ( .A(n43), .B(n41), .Z(n42) );
  XNOR U32 ( .A(n44), .B(n45), .Z(o[14]) );
  AND U33 ( .A(o[1]), .B(n46), .Z(n44) );
  XOR U34 ( .A(n47), .B(n45), .Z(n46) );
  XNOR U35 ( .A(n48), .B(n49), .Z(o[13]) );
  AND U36 ( .A(o[1]), .B(n50), .Z(n48) );
  XOR U37 ( .A(n51), .B(n49), .Z(n50) );
  XNOR U38 ( .A(n52), .B(n53), .Z(o[12]) );
  AND U39 ( .A(o[1]), .B(n54), .Z(n52) );
  XOR U40 ( .A(n55), .B(n53), .Z(n54) );
  XNOR U41 ( .A(n56), .B(n57), .Z(o[11]) );
  AND U42 ( .A(o[1]), .B(n58), .Z(n56) );
  XOR U43 ( .A(n59), .B(n57), .Z(n58) );
  XNOR U44 ( .A(n60), .B(n61), .Z(o[10]) );
  AND U45 ( .A(o[1]), .B(n62), .Z(n60) );
  XOR U46 ( .A(n63), .B(n61), .Z(n62) );
  XOR U47 ( .A(n64), .B(n65), .Z(o[0]) );
  AND U48 ( .A(o[1]), .B(n66), .Z(n65) );
  XOR U49 ( .A(n64), .B(n67), .Z(n66) );
  XOR U50 ( .A(n68), .B(n69), .Z(o[1]) );
  AND U51 ( .A(n70), .B(n71), .Z(n69) );
  XNOR U52 ( .A(n35), .B(n68), .Z(n71) );
  AND U53 ( .A(p_input[63]), .B(p_input[47]), .Z(n35) );
  XOR U54 ( .A(n68), .B(n34), .Z(n70) );
  AND U55 ( .A(p_input[15]), .B(p_input[31]), .Z(n34) );
  XOR U56 ( .A(n72), .B(n73), .Z(n68) );
  AND U57 ( .A(n74), .B(n75), .Z(n73) );
  XOR U58 ( .A(n72), .B(n39), .Z(n75) );
  XNOR U59 ( .A(p_input[46]), .B(n76), .Z(n39) );
  AND U60 ( .A(n67), .B(n77), .Z(n76) );
  XOR U61 ( .A(p_input[62]), .B(p_input[46]), .Z(n77) );
  XNOR U62 ( .A(n37), .B(n72), .Z(n74) );
  XOR U63 ( .A(n78), .B(n79), .Z(n37) );
  AND U64 ( .A(n64), .B(n80), .Z(n79) );
  XOR U65 ( .A(p_input[30]), .B(p_input[14]), .Z(n80) );
  XOR U66 ( .A(n81), .B(n82), .Z(n72) );
  AND U67 ( .A(n83), .B(n84), .Z(n82) );
  XOR U68 ( .A(n81), .B(n43), .Z(n84) );
  XNOR U69 ( .A(p_input[45]), .B(n85), .Z(n43) );
  AND U70 ( .A(n67), .B(n86), .Z(n85) );
  XOR U71 ( .A(p_input[61]), .B(p_input[45]), .Z(n86) );
  XNOR U72 ( .A(n41), .B(n81), .Z(n83) );
  XOR U73 ( .A(n87), .B(n88), .Z(n41) );
  AND U74 ( .A(n64), .B(n89), .Z(n88) );
  XOR U75 ( .A(p_input[29]), .B(p_input[13]), .Z(n89) );
  XOR U76 ( .A(n90), .B(n91), .Z(n81) );
  AND U77 ( .A(n92), .B(n93), .Z(n91) );
  XOR U78 ( .A(n90), .B(n47), .Z(n93) );
  XNOR U79 ( .A(p_input[44]), .B(n94), .Z(n47) );
  AND U80 ( .A(n67), .B(n95), .Z(n94) );
  XOR U81 ( .A(p_input[60]), .B(p_input[44]), .Z(n95) );
  XNOR U82 ( .A(n45), .B(n90), .Z(n92) );
  XOR U83 ( .A(n96), .B(n97), .Z(n45) );
  AND U84 ( .A(n64), .B(n98), .Z(n97) );
  XOR U85 ( .A(p_input[28]), .B(p_input[12]), .Z(n98) );
  XOR U86 ( .A(n99), .B(n100), .Z(n90) );
  AND U87 ( .A(n101), .B(n102), .Z(n100) );
  XOR U88 ( .A(n99), .B(n51), .Z(n102) );
  XNOR U89 ( .A(p_input[43]), .B(n103), .Z(n51) );
  AND U90 ( .A(n67), .B(n104), .Z(n103) );
  XOR U91 ( .A(p_input[59]), .B(p_input[43]), .Z(n104) );
  XNOR U92 ( .A(n49), .B(n99), .Z(n101) );
  XOR U93 ( .A(n105), .B(n106), .Z(n49) );
  AND U94 ( .A(n64), .B(n107), .Z(n106) );
  XOR U95 ( .A(p_input[27]), .B(p_input[11]), .Z(n107) );
  XOR U96 ( .A(n108), .B(n109), .Z(n99) );
  AND U97 ( .A(n110), .B(n111), .Z(n109) );
  XOR U98 ( .A(n108), .B(n55), .Z(n111) );
  XNOR U99 ( .A(p_input[42]), .B(n112), .Z(n55) );
  AND U100 ( .A(n67), .B(n113), .Z(n112) );
  XOR U101 ( .A(p_input[58]), .B(p_input[42]), .Z(n113) );
  XNOR U102 ( .A(n53), .B(n108), .Z(n110) );
  XOR U103 ( .A(n114), .B(n115), .Z(n53) );
  AND U104 ( .A(n64), .B(n116), .Z(n115) );
  XOR U105 ( .A(p_input[26]), .B(p_input[10]), .Z(n116) );
  XOR U106 ( .A(n117), .B(n118), .Z(n108) );
  AND U107 ( .A(n119), .B(n120), .Z(n118) );
  XOR U108 ( .A(n117), .B(n59), .Z(n120) );
  XNOR U109 ( .A(p_input[41]), .B(n121), .Z(n59) );
  AND U110 ( .A(n67), .B(n122), .Z(n121) );
  XOR U111 ( .A(p_input[57]), .B(p_input[41]), .Z(n122) );
  XNOR U112 ( .A(n57), .B(n117), .Z(n119) );
  XOR U113 ( .A(n123), .B(n124), .Z(n57) );
  AND U114 ( .A(n64), .B(n125), .Z(n124) );
  XOR U115 ( .A(p_input[9]), .B(p_input[25]), .Z(n125) );
  XOR U116 ( .A(n126), .B(n127), .Z(n117) );
  AND U117 ( .A(n128), .B(n129), .Z(n127) );
  XOR U118 ( .A(n126), .B(n63), .Z(n129) );
  XNOR U119 ( .A(p_input[40]), .B(n130), .Z(n63) );
  AND U120 ( .A(n67), .B(n131), .Z(n130) );
  XOR U121 ( .A(p_input[56]), .B(p_input[40]), .Z(n131) );
  XNOR U122 ( .A(n61), .B(n126), .Z(n128) );
  XOR U123 ( .A(n132), .B(n133), .Z(n61) );
  AND U124 ( .A(n64), .B(n134), .Z(n133) );
  XOR U125 ( .A(p_input[8]), .B(p_input[24]), .Z(n134) );
  XOR U126 ( .A(n135), .B(n136), .Z(n126) );
  AND U127 ( .A(n137), .B(n138), .Z(n136) );
  XOR U128 ( .A(n4), .B(n135), .Z(n138) );
  XNOR U129 ( .A(p_input[39]), .B(n139), .Z(n4) );
  AND U130 ( .A(n67), .B(n140), .Z(n139) );
  XOR U131 ( .A(p_input[55]), .B(p_input[39]), .Z(n140) );
  XNOR U132 ( .A(n135), .B(n2), .Z(n137) );
  XOR U133 ( .A(n141), .B(n142), .Z(n2) );
  AND U134 ( .A(n64), .B(n143), .Z(n142) );
  XOR U135 ( .A(p_input[7]), .B(p_input[23]), .Z(n143) );
  XOR U136 ( .A(n144), .B(n145), .Z(n135) );
  AND U137 ( .A(n146), .B(n147), .Z(n145) );
  XOR U138 ( .A(n144), .B(n8), .Z(n147) );
  XNOR U139 ( .A(p_input[38]), .B(n148), .Z(n8) );
  AND U140 ( .A(n67), .B(n149), .Z(n148) );
  XOR U141 ( .A(p_input[54]), .B(p_input[38]), .Z(n149) );
  XNOR U142 ( .A(n6), .B(n144), .Z(n146) );
  XOR U143 ( .A(n150), .B(n151), .Z(n6) );
  AND U144 ( .A(n64), .B(n152), .Z(n151) );
  XOR U145 ( .A(p_input[6]), .B(p_input[22]), .Z(n152) );
  XOR U146 ( .A(n153), .B(n154), .Z(n144) );
  AND U147 ( .A(n155), .B(n156), .Z(n154) );
  XOR U148 ( .A(n153), .B(n12), .Z(n156) );
  XNOR U149 ( .A(p_input[37]), .B(n157), .Z(n12) );
  AND U150 ( .A(n67), .B(n158), .Z(n157) );
  XOR U151 ( .A(p_input[53]), .B(p_input[37]), .Z(n158) );
  XNOR U152 ( .A(n10), .B(n153), .Z(n155) );
  XOR U153 ( .A(n159), .B(n160), .Z(n10) );
  AND U154 ( .A(n64), .B(n161), .Z(n160) );
  XOR U155 ( .A(p_input[5]), .B(p_input[21]), .Z(n161) );
  XOR U156 ( .A(n162), .B(n163), .Z(n153) );
  AND U157 ( .A(n164), .B(n165), .Z(n163) );
  XOR U158 ( .A(n162), .B(n16), .Z(n165) );
  XNOR U159 ( .A(p_input[36]), .B(n166), .Z(n16) );
  AND U160 ( .A(n67), .B(n167), .Z(n166) );
  XOR U161 ( .A(p_input[52]), .B(p_input[36]), .Z(n167) );
  XNOR U162 ( .A(n14), .B(n162), .Z(n164) );
  XOR U163 ( .A(n168), .B(n169), .Z(n14) );
  AND U164 ( .A(n64), .B(n170), .Z(n169) );
  XOR U165 ( .A(p_input[4]), .B(p_input[20]), .Z(n170) );
  XOR U166 ( .A(n171), .B(n172), .Z(n162) );
  AND U167 ( .A(n173), .B(n174), .Z(n172) );
  XOR U168 ( .A(n171), .B(n20), .Z(n174) );
  XNOR U169 ( .A(p_input[35]), .B(n175), .Z(n20) );
  AND U170 ( .A(n67), .B(n176), .Z(n175) );
  XOR U171 ( .A(p_input[51]), .B(p_input[35]), .Z(n176) );
  XNOR U172 ( .A(n18), .B(n171), .Z(n173) );
  XOR U173 ( .A(n177), .B(n178), .Z(n18) );
  AND U174 ( .A(n64), .B(n179), .Z(n178) );
  XOR U175 ( .A(p_input[3]), .B(p_input[19]), .Z(n179) );
  XOR U176 ( .A(n180), .B(n181), .Z(n171) );
  AND U177 ( .A(n182), .B(n183), .Z(n181) );
  XOR U178 ( .A(n180), .B(n24), .Z(n183) );
  XNOR U179 ( .A(p_input[34]), .B(n184), .Z(n24) );
  AND U180 ( .A(n67), .B(n185), .Z(n184) );
  XOR U181 ( .A(p_input[50]), .B(p_input[34]), .Z(n185) );
  XNOR U182 ( .A(n22), .B(n180), .Z(n182) );
  XOR U183 ( .A(n186), .B(n187), .Z(n22) );
  AND U184 ( .A(n64), .B(n188), .Z(n187) );
  XOR U185 ( .A(p_input[2]), .B(p_input[18]), .Z(n188) );
  XNOR U186 ( .A(n189), .B(n190), .Z(n180) );
  AND U187 ( .A(n191), .B(n192), .Z(n190) );
  XNOR U188 ( .A(n189), .B(n28), .Z(n192) );
  XNOR U189 ( .A(p_input[33]), .B(n193), .Z(n28) );
  AND U190 ( .A(n67), .B(n194), .Z(n193) );
  XNOR U191 ( .A(p_input[49]), .B(n195), .Z(n194) );
  IV U192 ( .A(p_input[33]), .Z(n195) );
  XOR U193 ( .A(n29), .B(n189), .Z(n191) );
  IV U194 ( .A(n26), .Z(n29) );
  XOR U195 ( .A(p_input[1]), .B(n196), .Z(n26) );
  AND U196 ( .A(n64), .B(n197), .Z(n196) );
  XOR U197 ( .A(p_input[1]), .B(p_input[17]), .Z(n197) );
  AND U198 ( .A(n31), .B(n33), .Z(n189) );
  XOR U199 ( .A(p_input[32]), .B(n198), .Z(n33) );
  AND U200 ( .A(n67), .B(n199), .Z(n198) );
  XOR U201 ( .A(p_input[48]), .B(p_input[32]), .Z(n199) );
  XOR U202 ( .A(n200), .B(n201), .Z(n67) );
  AND U203 ( .A(n202), .B(n203), .Z(n201) );
  XNOR U204 ( .A(p_input[63]), .B(n200), .Z(n203) );
  XOR U205 ( .A(n200), .B(p_input[47]), .Z(n202) );
  XOR U206 ( .A(n204), .B(n205), .Z(n200) );
  AND U207 ( .A(n206), .B(n207), .Z(n205) );
  XNOR U208 ( .A(p_input[62]), .B(n204), .Z(n207) );
  XOR U209 ( .A(n204), .B(p_input[46]), .Z(n206) );
  XOR U210 ( .A(n208), .B(n209), .Z(n204) );
  AND U211 ( .A(n210), .B(n211), .Z(n209) );
  XNOR U212 ( .A(p_input[61]), .B(n208), .Z(n211) );
  XOR U213 ( .A(n208), .B(p_input[45]), .Z(n210) );
  XOR U214 ( .A(n212), .B(n213), .Z(n208) );
  AND U215 ( .A(n214), .B(n215), .Z(n213) );
  XNOR U216 ( .A(p_input[60]), .B(n212), .Z(n215) );
  XOR U217 ( .A(n212), .B(p_input[44]), .Z(n214) );
  XOR U218 ( .A(n216), .B(n217), .Z(n212) );
  AND U219 ( .A(n218), .B(n219), .Z(n217) );
  XNOR U220 ( .A(p_input[59]), .B(n216), .Z(n219) );
  XOR U221 ( .A(n216), .B(p_input[43]), .Z(n218) );
  XOR U222 ( .A(n220), .B(n221), .Z(n216) );
  AND U223 ( .A(n222), .B(n223), .Z(n221) );
  XNOR U224 ( .A(p_input[58]), .B(n220), .Z(n223) );
  XOR U225 ( .A(n220), .B(p_input[42]), .Z(n222) );
  XOR U226 ( .A(n224), .B(n225), .Z(n220) );
  AND U227 ( .A(n226), .B(n227), .Z(n225) );
  XNOR U228 ( .A(p_input[57]), .B(n224), .Z(n227) );
  XOR U229 ( .A(n224), .B(p_input[41]), .Z(n226) );
  XOR U230 ( .A(n228), .B(n229), .Z(n224) );
  AND U231 ( .A(n230), .B(n231), .Z(n229) );
  XNOR U232 ( .A(p_input[56]), .B(n228), .Z(n231) );
  XOR U233 ( .A(n228), .B(p_input[40]), .Z(n230) );
  XOR U234 ( .A(n232), .B(n233), .Z(n228) );
  AND U235 ( .A(n234), .B(n235), .Z(n233) );
  XNOR U236 ( .A(p_input[55]), .B(n232), .Z(n235) );
  XOR U237 ( .A(n232), .B(p_input[39]), .Z(n234) );
  XOR U238 ( .A(n236), .B(n237), .Z(n232) );
  AND U239 ( .A(n238), .B(n239), .Z(n237) );
  XNOR U240 ( .A(p_input[54]), .B(n236), .Z(n239) );
  XOR U241 ( .A(n236), .B(p_input[38]), .Z(n238) );
  XOR U242 ( .A(n240), .B(n241), .Z(n236) );
  AND U243 ( .A(n242), .B(n243), .Z(n241) );
  XNOR U244 ( .A(p_input[53]), .B(n240), .Z(n243) );
  XOR U245 ( .A(n240), .B(p_input[37]), .Z(n242) );
  XOR U246 ( .A(n244), .B(n245), .Z(n240) );
  AND U247 ( .A(n246), .B(n247), .Z(n245) );
  XNOR U248 ( .A(p_input[52]), .B(n244), .Z(n247) );
  XOR U249 ( .A(n244), .B(p_input[36]), .Z(n246) );
  XOR U250 ( .A(n248), .B(n249), .Z(n244) );
  AND U251 ( .A(n250), .B(n251), .Z(n249) );
  XNOR U252 ( .A(p_input[51]), .B(n248), .Z(n251) );
  XOR U253 ( .A(n248), .B(p_input[35]), .Z(n250) );
  XOR U254 ( .A(n252), .B(n253), .Z(n248) );
  AND U255 ( .A(n254), .B(n255), .Z(n253) );
  XNOR U256 ( .A(p_input[50]), .B(n252), .Z(n255) );
  XOR U257 ( .A(n252), .B(p_input[34]), .Z(n254) );
  XNOR U258 ( .A(n256), .B(n257), .Z(n252) );
  AND U259 ( .A(n258), .B(n259), .Z(n257) );
  XOR U260 ( .A(p_input[49]), .B(n256), .Z(n259) );
  XNOR U261 ( .A(p_input[33]), .B(n256), .Z(n258) );
  AND U262 ( .A(p_input[48]), .B(n260), .Z(n256) );
  IV U263 ( .A(p_input[32]), .Z(n260) );
  XNOR U264 ( .A(p_input[0]), .B(n261), .Z(n31) );
  AND U265 ( .A(n64), .B(n262), .Z(n261) );
  XOR U266 ( .A(p_input[16]), .B(p_input[0]), .Z(n262) );
  XOR U267 ( .A(n263), .B(n264), .Z(n64) );
  AND U268 ( .A(n265), .B(n266), .Z(n264) );
  XNOR U269 ( .A(p_input[31]), .B(n263), .Z(n266) );
  XOR U270 ( .A(n263), .B(p_input[15]), .Z(n265) );
  XOR U271 ( .A(n267), .B(n268), .Z(n263) );
  AND U272 ( .A(n269), .B(n270), .Z(n268) );
  XNOR U273 ( .A(p_input[30]), .B(n267), .Z(n270) );
  XNOR U274 ( .A(n267), .B(n78), .Z(n269) );
  IV U275 ( .A(p_input[14]), .Z(n78) );
  XOR U276 ( .A(n271), .B(n272), .Z(n267) );
  AND U277 ( .A(n273), .B(n274), .Z(n272) );
  XNOR U278 ( .A(p_input[29]), .B(n271), .Z(n274) );
  XNOR U279 ( .A(n271), .B(n87), .Z(n273) );
  IV U280 ( .A(p_input[13]), .Z(n87) );
  XOR U281 ( .A(n275), .B(n276), .Z(n271) );
  AND U282 ( .A(n277), .B(n278), .Z(n276) );
  XNOR U283 ( .A(p_input[28]), .B(n275), .Z(n278) );
  XNOR U284 ( .A(n275), .B(n96), .Z(n277) );
  IV U285 ( .A(p_input[12]), .Z(n96) );
  XOR U286 ( .A(n279), .B(n280), .Z(n275) );
  AND U287 ( .A(n281), .B(n282), .Z(n280) );
  XNOR U288 ( .A(p_input[27]), .B(n279), .Z(n282) );
  XNOR U289 ( .A(n279), .B(n105), .Z(n281) );
  IV U290 ( .A(p_input[11]), .Z(n105) );
  XOR U291 ( .A(n283), .B(n284), .Z(n279) );
  AND U292 ( .A(n285), .B(n286), .Z(n284) );
  XNOR U293 ( .A(p_input[26]), .B(n283), .Z(n286) );
  XNOR U294 ( .A(n283), .B(n114), .Z(n285) );
  IV U295 ( .A(p_input[10]), .Z(n114) );
  XOR U296 ( .A(n287), .B(n288), .Z(n283) );
  AND U297 ( .A(n289), .B(n290), .Z(n288) );
  XNOR U298 ( .A(p_input[25]), .B(n287), .Z(n290) );
  XNOR U299 ( .A(n287), .B(n123), .Z(n289) );
  IV U300 ( .A(p_input[9]), .Z(n123) );
  XOR U301 ( .A(n291), .B(n292), .Z(n287) );
  AND U302 ( .A(n293), .B(n294), .Z(n292) );
  XNOR U303 ( .A(p_input[24]), .B(n291), .Z(n294) );
  XNOR U304 ( .A(n291), .B(n132), .Z(n293) );
  IV U305 ( .A(p_input[8]), .Z(n132) );
  XOR U306 ( .A(n295), .B(n296), .Z(n291) );
  AND U307 ( .A(n297), .B(n298), .Z(n296) );
  XNOR U308 ( .A(p_input[23]), .B(n295), .Z(n298) );
  XNOR U309 ( .A(n295), .B(n141), .Z(n297) );
  IV U310 ( .A(p_input[7]), .Z(n141) );
  XOR U311 ( .A(n299), .B(n300), .Z(n295) );
  AND U312 ( .A(n301), .B(n302), .Z(n300) );
  XNOR U313 ( .A(p_input[22]), .B(n299), .Z(n302) );
  XNOR U314 ( .A(n299), .B(n150), .Z(n301) );
  IV U315 ( .A(p_input[6]), .Z(n150) );
  XOR U316 ( .A(n303), .B(n304), .Z(n299) );
  AND U317 ( .A(n305), .B(n306), .Z(n304) );
  XNOR U318 ( .A(p_input[21]), .B(n303), .Z(n306) );
  XNOR U319 ( .A(n303), .B(n159), .Z(n305) );
  IV U320 ( .A(p_input[5]), .Z(n159) );
  XOR U321 ( .A(n307), .B(n308), .Z(n303) );
  AND U322 ( .A(n309), .B(n310), .Z(n308) );
  XNOR U323 ( .A(p_input[20]), .B(n307), .Z(n310) );
  XNOR U324 ( .A(n307), .B(n168), .Z(n309) );
  IV U325 ( .A(p_input[4]), .Z(n168) );
  XOR U326 ( .A(n311), .B(n312), .Z(n307) );
  AND U327 ( .A(n313), .B(n314), .Z(n312) );
  XNOR U328 ( .A(p_input[19]), .B(n311), .Z(n314) );
  XNOR U329 ( .A(n311), .B(n177), .Z(n313) );
  IV U330 ( .A(p_input[3]), .Z(n177) );
  XOR U331 ( .A(n315), .B(n316), .Z(n311) );
  AND U332 ( .A(n317), .B(n318), .Z(n316) );
  XNOR U333 ( .A(p_input[18]), .B(n315), .Z(n318) );
  XNOR U334 ( .A(n315), .B(n186), .Z(n317) );
  IV U335 ( .A(p_input[2]), .Z(n186) );
  XNOR U336 ( .A(n319), .B(n320), .Z(n315) );
  AND U337 ( .A(n321), .B(n322), .Z(n320) );
  XOR U338 ( .A(p_input[17]), .B(n319), .Z(n322) );
  XNOR U339 ( .A(p_input[1]), .B(n319), .Z(n321) );
  AND U340 ( .A(p_input[16]), .B(n323), .Z(n319) );
  IV U341 ( .A(p_input[0]), .Z(n323) );
endmodule

