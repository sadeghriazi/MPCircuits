
module knn_comb_BMR_W32_K2_N64 ( p_input, o );
  input [2079:0] p_input;
  output [63:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/min_val_out[0][16] , \knn_comb_/min_val_out[0][17] ,
         \knn_comb_/min_val_out[0][18] , \knn_comb_/min_val_out[0][19] ,
         \knn_comb_/min_val_out[0][20] , \knn_comb_/min_val_out[0][21] ,
         \knn_comb_/min_val_out[0][22] , \knn_comb_/min_val_out[0][23] ,
         \knn_comb_/min_val_out[0][24] , \knn_comb_/min_val_out[0][25] ,
         \knn_comb_/min_val_out[0][26] , \knn_comb_/min_val_out[0][27] ,
         \knn_comb_/min_val_out[0][28] , \knn_comb_/min_val_out[0][29] ,
         \knn_comb_/min_val_out[0][30] , \knn_comb_/min_val_out[0][31] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][31] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
         n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
         n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
         n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
         n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
         n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
         n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
         n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
         n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
         n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
         n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
         n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459,
         n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
         n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
         n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483,
         n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
         n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
         n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507,
         n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
         n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
         n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
         n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
         n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
         n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555,
         n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
         n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
         n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579,
         n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
         n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
         n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603,
         n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
         n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
         n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
         n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635,
         n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643,
         n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651,
         n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
         n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
         n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675,
         n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683,
         n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691,
         n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699,
         n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707,
         n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715,
         n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723,
         n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
         n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
         n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747,
         n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755,
         n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763,
         n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771,
         n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
         n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787,
         n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795,
         n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
         n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
         n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819,
         n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827,
         n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835,
         n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843,
         n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851,
         n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859,
         n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867,
         n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
         n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
         n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891,
         n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899,
         n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
         n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915,
         n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923,
         n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931,
         n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939,
         n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947,
         n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955,
         n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963,
         n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971,
         n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979,
         n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987,
         n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995,
         n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003,
         n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011,
         n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019,
         n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027,
         n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035,
         n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043,
         n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
         n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059,
         n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067,
         n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075,
         n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083,
         n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091,
         n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099,
         n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107,
         n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115,
         n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
         n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131,
         n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139,
         n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147,
         n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155,
         n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163,
         n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171,
         n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179,
         n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187,
         n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
         n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203,
         n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211,
         n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219,
         n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227,
         n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235,
         n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243,
         n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251,
         n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259,
         n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267,
         n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275,
         n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283,
         n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291,
         n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299,
         n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307,
         n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315,
         n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323,
         n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331,
         n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339,
         n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347,
         n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355,
         n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363,
         n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371,
         n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379,
         n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387,
         n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395,
         n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403,
         n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411,
         n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419,
         n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427,
         n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435,
         n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443,
         n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451,
         n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459,
         n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467,
         n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475,
         n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483,
         n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491,
         n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499,
         n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507,
         n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515,
         n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523,
         n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531,
         n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539,
         n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547,
         n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555,
         n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563,
         n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571,
         n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579,
         n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587,
         n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595,
         n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603,
         n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611,
         n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619,
         n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627,
         n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635,
         n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643,
         n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651,
         n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659,
         n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667,
         n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675,
         n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683,
         n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691,
         n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699,
         n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707,
         n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715,
         n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723,
         n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731,
         n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739,
         n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747,
         n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755,
         n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763,
         n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771,
         n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779,
         n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787,
         n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795,
         n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803,
         n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811,
         n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819,
         n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827,
         n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835,
         n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843,
         n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851,
         n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859,
         n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867,
         n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875,
         n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883,
         n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891,
         n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899,
         n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907,
         n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915,
         n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923,
         n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931,
         n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939,
         n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947,
         n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955,
         n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963,
         n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971,
         n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979,
         n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987,
         n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995,
         n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003,
         n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011,
         n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019,
         n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027,
         n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035,
         n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043,
         n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051,
         n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059,
         n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067,
         n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075,
         n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083,
         n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091,
         n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099,
         n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107,
         n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115,
         n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123,
         n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131,
         n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139,
         n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147,
         n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155,
         n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163,
         n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171,
         n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179,
         n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187,
         n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195,
         n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203,
         n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211,
         n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219,
         n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227,
         n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235,
         n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243,
         n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251,
         n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259,
         n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267,
         n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275,
         n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283,
         n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291,
         n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299,
         n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307,
         n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315,
         n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323,
         n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331,
         n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339,
         n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347,
         n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355,
         n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363,
         n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371,
         n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379,
         n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387,
         n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395,
         n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403,
         n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411,
         n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419,
         n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427,
         n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435,
         n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443,
         n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451,
         n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459,
         n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467,
         n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475,
         n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483,
         n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491,
         n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499,
         n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507,
         n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515,
         n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523,
         n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531,
         n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539,
         n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547,
         n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555,
         n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563,
         n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571,
         n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579,
         n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587,
         n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595,
         n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603,
         n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611,
         n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619,
         n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627,
         n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635,
         n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643,
         n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651,
         n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659,
         n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667,
         n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675,
         n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683,
         n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691,
         n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699,
         n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707,
         n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715,
         n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723,
         n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731,
         n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739,
         n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747,
         n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755,
         n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763,
         n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771,
         n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779,
         n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787,
         n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795,
         n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803,
         n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811,
         n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819,
         n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827,
         n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835,
         n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843,
         n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851,
         n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859,
         n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867,
         n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875,
         n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883,
         n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891,
         n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899,
         n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907,
         n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915,
         n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923,
         n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931,
         n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939,
         n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
         n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955,
         n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963,
         n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971,
         n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979,
         n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987,
         n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995,
         n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003,
         n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011,
         n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019,
         n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027,
         n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035,
         n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043,
         n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051,
         n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059,
         n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067,
         n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075,
         n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083,
         n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091,
         n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099,
         n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107,
         n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115,
         n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123,
         n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131,
         n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139,
         n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147,
         n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155,
         n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163,
         n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171,
         n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179,
         n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187,
         n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195,
         n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203,
         n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211,
         n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219,
         n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227,
         n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235,
         n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243,
         n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251,
         n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259,
         n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267,
         n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275,
         n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283,
         n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291,
         n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299,
         n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307,
         n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315,
         n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323,
         n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331,
         n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339,
         n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347,
         n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355,
         n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363,
         n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371,
         n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379,
         n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387,
         n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395,
         n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403,
         n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411,
         n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419,
         n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427,
         n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435,
         n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443,
         n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451,
         n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459,
         n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467,
         n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475,
         n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483,
         n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491,
         n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499,
         n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507,
         n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515,
         n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523,
         n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531,
         n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539,
         n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547,
         n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555,
         n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563,
         n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571,
         n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579,
         n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587,
         n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595,
         n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603,
         n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611,
         n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619,
         n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627,
         n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635,
         n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643,
         n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651,
         n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659,
         n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667,
         n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675,
         n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683,
         n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691,
         n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699,
         n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707,
         n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715,
         n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723,
         n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731,
         n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739,
         n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747,
         n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755,
         n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763,
         n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771,
         n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779,
         n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787,
         n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795,
         n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803,
         n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811,
         n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819,
         n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827,
         n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835,
         n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843,
         n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851,
         n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859,
         n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867,
         n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875,
         n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883,
         n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891,
         n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899,
         n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907,
         n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915,
         n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923,
         n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931,
         n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939,
         n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947,
         n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955,
         n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963,
         n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971,
         n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979,
         n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987,
         n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995,
         n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003,
         n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011,
         n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019,
         n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027,
         n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035,
         n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043,
         n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051,
         n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059,
         n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067,
         n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075,
         n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083,
         n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091,
         n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099,
         n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107,
         n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115,
         n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123,
         n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131,
         n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139,
         n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147,
         n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155,
         n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163,
         n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171,
         n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179,
         n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187,
         n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195,
         n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203,
         n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211,
         n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219,
         n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227,
         n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235,
         n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243,
         n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251,
         n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259,
         n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267,
         n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275,
         n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283,
         n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291,
         n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299,
         n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307,
         n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315,
         n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323,
         n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331,
         n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339,
         n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347,
         n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355,
         n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363,
         n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371,
         n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379,
         n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387,
         n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395,
         n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403,
         n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411,
         n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419,
         n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427,
         n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435,
         n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443,
         n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451,
         n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459,
         n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467,
         n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475,
         n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483,
         n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491,
         n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499,
         n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507,
         n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515,
         n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523,
         n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531,
         n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539,
         n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547,
         n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555,
         n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563,
         n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571,
         n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579,
         n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587,
         n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595,
         n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603,
         n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611,
         n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619,
         n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627,
         n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635,
         n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643,
         n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651,
         n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659,
         n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667,
         n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675,
         n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683,
         n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691,
         n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699,
         n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707,
         n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715,
         n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723,
         n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731,
         n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739,
         n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747,
         n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755,
         n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763,
         n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771,
         n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779,
         n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787,
         n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795,
         n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803,
         n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811,
         n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819,
         n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827,
         n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835,
         n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843,
         n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851,
         n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859,
         n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867,
         n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875,
         n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883,
         n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891,
         n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899,
         n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907,
         n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915,
         n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923,
         n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931,
         n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939,
         n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947,
         n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955,
         n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963,
         n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971,
         n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979,
         n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987,
         n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995,
         n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003,
         n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011,
         n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019,
         n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027,
         n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035,
         n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043,
         n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051,
         n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059,
         n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067,
         n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075,
         n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083,
         n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091,
         n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099,
         n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107,
         n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115,
         n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123,
         n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131,
         n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139,
         n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147,
         n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155,
         n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163,
         n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171,
         n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179,
         n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187,
         n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195,
         n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203,
         n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211,
         n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219,
         n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227,
         n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235,
         n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243,
         n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251,
         n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259,
         n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267,
         n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275,
         n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283,
         n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291,
         n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299,
         n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307,
         n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315,
         n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323,
         n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331,
         n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339,
         n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347,
         n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355,
         n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363,
         n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371,
         n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379,
         n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387,
         n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395,
         n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403,
         n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411,
         n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419,
         n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427,
         n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435,
         n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443,
         n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451,
         n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459,
         n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467,
         n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475,
         n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483,
         n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491,
         n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499,
         n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507,
         n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515,
         n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523,
         n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531,
         n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539,
         n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547,
         n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555,
         n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563,
         n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571,
         n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579,
         n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587,
         n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595,
         n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603,
         n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611,
         n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619,
         n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627,
         n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635,
         n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643,
         n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651,
         n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659,
         n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667,
         n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675,
         n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683,
         n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691,
         n26692, n26693, n26694, n26695, n26696, n26697, n26698, n26699,
         n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707,
         n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715,
         n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723,
         n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731,
         n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739,
         n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747,
         n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755,
         n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763,
         n26764, n26765, n26766, n26767, n26768, n26769, n26770, n26771,
         n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779,
         n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787,
         n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795,
         n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803,
         n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811,
         n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819,
         n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827,
         n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835,
         n26836, n26837, n26838, n26839, n26840, n26841, n26842, n26843,
         n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851,
         n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859,
         n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867,
         n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875,
         n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883,
         n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891,
         n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899,
         n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907,
         n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915,
         n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923,
         n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931,
         n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939,
         n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947,
         n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955,
         n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963,
         n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971,
         n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979,
         n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987,
         n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995,
         n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003,
         n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011,
         n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019,
         n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027,
         n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035,
         n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043,
         n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051,
         n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059,
         n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067,
         n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075,
         n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083,
         n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091,
         n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099,
         n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107,
         n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115,
         n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123,
         n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131,
         n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139,
         n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147,
         n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155,
         n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163,
         n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171,
         n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179,
         n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187,
         n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195,
         n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203,
         n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211,
         n27212, n27213, n27214, n27215, n27216, n27217, n27218, n27219,
         n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227,
         n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235,
         n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243,
         n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251,
         n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259,
         n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267,
         n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275,
         n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283,
         n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291,
         n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299,
         n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307,
         n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315,
         n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323,
         n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331,
         n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339,
         n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347,
         n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355,
         n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363,
         n27364, n27365, n27366, n27367, n27368, n27369, n27370, n27371,
         n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379,
         n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387,
         n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395,
         n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403,
         n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411,
         n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419,
         n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427,
         n27428, n27429, n27430, n27431, n27432, n27433, n27434, n27435,
         n27436, n27437, n27438, n27439, n27440, n27441, n27442, n27443,
         n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451,
         n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459,
         n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467,
         n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475,
         n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483,
         n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491,
         n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499,
         n27500, n27501, n27502, n27503, n27504, n27505, n27506, n27507,
         n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515,
         n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523,
         n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531,
         n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539,
         n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547,
         n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555,
         n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563,
         n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571,
         n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579,
         n27580, n27581, n27582, n27583, n27584, n27585, n27586, n27587,
         n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595,
         n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603,
         n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611,
         n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619,
         n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627,
         n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635,
         n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643,
         n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651,
         n27652, n27653, n27654, n27655, n27656, n27657, n27658, n27659,
         n27660, n27661, n27662, n27663, n27664, n27665, n27666, n27667,
         n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675,
         n27676, n27677, n27678, n27679, n27680, n27681, n27682, n27683,
         n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691,
         n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699,
         n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707,
         n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715,
         n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723,
         n27724, n27725, n27726, n27727, n27728, n27729, n27730, n27731,
         n27732, n27733, n27734, n27735, n27736, n27737, n27738, n27739,
         n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747,
         n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755,
         n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763,
         n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771,
         n27772, n27773, n27774, n27775, n27776, n27777, n27778, n27779,
         n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787,
         n27788, n27789, n27790, n27791, n27792, n27793, n27794, n27795,
         n27796, n27797, n27798, n27799, n27800, n27801, n27802, n27803,
         n27804, n27805, n27806, n27807, n27808, n27809, n27810, n27811,
         n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819,
         n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827,
         n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835,
         n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843,
         n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851,
         n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859,
         n27860, n27861, n27862, n27863, n27864, n27865, n27866, n27867,
         n27868, n27869, n27870, n27871, n27872, n27873, n27874, n27875,
         n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883,
         n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891,
         n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899,
         n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907,
         n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915,
         n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923,
         n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931,
         n27932, n27933, n27934, n27935, n27936, n27937, n27938, n27939,
         n27940, n27941, n27942, n27943, n27944, n27945, n27946, n27947,
         n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955,
         n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963,
         n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971,
         n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979,
         n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987,
         n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995,
         n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003,
         n28004, n28005, n28006, n28007, n28008, n28009, n28010, n28011,
         n28012, n28013, n28014, n28015, n28016, n28017, n28018, n28019,
         n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027,
         n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035,
         n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043,
         n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051,
         n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059,
         n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067,
         n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075,
         n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083,
         n28084, n28085, n28086, n28087, n28088, n28089, n28090, n28091,
         n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099,
         n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107,
         n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115,
         n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123,
         n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131,
         n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139,
         n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147,
         n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155,
         n28156, n28157, n28158, n28159, n28160, n28161, n28162, n28163,
         n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171,
         n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179,
         n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187,
         n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195,
         n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203,
         n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211,
         n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219,
         n28220, n28221, n28222, n28223, n28224, n28225, n28226, n28227,
         n28228, n28229, n28230, n28231, n28232, n28233, n28234, n28235,
         n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243,
         n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251,
         n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259,
         n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267,
         n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275,
         n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283,
         n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291,
         n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299,
         n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307,
         n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315,
         n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323,
         n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331,
         n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339,
         n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347,
         n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355,
         n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363,
         n28364, n28365, n28366, n28367, n28368, n28369, n28370, n28371,
         n28372, n28373, n28374, n28375, n28376, n28377, n28378, n28379,
         n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387,
         n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395,
         n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403,
         n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411,
         n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419,
         n28420, n28421, n28422, n28423, n28424, n28425, n28426, n28427,
         n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435,
         n28436, n28437, n28438, n28439, n28440, n28441, n28442, n28443,
         n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451,
         n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459,
         n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467,
         n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475,
         n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483,
         n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491,
         n28492, n28493, n28494, n28495, n28496, n28497, n28498, n28499,
         n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507,
         n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515,
         n28516, n28517, n28518, n28519, n28520, n28521, n28522, n28523,
         n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531,
         n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539,
         n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547,
         n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555,
         n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563,
         n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571,
         n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579,
         n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587,
         n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595,
         n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603,
         n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611,
         n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619,
         n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627,
         n28628, n28629, n28630, n28631, n28632, n28633, n28634, n28635,
         n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643,
         n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651,
         n28652, n28653, n28654, n28655, n28656, n28657, n28658, n28659,
         n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667,
         n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675,
         n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683,
         n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691,
         n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699,
         n28700, n28701, n28702, n28703, n28704, n28705, n28706, n28707,
         n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715,
         n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723,
         n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731,
         n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28739,
         n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747,
         n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755,
         n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763,
         n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771,
         n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779,
         n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787,
         n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795,
         n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803,
         n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811,
         n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819,
         n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827,
         n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835,
         n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843,
         n28844, n28845, n28846, n28847, n28848, n28849, n28850, n28851,
         n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859,
         n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867,
         n28868, n28869, n28870, n28871, n28872, n28873, n28874, n28875,
         n28876, n28877, n28878, n28879, n28880, n28881, n28882, n28883,
         n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891,
         n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899,
         n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907,
         n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915,
         n28916, n28917, n28918, n28919, n28920, n28921, n28922, n28923,
         n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931,
         n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939,
         n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947,
         n28948, n28949, n28950, n28951, n28952, n28953, n28954, n28955,
         n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963,
         n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971,
         n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979,
         n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987,
         n28988, n28989, n28990, n28991, n28992, n28993, n28994, n28995,
         n28996, n28997, n28998, n28999, n29000, n29001, n29002, n29003,
         n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011,
         n29012, n29013, n29014, n29015, n29016, n29017, n29018, n29019,
         n29020, n29021, n29022, n29023, n29024, n29025, n29026, n29027,
         n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035,
         n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043,
         n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051,
         n29052, n29053, n29054, n29055, n29056, n29057, n29058, n29059,
         n29060, n29061, n29062, n29063, n29064, n29065, n29066, n29067,
         n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075,
         n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083,
         n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091,
         n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099,
         n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107,
         n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115,
         n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123,
         n29124, n29125, n29126, n29127, n29128, n29129, n29130, n29131,
         n29132, n29133, n29134, n29135, n29136, n29137, n29138, n29139,
         n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147,
         n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155,
         n29156, n29157, n29158, n29159, n29160, n29161, n29162, n29163,
         n29164, n29165, n29166, n29167, n29168, n29169, n29170, n29171,
         n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179,
         n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187,
         n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195,
         n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203,
         n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211,
         n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219,
         n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227,
         n29228, n29229, n29230, n29231, n29232, n29233, n29234, n29235,
         n29236, n29237, n29238, n29239, n29240, n29241, n29242, n29243,
         n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251,
         n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259,
         n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267,
         n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275,
         n29276, n29277, n29278, n29279, n29280, n29281, n29282, n29283,
         n29284, n29285, n29286, n29287, n29288, n29289, n29290, n29291,
         n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299,
         n29300, n29301, n29302, n29303, n29304, n29305, n29306, n29307,
         n29308, n29309, n29310, n29311, n29312, n29313, n29314, n29315,
         n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323,
         n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331,
         n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339,
         n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347,
         n29348, n29349, n29350, n29351, n29352, n29353, n29354, n29355,
         n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363,
         n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371,
         n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379,
         n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387,
         n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395,
         n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403,
         n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411,
         n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29419,
         n29420, n29421, n29422, n29423, n29424, n29425, n29426, n29427,
         n29428, n29429, n29430, n29431, n29432, n29433, n29434, n29435,
         n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443,
         n29444, n29445, n29446, n29447, n29448, n29449, n29450, n29451,
         n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459,
         n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467,
         n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475,
         n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483,
         n29484, n29485, n29486, n29487, n29488, n29489, n29490, n29491,
         n29492, n29493, n29494, n29495, n29496, n29497, n29498, n29499,
         n29500, n29501, n29502, n29503, n29504, n29505, n29506, n29507,
         n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515,
         n29516, n29517, n29518, n29519, n29520, n29521, n29522, n29523,
         n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531,
         n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539,
         n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547,
         n29548, n29549, n29550, n29551, n29552, n29553, n29554, n29555,
         n29556, n29557, n29558, n29559, n29560, n29561, n29562, n29563,
         n29564, n29565, n29566, n29567, n29568, n29569, n29570, n29571,
         n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29579,
         n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587,
         n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595,
         n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603,
         n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611,
         n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619,
         n29620, n29621, n29622, n29623, n29624, n29625, n29626, n29627,
         n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635,
         n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643,
         n29644, n29645, n29646, n29647, n29648, n29649, n29650, n29651,
         n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659,
         n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667,
         n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675,
         n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683,
         n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691,
         n29692, n29693, n29694, n29695, n29696, n29697, n29698, n29699,
         n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707,
         n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715,
         n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723,
         n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731,
         n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739,
         n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747,
         n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755,
         n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763,
         n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771,
         n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779,
         n29780, n29781, n29782, n29783, n29784, n29785, n29786, n29787,
         n29788, n29789, n29790, n29791, n29792, n29793, n29794, n29795,
         n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803,
         n29804, n29805, n29806, n29807, n29808, n29809, n29810, n29811,
         n29812, n29813, n29814, n29815, n29816, n29817, n29818, n29819,
         n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827,
         n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835,
         n29836, n29837, n29838, n29839, n29840, n29841, n29842, n29843,
         n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851,
         n29852, n29853, n29854, n29855, n29856, n29857, n29858, n29859,
         n29860, n29861, n29862, n29863, n29864, n29865, n29866, n29867,
         n29868, n29869, n29870, n29871, n29872, n29873, n29874, n29875,
         n29876, n29877, n29878, n29879, n29880, n29881, n29882, n29883,
         n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891,
         n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899,
         n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907,
         n29908, n29909, n29910, n29911, n29912, n29913, n29914, n29915,
         n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923,
         n29924, n29925, n29926, n29927, n29928, n29929, n29930, n29931,
         n29932, n29933, n29934, n29935, n29936, n29937, n29938, n29939,
         n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947,
         n29948, n29949, n29950, n29951, n29952, n29953, n29954, n29955,
         n29956, n29957, n29958, n29959, n29960, n29961, n29962, n29963,
         n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971,
         n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979,
         n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987,
         n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995,
         n29996, n29997, n29998, n29999, n30000, n30001, n30002, n30003,
         n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011,
         n30012, n30013, n30014, n30015, n30016, n30017, n30018, n30019,
         n30020, n30021, n30022, n30023, n30024, n30025, n30026, n30027,
         n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035,
         n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043,
         n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051,
         n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059,
         n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067,
         n30068, n30069, n30070, n30071, n30072, n30073, n30074, n30075,
         n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083,
         n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091,
         n30092, n30093, n30094, n30095, n30096, n30097, n30098, n30099,
         n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107,
         n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115,
         n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123,
         n30124, n30125, n30126, n30127, n30128, n30129, n30130, n30131,
         n30132, n30133, n30134, n30135, n30136, n30137, n30138, n30139,
         n30140, n30141, n30142, n30143, n30144, n30145, n30146, n30147,
         n30148, n30149, n30150, n30151, n30152, n30153, n30154, n30155,
         n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163,
         n30164, n30165, n30166, n30167, n30168, n30169, n30170, n30171,
         n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179,
         n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187,
         n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195,
         n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203,
         n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211,
         n30212, n30213, n30214, n30215, n30216, n30217, n30218, n30219,
         n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227,
         n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235,
         n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243,
         n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251,
         n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259,
         n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267,
         n30268, n30269, n30270, n30271, n30272, n30273, n30274, n30275,
         n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283,
         n30284, n30285, n30286, n30287, n30288, n30289, n30290, n30291,
         n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299,
         n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307,
         n30308, n30309, n30310, n30311, n30312, n30313, n30314, n30315,
         n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323,
         n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331,
         n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339,
         n30340, n30341, n30342, n30343, n30344, n30345, n30346, n30347,
         n30348, n30349, n30350, n30351, n30352, n30353, n30354, n30355,
         n30356, n30357, n30358, n30359, n30360, n30361, n30362, n30363,
         n30364, n30365, n30366, n30367, n30368, n30369, n30370, n30371,
         n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379,
         n30380, n30381, n30382, n30383, n30384, n30385, n30386, n30387,
         n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395,
         n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403,
         n30404, n30405, n30406, n30407, n30408, n30409, n30410, n30411,
         n30412, n30413, n30414, n30415, n30416, n30417, n30418, n30419,
         n30420, n30421, n30422, n30423, n30424, n30425, n30426, n30427,
         n30428, n30429, n30430, n30431, n30432, n30433, n30434, n30435,
         n30436, n30437, n30438, n30439, n30440, n30441, n30442, n30443,
         n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451,
         n30452, n30453, n30454, n30455, n30456, n30457, n30458, n30459,
         n30460, n30461, n30462, n30463, n30464, n30465, n30466, n30467,
         n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475,
         n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483,
         n30484, n30485, n30486, n30487, n30488, n30489, n30490, n30491,
         n30492, n30493, n30494, n30495, n30496, n30497, n30498, n30499,
         n30500, n30501, n30502, n30503, n30504, n30505, n30506, n30507,
         n30508, n30509, n30510, n30511, n30512, n30513, n30514, n30515,
         n30516, n30517, n30518, n30519, n30520, n30521, n30522, n30523,
         n30524, n30525, n30526, n30527, n30528, n30529, n30530, n30531,
         n30532, n30533, n30534, n30535, n30536, n30537, n30538, n30539,
         n30540, n30541, n30542, n30543, n30544, n30545, n30546, n30547,
         n30548, n30549, n30550, n30551, n30552, n30553, n30554, n30555,
         n30556, n30557, n30558, n30559, n30560, n30561, n30562, n30563,
         n30564, n30565, n30566, n30567, n30568, n30569, n30570, n30571,
         n30572, n30573, n30574, n30575, n30576, n30577, n30578, n30579,
         n30580, n30581, n30582, n30583, n30584, n30585, n30586, n30587,
         n30588, n30589, n30590, n30591, n30592, n30593, n30594, n30595,
         n30596, n30597, n30598, n30599, n30600, n30601, n30602, n30603,
         n30604, n30605, n30606, n30607, n30608, n30609, n30610, n30611,
         n30612, n30613, n30614, n30615, n30616, n30617, n30618, n30619,
         n30620, n30621, n30622, n30623, n30624, n30625, n30626, n30627,
         n30628, n30629, n30630, n30631, n30632, n30633, n30634, n30635,
         n30636, n30637, n30638, n30639, n30640, n30641, n30642, n30643,
         n30644, n30645, n30646, n30647, n30648, n30649, n30650, n30651,
         n30652, n30653, n30654, n30655, n30656, n30657, n30658, n30659,
         n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667,
         n30668, n30669, n30670, n30671, n30672, n30673, n30674, n30675,
         n30676, n30677, n30678, n30679, n30680, n30681, n30682, n30683,
         n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691,
         n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699,
         n30700, n30701, n30702, n30703, n30704, n30705, n30706, n30707,
         n30708, n30709, n30710, n30711, n30712, n30713, n30714, n30715,
         n30716, n30717, n30718, n30719, n30720, n30721, n30722, n30723,
         n30724, n30725, n30726, n30727, n30728, n30729, n30730, n30731,
         n30732, n30733, n30734, n30735, n30736, n30737, n30738, n30739,
         n30740, n30741, n30742, n30743, n30744, n30745, n30746, n30747,
         n30748, n30749, n30750, n30751, n30752, n30753, n30754, n30755,
         n30756, n30757, n30758, n30759, n30760, n30761, n30762, n30763,
         n30764, n30765, n30766, n30767, n30768, n30769, n30770, n30771,
         n30772, n30773, n30774, n30775, n30776, n30777, n30778, n30779,
         n30780, n30781, n30782, n30783, n30784, n30785, n30786, n30787,
         n30788, n30789, n30790, n30791, n30792, n30793, n30794, n30795,
         n30796, n30797, n30798, n30799, n30800, n30801, n30802, n30803,
         n30804, n30805, n30806, n30807, n30808, n30809, n30810, n30811,
         n30812, n30813, n30814, n30815, n30816, n30817, n30818, n30819,
         n30820, n30821, n30822, n30823, n30824, n30825, n30826, n30827,
         n30828, n30829, n30830, n30831, n30832, n30833, n30834, n30835,
         n30836, n30837, n30838, n30839, n30840, n30841, n30842, n30843,
         n30844, n30845, n30846, n30847, n30848, n30849, n30850, n30851,
         n30852, n30853, n30854, n30855, n30856, n30857, n30858, n30859,
         n30860, n30861, n30862, n30863, n30864, n30865, n30866, n30867,
         n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30875,
         n30876, n30877, n30878, n30879, n30880, n30881, n30882, n30883,
         n30884, n30885, n30886, n30887, n30888, n30889, n30890, n30891,
         n30892, n30893, n30894, n30895, n30896, n30897, n30898, n30899,
         n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907,
         n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915,
         n30916, n30917, n30918, n30919, n30920, n30921, n30922, n30923,
         n30924, n30925, n30926, n30927, n30928, n30929, n30930, n30931,
         n30932, n30933, n30934, n30935, n30936, n30937, n30938, n30939,
         n30940, n30941, n30942, n30943, n30944, n30945, n30946, n30947,
         n30948, n30949, n30950, n30951, n30952, n30953, n30954, n30955,
         n30956, n30957, n30958, n30959, n30960, n30961, n30962, n30963,
         n30964, n30965, n30966, n30967, n30968, n30969, n30970, n30971,
         n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979,
         n30980, n30981, n30982, n30983, n30984, n30985, n30986, n30987,
         n30988, n30989, n30990, n30991, n30992, n30993, n30994, n30995,
         n30996, n30997, n30998, n30999, n31000, n31001, n31002, n31003,
         n31004, n31005, n31006, n31007, n31008, n31009, n31010, n31011,
         n31012, n31013, n31014, n31015, n31016, n31017, n31018, n31019,
         n31020, n31021, n31022, n31023, n31024, n31025, n31026, n31027,
         n31028, n31029, n31030, n31031, n31032, n31033, n31034, n31035,
         n31036, n31037, n31038, n31039, n31040, n31041, n31042, n31043,
         n31044, n31045, n31046, n31047, n31048, n31049, n31050, n31051,
         n31052, n31053, n31054, n31055, n31056, n31057, n31058, n31059,
         n31060, n31061, n31062, n31063, n31064, n31065, n31066, n31067,
         n31068, n31069, n31070, n31071, n31072, n31073, n31074, n31075,
         n31076, n31077, n31078, n31079, n31080, n31081, n31082, n31083,
         n31084, n31085, n31086, n31087, n31088, n31089, n31090, n31091,
         n31092, n31093, n31094, n31095, n31096, n31097, n31098, n31099,
         n31100, n31101, n31102, n31103, n31104, n31105, n31106, n31107,
         n31108, n31109, n31110, n31111, n31112, n31113, n31114, n31115,
         n31116, n31117, n31118, n31119, n31120, n31121, n31122, n31123,
         n31124, n31125, n31126, n31127, n31128, n31129, n31130, n31131,
         n31132, n31133, n31134, n31135, n31136, n31137, n31138, n31139,
         n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147,
         n31148, n31149, n31150, n31151, n31152, n31153, n31154, n31155,
         n31156, n31157, n31158, n31159, n31160, n31161, n31162, n31163,
         n31164, n31165, n31166, n31167, n31168, n31169, n31170, n31171,
         n31172, n31173, n31174, n31175, n31176, n31177, n31178, n31179,
         n31180, n31181, n31182, n31183, n31184, n31185, n31186, n31187,
         n31188, n31189, n31190, n31191, n31192, n31193, n31194, n31195,
         n31196, n31197, n31198, n31199, n31200, n31201, n31202, n31203,
         n31204, n31205, n31206, n31207, n31208, n31209, n31210, n31211,
         n31212, n31213, n31214, n31215, n31216, n31217, n31218, n31219,
         n31220, n31221, n31222, n31223, n31224, n31225, n31226, n31227,
         n31228, n31229, n31230, n31231, n31232, n31233, n31234, n31235,
         n31236, n31237, n31238, n31239, n31240, n31241, n31242, n31243,
         n31244, n31245, n31246, n31247, n31248, n31249, n31250, n31251,
         n31252, n31253, n31254, n31255, n31256, n31257, n31258, n31259,
         n31260, n31261, n31262, n31263, n31264, n31265, n31266, n31267,
         n31268, n31269, n31270, n31271, n31272, n31273, n31274, n31275,
         n31276, n31277, n31278, n31279, n31280, n31281, n31282, n31283,
         n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291,
         n31292, n31293, n31294, n31295, n31296, n31297, n31298, n31299,
         n31300, n31301, n31302, n31303, n31304, n31305, n31306, n31307,
         n31308, n31309, n31310, n31311, n31312, n31313, n31314, n31315,
         n31316, n31317, n31318, n31319, n31320, n31321, n31322, n31323,
         n31324, n31325, n31326, n31327, n31328, n31329, n31330, n31331,
         n31332, n31333, n31334, n31335, n31336, n31337, n31338, n31339,
         n31340, n31341, n31342, n31343, n31344, n31345, n31346, n31347,
         n31348, n31349, n31350, n31351, n31352, n31353, n31354, n31355,
         n31356, n31357, n31358, n31359, n31360, n31361, n31362, n31363,
         n31364, n31365, n31366, n31367, n31368, n31369, n31370, n31371,
         n31372, n31373, n31374, n31375, n31376, n31377, n31378, n31379,
         n31380, n31381, n31382, n31383, n31384, n31385, n31386, n31387,
         n31388, n31389, n31390, n31391, n31392, n31393, n31394, n31395,
         n31396, n31397, n31398, n31399, n31400, n31401, n31402, n31403,
         n31404, n31405, n31406, n31407, n31408, n31409, n31410, n31411,
         n31412, n31413, n31414, n31415, n31416, n31417, n31418, n31419,
         n31420, n31421, n31422, n31423, n31424, n31425, n31426, n31427,
         n31428, n31429, n31430, n31431, n31432, n31433, n31434, n31435,
         n31436, n31437, n31438, n31439, n31440, n31441, n31442, n31443,
         n31444, n31445, n31446, n31447, n31448, n31449, n31450, n31451,
         n31452, n31453, n31454, n31455, n31456, n31457, n31458, n31459,
         n31460, n31461, n31462, n31463, n31464, n31465, n31466, n31467,
         n31468, n31469, n31470, n31471, n31472, n31473, n31474, n31475,
         n31476, n31477, n31478, n31479, n31480, n31481, n31482, n31483,
         n31484, n31485, n31486, n31487, n31488, n31489, n31490, n31491,
         n31492, n31493, n31494, n31495, n31496, n31497, n31498, n31499,
         n31500, n31501, n31502, n31503, n31504, n31505, n31506, n31507,
         n31508, n31509, n31510, n31511, n31512, n31513, n31514, n31515,
         n31516, n31517, n31518, n31519, n31520, n31521, n31522, n31523,
         n31524, n31525, n31526, n31527, n31528, n31529, n31530, n31531,
         n31532, n31533, n31534, n31535, n31536, n31537, n31538, n31539,
         n31540, n31541, n31542, n31543, n31544, n31545, n31546, n31547,
         n31548, n31549, n31550, n31551, n31552, n31553, n31554, n31555,
         n31556, n31557, n31558, n31559, n31560, n31561, n31562, n31563,
         n31564, n31565, n31566, n31567, n31568, n31569, n31570, n31571,
         n31572, n31573, n31574, n31575, n31576, n31577, n31578, n31579,
         n31580, n31581, n31582, n31583, n31584, n31585, n31586, n31587,
         n31588, n31589, n31590, n31591, n31592, n31593, n31594, n31595,
         n31596, n31597, n31598, n31599, n31600, n31601, n31602, n31603,
         n31604, n31605, n31606, n31607, n31608, n31609, n31610, n31611,
         n31612, n31613, n31614, n31615, n31616, n31617, n31618, n31619,
         n31620, n31621, n31622, n31623, n31624, n31625, n31626, n31627,
         n31628, n31629, n31630, n31631, n31632, n31633, n31634, n31635,
         n31636, n31637, n31638, n31639, n31640, n31641, n31642, n31643,
         n31644, n31645, n31646, n31647, n31648, n31649, n31650, n31651,
         n31652, n31653, n31654, n31655, n31656, n31657, n31658, n31659,
         n31660, n31661, n31662, n31663, n31664, n31665, n31666, n31667,
         n31668, n31669, n31670, n31671, n31672, n31673, n31674, n31675,
         n31676, n31677, n31678, n31679, n31680, n31681, n31682, n31683,
         n31684, n31685, n31686, n31687, n31688, n31689, n31690, n31691,
         n31692, n31693, n31694, n31695, n31696, n31697, n31698, n31699,
         n31700, n31701, n31702, n31703, n31704, n31705, n31706, n31707,
         n31708, n31709, n31710, n31711, n31712, n31713, n31714, n31715,
         n31716, n31717, n31718, n31719, n31720, n31721, n31722, n31723,
         n31724, n31725, n31726, n31727, n31728, n31729, n31730, n31731,
         n31732, n31733, n31734, n31735, n31736, n31737, n31738, n31739,
         n31740, n31741, n31742, n31743, n31744, n31745, n31746, n31747,
         n31748, n31749, n31750, n31751, n31752, n31753, n31754, n31755,
         n31756, n31757, n31758, n31759, n31760, n31761, n31762, n31763,
         n31764, n31765, n31766, n31767, n31768, n31769, n31770, n31771,
         n31772, n31773, n31774, n31775, n31776, n31777, n31778, n31779,
         n31780, n31781, n31782, n31783, n31784, n31785, n31786, n31787,
         n31788, n31789, n31790, n31791, n31792, n31793, n31794, n31795,
         n31796, n31797, n31798, n31799, n31800, n31801, n31802, n31803,
         n31804, n31805, n31806, n31807, n31808, n31809, n31810, n31811,
         n31812, n31813, n31814, n31815, n31816, n31817, n31818, n31819,
         n31820, n31821, n31822, n31823, n31824, n31825, n31826, n31827,
         n31828, n31829, n31830, n31831, n31832, n31833, n31834, n31835,
         n31836, n31837, n31838, n31839, n31840, n31841, n31842, n31843,
         n31844, n31845, n31846, n31847, n31848, n31849, n31850, n31851,
         n31852, n31853, n31854, n31855, n31856, n31857, n31858, n31859,
         n31860, n31861, n31862, n31863, n31864, n31865, n31866, n31867,
         n31868, n31869, n31870, n31871, n31872, n31873, n31874, n31875,
         n31876, n31877, n31878, n31879, n31880, n31881, n31882, n31883,
         n31884, n31885, n31886, n31887, n31888, n31889, n31890, n31891,
         n31892, n31893, n31894, n31895, n31896, n31897, n31898, n31899,
         n31900, n31901, n31902, n31903, n31904, n31905, n31906, n31907,
         n31908, n31909, n31910, n31911, n31912, n31913, n31914, n31915,
         n31916, n31917, n31918, n31919, n31920, n31921, n31922, n31923,
         n31924, n31925, n31926, n31927, n31928, n31929, n31930, n31931,
         n31932, n31933, n31934, n31935, n31936, n31937, n31938, n31939,
         n31940, n31941, n31942, n31943, n31944, n31945, n31946, n31947,
         n31948, n31949, n31950, n31951, n31952, n31953, n31954, n31955,
         n31956, n31957, n31958, n31959, n31960, n31961, n31962, n31963,
         n31964, n31965, n31966, n31967, n31968, n31969, n31970, n31971,
         n31972, n31973, n31974, n31975, n31976, n31977, n31978, n31979,
         n31980, n31981, n31982, n31983, n31984, n31985, n31986, n31987,
         n31988, n31989, n31990, n31991, n31992, n31993, n31994, n31995,
         n31996, n31997, n31998, n31999, n32000, n32001, n32002, n32003,
         n32004, n32005, n32006, n32007, n32008, n32009, n32010, n32011,
         n32012, n32013, n32014, n32015, n32016, n32017, n32018, n32019,
         n32020, n32021, n32022, n32023, n32024, n32025, n32026, n32027,
         n32028, n32029, n32030, n32031, n32032, n32033, n32034, n32035,
         n32036, n32037, n32038, n32039, n32040, n32041, n32042, n32043,
         n32044, n32045, n32046, n32047, n32048, n32049, n32050, n32051,
         n32052, n32053, n32054, n32055, n32056, n32057, n32058, n32059,
         n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067,
         n32068, n32069, n32070, n32071, n32072, n32073, n32074, n32075,
         n32076, n32077, n32078, n32079, n32080, n32081, n32082, n32083,
         n32084, n32085, n32086, n32087, n32088, n32089, n32090, n32091,
         n32092, n32093, n32094, n32095, n32096, n32097, n32098, n32099,
         n32100, n32101, n32102, n32103, n32104, n32105, n32106, n32107,
         n32108, n32109, n32110, n32111, n32112, n32113, n32114, n32115,
         n32116, n32117, n32118, n32119, n32120, n32121, n32122, n32123,
         n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131,
         n32132, n32133, n32134, n32135, n32136, n32137, n32138, n32139,
         n32140, n32141, n32142, n32143, n32144, n32145, n32146, n32147,
         n32148, n32149, n32150, n32151, n32152, n32153, n32154, n32155,
         n32156, n32157, n32158, n32159, n32160, n32161, n32162, n32163,
         n32164, n32165, n32166, n32167, n32168, n32169, n32170, n32171,
         n32172, n32173, n32174, n32175, n32176, n32177, n32178, n32179,
         n32180, n32181, n32182, n32183, n32184, n32185, n32186, n32187,
         n32188, n32189, n32190, n32191, n32192, n32193, n32194, n32195,
         n32196, n32197, n32198, n32199, n32200, n32201, n32202, n32203,
         n32204, n32205, n32206, n32207, n32208, n32209, n32210, n32211,
         n32212, n32213, n32214, n32215, n32216, n32217, n32218, n32219,
         n32220, n32221, n32222, n32223, n32224, n32225, n32226, n32227,
         n32228, n32229, n32230, n32231, n32232, n32233, n32234, n32235,
         n32236, n32237, n32238, n32239, n32240, n32241, n32242, n32243,
         n32244, n32245, n32246, n32247, n32248, n32249, n32250, n32251,
         n32252, n32253, n32254, n32255, n32256, n32257, n32258, n32259,
         n32260, n32261, n32262, n32263, n32264, n32265, n32266, n32267,
         n32268, n32269, n32270, n32271, n32272, n32273, n32274, n32275,
         n32276, n32277, n32278, n32279, n32280, n32281, n32282, n32283,
         n32284, n32285, n32286, n32287, n32288, n32289, n32290, n32291,
         n32292, n32293, n32294, n32295, n32296, n32297, n32298, n32299,
         n32300, n32301, n32302, n32303, n32304, n32305, n32306, n32307,
         n32308, n32309, n32310, n32311, n32312, n32313, n32314, n32315,
         n32316, n32317, n32318, n32319, n32320, n32321, n32322, n32323,
         n32324, n32325, n32326, n32327, n32328, n32329, n32330, n32331,
         n32332, n32333, n32334, n32335, n32336, n32337, n32338, n32339,
         n32340, n32341, n32342, n32343, n32344, n32345, n32346, n32347,
         n32348, n32349, n32350, n32351, n32352, n32353, n32354, n32355,
         n32356, n32357, n32358, n32359, n32360, n32361, n32362, n32363,
         n32364, n32365, n32366, n32367, n32368, n32369, n32370, n32371,
         n32372, n32373, n32374, n32375, n32376, n32377, n32378, n32379,
         n32380, n32381, n32382, n32383, n32384, n32385, n32386, n32387,
         n32388, n32389, n32390, n32391, n32392, n32393, n32394, n32395,
         n32396, n32397, n32398, n32399, n32400, n32401, n32402, n32403,
         n32404, n32405, n32406, n32407, n32408, n32409, n32410, n32411,
         n32412, n32413, n32414, n32415, n32416, n32417, n32418, n32419,
         n32420, n32421, n32422, n32423, n32424, n32425, n32426, n32427,
         n32428, n32429, n32430, n32431, n32432, n32433, n32434, n32435,
         n32436, n32437, n32438, n32439, n32440, n32441, n32442, n32443,
         n32444, n32445, n32446, n32447, n32448, n32449, n32450, n32451,
         n32452, n32453, n32454, n32455, n32456, n32457, n32458, n32459,
         n32460, n32461, n32462, n32463, n32464, n32465, n32466, n32467,
         n32468, n32469, n32470, n32471, n32472, n32473, n32474, n32475,
         n32476, n32477, n32478, n32479, n32480, n32481, n32482, n32483,
         n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491,
         n32492, n32493, n32494, n32495, n32496, n32497, n32498, n32499,
         n32500, n32501, n32502, n32503, n32504, n32505, n32506, n32507,
         n32508, n32509, n32510, n32511, n32512, n32513, n32514, n32515,
         n32516, n32517, n32518, n32519, n32520, n32521, n32522, n32523,
         n32524, n32525, n32526, n32527, n32528, n32529, n32530, n32531,
         n32532, n32533, n32534, n32535, n32536, n32537, n32538, n32539,
         n32540, n32541, n32542, n32543, n32544, n32545, n32546, n32547,
         n32548, n32549, n32550, n32551, n32552, n32553, n32554, n32555,
         n32556, n32557, n32558, n32559, n32560, n32561, n32562, n32563,
         n32564, n32565, n32566, n32567, n32568, n32569, n32570, n32571,
         n32572, n32573, n32574, n32575, n32576, n32577, n32578, n32579,
         n32580, n32581, n32582, n32583, n32584, n32585, n32586, n32587,
         n32588, n32589, n32590, n32591, n32592, n32593, n32594, n32595,
         n32596, n32597, n32598, n32599, n32600, n32601, n32602, n32603,
         n32604, n32605, n32606, n32607, n32608, n32609, n32610, n32611,
         n32612, n32613, n32614, n32615, n32616, n32617, n32618, n32619,
         n32620, n32621, n32622, n32623, n32624, n32625, n32626, n32627,
         n32628, n32629, n32630, n32631, n32632, n32633, n32634, n32635,
         n32636, n32637, n32638, n32639, n32640, n32641, n32642, n32643,
         n32644, n32645, n32646, n32647, n32648, n32649, n32650, n32651,
         n32652, n32653, n32654, n32655, n32656, n32657, n32658, n32659,
         n32660, n32661, n32662, n32663, n32664, n32665, n32666, n32667,
         n32668, n32669, n32670, n32671, n32672, n32673, n32674, n32675,
         n32676, n32677, n32678, n32679, n32680, n32681, n32682, n32683,
         n32684, n32685, n32686, n32687, n32688, n32689, n32690, n32691,
         n32692, n32693, n32694, n32695, n32696, n32697, n32698, n32699,
         n32700, n32701, n32702, n32703, n32704, n32705, n32706, n32707,
         n32708, n32709, n32710, n32711, n32712, n32713, n32714, n32715,
         n32716, n32717, n32718, n32719, n32720, n32721, n32722, n32723,
         n32724, n32725, n32726, n32727, n32728, n32729, n32730, n32731,
         n32732, n32733, n32734, n32735, n32736, n32737, n32738, n32739,
         n32740, n32741, n32742, n32743, n32744, n32745, n32746, n32747,
         n32748, n32749, n32750, n32751, n32752, n32753, n32754, n32755,
         n32756, n32757, n32758, n32759, n32760, n32761, n32762, n32763,
         n32764, n32765, n32766, n32767, n32768, n32769, n32770, n32771,
         n32772, n32773, n32774, n32775, n32776, n32777, n32778, n32779,
         n32780, n32781, n32782, n32783, n32784, n32785, n32786, n32787,
         n32788, n32789, n32790, n32791, n32792, n32793, n32794, n32795,
         n32796, n32797, n32798, n32799, n32800, n32801, n32802, n32803,
         n32804, n32805, n32806, n32807, n32808, n32809, n32810, n32811,
         n32812, n32813, n32814, n32815, n32816, n32817, n32818, n32819,
         n32820, n32821, n32822, n32823, n32824, n32825, n32826, n32827,
         n32828, n32829, n32830, n32831, n32832, n32833, n32834, n32835,
         n32836, n32837, n32838, n32839, n32840, n32841, n32842, n32843,
         n32844, n32845, n32846, n32847, n32848, n32849, n32850, n32851,
         n32852, n32853, n32854, n32855, n32856, n32857, n32858, n32859,
         n32860, n32861, n32862, n32863, n32864, n32865, n32866, n32867,
         n32868, n32869, n32870, n32871, n32872, n32873, n32874, n32875,
         n32876, n32877, n32878, n32879, n32880, n32881, n32882, n32883,
         n32884, n32885, n32886, n32887, n32888, n32889, n32890, n32891,
         n32892, n32893, n32894, n32895, n32896, n32897, n32898, n32899,
         n32900, n32901, n32902, n32903, n32904, n32905, n32906, n32907,
         n32908, n32909, n32910, n32911, n32912, n32913, n32914, n32915,
         n32916, n32917, n32918, n32919, n32920, n32921, n32922, n32923,
         n32924, n32925, n32926, n32927, n32928, n32929, n32930, n32931,
         n32932, n32933, n32934, n32935, n32936, n32937, n32938, n32939,
         n32940, n32941, n32942, n32943, n32944, n32945, n32946, n32947,
         n32948, n32949, n32950, n32951, n32952, n32953, n32954, n32955,
         n32956, n32957, n32958, n32959, n32960, n32961, n32962, n32963,
         n32964, n32965, n32966, n32967, n32968, n32969, n32970, n32971,
         n32972, n32973, n32974, n32975, n32976, n32977, n32978, n32979,
         n32980, n32981, n32982, n32983, n32984, n32985, n32986, n32987,
         n32988, n32989, n32990, n32991, n32992, n32993, n32994, n32995,
         n32996, n32997, n32998, n32999, n33000, n33001, n33002, n33003,
         n33004, n33005, n33006, n33007, n33008, n33009, n33010, n33011,
         n33012, n33013, n33014, n33015, n33016, n33017, n33018, n33019,
         n33020, n33021, n33022, n33023, n33024, n33025, n33026, n33027,
         n33028, n33029, n33030, n33031, n33032, n33033, n33034, n33035,
         n33036, n33037, n33038, n33039, n33040, n33041, n33042, n33043,
         n33044, n33045, n33046, n33047, n33048, n33049, n33050, n33051,
         n33052, n33053, n33054, n33055, n33056, n33057, n33058, n33059,
         n33060, n33061, n33062, n33063, n33064, n33065, n33066, n33067,
         n33068, n33069, n33070, n33071, n33072, n33073, n33074, n33075,
         n33076, n33077, n33078, n33079, n33080, n33081, n33082, n33083,
         n33084, n33085, n33086, n33087, n33088, n33089, n33090, n33091,
         n33092, n33093, n33094, n33095, n33096, n33097, n33098, n33099,
         n33100, n33101, n33102, n33103, n33104, n33105, n33106, n33107,
         n33108, n33109, n33110, n33111, n33112, n33113, n33114, n33115,
         n33116, n33117, n33118, n33119, n33120, n33121, n33122, n33123,
         n33124, n33125, n33126, n33127, n33128, n33129, n33130, n33131,
         n33132, n33133, n33134, n33135, n33136, n33137, n33138, n33139,
         n33140, n33141, n33142, n33143, n33144, n33145, n33146, n33147,
         n33148, n33149, n33150, n33151, n33152, n33153, n33154, n33155,
         n33156, n33157, n33158, n33159, n33160, n33161, n33162, n33163,
         n33164, n33165, n33166, n33167, n33168, n33169, n33170, n33171,
         n33172, n33173, n33174, n33175, n33176, n33177, n33178, n33179,
         n33180, n33181, n33182, n33183, n33184, n33185, n33186, n33187,
         n33188, n33189, n33190, n33191, n33192, n33193, n33194, n33195,
         n33196, n33197, n33198, n33199, n33200, n33201, n33202, n33203,
         n33204, n33205, n33206, n33207, n33208, n33209, n33210, n33211,
         n33212, n33213, n33214, n33215, n33216, n33217, n33218, n33219,
         n33220, n33221, n33222, n33223, n33224, n33225, n33226, n33227,
         n33228, n33229, n33230, n33231, n33232, n33233, n33234, n33235,
         n33236, n33237, n33238, n33239, n33240, n33241, n33242, n33243,
         n33244, n33245, n33246, n33247, n33248, n33249, n33250, n33251,
         n33252, n33253, n33254, n33255, n33256, n33257, n33258, n33259,
         n33260, n33261, n33262, n33263, n33264, n33265, n33266, n33267,
         n33268, n33269, n33270, n33271, n33272, n33273, n33274, n33275,
         n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283,
         n33284, n33285, n33286, n33287, n33288, n33289, n33290, n33291,
         n33292, n33293, n33294, n33295, n33296, n33297, n33298, n33299,
         n33300, n33301, n33302, n33303, n33304, n33305, n33306, n33307,
         n33308, n33309, n33310, n33311, n33312, n33313, n33314, n33315,
         n33316, n33317, n33318, n33319, n33320, n33321, n33322, n33323,
         n33324, n33325, n33326, n33327, n33328, n33329, n33330, n33331,
         n33332, n33333, n33334, n33335, n33336, n33337, n33338, n33339,
         n33340, n33341, n33342, n33343, n33344, n33345, n33346, n33347,
         n33348, n33349, n33350, n33351, n33352, n33353, n33354, n33355,
         n33356, n33357, n33358, n33359, n33360, n33361, n33362, n33363,
         n33364, n33365, n33366, n33367, n33368, n33369, n33370, n33371,
         n33372, n33373, n33374, n33375, n33376, n33377, n33378, n33379,
         n33380, n33381, n33382, n33383, n33384, n33385, n33386, n33387,
         n33388, n33389, n33390, n33391, n33392, n33393, n33394, n33395,
         n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403,
         n33404, n33405, n33406, n33407, n33408, n33409, n33410, n33411,
         n33412, n33413, n33414, n33415, n33416, n33417, n33418, n33419,
         n33420, n33421, n33422, n33423, n33424, n33425, n33426, n33427,
         n33428, n33429, n33430, n33431, n33432, n33433, n33434, n33435,
         n33436, n33437, n33438, n33439, n33440, n33441, n33442, n33443,
         n33444, n33445, n33446, n33447, n33448, n33449, n33450, n33451,
         n33452, n33453, n33454, n33455, n33456, n33457, n33458, n33459,
         n33460, n33461, n33462, n33463, n33464, n33465, n33466, n33467,
         n33468, n33469, n33470, n33471, n33472, n33473, n33474, n33475,
         n33476, n33477, n33478, n33479, n33480, n33481, n33482, n33483,
         n33484, n33485, n33486, n33487, n33488, n33489, n33490, n33491,
         n33492, n33493, n33494, n33495, n33496, n33497, n33498, n33499,
         n33500, n33501, n33502, n33503, n33504, n33505, n33506, n33507,
         n33508, n33509, n33510, n33511, n33512, n33513, n33514, n33515,
         n33516, n33517, n33518, n33519, n33520, n33521, n33522, n33523,
         n33524, n33525, n33526, n33527, n33528, n33529, n33530, n33531,
         n33532, n33533, n33534, n33535, n33536, n33537, n33538, n33539,
         n33540, n33541, n33542, n33543, n33544, n33545, n33546, n33547,
         n33548, n33549, n33550, n33551, n33552, n33553, n33554, n33555,
         n33556, n33557, n33558, n33559, n33560, n33561, n33562, n33563,
         n33564, n33565, n33566, n33567, n33568, n33569, n33570, n33571,
         n33572, n33573, n33574, n33575, n33576, n33577, n33578, n33579,
         n33580, n33581, n33582, n33583, n33584, n33585, n33586, n33587,
         n33588, n33589, n33590, n33591, n33592, n33593, n33594, n33595,
         n33596, n33597, n33598, n33599, n33600, n33601, n33602, n33603,
         n33604, n33605, n33606, n33607, n33608, n33609, n33610, n33611,
         n33612, n33613, n33614, n33615, n33616, n33617, n33618, n33619,
         n33620, n33621, n33622, n33623, n33624, n33625, n33626, n33627,
         n33628, n33629, n33630, n33631, n33632, n33633, n33634, n33635,
         n33636, n33637, n33638, n33639, n33640, n33641, n33642, n33643,
         n33644, n33645, n33646, n33647, n33648, n33649, n33650, n33651,
         n33652, n33653, n33654, n33655, n33656, n33657, n33658, n33659,
         n33660, n33661, n33662, n33663, n33664, n33665, n33666, n33667,
         n33668, n33669, n33670, n33671, n33672, n33673, n33674, n33675,
         n33676, n33677, n33678, n33679, n33680, n33681, n33682, n33683,
         n33684, n33685, n33686, n33687, n33688, n33689, n33690, n33691,
         n33692, n33693, n33694, n33695, n33696, n33697, n33698, n33699,
         n33700, n33701, n33702, n33703, n33704, n33705, n33706, n33707,
         n33708, n33709, n33710, n33711, n33712, n33713, n33714, n33715,
         n33716, n33717, n33718, n33719, n33720, n33721, n33722, n33723,
         n33724, n33725, n33726, n33727, n33728, n33729, n33730, n33731,
         n33732, n33733, n33734, n33735, n33736, n33737, n33738, n33739,
         n33740, n33741, n33742, n33743, n33744, n33745, n33746, n33747,
         n33748, n33749, n33750, n33751, n33752, n33753, n33754, n33755,
         n33756, n33757, n33758, n33759, n33760, n33761, n33762, n33763,
         n33764, n33765, n33766, n33767, n33768, n33769, n33770, n33771,
         n33772, n33773, n33774, n33775, n33776, n33777, n33778, n33779,
         n33780, n33781, n33782, n33783, n33784, n33785, n33786, n33787,
         n33788, n33789, n33790, n33791, n33792, n33793, n33794, n33795,
         n33796, n33797, n33798, n33799, n33800, n33801, n33802, n33803,
         n33804, n33805, n33806, n33807, n33808, n33809, n33810, n33811,
         n33812, n33813, n33814, n33815, n33816, n33817, n33818, n33819,
         n33820, n33821, n33822, n33823, n33824, n33825, n33826, n33827,
         n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835,
         n33836, n33837, n33838, n33839, n33840, n33841, n33842, n33843,
         n33844, n33845, n33846, n33847, n33848, n33849, n33850, n33851,
         n33852, n33853, n33854, n33855, n33856, n33857, n33858, n33859,
         n33860, n33861, n33862, n33863, n33864, n33865, n33866, n33867,
         n33868, n33869, n33870, n33871, n33872, n33873, n33874, n33875,
         n33876, n33877, n33878, n33879, n33880, n33881, n33882, n33883,
         n33884, n33885, n33886, n33887, n33888, n33889, n33890, n33891,
         n33892, n33893, n33894, n33895, n33896, n33897, n33898, n33899,
         n33900, n33901, n33902, n33903, n33904, n33905, n33906, n33907,
         n33908, n33909, n33910, n33911, n33912, n33913, n33914, n33915,
         n33916, n33917, n33918, n33919, n33920, n33921, n33922, n33923,
         n33924, n33925, n33926, n33927, n33928, n33929, n33930, n33931,
         n33932, n33933, n33934, n33935, n33936, n33937, n33938, n33939,
         n33940, n33941, n33942, n33943, n33944, n33945, n33946, n33947,
         n33948, n33949, n33950, n33951, n33952, n33953, n33954, n33955,
         n33956, n33957, n33958, n33959, n33960, n33961, n33962, n33963,
         n33964, n33965, n33966, n33967, n33968, n33969, n33970, n33971,
         n33972, n33973, n33974, n33975, n33976, n33977, n33978, n33979,
         n33980, n33981, n33982, n33983, n33984, n33985, n33986, n33987,
         n33988, n33989, n33990, n33991, n33992, n33993, n33994, n33995,
         n33996, n33997, n33998, n33999, n34000, n34001, n34002, n34003,
         n34004, n34005, n34006, n34007, n34008, n34009, n34010, n34011,
         n34012, n34013, n34014, n34015, n34016, n34017, n34018, n34019,
         n34020, n34021, n34022, n34023, n34024, n34025, n34026, n34027,
         n34028, n34029, n34030, n34031, n34032, n34033, n34034, n34035,
         n34036, n34037, n34038, n34039, n34040, n34041, n34042, n34043,
         n34044, n34045, n34046, n34047, n34048, n34049, n34050, n34051,
         n34052, n34053, n34054, n34055, n34056, n34057, n34058, n34059,
         n34060, n34061, n34062, n34063, n34064, n34065, n34066, n34067,
         n34068, n34069, n34070, n34071, n34072, n34073, n34074, n34075,
         n34076, n34077, n34078, n34079, n34080, n34081, n34082, n34083,
         n34084, n34085, n34086, n34087, n34088, n34089, n34090, n34091,
         n34092, n34093, n34094, n34095, n34096, n34097, n34098, n34099,
         n34100, n34101, n34102, n34103, n34104, n34105, n34106, n34107,
         n34108, n34109, n34110, n34111, n34112, n34113, n34114, n34115,
         n34116, n34117, n34118, n34119, n34120, n34121, n34122, n34123,
         n34124, n34125, n34126, n34127, n34128, n34129, n34130, n34131,
         n34132, n34133, n34134, n34135, n34136, n34137, n34138, n34139,
         n34140, n34141, n34142, n34143, n34144, n34145, n34146, n34147,
         n34148;
  assign \knn_comb_/min_val_out[0][0]  = p_input[2016];
  assign \knn_comb_/min_val_out[0][1]  = p_input[2017];
  assign \knn_comb_/min_val_out[0][2]  = p_input[2018];
  assign \knn_comb_/min_val_out[0][3]  = p_input[2019];
  assign \knn_comb_/min_val_out[0][4]  = p_input[2020];
  assign \knn_comb_/min_val_out[0][5]  = p_input[2021];
  assign \knn_comb_/min_val_out[0][6]  = p_input[2022];
  assign \knn_comb_/min_val_out[0][7]  = p_input[2023];
  assign \knn_comb_/min_val_out[0][8]  = p_input[2024];
  assign \knn_comb_/min_val_out[0][9]  = p_input[2025];
  assign \knn_comb_/min_val_out[0][10]  = p_input[2026];
  assign \knn_comb_/min_val_out[0][11]  = p_input[2027];
  assign \knn_comb_/min_val_out[0][12]  = p_input[2028];
  assign \knn_comb_/min_val_out[0][13]  = p_input[2029];
  assign \knn_comb_/min_val_out[0][14]  = p_input[2030];
  assign \knn_comb_/min_val_out[0][15]  = p_input[2031];
  assign \knn_comb_/min_val_out[0][16]  = p_input[2032];
  assign \knn_comb_/min_val_out[0][17]  = p_input[2033];
  assign \knn_comb_/min_val_out[0][18]  = p_input[2034];
  assign \knn_comb_/min_val_out[0][19]  = p_input[2035];
  assign \knn_comb_/min_val_out[0][20]  = p_input[2036];
  assign \knn_comb_/min_val_out[0][21]  = p_input[2037];
  assign \knn_comb_/min_val_out[0][22]  = p_input[2038];
  assign \knn_comb_/min_val_out[0][23]  = p_input[2039];
  assign \knn_comb_/min_val_out[0][24]  = p_input[2040];
  assign \knn_comb_/min_val_out[0][25]  = p_input[2041];
  assign \knn_comb_/min_val_out[0][26]  = p_input[2042];
  assign \knn_comb_/min_val_out[0][27]  = p_input[2043];
  assign \knn_comb_/min_val_out[0][28]  = p_input[2044];
  assign \knn_comb_/min_val_out[0][29]  = p_input[2045];
  assign \knn_comb_/min_val_out[0][30]  = p_input[2046];
  assign \knn_comb_/min_val_out[0][31]  = p_input[2047];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][0]  = p_input[1984];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][1]  = p_input[1985];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][2]  = p_input[1986];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][3]  = p_input[1987];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][4]  = p_input[1988];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][5]  = p_input[1989];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][6]  = p_input[1990];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][7]  = p_input[1991];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][8]  = p_input[1992];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][9]  = p_input[1993];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][10]  = p_input[1994];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][11]  = p_input[1995];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][12]  = p_input[1996];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][13]  = p_input[1997];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][14]  = p_input[1998];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][15]  = p_input[1999];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][16]  = p_input[2000];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][17]  = p_input[2001];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][18]  = p_input[2002];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][19]  = p_input[2003];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][20]  = p_input[2004];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][21]  = p_input[2005];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][22]  = p_input[2006];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][23]  = p_input[2007];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][24]  = p_input[2008];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][25]  = p_input[2009];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][26]  = p_input[2010];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][27]  = p_input[2011];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][28]  = p_input[2012];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][29]  = p_input[2013];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][30]  = p_input[2014];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][31]  = p_input[2015];

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  XOR U2 ( .A(n3), .B(n4), .Z(o[8]) );
  XOR U3 ( .A(n5), .B(n6), .Z(o[7]) );
  XOR U4 ( .A(n7), .B(n8), .Z(o[6]) );
  XOR U5 ( .A(n9), .B(n10), .Z(o[63]) );
  XOR U6 ( .A(n11), .B(n12), .Z(o[62]) );
  XOR U7 ( .A(n13), .B(n14), .Z(o[61]) );
  XOR U8 ( .A(n15), .B(n16), .Z(o[60]) );
  XOR U9 ( .A(n17), .B(n18), .Z(o[5]) );
  XOR U10 ( .A(n19), .B(n20), .Z(o[59]) );
  XOR U11 ( .A(n21), .B(n22), .Z(o[58]) );
  XOR U12 ( .A(n23), .B(n24), .Z(o[57]) );
  XOR U13 ( .A(n25), .B(n26), .Z(o[56]) );
  XOR U14 ( .A(n27), .B(n28), .Z(o[55]) );
  XOR U15 ( .A(n29), .B(n30), .Z(o[54]) );
  XOR U16 ( .A(n31), .B(n32), .Z(o[53]) );
  XOR U17 ( .A(n33), .B(n34), .Z(o[52]) );
  XOR U18 ( .A(n35), .B(n36), .Z(o[51]) );
  XOR U19 ( .A(n37), .B(n38), .Z(o[50]) );
  XOR U20 ( .A(n39), .B(n40), .Z(o[4]) );
  XOR U21 ( .A(n41), .B(n42), .Z(o[49]) );
  XOR U22 ( .A(n43), .B(n44), .Z(o[48]) );
  XOR U23 ( .A(n45), .B(n46), .Z(o[47]) );
  XOR U24 ( .A(n47), .B(n48), .Z(o[46]) );
  XOR U25 ( .A(n49), .B(n50), .Z(o[45]) );
  XOR U26 ( .A(n51), .B(n52), .Z(o[44]) );
  XOR U27 ( .A(n53), .B(n54), .Z(o[43]) );
  XOR U28 ( .A(n55), .B(n56), .Z(o[42]) );
  XOR U29 ( .A(n1), .B(n57), .Z(o[41]) );
  AND U30 ( .A(n58), .B(n59), .Z(n1) );
  XOR U31 ( .A(n2), .B(n57), .Z(n59) );
  XOR U32 ( .A(n60), .B(n61), .Z(n57) );
  AND U33 ( .A(n62), .B(n63), .Z(n61) );
  XOR U34 ( .A(p_input[9]), .B(n60), .Z(n63) );
  XOR U35 ( .A(n64), .B(n65), .Z(n60) );
  AND U36 ( .A(n66), .B(n67), .Z(n65) );
  XOR U37 ( .A(n68), .B(n69), .Z(n2) );
  AND U38 ( .A(n70), .B(n67), .Z(n69) );
  XNOR U39 ( .A(n71), .B(n64), .Z(n67) );
  XOR U40 ( .A(n72), .B(n73), .Z(n64) );
  AND U41 ( .A(n74), .B(n75), .Z(n73) );
  XOR U42 ( .A(p_input[41]), .B(n72), .Z(n75) );
  XOR U43 ( .A(n76), .B(n77), .Z(n72) );
  AND U44 ( .A(n78), .B(n79), .Z(n77) );
  IV U45 ( .A(n68), .Z(n71) );
  XNOR U46 ( .A(n80), .B(n81), .Z(n68) );
  AND U47 ( .A(n82), .B(n79), .Z(n81) );
  XNOR U48 ( .A(n80), .B(n76), .Z(n79) );
  XOR U49 ( .A(n83), .B(n84), .Z(n76) );
  AND U50 ( .A(n85), .B(n86), .Z(n84) );
  XOR U51 ( .A(p_input[73]), .B(n83), .Z(n86) );
  XOR U52 ( .A(n87), .B(n88), .Z(n83) );
  AND U53 ( .A(n89), .B(n90), .Z(n88) );
  XOR U54 ( .A(n91), .B(n92), .Z(n80) );
  AND U55 ( .A(n93), .B(n90), .Z(n92) );
  XNOR U56 ( .A(n91), .B(n87), .Z(n90) );
  XOR U57 ( .A(n94), .B(n95), .Z(n87) );
  AND U58 ( .A(n96), .B(n97), .Z(n95) );
  XOR U59 ( .A(p_input[105]), .B(n94), .Z(n97) );
  XOR U60 ( .A(n98), .B(n99), .Z(n94) );
  AND U61 ( .A(n100), .B(n101), .Z(n99) );
  XOR U62 ( .A(n102), .B(n103), .Z(n91) );
  AND U63 ( .A(n104), .B(n101), .Z(n103) );
  XNOR U64 ( .A(n102), .B(n98), .Z(n101) );
  XOR U65 ( .A(n105), .B(n106), .Z(n98) );
  AND U66 ( .A(n107), .B(n108), .Z(n106) );
  XOR U67 ( .A(p_input[137]), .B(n105), .Z(n108) );
  XOR U68 ( .A(n109), .B(n110), .Z(n105) );
  AND U69 ( .A(n111), .B(n112), .Z(n110) );
  XOR U70 ( .A(n113), .B(n114), .Z(n102) );
  AND U71 ( .A(n115), .B(n112), .Z(n114) );
  XNOR U72 ( .A(n113), .B(n109), .Z(n112) );
  XOR U73 ( .A(n116), .B(n117), .Z(n109) );
  AND U74 ( .A(n118), .B(n119), .Z(n117) );
  XOR U75 ( .A(p_input[169]), .B(n116), .Z(n119) );
  XOR U76 ( .A(n120), .B(n121), .Z(n116) );
  AND U77 ( .A(n122), .B(n123), .Z(n121) );
  XOR U78 ( .A(n124), .B(n125), .Z(n113) );
  AND U79 ( .A(n126), .B(n123), .Z(n125) );
  XNOR U80 ( .A(n124), .B(n120), .Z(n123) );
  XOR U81 ( .A(n127), .B(n128), .Z(n120) );
  AND U82 ( .A(n129), .B(n130), .Z(n128) );
  XOR U83 ( .A(p_input[201]), .B(n127), .Z(n130) );
  XOR U84 ( .A(n131), .B(n132), .Z(n127) );
  AND U85 ( .A(n133), .B(n134), .Z(n132) );
  XOR U86 ( .A(n135), .B(n136), .Z(n124) );
  AND U87 ( .A(n137), .B(n134), .Z(n136) );
  XNOR U88 ( .A(n135), .B(n131), .Z(n134) );
  XOR U89 ( .A(n138), .B(n139), .Z(n131) );
  AND U90 ( .A(n140), .B(n141), .Z(n139) );
  XOR U91 ( .A(p_input[233]), .B(n138), .Z(n141) );
  XOR U92 ( .A(n142), .B(n143), .Z(n138) );
  AND U93 ( .A(n144), .B(n145), .Z(n143) );
  XOR U94 ( .A(n146), .B(n147), .Z(n135) );
  AND U95 ( .A(n148), .B(n145), .Z(n147) );
  XNOR U96 ( .A(n146), .B(n142), .Z(n145) );
  XOR U97 ( .A(n149), .B(n150), .Z(n142) );
  AND U98 ( .A(n151), .B(n152), .Z(n150) );
  XOR U99 ( .A(p_input[265]), .B(n149), .Z(n152) );
  XOR U100 ( .A(n153), .B(n154), .Z(n149) );
  AND U101 ( .A(n155), .B(n156), .Z(n154) );
  XOR U102 ( .A(n157), .B(n158), .Z(n146) );
  AND U103 ( .A(n159), .B(n156), .Z(n158) );
  XNOR U104 ( .A(n157), .B(n153), .Z(n156) );
  XOR U105 ( .A(n160), .B(n161), .Z(n153) );
  AND U106 ( .A(n162), .B(n163), .Z(n161) );
  XOR U107 ( .A(p_input[297]), .B(n160), .Z(n163) );
  XOR U108 ( .A(n164), .B(n165), .Z(n160) );
  AND U109 ( .A(n166), .B(n167), .Z(n165) );
  XOR U110 ( .A(n168), .B(n169), .Z(n157) );
  AND U111 ( .A(n170), .B(n167), .Z(n169) );
  XNOR U112 ( .A(n168), .B(n164), .Z(n167) );
  XOR U113 ( .A(n171), .B(n172), .Z(n164) );
  AND U114 ( .A(n173), .B(n174), .Z(n172) );
  XOR U115 ( .A(p_input[329]), .B(n171), .Z(n174) );
  XOR U116 ( .A(n175), .B(n176), .Z(n171) );
  AND U117 ( .A(n177), .B(n178), .Z(n176) );
  XOR U118 ( .A(n179), .B(n180), .Z(n168) );
  AND U119 ( .A(n181), .B(n178), .Z(n180) );
  XNOR U120 ( .A(n179), .B(n175), .Z(n178) );
  XOR U121 ( .A(n182), .B(n183), .Z(n175) );
  AND U122 ( .A(n184), .B(n185), .Z(n183) );
  XOR U123 ( .A(p_input[361]), .B(n182), .Z(n185) );
  XOR U124 ( .A(n186), .B(n187), .Z(n182) );
  AND U125 ( .A(n188), .B(n189), .Z(n187) );
  XOR U126 ( .A(n190), .B(n191), .Z(n179) );
  AND U127 ( .A(n192), .B(n189), .Z(n191) );
  XNOR U128 ( .A(n190), .B(n186), .Z(n189) );
  XOR U129 ( .A(n193), .B(n194), .Z(n186) );
  AND U130 ( .A(n195), .B(n196), .Z(n194) );
  XOR U131 ( .A(p_input[393]), .B(n193), .Z(n196) );
  XOR U132 ( .A(n197), .B(n198), .Z(n193) );
  AND U133 ( .A(n199), .B(n200), .Z(n198) );
  XOR U134 ( .A(n201), .B(n202), .Z(n190) );
  AND U135 ( .A(n203), .B(n200), .Z(n202) );
  XNOR U136 ( .A(n201), .B(n197), .Z(n200) );
  XOR U137 ( .A(n204), .B(n205), .Z(n197) );
  AND U138 ( .A(n206), .B(n207), .Z(n205) );
  XOR U139 ( .A(p_input[425]), .B(n204), .Z(n207) );
  XOR U140 ( .A(n208), .B(n209), .Z(n204) );
  AND U141 ( .A(n210), .B(n211), .Z(n209) );
  XOR U142 ( .A(n212), .B(n213), .Z(n201) );
  AND U143 ( .A(n214), .B(n211), .Z(n213) );
  XNOR U144 ( .A(n212), .B(n208), .Z(n211) );
  XOR U145 ( .A(n215), .B(n216), .Z(n208) );
  AND U146 ( .A(n217), .B(n218), .Z(n216) );
  XOR U147 ( .A(p_input[457]), .B(n215), .Z(n218) );
  XOR U148 ( .A(n219), .B(n220), .Z(n215) );
  AND U149 ( .A(n221), .B(n222), .Z(n220) );
  XOR U150 ( .A(n223), .B(n224), .Z(n212) );
  AND U151 ( .A(n225), .B(n222), .Z(n224) );
  XNOR U152 ( .A(n223), .B(n219), .Z(n222) );
  XOR U153 ( .A(n226), .B(n227), .Z(n219) );
  AND U154 ( .A(n228), .B(n229), .Z(n227) );
  XOR U155 ( .A(p_input[489]), .B(n226), .Z(n229) );
  XOR U156 ( .A(n230), .B(n231), .Z(n226) );
  AND U157 ( .A(n232), .B(n233), .Z(n231) );
  XOR U158 ( .A(n234), .B(n235), .Z(n223) );
  AND U159 ( .A(n236), .B(n233), .Z(n235) );
  XNOR U160 ( .A(n234), .B(n230), .Z(n233) );
  XOR U161 ( .A(n237), .B(n238), .Z(n230) );
  AND U162 ( .A(n239), .B(n240), .Z(n238) );
  XOR U163 ( .A(p_input[521]), .B(n237), .Z(n240) );
  XOR U164 ( .A(n241), .B(n242), .Z(n237) );
  AND U165 ( .A(n243), .B(n244), .Z(n242) );
  XOR U166 ( .A(n245), .B(n246), .Z(n234) );
  AND U167 ( .A(n247), .B(n244), .Z(n246) );
  XNOR U168 ( .A(n245), .B(n241), .Z(n244) );
  XOR U169 ( .A(n248), .B(n249), .Z(n241) );
  AND U170 ( .A(n250), .B(n251), .Z(n249) );
  XOR U171 ( .A(p_input[553]), .B(n248), .Z(n251) );
  XOR U172 ( .A(n252), .B(n253), .Z(n248) );
  AND U173 ( .A(n254), .B(n255), .Z(n253) );
  XOR U174 ( .A(n256), .B(n257), .Z(n245) );
  AND U175 ( .A(n258), .B(n255), .Z(n257) );
  XNOR U176 ( .A(n256), .B(n252), .Z(n255) );
  XOR U177 ( .A(n259), .B(n260), .Z(n252) );
  AND U178 ( .A(n261), .B(n262), .Z(n260) );
  XOR U179 ( .A(p_input[585]), .B(n259), .Z(n262) );
  XOR U180 ( .A(n263), .B(n264), .Z(n259) );
  AND U181 ( .A(n265), .B(n266), .Z(n264) );
  XOR U182 ( .A(n267), .B(n268), .Z(n256) );
  AND U183 ( .A(n269), .B(n266), .Z(n268) );
  XNOR U184 ( .A(n267), .B(n263), .Z(n266) );
  XOR U185 ( .A(n270), .B(n271), .Z(n263) );
  AND U186 ( .A(n272), .B(n273), .Z(n271) );
  XOR U187 ( .A(p_input[617]), .B(n270), .Z(n273) );
  XOR U188 ( .A(n274), .B(n275), .Z(n270) );
  AND U189 ( .A(n276), .B(n277), .Z(n275) );
  XOR U190 ( .A(n278), .B(n279), .Z(n267) );
  AND U191 ( .A(n280), .B(n277), .Z(n279) );
  XNOR U192 ( .A(n278), .B(n274), .Z(n277) );
  XOR U193 ( .A(n281), .B(n282), .Z(n274) );
  AND U194 ( .A(n283), .B(n284), .Z(n282) );
  XOR U195 ( .A(p_input[649]), .B(n281), .Z(n284) );
  XOR U196 ( .A(n285), .B(n286), .Z(n281) );
  AND U197 ( .A(n287), .B(n288), .Z(n286) );
  XOR U198 ( .A(n289), .B(n290), .Z(n278) );
  AND U199 ( .A(n291), .B(n288), .Z(n290) );
  XNOR U200 ( .A(n289), .B(n285), .Z(n288) );
  XOR U201 ( .A(n292), .B(n293), .Z(n285) );
  AND U202 ( .A(n294), .B(n295), .Z(n293) );
  XOR U203 ( .A(p_input[681]), .B(n292), .Z(n295) );
  XOR U204 ( .A(n296), .B(n297), .Z(n292) );
  AND U205 ( .A(n298), .B(n299), .Z(n297) );
  XOR U206 ( .A(n300), .B(n301), .Z(n289) );
  AND U207 ( .A(n302), .B(n299), .Z(n301) );
  XNOR U208 ( .A(n300), .B(n296), .Z(n299) );
  XOR U209 ( .A(n303), .B(n304), .Z(n296) );
  AND U210 ( .A(n305), .B(n306), .Z(n304) );
  XOR U211 ( .A(p_input[713]), .B(n303), .Z(n306) );
  XOR U212 ( .A(n307), .B(n308), .Z(n303) );
  AND U213 ( .A(n309), .B(n310), .Z(n308) );
  XOR U214 ( .A(n311), .B(n312), .Z(n300) );
  AND U215 ( .A(n313), .B(n310), .Z(n312) );
  XNOR U216 ( .A(n311), .B(n307), .Z(n310) );
  XOR U217 ( .A(n314), .B(n315), .Z(n307) );
  AND U218 ( .A(n316), .B(n317), .Z(n315) );
  XOR U219 ( .A(p_input[745]), .B(n314), .Z(n317) );
  XOR U220 ( .A(n318), .B(n319), .Z(n314) );
  AND U221 ( .A(n320), .B(n321), .Z(n319) );
  XOR U222 ( .A(n322), .B(n323), .Z(n311) );
  AND U223 ( .A(n324), .B(n321), .Z(n323) );
  XNOR U224 ( .A(n322), .B(n318), .Z(n321) );
  XOR U225 ( .A(n325), .B(n326), .Z(n318) );
  AND U226 ( .A(n327), .B(n328), .Z(n326) );
  XOR U227 ( .A(p_input[777]), .B(n325), .Z(n328) );
  XOR U228 ( .A(n329), .B(n330), .Z(n325) );
  AND U229 ( .A(n331), .B(n332), .Z(n330) );
  XOR U230 ( .A(n333), .B(n334), .Z(n322) );
  AND U231 ( .A(n335), .B(n332), .Z(n334) );
  XNOR U232 ( .A(n333), .B(n329), .Z(n332) );
  XOR U233 ( .A(n336), .B(n337), .Z(n329) );
  AND U234 ( .A(n338), .B(n339), .Z(n337) );
  XOR U235 ( .A(p_input[809]), .B(n336), .Z(n339) );
  XOR U236 ( .A(n340), .B(n341), .Z(n336) );
  AND U237 ( .A(n342), .B(n343), .Z(n341) );
  XOR U238 ( .A(n344), .B(n345), .Z(n333) );
  AND U239 ( .A(n346), .B(n343), .Z(n345) );
  XNOR U240 ( .A(n344), .B(n340), .Z(n343) );
  XOR U241 ( .A(n347), .B(n348), .Z(n340) );
  AND U242 ( .A(n349), .B(n350), .Z(n348) );
  XOR U243 ( .A(p_input[841]), .B(n347), .Z(n350) );
  XOR U244 ( .A(n351), .B(n352), .Z(n347) );
  AND U245 ( .A(n353), .B(n354), .Z(n352) );
  XOR U246 ( .A(n355), .B(n356), .Z(n344) );
  AND U247 ( .A(n357), .B(n354), .Z(n356) );
  XNOR U248 ( .A(n355), .B(n351), .Z(n354) );
  XOR U249 ( .A(n358), .B(n359), .Z(n351) );
  AND U250 ( .A(n360), .B(n361), .Z(n359) );
  XOR U251 ( .A(p_input[873]), .B(n358), .Z(n361) );
  XOR U252 ( .A(n362), .B(n363), .Z(n358) );
  AND U253 ( .A(n364), .B(n365), .Z(n363) );
  XOR U254 ( .A(n366), .B(n367), .Z(n355) );
  AND U255 ( .A(n368), .B(n365), .Z(n367) );
  XNOR U256 ( .A(n366), .B(n362), .Z(n365) );
  XOR U257 ( .A(n369), .B(n370), .Z(n362) );
  AND U258 ( .A(n371), .B(n372), .Z(n370) );
  XOR U259 ( .A(p_input[905]), .B(n369), .Z(n372) );
  XOR U260 ( .A(n373), .B(n374), .Z(n369) );
  AND U261 ( .A(n375), .B(n376), .Z(n374) );
  XOR U262 ( .A(n377), .B(n378), .Z(n366) );
  AND U263 ( .A(n379), .B(n376), .Z(n378) );
  XNOR U264 ( .A(n377), .B(n373), .Z(n376) );
  XOR U265 ( .A(n380), .B(n381), .Z(n373) );
  AND U266 ( .A(n382), .B(n383), .Z(n381) );
  XOR U267 ( .A(p_input[937]), .B(n380), .Z(n383) );
  XOR U268 ( .A(n384), .B(n385), .Z(n380) );
  AND U269 ( .A(n386), .B(n387), .Z(n385) );
  XOR U270 ( .A(n388), .B(n389), .Z(n377) );
  AND U271 ( .A(n390), .B(n387), .Z(n389) );
  XNOR U272 ( .A(n388), .B(n384), .Z(n387) );
  XOR U273 ( .A(n391), .B(n392), .Z(n384) );
  AND U274 ( .A(n393), .B(n394), .Z(n392) );
  XOR U275 ( .A(p_input[969]), .B(n391), .Z(n394) );
  XOR U276 ( .A(n395), .B(n396), .Z(n391) );
  AND U277 ( .A(n397), .B(n398), .Z(n396) );
  XOR U278 ( .A(n399), .B(n400), .Z(n388) );
  AND U279 ( .A(n401), .B(n398), .Z(n400) );
  XNOR U280 ( .A(n399), .B(n395), .Z(n398) );
  XOR U281 ( .A(n402), .B(n403), .Z(n395) );
  AND U282 ( .A(n404), .B(n405), .Z(n403) );
  XOR U283 ( .A(p_input[1001]), .B(n402), .Z(n405) );
  XOR U284 ( .A(n406), .B(n407), .Z(n402) );
  AND U285 ( .A(n408), .B(n409), .Z(n407) );
  XOR U286 ( .A(n410), .B(n411), .Z(n399) );
  AND U287 ( .A(n412), .B(n409), .Z(n411) );
  XNOR U288 ( .A(n410), .B(n406), .Z(n409) );
  XOR U289 ( .A(n413), .B(n414), .Z(n406) );
  AND U290 ( .A(n415), .B(n416), .Z(n414) );
  XOR U291 ( .A(p_input[1033]), .B(n413), .Z(n416) );
  XOR U292 ( .A(n417), .B(n418), .Z(n413) );
  AND U293 ( .A(n419), .B(n420), .Z(n418) );
  XOR U294 ( .A(n421), .B(n422), .Z(n410) );
  AND U295 ( .A(n423), .B(n420), .Z(n422) );
  XNOR U296 ( .A(n421), .B(n417), .Z(n420) );
  XOR U297 ( .A(n424), .B(n425), .Z(n417) );
  AND U298 ( .A(n426), .B(n427), .Z(n425) );
  XOR U299 ( .A(p_input[1065]), .B(n424), .Z(n427) );
  XOR U300 ( .A(n428), .B(n429), .Z(n424) );
  AND U301 ( .A(n430), .B(n431), .Z(n429) );
  XOR U302 ( .A(n432), .B(n433), .Z(n421) );
  AND U303 ( .A(n434), .B(n431), .Z(n433) );
  XNOR U304 ( .A(n432), .B(n428), .Z(n431) );
  XOR U305 ( .A(n435), .B(n436), .Z(n428) );
  AND U306 ( .A(n437), .B(n438), .Z(n436) );
  XOR U307 ( .A(p_input[1097]), .B(n435), .Z(n438) );
  XOR U308 ( .A(n439), .B(n440), .Z(n435) );
  AND U309 ( .A(n441), .B(n442), .Z(n440) );
  XOR U310 ( .A(n443), .B(n444), .Z(n432) );
  AND U311 ( .A(n445), .B(n442), .Z(n444) );
  XNOR U312 ( .A(n443), .B(n439), .Z(n442) );
  XOR U313 ( .A(n446), .B(n447), .Z(n439) );
  AND U314 ( .A(n448), .B(n449), .Z(n447) );
  XOR U315 ( .A(p_input[1129]), .B(n446), .Z(n449) );
  XOR U316 ( .A(n450), .B(n451), .Z(n446) );
  AND U317 ( .A(n452), .B(n453), .Z(n451) );
  XOR U318 ( .A(n454), .B(n455), .Z(n443) );
  AND U319 ( .A(n456), .B(n453), .Z(n455) );
  XNOR U320 ( .A(n454), .B(n450), .Z(n453) );
  XOR U321 ( .A(n457), .B(n458), .Z(n450) );
  AND U322 ( .A(n459), .B(n460), .Z(n458) );
  XOR U323 ( .A(p_input[1161]), .B(n457), .Z(n460) );
  XOR U324 ( .A(n461), .B(n462), .Z(n457) );
  AND U325 ( .A(n463), .B(n464), .Z(n462) );
  XOR U326 ( .A(n465), .B(n466), .Z(n454) );
  AND U327 ( .A(n467), .B(n464), .Z(n466) );
  XNOR U328 ( .A(n465), .B(n461), .Z(n464) );
  XOR U329 ( .A(n468), .B(n469), .Z(n461) );
  AND U330 ( .A(n470), .B(n471), .Z(n469) );
  XOR U331 ( .A(p_input[1193]), .B(n468), .Z(n471) );
  XOR U332 ( .A(n472), .B(n473), .Z(n468) );
  AND U333 ( .A(n474), .B(n475), .Z(n473) );
  XOR U334 ( .A(n476), .B(n477), .Z(n465) );
  AND U335 ( .A(n478), .B(n475), .Z(n477) );
  XNOR U336 ( .A(n476), .B(n472), .Z(n475) );
  XOR U337 ( .A(n479), .B(n480), .Z(n472) );
  AND U338 ( .A(n481), .B(n482), .Z(n480) );
  XOR U339 ( .A(p_input[1225]), .B(n479), .Z(n482) );
  XOR U340 ( .A(n483), .B(n484), .Z(n479) );
  AND U341 ( .A(n485), .B(n486), .Z(n484) );
  XOR U342 ( .A(n487), .B(n488), .Z(n476) );
  AND U343 ( .A(n489), .B(n486), .Z(n488) );
  XNOR U344 ( .A(n487), .B(n483), .Z(n486) );
  XOR U345 ( .A(n490), .B(n491), .Z(n483) );
  AND U346 ( .A(n492), .B(n493), .Z(n491) );
  XOR U347 ( .A(p_input[1257]), .B(n490), .Z(n493) );
  XOR U348 ( .A(n494), .B(n495), .Z(n490) );
  AND U349 ( .A(n496), .B(n497), .Z(n495) );
  XOR U350 ( .A(n498), .B(n499), .Z(n487) );
  AND U351 ( .A(n500), .B(n497), .Z(n499) );
  XNOR U352 ( .A(n498), .B(n494), .Z(n497) );
  XOR U353 ( .A(n501), .B(n502), .Z(n494) );
  AND U354 ( .A(n503), .B(n504), .Z(n502) );
  XOR U355 ( .A(p_input[1289]), .B(n501), .Z(n504) );
  XOR U356 ( .A(n505), .B(n506), .Z(n501) );
  AND U357 ( .A(n507), .B(n508), .Z(n506) );
  XOR U358 ( .A(n509), .B(n510), .Z(n498) );
  AND U359 ( .A(n511), .B(n508), .Z(n510) );
  XNOR U360 ( .A(n509), .B(n505), .Z(n508) );
  XOR U361 ( .A(n512), .B(n513), .Z(n505) );
  AND U362 ( .A(n514), .B(n515), .Z(n513) );
  XOR U363 ( .A(p_input[1321]), .B(n512), .Z(n515) );
  XOR U364 ( .A(n516), .B(n517), .Z(n512) );
  AND U365 ( .A(n518), .B(n519), .Z(n517) );
  XOR U366 ( .A(n520), .B(n521), .Z(n509) );
  AND U367 ( .A(n522), .B(n519), .Z(n521) );
  XNOR U368 ( .A(n520), .B(n516), .Z(n519) );
  XOR U369 ( .A(n523), .B(n524), .Z(n516) );
  AND U370 ( .A(n525), .B(n526), .Z(n524) );
  XOR U371 ( .A(p_input[1353]), .B(n523), .Z(n526) );
  XOR U372 ( .A(n527), .B(n528), .Z(n523) );
  AND U373 ( .A(n529), .B(n530), .Z(n528) );
  XOR U374 ( .A(n531), .B(n532), .Z(n520) );
  AND U375 ( .A(n533), .B(n530), .Z(n532) );
  XNOR U376 ( .A(n531), .B(n527), .Z(n530) );
  XOR U377 ( .A(n534), .B(n535), .Z(n527) );
  AND U378 ( .A(n536), .B(n537), .Z(n535) );
  XOR U379 ( .A(p_input[1385]), .B(n534), .Z(n537) );
  XOR U380 ( .A(n538), .B(n539), .Z(n534) );
  AND U381 ( .A(n540), .B(n541), .Z(n539) );
  XOR U382 ( .A(n542), .B(n543), .Z(n531) );
  AND U383 ( .A(n544), .B(n541), .Z(n543) );
  XNOR U384 ( .A(n542), .B(n538), .Z(n541) );
  XOR U385 ( .A(n545), .B(n546), .Z(n538) );
  AND U386 ( .A(n547), .B(n548), .Z(n546) );
  XOR U387 ( .A(p_input[1417]), .B(n545), .Z(n548) );
  XOR U388 ( .A(n549), .B(n550), .Z(n545) );
  AND U389 ( .A(n551), .B(n552), .Z(n550) );
  XOR U390 ( .A(n553), .B(n554), .Z(n542) );
  AND U391 ( .A(n555), .B(n552), .Z(n554) );
  XNOR U392 ( .A(n553), .B(n549), .Z(n552) );
  XOR U393 ( .A(n556), .B(n557), .Z(n549) );
  AND U394 ( .A(n558), .B(n559), .Z(n557) );
  XOR U395 ( .A(p_input[1449]), .B(n556), .Z(n559) );
  XOR U396 ( .A(n560), .B(n561), .Z(n556) );
  AND U397 ( .A(n562), .B(n563), .Z(n561) );
  XOR U398 ( .A(n564), .B(n565), .Z(n553) );
  AND U399 ( .A(n566), .B(n563), .Z(n565) );
  XNOR U400 ( .A(n564), .B(n560), .Z(n563) );
  XOR U401 ( .A(n567), .B(n568), .Z(n560) );
  AND U402 ( .A(n569), .B(n570), .Z(n568) );
  XOR U403 ( .A(p_input[1481]), .B(n567), .Z(n570) );
  XOR U404 ( .A(n571), .B(n572), .Z(n567) );
  AND U405 ( .A(n573), .B(n574), .Z(n572) );
  XOR U406 ( .A(n575), .B(n576), .Z(n564) );
  AND U407 ( .A(n577), .B(n574), .Z(n576) );
  XNOR U408 ( .A(n575), .B(n571), .Z(n574) );
  XOR U409 ( .A(n578), .B(n579), .Z(n571) );
  AND U410 ( .A(n580), .B(n581), .Z(n579) );
  XOR U411 ( .A(p_input[1513]), .B(n578), .Z(n581) );
  XOR U412 ( .A(n582), .B(n583), .Z(n578) );
  AND U413 ( .A(n584), .B(n585), .Z(n583) );
  XOR U414 ( .A(n586), .B(n587), .Z(n575) );
  AND U415 ( .A(n588), .B(n585), .Z(n587) );
  XNOR U416 ( .A(n586), .B(n582), .Z(n585) );
  XOR U417 ( .A(n589), .B(n590), .Z(n582) );
  AND U418 ( .A(n591), .B(n592), .Z(n590) );
  XOR U419 ( .A(p_input[1545]), .B(n589), .Z(n592) );
  XOR U420 ( .A(n593), .B(n594), .Z(n589) );
  AND U421 ( .A(n595), .B(n596), .Z(n594) );
  XOR U422 ( .A(n597), .B(n598), .Z(n586) );
  AND U423 ( .A(n599), .B(n596), .Z(n598) );
  XNOR U424 ( .A(n597), .B(n593), .Z(n596) );
  XOR U425 ( .A(n600), .B(n601), .Z(n593) );
  AND U426 ( .A(n602), .B(n603), .Z(n601) );
  XOR U427 ( .A(p_input[1577]), .B(n600), .Z(n603) );
  XOR U428 ( .A(n604), .B(n605), .Z(n600) );
  AND U429 ( .A(n606), .B(n607), .Z(n605) );
  XOR U430 ( .A(n608), .B(n609), .Z(n597) );
  AND U431 ( .A(n610), .B(n607), .Z(n609) );
  XNOR U432 ( .A(n608), .B(n604), .Z(n607) );
  XOR U433 ( .A(n611), .B(n612), .Z(n604) );
  AND U434 ( .A(n613), .B(n614), .Z(n612) );
  XOR U435 ( .A(p_input[1609]), .B(n611), .Z(n614) );
  XOR U436 ( .A(n615), .B(n616), .Z(n611) );
  AND U437 ( .A(n617), .B(n618), .Z(n616) );
  XOR U438 ( .A(n619), .B(n620), .Z(n608) );
  AND U439 ( .A(n621), .B(n618), .Z(n620) );
  XNOR U440 ( .A(n619), .B(n615), .Z(n618) );
  XOR U441 ( .A(n622), .B(n623), .Z(n615) );
  AND U442 ( .A(n624), .B(n625), .Z(n623) );
  XOR U443 ( .A(p_input[1641]), .B(n622), .Z(n625) );
  XOR U444 ( .A(n626), .B(n627), .Z(n622) );
  AND U445 ( .A(n628), .B(n629), .Z(n627) );
  XOR U446 ( .A(n630), .B(n631), .Z(n619) );
  AND U447 ( .A(n632), .B(n629), .Z(n631) );
  XNOR U448 ( .A(n630), .B(n626), .Z(n629) );
  XOR U449 ( .A(n633), .B(n634), .Z(n626) );
  AND U450 ( .A(n635), .B(n636), .Z(n634) );
  XOR U451 ( .A(p_input[1673]), .B(n633), .Z(n636) );
  XOR U452 ( .A(n637), .B(n638), .Z(n633) );
  AND U453 ( .A(n639), .B(n640), .Z(n638) );
  XOR U454 ( .A(n641), .B(n642), .Z(n630) );
  AND U455 ( .A(n643), .B(n640), .Z(n642) );
  XNOR U456 ( .A(n641), .B(n637), .Z(n640) );
  XOR U457 ( .A(n644), .B(n645), .Z(n637) );
  AND U458 ( .A(n646), .B(n647), .Z(n645) );
  XOR U459 ( .A(p_input[1705]), .B(n644), .Z(n647) );
  XOR U460 ( .A(n648), .B(n649), .Z(n644) );
  AND U461 ( .A(n650), .B(n651), .Z(n649) );
  XOR U462 ( .A(n652), .B(n653), .Z(n641) );
  AND U463 ( .A(n654), .B(n651), .Z(n653) );
  XNOR U464 ( .A(n652), .B(n648), .Z(n651) );
  XOR U465 ( .A(n655), .B(n656), .Z(n648) );
  AND U466 ( .A(n657), .B(n658), .Z(n656) );
  XOR U467 ( .A(p_input[1737]), .B(n655), .Z(n658) );
  XOR U468 ( .A(n659), .B(n660), .Z(n655) );
  AND U469 ( .A(n661), .B(n662), .Z(n660) );
  XOR U470 ( .A(n663), .B(n664), .Z(n652) );
  AND U471 ( .A(n665), .B(n662), .Z(n664) );
  XNOR U472 ( .A(n663), .B(n659), .Z(n662) );
  XOR U473 ( .A(n666), .B(n667), .Z(n659) );
  AND U474 ( .A(n668), .B(n669), .Z(n667) );
  XOR U475 ( .A(p_input[1769]), .B(n666), .Z(n669) );
  XOR U476 ( .A(n670), .B(n671), .Z(n666) );
  AND U477 ( .A(n672), .B(n673), .Z(n671) );
  XOR U478 ( .A(n674), .B(n675), .Z(n663) );
  AND U479 ( .A(n676), .B(n673), .Z(n675) );
  XNOR U480 ( .A(n674), .B(n670), .Z(n673) );
  XOR U481 ( .A(n677), .B(n678), .Z(n670) );
  AND U482 ( .A(n679), .B(n680), .Z(n678) );
  XOR U483 ( .A(p_input[1801]), .B(n677), .Z(n680) );
  XOR U484 ( .A(n681), .B(n682), .Z(n677) );
  AND U485 ( .A(n683), .B(n684), .Z(n682) );
  XOR U486 ( .A(n685), .B(n686), .Z(n674) );
  AND U487 ( .A(n687), .B(n684), .Z(n686) );
  XNOR U488 ( .A(n685), .B(n681), .Z(n684) );
  XOR U489 ( .A(n688), .B(n689), .Z(n681) );
  AND U490 ( .A(n690), .B(n691), .Z(n689) );
  XOR U491 ( .A(p_input[1833]), .B(n688), .Z(n691) );
  XOR U492 ( .A(n692), .B(n693), .Z(n688) );
  AND U493 ( .A(n694), .B(n695), .Z(n693) );
  XOR U494 ( .A(n696), .B(n697), .Z(n685) );
  AND U495 ( .A(n698), .B(n695), .Z(n697) );
  XNOR U496 ( .A(n696), .B(n692), .Z(n695) );
  XOR U497 ( .A(n699), .B(n700), .Z(n692) );
  AND U498 ( .A(n701), .B(n702), .Z(n700) );
  XOR U499 ( .A(p_input[1865]), .B(n699), .Z(n702) );
  XOR U500 ( .A(n703), .B(n704), .Z(n699) );
  AND U501 ( .A(n705), .B(n706), .Z(n704) );
  XOR U502 ( .A(n707), .B(n708), .Z(n696) );
  AND U503 ( .A(n709), .B(n706), .Z(n708) );
  XNOR U504 ( .A(n707), .B(n703), .Z(n706) );
  XOR U505 ( .A(n710), .B(n711), .Z(n703) );
  AND U506 ( .A(n712), .B(n713), .Z(n711) );
  XOR U507 ( .A(p_input[1897]), .B(n710), .Z(n713) );
  XOR U508 ( .A(n714), .B(n715), .Z(n710) );
  AND U509 ( .A(n716), .B(n717), .Z(n715) );
  XOR U510 ( .A(n718), .B(n719), .Z(n707) );
  AND U511 ( .A(n720), .B(n717), .Z(n719) );
  XNOR U512 ( .A(n718), .B(n714), .Z(n717) );
  XOR U513 ( .A(n721), .B(n722), .Z(n714) );
  AND U514 ( .A(n723), .B(n724), .Z(n722) );
  XOR U515 ( .A(p_input[1929]), .B(n721), .Z(n724) );
  XOR U516 ( .A(n725), .B(n726), .Z(n721) );
  AND U517 ( .A(n727), .B(n728), .Z(n726) );
  XOR U518 ( .A(n729), .B(n730), .Z(n718) );
  AND U519 ( .A(n731), .B(n728), .Z(n730) );
  XNOR U520 ( .A(n729), .B(n725), .Z(n728) );
  XOR U521 ( .A(n732), .B(n733), .Z(n725) );
  AND U522 ( .A(n734), .B(n735), .Z(n733) );
  XOR U523 ( .A(p_input[1961]), .B(n732), .Z(n735) );
  XNOR U524 ( .A(n736), .B(n737), .Z(n732) );
  AND U525 ( .A(n738), .B(n739), .Z(n737) );
  XNOR U526 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n740), .Z(n729) );
  AND U527 ( .A(n741), .B(n739), .Z(n740) );
  XOR U528 ( .A(n742), .B(n736), .Z(n739) );
  XOR U529 ( .A(n3), .B(n743), .Z(o[40]) );
  AND U530 ( .A(n58), .B(n744), .Z(n3) );
  XOR U531 ( .A(n4), .B(n743), .Z(n744) );
  XOR U532 ( .A(n745), .B(n746), .Z(n743) );
  AND U533 ( .A(n62), .B(n747), .Z(n746) );
  XOR U534 ( .A(p_input[8]), .B(n745), .Z(n747) );
  XOR U535 ( .A(n748), .B(n749), .Z(n745) );
  AND U536 ( .A(n66), .B(n750), .Z(n749) );
  XOR U537 ( .A(n751), .B(n752), .Z(n4) );
  AND U538 ( .A(n70), .B(n750), .Z(n752) );
  XNOR U539 ( .A(n753), .B(n748), .Z(n750) );
  XOR U540 ( .A(n754), .B(n755), .Z(n748) );
  AND U541 ( .A(n74), .B(n756), .Z(n755) );
  XOR U542 ( .A(p_input[40]), .B(n754), .Z(n756) );
  XOR U543 ( .A(n757), .B(n758), .Z(n754) );
  AND U544 ( .A(n78), .B(n759), .Z(n758) );
  IV U545 ( .A(n751), .Z(n753) );
  XNOR U546 ( .A(n760), .B(n761), .Z(n751) );
  AND U547 ( .A(n82), .B(n759), .Z(n761) );
  XNOR U548 ( .A(n760), .B(n757), .Z(n759) );
  XOR U549 ( .A(n762), .B(n763), .Z(n757) );
  AND U550 ( .A(n85), .B(n764), .Z(n763) );
  XOR U551 ( .A(p_input[72]), .B(n762), .Z(n764) );
  XOR U552 ( .A(n765), .B(n766), .Z(n762) );
  AND U553 ( .A(n89), .B(n767), .Z(n766) );
  XOR U554 ( .A(n768), .B(n769), .Z(n760) );
  AND U555 ( .A(n93), .B(n767), .Z(n769) );
  XNOR U556 ( .A(n768), .B(n765), .Z(n767) );
  XOR U557 ( .A(n770), .B(n771), .Z(n765) );
  AND U558 ( .A(n96), .B(n772), .Z(n771) );
  XOR U559 ( .A(p_input[104]), .B(n770), .Z(n772) );
  XOR U560 ( .A(n773), .B(n774), .Z(n770) );
  AND U561 ( .A(n100), .B(n775), .Z(n774) );
  XOR U562 ( .A(n776), .B(n777), .Z(n768) );
  AND U563 ( .A(n104), .B(n775), .Z(n777) );
  XNOR U564 ( .A(n776), .B(n773), .Z(n775) );
  XOR U565 ( .A(n778), .B(n779), .Z(n773) );
  AND U566 ( .A(n107), .B(n780), .Z(n779) );
  XOR U567 ( .A(p_input[136]), .B(n778), .Z(n780) );
  XOR U568 ( .A(n781), .B(n782), .Z(n778) );
  AND U569 ( .A(n111), .B(n783), .Z(n782) );
  XOR U570 ( .A(n784), .B(n785), .Z(n776) );
  AND U571 ( .A(n115), .B(n783), .Z(n785) );
  XNOR U572 ( .A(n784), .B(n781), .Z(n783) );
  XOR U573 ( .A(n786), .B(n787), .Z(n781) );
  AND U574 ( .A(n118), .B(n788), .Z(n787) );
  XOR U575 ( .A(p_input[168]), .B(n786), .Z(n788) );
  XOR U576 ( .A(n789), .B(n790), .Z(n786) );
  AND U577 ( .A(n122), .B(n791), .Z(n790) );
  XOR U578 ( .A(n792), .B(n793), .Z(n784) );
  AND U579 ( .A(n126), .B(n791), .Z(n793) );
  XNOR U580 ( .A(n792), .B(n789), .Z(n791) );
  XOR U581 ( .A(n794), .B(n795), .Z(n789) );
  AND U582 ( .A(n129), .B(n796), .Z(n795) );
  XOR U583 ( .A(p_input[200]), .B(n794), .Z(n796) );
  XOR U584 ( .A(n797), .B(n798), .Z(n794) );
  AND U585 ( .A(n133), .B(n799), .Z(n798) );
  XOR U586 ( .A(n800), .B(n801), .Z(n792) );
  AND U587 ( .A(n137), .B(n799), .Z(n801) );
  XNOR U588 ( .A(n800), .B(n797), .Z(n799) );
  XOR U589 ( .A(n802), .B(n803), .Z(n797) );
  AND U590 ( .A(n140), .B(n804), .Z(n803) );
  XOR U591 ( .A(p_input[232]), .B(n802), .Z(n804) );
  XOR U592 ( .A(n805), .B(n806), .Z(n802) );
  AND U593 ( .A(n144), .B(n807), .Z(n806) );
  XOR U594 ( .A(n808), .B(n809), .Z(n800) );
  AND U595 ( .A(n148), .B(n807), .Z(n809) );
  XNOR U596 ( .A(n808), .B(n805), .Z(n807) );
  XOR U597 ( .A(n810), .B(n811), .Z(n805) );
  AND U598 ( .A(n151), .B(n812), .Z(n811) );
  XOR U599 ( .A(p_input[264]), .B(n810), .Z(n812) );
  XOR U600 ( .A(n813), .B(n814), .Z(n810) );
  AND U601 ( .A(n155), .B(n815), .Z(n814) );
  XOR U602 ( .A(n816), .B(n817), .Z(n808) );
  AND U603 ( .A(n159), .B(n815), .Z(n817) );
  XNOR U604 ( .A(n816), .B(n813), .Z(n815) );
  XOR U605 ( .A(n818), .B(n819), .Z(n813) );
  AND U606 ( .A(n162), .B(n820), .Z(n819) );
  XOR U607 ( .A(p_input[296]), .B(n818), .Z(n820) );
  XOR U608 ( .A(n821), .B(n822), .Z(n818) );
  AND U609 ( .A(n166), .B(n823), .Z(n822) );
  XOR U610 ( .A(n824), .B(n825), .Z(n816) );
  AND U611 ( .A(n170), .B(n823), .Z(n825) );
  XNOR U612 ( .A(n824), .B(n821), .Z(n823) );
  XOR U613 ( .A(n826), .B(n827), .Z(n821) );
  AND U614 ( .A(n173), .B(n828), .Z(n827) );
  XOR U615 ( .A(p_input[328]), .B(n826), .Z(n828) );
  XOR U616 ( .A(n829), .B(n830), .Z(n826) );
  AND U617 ( .A(n177), .B(n831), .Z(n830) );
  XOR U618 ( .A(n832), .B(n833), .Z(n824) );
  AND U619 ( .A(n181), .B(n831), .Z(n833) );
  XNOR U620 ( .A(n832), .B(n829), .Z(n831) );
  XOR U621 ( .A(n834), .B(n835), .Z(n829) );
  AND U622 ( .A(n184), .B(n836), .Z(n835) );
  XOR U623 ( .A(p_input[360]), .B(n834), .Z(n836) );
  XOR U624 ( .A(n837), .B(n838), .Z(n834) );
  AND U625 ( .A(n188), .B(n839), .Z(n838) );
  XOR U626 ( .A(n840), .B(n841), .Z(n832) );
  AND U627 ( .A(n192), .B(n839), .Z(n841) );
  XNOR U628 ( .A(n840), .B(n837), .Z(n839) );
  XOR U629 ( .A(n842), .B(n843), .Z(n837) );
  AND U630 ( .A(n195), .B(n844), .Z(n843) );
  XOR U631 ( .A(p_input[392]), .B(n842), .Z(n844) );
  XOR U632 ( .A(n845), .B(n846), .Z(n842) );
  AND U633 ( .A(n199), .B(n847), .Z(n846) );
  XOR U634 ( .A(n848), .B(n849), .Z(n840) );
  AND U635 ( .A(n203), .B(n847), .Z(n849) );
  XNOR U636 ( .A(n848), .B(n845), .Z(n847) );
  XOR U637 ( .A(n850), .B(n851), .Z(n845) );
  AND U638 ( .A(n206), .B(n852), .Z(n851) );
  XOR U639 ( .A(p_input[424]), .B(n850), .Z(n852) );
  XOR U640 ( .A(n853), .B(n854), .Z(n850) );
  AND U641 ( .A(n210), .B(n855), .Z(n854) );
  XOR U642 ( .A(n856), .B(n857), .Z(n848) );
  AND U643 ( .A(n214), .B(n855), .Z(n857) );
  XNOR U644 ( .A(n856), .B(n853), .Z(n855) );
  XOR U645 ( .A(n858), .B(n859), .Z(n853) );
  AND U646 ( .A(n217), .B(n860), .Z(n859) );
  XOR U647 ( .A(p_input[456]), .B(n858), .Z(n860) );
  XOR U648 ( .A(n861), .B(n862), .Z(n858) );
  AND U649 ( .A(n221), .B(n863), .Z(n862) );
  XOR U650 ( .A(n864), .B(n865), .Z(n856) );
  AND U651 ( .A(n225), .B(n863), .Z(n865) );
  XNOR U652 ( .A(n864), .B(n861), .Z(n863) );
  XOR U653 ( .A(n866), .B(n867), .Z(n861) );
  AND U654 ( .A(n228), .B(n868), .Z(n867) );
  XOR U655 ( .A(p_input[488]), .B(n866), .Z(n868) );
  XOR U656 ( .A(n869), .B(n870), .Z(n866) );
  AND U657 ( .A(n232), .B(n871), .Z(n870) );
  XOR U658 ( .A(n872), .B(n873), .Z(n864) );
  AND U659 ( .A(n236), .B(n871), .Z(n873) );
  XNOR U660 ( .A(n872), .B(n869), .Z(n871) );
  XOR U661 ( .A(n874), .B(n875), .Z(n869) );
  AND U662 ( .A(n239), .B(n876), .Z(n875) );
  XOR U663 ( .A(p_input[520]), .B(n874), .Z(n876) );
  XOR U664 ( .A(n877), .B(n878), .Z(n874) );
  AND U665 ( .A(n243), .B(n879), .Z(n878) );
  XOR U666 ( .A(n880), .B(n881), .Z(n872) );
  AND U667 ( .A(n247), .B(n879), .Z(n881) );
  XNOR U668 ( .A(n880), .B(n877), .Z(n879) );
  XOR U669 ( .A(n882), .B(n883), .Z(n877) );
  AND U670 ( .A(n250), .B(n884), .Z(n883) );
  XOR U671 ( .A(p_input[552]), .B(n882), .Z(n884) );
  XOR U672 ( .A(n885), .B(n886), .Z(n882) );
  AND U673 ( .A(n254), .B(n887), .Z(n886) );
  XOR U674 ( .A(n888), .B(n889), .Z(n880) );
  AND U675 ( .A(n258), .B(n887), .Z(n889) );
  XNOR U676 ( .A(n888), .B(n885), .Z(n887) );
  XOR U677 ( .A(n890), .B(n891), .Z(n885) );
  AND U678 ( .A(n261), .B(n892), .Z(n891) );
  XOR U679 ( .A(p_input[584]), .B(n890), .Z(n892) );
  XOR U680 ( .A(n893), .B(n894), .Z(n890) );
  AND U681 ( .A(n265), .B(n895), .Z(n894) );
  XOR U682 ( .A(n896), .B(n897), .Z(n888) );
  AND U683 ( .A(n269), .B(n895), .Z(n897) );
  XNOR U684 ( .A(n896), .B(n893), .Z(n895) );
  XOR U685 ( .A(n898), .B(n899), .Z(n893) );
  AND U686 ( .A(n272), .B(n900), .Z(n899) );
  XOR U687 ( .A(p_input[616]), .B(n898), .Z(n900) );
  XOR U688 ( .A(n901), .B(n902), .Z(n898) );
  AND U689 ( .A(n276), .B(n903), .Z(n902) );
  XOR U690 ( .A(n904), .B(n905), .Z(n896) );
  AND U691 ( .A(n280), .B(n903), .Z(n905) );
  XNOR U692 ( .A(n904), .B(n901), .Z(n903) );
  XOR U693 ( .A(n906), .B(n907), .Z(n901) );
  AND U694 ( .A(n283), .B(n908), .Z(n907) );
  XOR U695 ( .A(p_input[648]), .B(n906), .Z(n908) );
  XOR U696 ( .A(n909), .B(n910), .Z(n906) );
  AND U697 ( .A(n287), .B(n911), .Z(n910) );
  XOR U698 ( .A(n912), .B(n913), .Z(n904) );
  AND U699 ( .A(n291), .B(n911), .Z(n913) );
  XNOR U700 ( .A(n912), .B(n909), .Z(n911) );
  XOR U701 ( .A(n914), .B(n915), .Z(n909) );
  AND U702 ( .A(n294), .B(n916), .Z(n915) );
  XOR U703 ( .A(p_input[680]), .B(n914), .Z(n916) );
  XOR U704 ( .A(n917), .B(n918), .Z(n914) );
  AND U705 ( .A(n298), .B(n919), .Z(n918) );
  XOR U706 ( .A(n920), .B(n921), .Z(n912) );
  AND U707 ( .A(n302), .B(n919), .Z(n921) );
  XNOR U708 ( .A(n920), .B(n917), .Z(n919) );
  XOR U709 ( .A(n922), .B(n923), .Z(n917) );
  AND U710 ( .A(n305), .B(n924), .Z(n923) );
  XOR U711 ( .A(p_input[712]), .B(n922), .Z(n924) );
  XOR U712 ( .A(n925), .B(n926), .Z(n922) );
  AND U713 ( .A(n309), .B(n927), .Z(n926) );
  XOR U714 ( .A(n928), .B(n929), .Z(n920) );
  AND U715 ( .A(n313), .B(n927), .Z(n929) );
  XNOR U716 ( .A(n928), .B(n925), .Z(n927) );
  XOR U717 ( .A(n930), .B(n931), .Z(n925) );
  AND U718 ( .A(n316), .B(n932), .Z(n931) );
  XOR U719 ( .A(p_input[744]), .B(n930), .Z(n932) );
  XOR U720 ( .A(n933), .B(n934), .Z(n930) );
  AND U721 ( .A(n320), .B(n935), .Z(n934) );
  XOR U722 ( .A(n936), .B(n937), .Z(n928) );
  AND U723 ( .A(n324), .B(n935), .Z(n937) );
  XNOR U724 ( .A(n936), .B(n933), .Z(n935) );
  XOR U725 ( .A(n938), .B(n939), .Z(n933) );
  AND U726 ( .A(n327), .B(n940), .Z(n939) );
  XOR U727 ( .A(p_input[776]), .B(n938), .Z(n940) );
  XOR U728 ( .A(n941), .B(n942), .Z(n938) );
  AND U729 ( .A(n331), .B(n943), .Z(n942) );
  XOR U730 ( .A(n944), .B(n945), .Z(n936) );
  AND U731 ( .A(n335), .B(n943), .Z(n945) );
  XNOR U732 ( .A(n944), .B(n941), .Z(n943) );
  XOR U733 ( .A(n946), .B(n947), .Z(n941) );
  AND U734 ( .A(n338), .B(n948), .Z(n947) );
  XOR U735 ( .A(p_input[808]), .B(n946), .Z(n948) );
  XOR U736 ( .A(n949), .B(n950), .Z(n946) );
  AND U737 ( .A(n342), .B(n951), .Z(n950) );
  XOR U738 ( .A(n952), .B(n953), .Z(n944) );
  AND U739 ( .A(n346), .B(n951), .Z(n953) );
  XNOR U740 ( .A(n952), .B(n949), .Z(n951) );
  XOR U741 ( .A(n954), .B(n955), .Z(n949) );
  AND U742 ( .A(n349), .B(n956), .Z(n955) );
  XOR U743 ( .A(p_input[840]), .B(n954), .Z(n956) );
  XOR U744 ( .A(n957), .B(n958), .Z(n954) );
  AND U745 ( .A(n353), .B(n959), .Z(n958) );
  XOR U746 ( .A(n960), .B(n961), .Z(n952) );
  AND U747 ( .A(n357), .B(n959), .Z(n961) );
  XNOR U748 ( .A(n960), .B(n957), .Z(n959) );
  XOR U749 ( .A(n962), .B(n963), .Z(n957) );
  AND U750 ( .A(n360), .B(n964), .Z(n963) );
  XOR U751 ( .A(p_input[872]), .B(n962), .Z(n964) );
  XOR U752 ( .A(n965), .B(n966), .Z(n962) );
  AND U753 ( .A(n364), .B(n967), .Z(n966) );
  XOR U754 ( .A(n968), .B(n969), .Z(n960) );
  AND U755 ( .A(n368), .B(n967), .Z(n969) );
  XNOR U756 ( .A(n968), .B(n965), .Z(n967) );
  XOR U757 ( .A(n970), .B(n971), .Z(n965) );
  AND U758 ( .A(n371), .B(n972), .Z(n971) );
  XOR U759 ( .A(p_input[904]), .B(n970), .Z(n972) );
  XOR U760 ( .A(n973), .B(n974), .Z(n970) );
  AND U761 ( .A(n375), .B(n975), .Z(n974) );
  XOR U762 ( .A(n976), .B(n977), .Z(n968) );
  AND U763 ( .A(n379), .B(n975), .Z(n977) );
  XNOR U764 ( .A(n976), .B(n973), .Z(n975) );
  XOR U765 ( .A(n978), .B(n979), .Z(n973) );
  AND U766 ( .A(n382), .B(n980), .Z(n979) );
  XOR U767 ( .A(p_input[936]), .B(n978), .Z(n980) );
  XOR U768 ( .A(n981), .B(n982), .Z(n978) );
  AND U769 ( .A(n386), .B(n983), .Z(n982) );
  XOR U770 ( .A(n984), .B(n985), .Z(n976) );
  AND U771 ( .A(n390), .B(n983), .Z(n985) );
  XNOR U772 ( .A(n984), .B(n981), .Z(n983) );
  XOR U773 ( .A(n986), .B(n987), .Z(n981) );
  AND U774 ( .A(n393), .B(n988), .Z(n987) );
  XOR U775 ( .A(p_input[968]), .B(n986), .Z(n988) );
  XOR U776 ( .A(n989), .B(n990), .Z(n986) );
  AND U777 ( .A(n397), .B(n991), .Z(n990) );
  XOR U778 ( .A(n992), .B(n993), .Z(n984) );
  AND U779 ( .A(n401), .B(n991), .Z(n993) );
  XNOR U780 ( .A(n992), .B(n989), .Z(n991) );
  XOR U781 ( .A(n994), .B(n995), .Z(n989) );
  AND U782 ( .A(n404), .B(n996), .Z(n995) );
  XOR U783 ( .A(p_input[1000]), .B(n994), .Z(n996) );
  XOR U784 ( .A(n997), .B(n998), .Z(n994) );
  AND U785 ( .A(n408), .B(n999), .Z(n998) );
  XOR U786 ( .A(n1000), .B(n1001), .Z(n992) );
  AND U787 ( .A(n412), .B(n999), .Z(n1001) );
  XNOR U788 ( .A(n1000), .B(n997), .Z(n999) );
  XOR U789 ( .A(n1002), .B(n1003), .Z(n997) );
  AND U790 ( .A(n415), .B(n1004), .Z(n1003) );
  XOR U791 ( .A(p_input[1032]), .B(n1002), .Z(n1004) );
  XOR U792 ( .A(n1005), .B(n1006), .Z(n1002) );
  AND U793 ( .A(n419), .B(n1007), .Z(n1006) );
  XOR U794 ( .A(n1008), .B(n1009), .Z(n1000) );
  AND U795 ( .A(n423), .B(n1007), .Z(n1009) );
  XNOR U796 ( .A(n1008), .B(n1005), .Z(n1007) );
  XOR U797 ( .A(n1010), .B(n1011), .Z(n1005) );
  AND U798 ( .A(n426), .B(n1012), .Z(n1011) );
  XOR U799 ( .A(p_input[1064]), .B(n1010), .Z(n1012) );
  XOR U800 ( .A(n1013), .B(n1014), .Z(n1010) );
  AND U801 ( .A(n430), .B(n1015), .Z(n1014) );
  XOR U802 ( .A(n1016), .B(n1017), .Z(n1008) );
  AND U803 ( .A(n434), .B(n1015), .Z(n1017) );
  XNOR U804 ( .A(n1016), .B(n1013), .Z(n1015) );
  XOR U805 ( .A(n1018), .B(n1019), .Z(n1013) );
  AND U806 ( .A(n437), .B(n1020), .Z(n1019) );
  XOR U807 ( .A(p_input[1096]), .B(n1018), .Z(n1020) );
  XOR U808 ( .A(n1021), .B(n1022), .Z(n1018) );
  AND U809 ( .A(n441), .B(n1023), .Z(n1022) );
  XOR U810 ( .A(n1024), .B(n1025), .Z(n1016) );
  AND U811 ( .A(n445), .B(n1023), .Z(n1025) );
  XNOR U812 ( .A(n1024), .B(n1021), .Z(n1023) );
  XOR U813 ( .A(n1026), .B(n1027), .Z(n1021) );
  AND U814 ( .A(n448), .B(n1028), .Z(n1027) );
  XOR U815 ( .A(p_input[1128]), .B(n1026), .Z(n1028) );
  XOR U816 ( .A(n1029), .B(n1030), .Z(n1026) );
  AND U817 ( .A(n452), .B(n1031), .Z(n1030) );
  XOR U818 ( .A(n1032), .B(n1033), .Z(n1024) );
  AND U819 ( .A(n456), .B(n1031), .Z(n1033) );
  XNOR U820 ( .A(n1032), .B(n1029), .Z(n1031) );
  XOR U821 ( .A(n1034), .B(n1035), .Z(n1029) );
  AND U822 ( .A(n459), .B(n1036), .Z(n1035) );
  XOR U823 ( .A(p_input[1160]), .B(n1034), .Z(n1036) );
  XOR U824 ( .A(n1037), .B(n1038), .Z(n1034) );
  AND U825 ( .A(n463), .B(n1039), .Z(n1038) );
  XOR U826 ( .A(n1040), .B(n1041), .Z(n1032) );
  AND U827 ( .A(n467), .B(n1039), .Z(n1041) );
  XNOR U828 ( .A(n1040), .B(n1037), .Z(n1039) );
  XOR U829 ( .A(n1042), .B(n1043), .Z(n1037) );
  AND U830 ( .A(n470), .B(n1044), .Z(n1043) );
  XOR U831 ( .A(p_input[1192]), .B(n1042), .Z(n1044) );
  XOR U832 ( .A(n1045), .B(n1046), .Z(n1042) );
  AND U833 ( .A(n474), .B(n1047), .Z(n1046) );
  XOR U834 ( .A(n1048), .B(n1049), .Z(n1040) );
  AND U835 ( .A(n478), .B(n1047), .Z(n1049) );
  XNOR U836 ( .A(n1048), .B(n1045), .Z(n1047) );
  XOR U837 ( .A(n1050), .B(n1051), .Z(n1045) );
  AND U838 ( .A(n481), .B(n1052), .Z(n1051) );
  XOR U839 ( .A(p_input[1224]), .B(n1050), .Z(n1052) );
  XOR U840 ( .A(n1053), .B(n1054), .Z(n1050) );
  AND U841 ( .A(n485), .B(n1055), .Z(n1054) );
  XOR U842 ( .A(n1056), .B(n1057), .Z(n1048) );
  AND U843 ( .A(n489), .B(n1055), .Z(n1057) );
  XNOR U844 ( .A(n1056), .B(n1053), .Z(n1055) );
  XOR U845 ( .A(n1058), .B(n1059), .Z(n1053) );
  AND U846 ( .A(n492), .B(n1060), .Z(n1059) );
  XOR U847 ( .A(p_input[1256]), .B(n1058), .Z(n1060) );
  XOR U848 ( .A(n1061), .B(n1062), .Z(n1058) );
  AND U849 ( .A(n496), .B(n1063), .Z(n1062) );
  XOR U850 ( .A(n1064), .B(n1065), .Z(n1056) );
  AND U851 ( .A(n500), .B(n1063), .Z(n1065) );
  XNOR U852 ( .A(n1064), .B(n1061), .Z(n1063) );
  XOR U853 ( .A(n1066), .B(n1067), .Z(n1061) );
  AND U854 ( .A(n503), .B(n1068), .Z(n1067) );
  XOR U855 ( .A(p_input[1288]), .B(n1066), .Z(n1068) );
  XOR U856 ( .A(n1069), .B(n1070), .Z(n1066) );
  AND U857 ( .A(n507), .B(n1071), .Z(n1070) );
  XOR U858 ( .A(n1072), .B(n1073), .Z(n1064) );
  AND U859 ( .A(n511), .B(n1071), .Z(n1073) );
  XNOR U860 ( .A(n1072), .B(n1069), .Z(n1071) );
  XOR U861 ( .A(n1074), .B(n1075), .Z(n1069) );
  AND U862 ( .A(n514), .B(n1076), .Z(n1075) );
  XOR U863 ( .A(p_input[1320]), .B(n1074), .Z(n1076) );
  XOR U864 ( .A(n1077), .B(n1078), .Z(n1074) );
  AND U865 ( .A(n518), .B(n1079), .Z(n1078) );
  XOR U866 ( .A(n1080), .B(n1081), .Z(n1072) );
  AND U867 ( .A(n522), .B(n1079), .Z(n1081) );
  XNOR U868 ( .A(n1080), .B(n1077), .Z(n1079) );
  XOR U869 ( .A(n1082), .B(n1083), .Z(n1077) );
  AND U870 ( .A(n525), .B(n1084), .Z(n1083) );
  XOR U871 ( .A(p_input[1352]), .B(n1082), .Z(n1084) );
  XOR U872 ( .A(n1085), .B(n1086), .Z(n1082) );
  AND U873 ( .A(n529), .B(n1087), .Z(n1086) );
  XOR U874 ( .A(n1088), .B(n1089), .Z(n1080) );
  AND U875 ( .A(n533), .B(n1087), .Z(n1089) );
  XNOR U876 ( .A(n1088), .B(n1085), .Z(n1087) );
  XOR U877 ( .A(n1090), .B(n1091), .Z(n1085) );
  AND U878 ( .A(n536), .B(n1092), .Z(n1091) );
  XOR U879 ( .A(p_input[1384]), .B(n1090), .Z(n1092) );
  XOR U880 ( .A(n1093), .B(n1094), .Z(n1090) );
  AND U881 ( .A(n540), .B(n1095), .Z(n1094) );
  XOR U882 ( .A(n1096), .B(n1097), .Z(n1088) );
  AND U883 ( .A(n544), .B(n1095), .Z(n1097) );
  XNOR U884 ( .A(n1096), .B(n1093), .Z(n1095) );
  XOR U885 ( .A(n1098), .B(n1099), .Z(n1093) );
  AND U886 ( .A(n547), .B(n1100), .Z(n1099) );
  XOR U887 ( .A(p_input[1416]), .B(n1098), .Z(n1100) );
  XOR U888 ( .A(n1101), .B(n1102), .Z(n1098) );
  AND U889 ( .A(n551), .B(n1103), .Z(n1102) );
  XOR U890 ( .A(n1104), .B(n1105), .Z(n1096) );
  AND U891 ( .A(n555), .B(n1103), .Z(n1105) );
  XNOR U892 ( .A(n1104), .B(n1101), .Z(n1103) );
  XOR U893 ( .A(n1106), .B(n1107), .Z(n1101) );
  AND U894 ( .A(n558), .B(n1108), .Z(n1107) );
  XOR U895 ( .A(p_input[1448]), .B(n1106), .Z(n1108) );
  XOR U896 ( .A(n1109), .B(n1110), .Z(n1106) );
  AND U897 ( .A(n562), .B(n1111), .Z(n1110) );
  XOR U898 ( .A(n1112), .B(n1113), .Z(n1104) );
  AND U899 ( .A(n566), .B(n1111), .Z(n1113) );
  XNOR U900 ( .A(n1112), .B(n1109), .Z(n1111) );
  XOR U901 ( .A(n1114), .B(n1115), .Z(n1109) );
  AND U902 ( .A(n569), .B(n1116), .Z(n1115) );
  XOR U903 ( .A(p_input[1480]), .B(n1114), .Z(n1116) );
  XOR U904 ( .A(n1117), .B(n1118), .Z(n1114) );
  AND U905 ( .A(n573), .B(n1119), .Z(n1118) );
  XOR U906 ( .A(n1120), .B(n1121), .Z(n1112) );
  AND U907 ( .A(n577), .B(n1119), .Z(n1121) );
  XNOR U908 ( .A(n1120), .B(n1117), .Z(n1119) );
  XOR U909 ( .A(n1122), .B(n1123), .Z(n1117) );
  AND U910 ( .A(n580), .B(n1124), .Z(n1123) );
  XOR U911 ( .A(p_input[1512]), .B(n1122), .Z(n1124) );
  XOR U912 ( .A(n1125), .B(n1126), .Z(n1122) );
  AND U913 ( .A(n584), .B(n1127), .Z(n1126) );
  XOR U914 ( .A(n1128), .B(n1129), .Z(n1120) );
  AND U915 ( .A(n588), .B(n1127), .Z(n1129) );
  XNOR U916 ( .A(n1128), .B(n1125), .Z(n1127) );
  XOR U917 ( .A(n1130), .B(n1131), .Z(n1125) );
  AND U918 ( .A(n591), .B(n1132), .Z(n1131) );
  XOR U919 ( .A(p_input[1544]), .B(n1130), .Z(n1132) );
  XOR U920 ( .A(n1133), .B(n1134), .Z(n1130) );
  AND U921 ( .A(n595), .B(n1135), .Z(n1134) );
  XOR U922 ( .A(n1136), .B(n1137), .Z(n1128) );
  AND U923 ( .A(n599), .B(n1135), .Z(n1137) );
  XNOR U924 ( .A(n1136), .B(n1133), .Z(n1135) );
  XOR U925 ( .A(n1138), .B(n1139), .Z(n1133) );
  AND U926 ( .A(n602), .B(n1140), .Z(n1139) );
  XOR U927 ( .A(p_input[1576]), .B(n1138), .Z(n1140) );
  XOR U928 ( .A(n1141), .B(n1142), .Z(n1138) );
  AND U929 ( .A(n606), .B(n1143), .Z(n1142) );
  XOR U930 ( .A(n1144), .B(n1145), .Z(n1136) );
  AND U931 ( .A(n610), .B(n1143), .Z(n1145) );
  XNOR U932 ( .A(n1144), .B(n1141), .Z(n1143) );
  XOR U933 ( .A(n1146), .B(n1147), .Z(n1141) );
  AND U934 ( .A(n613), .B(n1148), .Z(n1147) );
  XOR U935 ( .A(p_input[1608]), .B(n1146), .Z(n1148) );
  XOR U936 ( .A(n1149), .B(n1150), .Z(n1146) );
  AND U937 ( .A(n617), .B(n1151), .Z(n1150) );
  XOR U938 ( .A(n1152), .B(n1153), .Z(n1144) );
  AND U939 ( .A(n621), .B(n1151), .Z(n1153) );
  XNOR U940 ( .A(n1152), .B(n1149), .Z(n1151) );
  XOR U941 ( .A(n1154), .B(n1155), .Z(n1149) );
  AND U942 ( .A(n624), .B(n1156), .Z(n1155) );
  XOR U943 ( .A(p_input[1640]), .B(n1154), .Z(n1156) );
  XOR U944 ( .A(n1157), .B(n1158), .Z(n1154) );
  AND U945 ( .A(n628), .B(n1159), .Z(n1158) );
  XOR U946 ( .A(n1160), .B(n1161), .Z(n1152) );
  AND U947 ( .A(n632), .B(n1159), .Z(n1161) );
  XNOR U948 ( .A(n1160), .B(n1157), .Z(n1159) );
  XOR U949 ( .A(n1162), .B(n1163), .Z(n1157) );
  AND U950 ( .A(n635), .B(n1164), .Z(n1163) );
  XOR U951 ( .A(p_input[1672]), .B(n1162), .Z(n1164) );
  XOR U952 ( .A(n1165), .B(n1166), .Z(n1162) );
  AND U953 ( .A(n639), .B(n1167), .Z(n1166) );
  XOR U954 ( .A(n1168), .B(n1169), .Z(n1160) );
  AND U955 ( .A(n643), .B(n1167), .Z(n1169) );
  XNOR U956 ( .A(n1168), .B(n1165), .Z(n1167) );
  XOR U957 ( .A(n1170), .B(n1171), .Z(n1165) );
  AND U958 ( .A(n646), .B(n1172), .Z(n1171) );
  XOR U959 ( .A(p_input[1704]), .B(n1170), .Z(n1172) );
  XOR U960 ( .A(n1173), .B(n1174), .Z(n1170) );
  AND U961 ( .A(n650), .B(n1175), .Z(n1174) );
  XOR U962 ( .A(n1176), .B(n1177), .Z(n1168) );
  AND U963 ( .A(n654), .B(n1175), .Z(n1177) );
  XNOR U964 ( .A(n1176), .B(n1173), .Z(n1175) );
  XOR U965 ( .A(n1178), .B(n1179), .Z(n1173) );
  AND U966 ( .A(n657), .B(n1180), .Z(n1179) );
  XOR U967 ( .A(p_input[1736]), .B(n1178), .Z(n1180) );
  XOR U968 ( .A(n1181), .B(n1182), .Z(n1178) );
  AND U969 ( .A(n661), .B(n1183), .Z(n1182) );
  XOR U970 ( .A(n1184), .B(n1185), .Z(n1176) );
  AND U971 ( .A(n665), .B(n1183), .Z(n1185) );
  XNOR U972 ( .A(n1184), .B(n1181), .Z(n1183) );
  XOR U973 ( .A(n1186), .B(n1187), .Z(n1181) );
  AND U974 ( .A(n668), .B(n1188), .Z(n1187) );
  XOR U975 ( .A(p_input[1768]), .B(n1186), .Z(n1188) );
  XOR U976 ( .A(n1189), .B(n1190), .Z(n1186) );
  AND U977 ( .A(n672), .B(n1191), .Z(n1190) );
  XOR U978 ( .A(n1192), .B(n1193), .Z(n1184) );
  AND U979 ( .A(n676), .B(n1191), .Z(n1193) );
  XNOR U980 ( .A(n1192), .B(n1189), .Z(n1191) );
  XOR U981 ( .A(n1194), .B(n1195), .Z(n1189) );
  AND U982 ( .A(n679), .B(n1196), .Z(n1195) );
  XOR U983 ( .A(p_input[1800]), .B(n1194), .Z(n1196) );
  XOR U984 ( .A(n1197), .B(n1198), .Z(n1194) );
  AND U985 ( .A(n683), .B(n1199), .Z(n1198) );
  XOR U986 ( .A(n1200), .B(n1201), .Z(n1192) );
  AND U987 ( .A(n687), .B(n1199), .Z(n1201) );
  XNOR U988 ( .A(n1200), .B(n1197), .Z(n1199) );
  XOR U989 ( .A(n1202), .B(n1203), .Z(n1197) );
  AND U990 ( .A(n690), .B(n1204), .Z(n1203) );
  XOR U991 ( .A(p_input[1832]), .B(n1202), .Z(n1204) );
  XOR U992 ( .A(n1205), .B(n1206), .Z(n1202) );
  AND U993 ( .A(n694), .B(n1207), .Z(n1206) );
  XOR U994 ( .A(n1208), .B(n1209), .Z(n1200) );
  AND U995 ( .A(n698), .B(n1207), .Z(n1209) );
  XNOR U996 ( .A(n1208), .B(n1205), .Z(n1207) );
  XOR U997 ( .A(n1210), .B(n1211), .Z(n1205) );
  AND U998 ( .A(n701), .B(n1212), .Z(n1211) );
  XOR U999 ( .A(p_input[1864]), .B(n1210), .Z(n1212) );
  XOR U1000 ( .A(n1213), .B(n1214), .Z(n1210) );
  AND U1001 ( .A(n705), .B(n1215), .Z(n1214) );
  XOR U1002 ( .A(n1216), .B(n1217), .Z(n1208) );
  AND U1003 ( .A(n709), .B(n1215), .Z(n1217) );
  XNOR U1004 ( .A(n1216), .B(n1213), .Z(n1215) );
  XOR U1005 ( .A(n1218), .B(n1219), .Z(n1213) );
  AND U1006 ( .A(n712), .B(n1220), .Z(n1219) );
  XOR U1007 ( .A(p_input[1896]), .B(n1218), .Z(n1220) );
  XOR U1008 ( .A(n1221), .B(n1222), .Z(n1218) );
  AND U1009 ( .A(n716), .B(n1223), .Z(n1222) );
  XOR U1010 ( .A(n1224), .B(n1225), .Z(n1216) );
  AND U1011 ( .A(n720), .B(n1223), .Z(n1225) );
  XNOR U1012 ( .A(n1224), .B(n1221), .Z(n1223) );
  XOR U1013 ( .A(n1226), .B(n1227), .Z(n1221) );
  AND U1014 ( .A(n723), .B(n1228), .Z(n1227) );
  XOR U1015 ( .A(p_input[1928]), .B(n1226), .Z(n1228) );
  XOR U1016 ( .A(n1229), .B(n1230), .Z(n1226) );
  AND U1017 ( .A(n727), .B(n1231), .Z(n1230) );
  XOR U1018 ( .A(n1232), .B(n1233), .Z(n1224) );
  AND U1019 ( .A(n731), .B(n1231), .Z(n1233) );
  XNOR U1020 ( .A(n1232), .B(n1229), .Z(n1231) );
  XOR U1021 ( .A(n1234), .B(n1235), .Z(n1229) );
  AND U1022 ( .A(n734), .B(n1236), .Z(n1235) );
  XOR U1023 ( .A(p_input[1960]), .B(n1234), .Z(n1236) );
  XNOR U1024 ( .A(n1237), .B(n1238), .Z(n1234) );
  AND U1025 ( .A(n738), .B(n1239), .Z(n1238) );
  XNOR U1026 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n1240), .Z(n1232) );
  AND U1027 ( .A(n741), .B(n1239), .Z(n1240) );
  XOR U1028 ( .A(n1241), .B(n1237), .Z(n1239) );
  IV U1029 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .Z(n1237) );
  IV U1030 ( .A(\knn_comb_/min_val_out[0][8] ), .Z(n1241) );
  XOR U1031 ( .A(n1242), .B(n1243), .Z(o[3]) );
  XOR U1032 ( .A(n5), .B(n1244), .Z(o[39]) );
  AND U1033 ( .A(n58), .B(n1245), .Z(n5) );
  XOR U1034 ( .A(n6), .B(n1244), .Z(n1245) );
  XOR U1035 ( .A(n1246), .B(n1247), .Z(n1244) );
  AND U1036 ( .A(n62), .B(n1248), .Z(n1247) );
  XOR U1037 ( .A(p_input[7]), .B(n1246), .Z(n1248) );
  XOR U1038 ( .A(n1249), .B(n1250), .Z(n1246) );
  AND U1039 ( .A(n66), .B(n1251), .Z(n1250) );
  XOR U1040 ( .A(n1252), .B(n1253), .Z(n6) );
  AND U1041 ( .A(n70), .B(n1251), .Z(n1253) );
  XNOR U1042 ( .A(n1254), .B(n1249), .Z(n1251) );
  XOR U1043 ( .A(n1255), .B(n1256), .Z(n1249) );
  AND U1044 ( .A(n74), .B(n1257), .Z(n1256) );
  XOR U1045 ( .A(p_input[39]), .B(n1255), .Z(n1257) );
  XOR U1046 ( .A(n1258), .B(n1259), .Z(n1255) );
  AND U1047 ( .A(n78), .B(n1260), .Z(n1259) );
  IV U1048 ( .A(n1252), .Z(n1254) );
  XNOR U1049 ( .A(n1261), .B(n1262), .Z(n1252) );
  AND U1050 ( .A(n82), .B(n1260), .Z(n1262) );
  XNOR U1051 ( .A(n1261), .B(n1258), .Z(n1260) );
  XOR U1052 ( .A(n1263), .B(n1264), .Z(n1258) );
  AND U1053 ( .A(n85), .B(n1265), .Z(n1264) );
  XOR U1054 ( .A(p_input[71]), .B(n1263), .Z(n1265) );
  XOR U1055 ( .A(n1266), .B(n1267), .Z(n1263) );
  AND U1056 ( .A(n89), .B(n1268), .Z(n1267) );
  XOR U1057 ( .A(n1269), .B(n1270), .Z(n1261) );
  AND U1058 ( .A(n93), .B(n1268), .Z(n1270) );
  XNOR U1059 ( .A(n1269), .B(n1266), .Z(n1268) );
  XOR U1060 ( .A(n1271), .B(n1272), .Z(n1266) );
  AND U1061 ( .A(n96), .B(n1273), .Z(n1272) );
  XOR U1062 ( .A(p_input[103]), .B(n1271), .Z(n1273) );
  XOR U1063 ( .A(n1274), .B(n1275), .Z(n1271) );
  AND U1064 ( .A(n100), .B(n1276), .Z(n1275) );
  XOR U1065 ( .A(n1277), .B(n1278), .Z(n1269) );
  AND U1066 ( .A(n104), .B(n1276), .Z(n1278) );
  XNOR U1067 ( .A(n1277), .B(n1274), .Z(n1276) );
  XOR U1068 ( .A(n1279), .B(n1280), .Z(n1274) );
  AND U1069 ( .A(n107), .B(n1281), .Z(n1280) );
  XOR U1070 ( .A(p_input[135]), .B(n1279), .Z(n1281) );
  XOR U1071 ( .A(n1282), .B(n1283), .Z(n1279) );
  AND U1072 ( .A(n111), .B(n1284), .Z(n1283) );
  XOR U1073 ( .A(n1285), .B(n1286), .Z(n1277) );
  AND U1074 ( .A(n115), .B(n1284), .Z(n1286) );
  XNOR U1075 ( .A(n1285), .B(n1282), .Z(n1284) );
  XOR U1076 ( .A(n1287), .B(n1288), .Z(n1282) );
  AND U1077 ( .A(n118), .B(n1289), .Z(n1288) );
  XOR U1078 ( .A(p_input[167]), .B(n1287), .Z(n1289) );
  XOR U1079 ( .A(n1290), .B(n1291), .Z(n1287) );
  AND U1080 ( .A(n122), .B(n1292), .Z(n1291) );
  XOR U1081 ( .A(n1293), .B(n1294), .Z(n1285) );
  AND U1082 ( .A(n126), .B(n1292), .Z(n1294) );
  XNOR U1083 ( .A(n1293), .B(n1290), .Z(n1292) );
  XOR U1084 ( .A(n1295), .B(n1296), .Z(n1290) );
  AND U1085 ( .A(n129), .B(n1297), .Z(n1296) );
  XOR U1086 ( .A(p_input[199]), .B(n1295), .Z(n1297) );
  XOR U1087 ( .A(n1298), .B(n1299), .Z(n1295) );
  AND U1088 ( .A(n133), .B(n1300), .Z(n1299) );
  XOR U1089 ( .A(n1301), .B(n1302), .Z(n1293) );
  AND U1090 ( .A(n137), .B(n1300), .Z(n1302) );
  XNOR U1091 ( .A(n1301), .B(n1298), .Z(n1300) );
  XOR U1092 ( .A(n1303), .B(n1304), .Z(n1298) );
  AND U1093 ( .A(n140), .B(n1305), .Z(n1304) );
  XOR U1094 ( .A(p_input[231]), .B(n1303), .Z(n1305) );
  XOR U1095 ( .A(n1306), .B(n1307), .Z(n1303) );
  AND U1096 ( .A(n144), .B(n1308), .Z(n1307) );
  XOR U1097 ( .A(n1309), .B(n1310), .Z(n1301) );
  AND U1098 ( .A(n148), .B(n1308), .Z(n1310) );
  XNOR U1099 ( .A(n1309), .B(n1306), .Z(n1308) );
  XOR U1100 ( .A(n1311), .B(n1312), .Z(n1306) );
  AND U1101 ( .A(n151), .B(n1313), .Z(n1312) );
  XOR U1102 ( .A(p_input[263]), .B(n1311), .Z(n1313) );
  XOR U1103 ( .A(n1314), .B(n1315), .Z(n1311) );
  AND U1104 ( .A(n155), .B(n1316), .Z(n1315) );
  XOR U1105 ( .A(n1317), .B(n1318), .Z(n1309) );
  AND U1106 ( .A(n159), .B(n1316), .Z(n1318) );
  XNOR U1107 ( .A(n1317), .B(n1314), .Z(n1316) );
  XOR U1108 ( .A(n1319), .B(n1320), .Z(n1314) );
  AND U1109 ( .A(n162), .B(n1321), .Z(n1320) );
  XOR U1110 ( .A(p_input[295]), .B(n1319), .Z(n1321) );
  XOR U1111 ( .A(n1322), .B(n1323), .Z(n1319) );
  AND U1112 ( .A(n166), .B(n1324), .Z(n1323) );
  XOR U1113 ( .A(n1325), .B(n1326), .Z(n1317) );
  AND U1114 ( .A(n170), .B(n1324), .Z(n1326) );
  XNOR U1115 ( .A(n1325), .B(n1322), .Z(n1324) );
  XOR U1116 ( .A(n1327), .B(n1328), .Z(n1322) );
  AND U1117 ( .A(n173), .B(n1329), .Z(n1328) );
  XOR U1118 ( .A(p_input[327]), .B(n1327), .Z(n1329) );
  XOR U1119 ( .A(n1330), .B(n1331), .Z(n1327) );
  AND U1120 ( .A(n177), .B(n1332), .Z(n1331) );
  XOR U1121 ( .A(n1333), .B(n1334), .Z(n1325) );
  AND U1122 ( .A(n181), .B(n1332), .Z(n1334) );
  XNOR U1123 ( .A(n1333), .B(n1330), .Z(n1332) );
  XOR U1124 ( .A(n1335), .B(n1336), .Z(n1330) );
  AND U1125 ( .A(n184), .B(n1337), .Z(n1336) );
  XOR U1126 ( .A(p_input[359]), .B(n1335), .Z(n1337) );
  XOR U1127 ( .A(n1338), .B(n1339), .Z(n1335) );
  AND U1128 ( .A(n188), .B(n1340), .Z(n1339) );
  XOR U1129 ( .A(n1341), .B(n1342), .Z(n1333) );
  AND U1130 ( .A(n192), .B(n1340), .Z(n1342) );
  XNOR U1131 ( .A(n1341), .B(n1338), .Z(n1340) );
  XOR U1132 ( .A(n1343), .B(n1344), .Z(n1338) );
  AND U1133 ( .A(n195), .B(n1345), .Z(n1344) );
  XOR U1134 ( .A(p_input[391]), .B(n1343), .Z(n1345) );
  XOR U1135 ( .A(n1346), .B(n1347), .Z(n1343) );
  AND U1136 ( .A(n199), .B(n1348), .Z(n1347) );
  XOR U1137 ( .A(n1349), .B(n1350), .Z(n1341) );
  AND U1138 ( .A(n203), .B(n1348), .Z(n1350) );
  XNOR U1139 ( .A(n1349), .B(n1346), .Z(n1348) );
  XOR U1140 ( .A(n1351), .B(n1352), .Z(n1346) );
  AND U1141 ( .A(n206), .B(n1353), .Z(n1352) );
  XOR U1142 ( .A(p_input[423]), .B(n1351), .Z(n1353) );
  XOR U1143 ( .A(n1354), .B(n1355), .Z(n1351) );
  AND U1144 ( .A(n210), .B(n1356), .Z(n1355) );
  XOR U1145 ( .A(n1357), .B(n1358), .Z(n1349) );
  AND U1146 ( .A(n214), .B(n1356), .Z(n1358) );
  XNOR U1147 ( .A(n1357), .B(n1354), .Z(n1356) );
  XOR U1148 ( .A(n1359), .B(n1360), .Z(n1354) );
  AND U1149 ( .A(n217), .B(n1361), .Z(n1360) );
  XOR U1150 ( .A(p_input[455]), .B(n1359), .Z(n1361) );
  XOR U1151 ( .A(n1362), .B(n1363), .Z(n1359) );
  AND U1152 ( .A(n221), .B(n1364), .Z(n1363) );
  XOR U1153 ( .A(n1365), .B(n1366), .Z(n1357) );
  AND U1154 ( .A(n225), .B(n1364), .Z(n1366) );
  XNOR U1155 ( .A(n1365), .B(n1362), .Z(n1364) );
  XOR U1156 ( .A(n1367), .B(n1368), .Z(n1362) );
  AND U1157 ( .A(n228), .B(n1369), .Z(n1368) );
  XOR U1158 ( .A(p_input[487]), .B(n1367), .Z(n1369) );
  XOR U1159 ( .A(n1370), .B(n1371), .Z(n1367) );
  AND U1160 ( .A(n232), .B(n1372), .Z(n1371) );
  XOR U1161 ( .A(n1373), .B(n1374), .Z(n1365) );
  AND U1162 ( .A(n236), .B(n1372), .Z(n1374) );
  XNOR U1163 ( .A(n1373), .B(n1370), .Z(n1372) );
  XOR U1164 ( .A(n1375), .B(n1376), .Z(n1370) );
  AND U1165 ( .A(n239), .B(n1377), .Z(n1376) );
  XOR U1166 ( .A(p_input[519]), .B(n1375), .Z(n1377) );
  XOR U1167 ( .A(n1378), .B(n1379), .Z(n1375) );
  AND U1168 ( .A(n243), .B(n1380), .Z(n1379) );
  XOR U1169 ( .A(n1381), .B(n1382), .Z(n1373) );
  AND U1170 ( .A(n247), .B(n1380), .Z(n1382) );
  XNOR U1171 ( .A(n1381), .B(n1378), .Z(n1380) );
  XOR U1172 ( .A(n1383), .B(n1384), .Z(n1378) );
  AND U1173 ( .A(n250), .B(n1385), .Z(n1384) );
  XOR U1174 ( .A(p_input[551]), .B(n1383), .Z(n1385) );
  XOR U1175 ( .A(n1386), .B(n1387), .Z(n1383) );
  AND U1176 ( .A(n254), .B(n1388), .Z(n1387) );
  XOR U1177 ( .A(n1389), .B(n1390), .Z(n1381) );
  AND U1178 ( .A(n258), .B(n1388), .Z(n1390) );
  XNOR U1179 ( .A(n1389), .B(n1386), .Z(n1388) );
  XOR U1180 ( .A(n1391), .B(n1392), .Z(n1386) );
  AND U1181 ( .A(n261), .B(n1393), .Z(n1392) );
  XOR U1182 ( .A(p_input[583]), .B(n1391), .Z(n1393) );
  XOR U1183 ( .A(n1394), .B(n1395), .Z(n1391) );
  AND U1184 ( .A(n265), .B(n1396), .Z(n1395) );
  XOR U1185 ( .A(n1397), .B(n1398), .Z(n1389) );
  AND U1186 ( .A(n269), .B(n1396), .Z(n1398) );
  XNOR U1187 ( .A(n1397), .B(n1394), .Z(n1396) );
  XOR U1188 ( .A(n1399), .B(n1400), .Z(n1394) );
  AND U1189 ( .A(n272), .B(n1401), .Z(n1400) );
  XOR U1190 ( .A(p_input[615]), .B(n1399), .Z(n1401) );
  XOR U1191 ( .A(n1402), .B(n1403), .Z(n1399) );
  AND U1192 ( .A(n276), .B(n1404), .Z(n1403) );
  XOR U1193 ( .A(n1405), .B(n1406), .Z(n1397) );
  AND U1194 ( .A(n280), .B(n1404), .Z(n1406) );
  XNOR U1195 ( .A(n1405), .B(n1402), .Z(n1404) );
  XOR U1196 ( .A(n1407), .B(n1408), .Z(n1402) );
  AND U1197 ( .A(n283), .B(n1409), .Z(n1408) );
  XOR U1198 ( .A(p_input[647]), .B(n1407), .Z(n1409) );
  XOR U1199 ( .A(n1410), .B(n1411), .Z(n1407) );
  AND U1200 ( .A(n287), .B(n1412), .Z(n1411) );
  XOR U1201 ( .A(n1413), .B(n1414), .Z(n1405) );
  AND U1202 ( .A(n291), .B(n1412), .Z(n1414) );
  XNOR U1203 ( .A(n1413), .B(n1410), .Z(n1412) );
  XOR U1204 ( .A(n1415), .B(n1416), .Z(n1410) );
  AND U1205 ( .A(n294), .B(n1417), .Z(n1416) );
  XOR U1206 ( .A(p_input[679]), .B(n1415), .Z(n1417) );
  XOR U1207 ( .A(n1418), .B(n1419), .Z(n1415) );
  AND U1208 ( .A(n298), .B(n1420), .Z(n1419) );
  XOR U1209 ( .A(n1421), .B(n1422), .Z(n1413) );
  AND U1210 ( .A(n302), .B(n1420), .Z(n1422) );
  XNOR U1211 ( .A(n1421), .B(n1418), .Z(n1420) );
  XOR U1212 ( .A(n1423), .B(n1424), .Z(n1418) );
  AND U1213 ( .A(n305), .B(n1425), .Z(n1424) );
  XOR U1214 ( .A(p_input[711]), .B(n1423), .Z(n1425) );
  XOR U1215 ( .A(n1426), .B(n1427), .Z(n1423) );
  AND U1216 ( .A(n309), .B(n1428), .Z(n1427) );
  XOR U1217 ( .A(n1429), .B(n1430), .Z(n1421) );
  AND U1218 ( .A(n313), .B(n1428), .Z(n1430) );
  XNOR U1219 ( .A(n1429), .B(n1426), .Z(n1428) );
  XOR U1220 ( .A(n1431), .B(n1432), .Z(n1426) );
  AND U1221 ( .A(n316), .B(n1433), .Z(n1432) );
  XOR U1222 ( .A(p_input[743]), .B(n1431), .Z(n1433) );
  XOR U1223 ( .A(n1434), .B(n1435), .Z(n1431) );
  AND U1224 ( .A(n320), .B(n1436), .Z(n1435) );
  XOR U1225 ( .A(n1437), .B(n1438), .Z(n1429) );
  AND U1226 ( .A(n324), .B(n1436), .Z(n1438) );
  XNOR U1227 ( .A(n1437), .B(n1434), .Z(n1436) );
  XOR U1228 ( .A(n1439), .B(n1440), .Z(n1434) );
  AND U1229 ( .A(n327), .B(n1441), .Z(n1440) );
  XOR U1230 ( .A(p_input[775]), .B(n1439), .Z(n1441) );
  XOR U1231 ( .A(n1442), .B(n1443), .Z(n1439) );
  AND U1232 ( .A(n331), .B(n1444), .Z(n1443) );
  XOR U1233 ( .A(n1445), .B(n1446), .Z(n1437) );
  AND U1234 ( .A(n335), .B(n1444), .Z(n1446) );
  XNOR U1235 ( .A(n1445), .B(n1442), .Z(n1444) );
  XOR U1236 ( .A(n1447), .B(n1448), .Z(n1442) );
  AND U1237 ( .A(n338), .B(n1449), .Z(n1448) );
  XOR U1238 ( .A(p_input[807]), .B(n1447), .Z(n1449) );
  XOR U1239 ( .A(n1450), .B(n1451), .Z(n1447) );
  AND U1240 ( .A(n342), .B(n1452), .Z(n1451) );
  XOR U1241 ( .A(n1453), .B(n1454), .Z(n1445) );
  AND U1242 ( .A(n346), .B(n1452), .Z(n1454) );
  XNOR U1243 ( .A(n1453), .B(n1450), .Z(n1452) );
  XOR U1244 ( .A(n1455), .B(n1456), .Z(n1450) );
  AND U1245 ( .A(n349), .B(n1457), .Z(n1456) );
  XOR U1246 ( .A(p_input[839]), .B(n1455), .Z(n1457) );
  XOR U1247 ( .A(n1458), .B(n1459), .Z(n1455) );
  AND U1248 ( .A(n353), .B(n1460), .Z(n1459) );
  XOR U1249 ( .A(n1461), .B(n1462), .Z(n1453) );
  AND U1250 ( .A(n357), .B(n1460), .Z(n1462) );
  XNOR U1251 ( .A(n1461), .B(n1458), .Z(n1460) );
  XOR U1252 ( .A(n1463), .B(n1464), .Z(n1458) );
  AND U1253 ( .A(n360), .B(n1465), .Z(n1464) );
  XOR U1254 ( .A(p_input[871]), .B(n1463), .Z(n1465) );
  XOR U1255 ( .A(n1466), .B(n1467), .Z(n1463) );
  AND U1256 ( .A(n364), .B(n1468), .Z(n1467) );
  XOR U1257 ( .A(n1469), .B(n1470), .Z(n1461) );
  AND U1258 ( .A(n368), .B(n1468), .Z(n1470) );
  XNOR U1259 ( .A(n1469), .B(n1466), .Z(n1468) );
  XOR U1260 ( .A(n1471), .B(n1472), .Z(n1466) );
  AND U1261 ( .A(n371), .B(n1473), .Z(n1472) );
  XOR U1262 ( .A(p_input[903]), .B(n1471), .Z(n1473) );
  XOR U1263 ( .A(n1474), .B(n1475), .Z(n1471) );
  AND U1264 ( .A(n375), .B(n1476), .Z(n1475) );
  XOR U1265 ( .A(n1477), .B(n1478), .Z(n1469) );
  AND U1266 ( .A(n379), .B(n1476), .Z(n1478) );
  XNOR U1267 ( .A(n1477), .B(n1474), .Z(n1476) );
  XOR U1268 ( .A(n1479), .B(n1480), .Z(n1474) );
  AND U1269 ( .A(n382), .B(n1481), .Z(n1480) );
  XOR U1270 ( .A(p_input[935]), .B(n1479), .Z(n1481) );
  XOR U1271 ( .A(n1482), .B(n1483), .Z(n1479) );
  AND U1272 ( .A(n386), .B(n1484), .Z(n1483) );
  XOR U1273 ( .A(n1485), .B(n1486), .Z(n1477) );
  AND U1274 ( .A(n390), .B(n1484), .Z(n1486) );
  XNOR U1275 ( .A(n1485), .B(n1482), .Z(n1484) );
  XOR U1276 ( .A(n1487), .B(n1488), .Z(n1482) );
  AND U1277 ( .A(n393), .B(n1489), .Z(n1488) );
  XOR U1278 ( .A(p_input[967]), .B(n1487), .Z(n1489) );
  XOR U1279 ( .A(n1490), .B(n1491), .Z(n1487) );
  AND U1280 ( .A(n397), .B(n1492), .Z(n1491) );
  XOR U1281 ( .A(n1493), .B(n1494), .Z(n1485) );
  AND U1282 ( .A(n401), .B(n1492), .Z(n1494) );
  XNOR U1283 ( .A(n1493), .B(n1490), .Z(n1492) );
  XOR U1284 ( .A(n1495), .B(n1496), .Z(n1490) );
  AND U1285 ( .A(n404), .B(n1497), .Z(n1496) );
  XOR U1286 ( .A(p_input[999]), .B(n1495), .Z(n1497) );
  XOR U1287 ( .A(n1498), .B(n1499), .Z(n1495) );
  AND U1288 ( .A(n408), .B(n1500), .Z(n1499) );
  XOR U1289 ( .A(n1501), .B(n1502), .Z(n1493) );
  AND U1290 ( .A(n412), .B(n1500), .Z(n1502) );
  XNOR U1291 ( .A(n1501), .B(n1498), .Z(n1500) );
  XOR U1292 ( .A(n1503), .B(n1504), .Z(n1498) );
  AND U1293 ( .A(n415), .B(n1505), .Z(n1504) );
  XOR U1294 ( .A(p_input[1031]), .B(n1503), .Z(n1505) );
  XOR U1295 ( .A(n1506), .B(n1507), .Z(n1503) );
  AND U1296 ( .A(n419), .B(n1508), .Z(n1507) );
  XOR U1297 ( .A(n1509), .B(n1510), .Z(n1501) );
  AND U1298 ( .A(n423), .B(n1508), .Z(n1510) );
  XNOR U1299 ( .A(n1509), .B(n1506), .Z(n1508) );
  XOR U1300 ( .A(n1511), .B(n1512), .Z(n1506) );
  AND U1301 ( .A(n426), .B(n1513), .Z(n1512) );
  XOR U1302 ( .A(p_input[1063]), .B(n1511), .Z(n1513) );
  XOR U1303 ( .A(n1514), .B(n1515), .Z(n1511) );
  AND U1304 ( .A(n430), .B(n1516), .Z(n1515) );
  XOR U1305 ( .A(n1517), .B(n1518), .Z(n1509) );
  AND U1306 ( .A(n434), .B(n1516), .Z(n1518) );
  XNOR U1307 ( .A(n1517), .B(n1514), .Z(n1516) );
  XOR U1308 ( .A(n1519), .B(n1520), .Z(n1514) );
  AND U1309 ( .A(n437), .B(n1521), .Z(n1520) );
  XOR U1310 ( .A(p_input[1095]), .B(n1519), .Z(n1521) );
  XOR U1311 ( .A(n1522), .B(n1523), .Z(n1519) );
  AND U1312 ( .A(n441), .B(n1524), .Z(n1523) );
  XOR U1313 ( .A(n1525), .B(n1526), .Z(n1517) );
  AND U1314 ( .A(n445), .B(n1524), .Z(n1526) );
  XNOR U1315 ( .A(n1525), .B(n1522), .Z(n1524) );
  XOR U1316 ( .A(n1527), .B(n1528), .Z(n1522) );
  AND U1317 ( .A(n448), .B(n1529), .Z(n1528) );
  XOR U1318 ( .A(p_input[1127]), .B(n1527), .Z(n1529) );
  XOR U1319 ( .A(n1530), .B(n1531), .Z(n1527) );
  AND U1320 ( .A(n452), .B(n1532), .Z(n1531) );
  XOR U1321 ( .A(n1533), .B(n1534), .Z(n1525) );
  AND U1322 ( .A(n456), .B(n1532), .Z(n1534) );
  XNOR U1323 ( .A(n1533), .B(n1530), .Z(n1532) );
  XOR U1324 ( .A(n1535), .B(n1536), .Z(n1530) );
  AND U1325 ( .A(n459), .B(n1537), .Z(n1536) );
  XOR U1326 ( .A(p_input[1159]), .B(n1535), .Z(n1537) );
  XOR U1327 ( .A(n1538), .B(n1539), .Z(n1535) );
  AND U1328 ( .A(n463), .B(n1540), .Z(n1539) );
  XOR U1329 ( .A(n1541), .B(n1542), .Z(n1533) );
  AND U1330 ( .A(n467), .B(n1540), .Z(n1542) );
  XNOR U1331 ( .A(n1541), .B(n1538), .Z(n1540) );
  XOR U1332 ( .A(n1543), .B(n1544), .Z(n1538) );
  AND U1333 ( .A(n470), .B(n1545), .Z(n1544) );
  XOR U1334 ( .A(p_input[1191]), .B(n1543), .Z(n1545) );
  XOR U1335 ( .A(n1546), .B(n1547), .Z(n1543) );
  AND U1336 ( .A(n474), .B(n1548), .Z(n1547) );
  XOR U1337 ( .A(n1549), .B(n1550), .Z(n1541) );
  AND U1338 ( .A(n478), .B(n1548), .Z(n1550) );
  XNOR U1339 ( .A(n1549), .B(n1546), .Z(n1548) );
  XOR U1340 ( .A(n1551), .B(n1552), .Z(n1546) );
  AND U1341 ( .A(n481), .B(n1553), .Z(n1552) );
  XOR U1342 ( .A(p_input[1223]), .B(n1551), .Z(n1553) );
  XOR U1343 ( .A(n1554), .B(n1555), .Z(n1551) );
  AND U1344 ( .A(n485), .B(n1556), .Z(n1555) );
  XOR U1345 ( .A(n1557), .B(n1558), .Z(n1549) );
  AND U1346 ( .A(n489), .B(n1556), .Z(n1558) );
  XNOR U1347 ( .A(n1557), .B(n1554), .Z(n1556) );
  XOR U1348 ( .A(n1559), .B(n1560), .Z(n1554) );
  AND U1349 ( .A(n492), .B(n1561), .Z(n1560) );
  XOR U1350 ( .A(p_input[1255]), .B(n1559), .Z(n1561) );
  XOR U1351 ( .A(n1562), .B(n1563), .Z(n1559) );
  AND U1352 ( .A(n496), .B(n1564), .Z(n1563) );
  XOR U1353 ( .A(n1565), .B(n1566), .Z(n1557) );
  AND U1354 ( .A(n500), .B(n1564), .Z(n1566) );
  XNOR U1355 ( .A(n1565), .B(n1562), .Z(n1564) );
  XOR U1356 ( .A(n1567), .B(n1568), .Z(n1562) );
  AND U1357 ( .A(n503), .B(n1569), .Z(n1568) );
  XOR U1358 ( .A(p_input[1287]), .B(n1567), .Z(n1569) );
  XOR U1359 ( .A(n1570), .B(n1571), .Z(n1567) );
  AND U1360 ( .A(n507), .B(n1572), .Z(n1571) );
  XOR U1361 ( .A(n1573), .B(n1574), .Z(n1565) );
  AND U1362 ( .A(n511), .B(n1572), .Z(n1574) );
  XNOR U1363 ( .A(n1573), .B(n1570), .Z(n1572) );
  XOR U1364 ( .A(n1575), .B(n1576), .Z(n1570) );
  AND U1365 ( .A(n514), .B(n1577), .Z(n1576) );
  XOR U1366 ( .A(p_input[1319]), .B(n1575), .Z(n1577) );
  XOR U1367 ( .A(n1578), .B(n1579), .Z(n1575) );
  AND U1368 ( .A(n518), .B(n1580), .Z(n1579) );
  XOR U1369 ( .A(n1581), .B(n1582), .Z(n1573) );
  AND U1370 ( .A(n522), .B(n1580), .Z(n1582) );
  XNOR U1371 ( .A(n1581), .B(n1578), .Z(n1580) );
  XOR U1372 ( .A(n1583), .B(n1584), .Z(n1578) );
  AND U1373 ( .A(n525), .B(n1585), .Z(n1584) );
  XOR U1374 ( .A(p_input[1351]), .B(n1583), .Z(n1585) );
  XOR U1375 ( .A(n1586), .B(n1587), .Z(n1583) );
  AND U1376 ( .A(n529), .B(n1588), .Z(n1587) );
  XOR U1377 ( .A(n1589), .B(n1590), .Z(n1581) );
  AND U1378 ( .A(n533), .B(n1588), .Z(n1590) );
  XNOR U1379 ( .A(n1589), .B(n1586), .Z(n1588) );
  XOR U1380 ( .A(n1591), .B(n1592), .Z(n1586) );
  AND U1381 ( .A(n536), .B(n1593), .Z(n1592) );
  XOR U1382 ( .A(p_input[1383]), .B(n1591), .Z(n1593) );
  XOR U1383 ( .A(n1594), .B(n1595), .Z(n1591) );
  AND U1384 ( .A(n540), .B(n1596), .Z(n1595) );
  XOR U1385 ( .A(n1597), .B(n1598), .Z(n1589) );
  AND U1386 ( .A(n544), .B(n1596), .Z(n1598) );
  XNOR U1387 ( .A(n1597), .B(n1594), .Z(n1596) );
  XOR U1388 ( .A(n1599), .B(n1600), .Z(n1594) );
  AND U1389 ( .A(n547), .B(n1601), .Z(n1600) );
  XOR U1390 ( .A(p_input[1415]), .B(n1599), .Z(n1601) );
  XOR U1391 ( .A(n1602), .B(n1603), .Z(n1599) );
  AND U1392 ( .A(n551), .B(n1604), .Z(n1603) );
  XOR U1393 ( .A(n1605), .B(n1606), .Z(n1597) );
  AND U1394 ( .A(n555), .B(n1604), .Z(n1606) );
  XNOR U1395 ( .A(n1605), .B(n1602), .Z(n1604) );
  XOR U1396 ( .A(n1607), .B(n1608), .Z(n1602) );
  AND U1397 ( .A(n558), .B(n1609), .Z(n1608) );
  XOR U1398 ( .A(p_input[1447]), .B(n1607), .Z(n1609) );
  XOR U1399 ( .A(n1610), .B(n1611), .Z(n1607) );
  AND U1400 ( .A(n562), .B(n1612), .Z(n1611) );
  XOR U1401 ( .A(n1613), .B(n1614), .Z(n1605) );
  AND U1402 ( .A(n566), .B(n1612), .Z(n1614) );
  XNOR U1403 ( .A(n1613), .B(n1610), .Z(n1612) );
  XOR U1404 ( .A(n1615), .B(n1616), .Z(n1610) );
  AND U1405 ( .A(n569), .B(n1617), .Z(n1616) );
  XOR U1406 ( .A(p_input[1479]), .B(n1615), .Z(n1617) );
  XOR U1407 ( .A(n1618), .B(n1619), .Z(n1615) );
  AND U1408 ( .A(n573), .B(n1620), .Z(n1619) );
  XOR U1409 ( .A(n1621), .B(n1622), .Z(n1613) );
  AND U1410 ( .A(n577), .B(n1620), .Z(n1622) );
  XNOR U1411 ( .A(n1621), .B(n1618), .Z(n1620) );
  XOR U1412 ( .A(n1623), .B(n1624), .Z(n1618) );
  AND U1413 ( .A(n580), .B(n1625), .Z(n1624) );
  XOR U1414 ( .A(p_input[1511]), .B(n1623), .Z(n1625) );
  XOR U1415 ( .A(n1626), .B(n1627), .Z(n1623) );
  AND U1416 ( .A(n584), .B(n1628), .Z(n1627) );
  XOR U1417 ( .A(n1629), .B(n1630), .Z(n1621) );
  AND U1418 ( .A(n588), .B(n1628), .Z(n1630) );
  XNOR U1419 ( .A(n1629), .B(n1626), .Z(n1628) );
  XOR U1420 ( .A(n1631), .B(n1632), .Z(n1626) );
  AND U1421 ( .A(n591), .B(n1633), .Z(n1632) );
  XOR U1422 ( .A(p_input[1543]), .B(n1631), .Z(n1633) );
  XOR U1423 ( .A(n1634), .B(n1635), .Z(n1631) );
  AND U1424 ( .A(n595), .B(n1636), .Z(n1635) );
  XOR U1425 ( .A(n1637), .B(n1638), .Z(n1629) );
  AND U1426 ( .A(n599), .B(n1636), .Z(n1638) );
  XNOR U1427 ( .A(n1637), .B(n1634), .Z(n1636) );
  XOR U1428 ( .A(n1639), .B(n1640), .Z(n1634) );
  AND U1429 ( .A(n602), .B(n1641), .Z(n1640) );
  XOR U1430 ( .A(p_input[1575]), .B(n1639), .Z(n1641) );
  XOR U1431 ( .A(n1642), .B(n1643), .Z(n1639) );
  AND U1432 ( .A(n606), .B(n1644), .Z(n1643) );
  XOR U1433 ( .A(n1645), .B(n1646), .Z(n1637) );
  AND U1434 ( .A(n610), .B(n1644), .Z(n1646) );
  XNOR U1435 ( .A(n1645), .B(n1642), .Z(n1644) );
  XOR U1436 ( .A(n1647), .B(n1648), .Z(n1642) );
  AND U1437 ( .A(n613), .B(n1649), .Z(n1648) );
  XOR U1438 ( .A(p_input[1607]), .B(n1647), .Z(n1649) );
  XOR U1439 ( .A(n1650), .B(n1651), .Z(n1647) );
  AND U1440 ( .A(n617), .B(n1652), .Z(n1651) );
  XOR U1441 ( .A(n1653), .B(n1654), .Z(n1645) );
  AND U1442 ( .A(n621), .B(n1652), .Z(n1654) );
  XNOR U1443 ( .A(n1653), .B(n1650), .Z(n1652) );
  XOR U1444 ( .A(n1655), .B(n1656), .Z(n1650) );
  AND U1445 ( .A(n624), .B(n1657), .Z(n1656) );
  XOR U1446 ( .A(p_input[1639]), .B(n1655), .Z(n1657) );
  XOR U1447 ( .A(n1658), .B(n1659), .Z(n1655) );
  AND U1448 ( .A(n628), .B(n1660), .Z(n1659) );
  XOR U1449 ( .A(n1661), .B(n1662), .Z(n1653) );
  AND U1450 ( .A(n632), .B(n1660), .Z(n1662) );
  XNOR U1451 ( .A(n1661), .B(n1658), .Z(n1660) );
  XOR U1452 ( .A(n1663), .B(n1664), .Z(n1658) );
  AND U1453 ( .A(n635), .B(n1665), .Z(n1664) );
  XOR U1454 ( .A(p_input[1671]), .B(n1663), .Z(n1665) );
  XOR U1455 ( .A(n1666), .B(n1667), .Z(n1663) );
  AND U1456 ( .A(n639), .B(n1668), .Z(n1667) );
  XOR U1457 ( .A(n1669), .B(n1670), .Z(n1661) );
  AND U1458 ( .A(n643), .B(n1668), .Z(n1670) );
  XNOR U1459 ( .A(n1669), .B(n1666), .Z(n1668) );
  XOR U1460 ( .A(n1671), .B(n1672), .Z(n1666) );
  AND U1461 ( .A(n646), .B(n1673), .Z(n1672) );
  XOR U1462 ( .A(p_input[1703]), .B(n1671), .Z(n1673) );
  XOR U1463 ( .A(n1674), .B(n1675), .Z(n1671) );
  AND U1464 ( .A(n650), .B(n1676), .Z(n1675) );
  XOR U1465 ( .A(n1677), .B(n1678), .Z(n1669) );
  AND U1466 ( .A(n654), .B(n1676), .Z(n1678) );
  XNOR U1467 ( .A(n1677), .B(n1674), .Z(n1676) );
  XOR U1468 ( .A(n1679), .B(n1680), .Z(n1674) );
  AND U1469 ( .A(n657), .B(n1681), .Z(n1680) );
  XOR U1470 ( .A(p_input[1735]), .B(n1679), .Z(n1681) );
  XOR U1471 ( .A(n1682), .B(n1683), .Z(n1679) );
  AND U1472 ( .A(n661), .B(n1684), .Z(n1683) );
  XOR U1473 ( .A(n1685), .B(n1686), .Z(n1677) );
  AND U1474 ( .A(n665), .B(n1684), .Z(n1686) );
  XNOR U1475 ( .A(n1685), .B(n1682), .Z(n1684) );
  XOR U1476 ( .A(n1687), .B(n1688), .Z(n1682) );
  AND U1477 ( .A(n668), .B(n1689), .Z(n1688) );
  XOR U1478 ( .A(p_input[1767]), .B(n1687), .Z(n1689) );
  XOR U1479 ( .A(n1690), .B(n1691), .Z(n1687) );
  AND U1480 ( .A(n672), .B(n1692), .Z(n1691) );
  XOR U1481 ( .A(n1693), .B(n1694), .Z(n1685) );
  AND U1482 ( .A(n676), .B(n1692), .Z(n1694) );
  XNOR U1483 ( .A(n1693), .B(n1690), .Z(n1692) );
  XOR U1484 ( .A(n1695), .B(n1696), .Z(n1690) );
  AND U1485 ( .A(n679), .B(n1697), .Z(n1696) );
  XOR U1486 ( .A(p_input[1799]), .B(n1695), .Z(n1697) );
  XOR U1487 ( .A(n1698), .B(n1699), .Z(n1695) );
  AND U1488 ( .A(n683), .B(n1700), .Z(n1699) );
  XOR U1489 ( .A(n1701), .B(n1702), .Z(n1693) );
  AND U1490 ( .A(n687), .B(n1700), .Z(n1702) );
  XNOR U1491 ( .A(n1701), .B(n1698), .Z(n1700) );
  XOR U1492 ( .A(n1703), .B(n1704), .Z(n1698) );
  AND U1493 ( .A(n690), .B(n1705), .Z(n1704) );
  XOR U1494 ( .A(p_input[1831]), .B(n1703), .Z(n1705) );
  XOR U1495 ( .A(n1706), .B(n1707), .Z(n1703) );
  AND U1496 ( .A(n694), .B(n1708), .Z(n1707) );
  XOR U1497 ( .A(n1709), .B(n1710), .Z(n1701) );
  AND U1498 ( .A(n698), .B(n1708), .Z(n1710) );
  XNOR U1499 ( .A(n1709), .B(n1706), .Z(n1708) );
  XOR U1500 ( .A(n1711), .B(n1712), .Z(n1706) );
  AND U1501 ( .A(n701), .B(n1713), .Z(n1712) );
  XOR U1502 ( .A(p_input[1863]), .B(n1711), .Z(n1713) );
  XOR U1503 ( .A(n1714), .B(n1715), .Z(n1711) );
  AND U1504 ( .A(n705), .B(n1716), .Z(n1715) );
  XOR U1505 ( .A(n1717), .B(n1718), .Z(n1709) );
  AND U1506 ( .A(n709), .B(n1716), .Z(n1718) );
  XNOR U1507 ( .A(n1717), .B(n1714), .Z(n1716) );
  XOR U1508 ( .A(n1719), .B(n1720), .Z(n1714) );
  AND U1509 ( .A(n712), .B(n1721), .Z(n1720) );
  XOR U1510 ( .A(p_input[1895]), .B(n1719), .Z(n1721) );
  XOR U1511 ( .A(n1722), .B(n1723), .Z(n1719) );
  AND U1512 ( .A(n716), .B(n1724), .Z(n1723) );
  XOR U1513 ( .A(n1725), .B(n1726), .Z(n1717) );
  AND U1514 ( .A(n720), .B(n1724), .Z(n1726) );
  XNOR U1515 ( .A(n1725), .B(n1722), .Z(n1724) );
  XOR U1516 ( .A(n1727), .B(n1728), .Z(n1722) );
  AND U1517 ( .A(n723), .B(n1729), .Z(n1728) );
  XOR U1518 ( .A(p_input[1927]), .B(n1727), .Z(n1729) );
  XOR U1519 ( .A(n1730), .B(n1731), .Z(n1727) );
  AND U1520 ( .A(n727), .B(n1732), .Z(n1731) );
  XOR U1521 ( .A(n1733), .B(n1734), .Z(n1725) );
  AND U1522 ( .A(n731), .B(n1732), .Z(n1734) );
  XNOR U1523 ( .A(n1733), .B(n1730), .Z(n1732) );
  XOR U1524 ( .A(n1735), .B(n1736), .Z(n1730) );
  AND U1525 ( .A(n734), .B(n1737), .Z(n1736) );
  XOR U1526 ( .A(p_input[1959]), .B(n1735), .Z(n1737) );
  XNOR U1527 ( .A(n1738), .B(n1739), .Z(n1735) );
  AND U1528 ( .A(n738), .B(n1740), .Z(n1739) );
  XNOR U1529 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n1741), .Z(n1733) );
  AND U1530 ( .A(n741), .B(n1740), .Z(n1741) );
  XOR U1531 ( .A(n1742), .B(n1738), .Z(n1740) );
  XOR U1532 ( .A(n7), .B(n1743), .Z(o[38]) );
  AND U1533 ( .A(n58), .B(n1744), .Z(n7) );
  XOR U1534 ( .A(n8), .B(n1743), .Z(n1744) );
  XOR U1535 ( .A(n1745), .B(n1746), .Z(n1743) );
  AND U1536 ( .A(n62), .B(n1747), .Z(n1746) );
  XOR U1537 ( .A(p_input[6]), .B(n1745), .Z(n1747) );
  XOR U1538 ( .A(n1748), .B(n1749), .Z(n1745) );
  AND U1539 ( .A(n66), .B(n1750), .Z(n1749) );
  XOR U1540 ( .A(n1751), .B(n1752), .Z(n8) );
  AND U1541 ( .A(n70), .B(n1750), .Z(n1752) );
  XNOR U1542 ( .A(n1753), .B(n1748), .Z(n1750) );
  XOR U1543 ( .A(n1754), .B(n1755), .Z(n1748) );
  AND U1544 ( .A(n74), .B(n1756), .Z(n1755) );
  XOR U1545 ( .A(p_input[38]), .B(n1754), .Z(n1756) );
  XOR U1546 ( .A(n1757), .B(n1758), .Z(n1754) );
  AND U1547 ( .A(n78), .B(n1759), .Z(n1758) );
  IV U1548 ( .A(n1751), .Z(n1753) );
  XNOR U1549 ( .A(n1760), .B(n1761), .Z(n1751) );
  AND U1550 ( .A(n82), .B(n1759), .Z(n1761) );
  XNOR U1551 ( .A(n1760), .B(n1757), .Z(n1759) );
  XOR U1552 ( .A(n1762), .B(n1763), .Z(n1757) );
  AND U1553 ( .A(n85), .B(n1764), .Z(n1763) );
  XOR U1554 ( .A(p_input[70]), .B(n1762), .Z(n1764) );
  XOR U1555 ( .A(n1765), .B(n1766), .Z(n1762) );
  AND U1556 ( .A(n89), .B(n1767), .Z(n1766) );
  XOR U1557 ( .A(n1768), .B(n1769), .Z(n1760) );
  AND U1558 ( .A(n93), .B(n1767), .Z(n1769) );
  XNOR U1559 ( .A(n1768), .B(n1765), .Z(n1767) );
  XOR U1560 ( .A(n1770), .B(n1771), .Z(n1765) );
  AND U1561 ( .A(n96), .B(n1772), .Z(n1771) );
  XOR U1562 ( .A(p_input[102]), .B(n1770), .Z(n1772) );
  XOR U1563 ( .A(n1773), .B(n1774), .Z(n1770) );
  AND U1564 ( .A(n100), .B(n1775), .Z(n1774) );
  XOR U1565 ( .A(n1776), .B(n1777), .Z(n1768) );
  AND U1566 ( .A(n104), .B(n1775), .Z(n1777) );
  XNOR U1567 ( .A(n1776), .B(n1773), .Z(n1775) );
  XOR U1568 ( .A(n1778), .B(n1779), .Z(n1773) );
  AND U1569 ( .A(n107), .B(n1780), .Z(n1779) );
  XOR U1570 ( .A(p_input[134]), .B(n1778), .Z(n1780) );
  XOR U1571 ( .A(n1781), .B(n1782), .Z(n1778) );
  AND U1572 ( .A(n111), .B(n1783), .Z(n1782) );
  XOR U1573 ( .A(n1784), .B(n1785), .Z(n1776) );
  AND U1574 ( .A(n115), .B(n1783), .Z(n1785) );
  XNOR U1575 ( .A(n1784), .B(n1781), .Z(n1783) );
  XOR U1576 ( .A(n1786), .B(n1787), .Z(n1781) );
  AND U1577 ( .A(n118), .B(n1788), .Z(n1787) );
  XOR U1578 ( .A(p_input[166]), .B(n1786), .Z(n1788) );
  XOR U1579 ( .A(n1789), .B(n1790), .Z(n1786) );
  AND U1580 ( .A(n122), .B(n1791), .Z(n1790) );
  XOR U1581 ( .A(n1792), .B(n1793), .Z(n1784) );
  AND U1582 ( .A(n126), .B(n1791), .Z(n1793) );
  XNOR U1583 ( .A(n1792), .B(n1789), .Z(n1791) );
  XOR U1584 ( .A(n1794), .B(n1795), .Z(n1789) );
  AND U1585 ( .A(n129), .B(n1796), .Z(n1795) );
  XOR U1586 ( .A(p_input[198]), .B(n1794), .Z(n1796) );
  XOR U1587 ( .A(n1797), .B(n1798), .Z(n1794) );
  AND U1588 ( .A(n133), .B(n1799), .Z(n1798) );
  XOR U1589 ( .A(n1800), .B(n1801), .Z(n1792) );
  AND U1590 ( .A(n137), .B(n1799), .Z(n1801) );
  XNOR U1591 ( .A(n1800), .B(n1797), .Z(n1799) );
  XOR U1592 ( .A(n1802), .B(n1803), .Z(n1797) );
  AND U1593 ( .A(n140), .B(n1804), .Z(n1803) );
  XOR U1594 ( .A(p_input[230]), .B(n1802), .Z(n1804) );
  XOR U1595 ( .A(n1805), .B(n1806), .Z(n1802) );
  AND U1596 ( .A(n144), .B(n1807), .Z(n1806) );
  XOR U1597 ( .A(n1808), .B(n1809), .Z(n1800) );
  AND U1598 ( .A(n148), .B(n1807), .Z(n1809) );
  XNOR U1599 ( .A(n1808), .B(n1805), .Z(n1807) );
  XOR U1600 ( .A(n1810), .B(n1811), .Z(n1805) );
  AND U1601 ( .A(n151), .B(n1812), .Z(n1811) );
  XOR U1602 ( .A(p_input[262]), .B(n1810), .Z(n1812) );
  XOR U1603 ( .A(n1813), .B(n1814), .Z(n1810) );
  AND U1604 ( .A(n155), .B(n1815), .Z(n1814) );
  XOR U1605 ( .A(n1816), .B(n1817), .Z(n1808) );
  AND U1606 ( .A(n159), .B(n1815), .Z(n1817) );
  XNOR U1607 ( .A(n1816), .B(n1813), .Z(n1815) );
  XOR U1608 ( .A(n1818), .B(n1819), .Z(n1813) );
  AND U1609 ( .A(n162), .B(n1820), .Z(n1819) );
  XOR U1610 ( .A(p_input[294]), .B(n1818), .Z(n1820) );
  XOR U1611 ( .A(n1821), .B(n1822), .Z(n1818) );
  AND U1612 ( .A(n166), .B(n1823), .Z(n1822) );
  XOR U1613 ( .A(n1824), .B(n1825), .Z(n1816) );
  AND U1614 ( .A(n170), .B(n1823), .Z(n1825) );
  XNOR U1615 ( .A(n1824), .B(n1821), .Z(n1823) );
  XOR U1616 ( .A(n1826), .B(n1827), .Z(n1821) );
  AND U1617 ( .A(n173), .B(n1828), .Z(n1827) );
  XOR U1618 ( .A(p_input[326]), .B(n1826), .Z(n1828) );
  XOR U1619 ( .A(n1829), .B(n1830), .Z(n1826) );
  AND U1620 ( .A(n177), .B(n1831), .Z(n1830) );
  XOR U1621 ( .A(n1832), .B(n1833), .Z(n1824) );
  AND U1622 ( .A(n181), .B(n1831), .Z(n1833) );
  XNOR U1623 ( .A(n1832), .B(n1829), .Z(n1831) );
  XOR U1624 ( .A(n1834), .B(n1835), .Z(n1829) );
  AND U1625 ( .A(n184), .B(n1836), .Z(n1835) );
  XOR U1626 ( .A(p_input[358]), .B(n1834), .Z(n1836) );
  XOR U1627 ( .A(n1837), .B(n1838), .Z(n1834) );
  AND U1628 ( .A(n188), .B(n1839), .Z(n1838) );
  XOR U1629 ( .A(n1840), .B(n1841), .Z(n1832) );
  AND U1630 ( .A(n192), .B(n1839), .Z(n1841) );
  XNOR U1631 ( .A(n1840), .B(n1837), .Z(n1839) );
  XOR U1632 ( .A(n1842), .B(n1843), .Z(n1837) );
  AND U1633 ( .A(n195), .B(n1844), .Z(n1843) );
  XOR U1634 ( .A(p_input[390]), .B(n1842), .Z(n1844) );
  XOR U1635 ( .A(n1845), .B(n1846), .Z(n1842) );
  AND U1636 ( .A(n199), .B(n1847), .Z(n1846) );
  XOR U1637 ( .A(n1848), .B(n1849), .Z(n1840) );
  AND U1638 ( .A(n203), .B(n1847), .Z(n1849) );
  XNOR U1639 ( .A(n1848), .B(n1845), .Z(n1847) );
  XOR U1640 ( .A(n1850), .B(n1851), .Z(n1845) );
  AND U1641 ( .A(n206), .B(n1852), .Z(n1851) );
  XOR U1642 ( .A(p_input[422]), .B(n1850), .Z(n1852) );
  XOR U1643 ( .A(n1853), .B(n1854), .Z(n1850) );
  AND U1644 ( .A(n210), .B(n1855), .Z(n1854) );
  XOR U1645 ( .A(n1856), .B(n1857), .Z(n1848) );
  AND U1646 ( .A(n214), .B(n1855), .Z(n1857) );
  XNOR U1647 ( .A(n1856), .B(n1853), .Z(n1855) );
  XOR U1648 ( .A(n1858), .B(n1859), .Z(n1853) );
  AND U1649 ( .A(n217), .B(n1860), .Z(n1859) );
  XOR U1650 ( .A(p_input[454]), .B(n1858), .Z(n1860) );
  XOR U1651 ( .A(n1861), .B(n1862), .Z(n1858) );
  AND U1652 ( .A(n221), .B(n1863), .Z(n1862) );
  XOR U1653 ( .A(n1864), .B(n1865), .Z(n1856) );
  AND U1654 ( .A(n225), .B(n1863), .Z(n1865) );
  XNOR U1655 ( .A(n1864), .B(n1861), .Z(n1863) );
  XOR U1656 ( .A(n1866), .B(n1867), .Z(n1861) );
  AND U1657 ( .A(n228), .B(n1868), .Z(n1867) );
  XOR U1658 ( .A(p_input[486]), .B(n1866), .Z(n1868) );
  XOR U1659 ( .A(n1869), .B(n1870), .Z(n1866) );
  AND U1660 ( .A(n232), .B(n1871), .Z(n1870) );
  XOR U1661 ( .A(n1872), .B(n1873), .Z(n1864) );
  AND U1662 ( .A(n236), .B(n1871), .Z(n1873) );
  XNOR U1663 ( .A(n1872), .B(n1869), .Z(n1871) );
  XOR U1664 ( .A(n1874), .B(n1875), .Z(n1869) );
  AND U1665 ( .A(n239), .B(n1876), .Z(n1875) );
  XOR U1666 ( .A(p_input[518]), .B(n1874), .Z(n1876) );
  XOR U1667 ( .A(n1877), .B(n1878), .Z(n1874) );
  AND U1668 ( .A(n243), .B(n1879), .Z(n1878) );
  XOR U1669 ( .A(n1880), .B(n1881), .Z(n1872) );
  AND U1670 ( .A(n247), .B(n1879), .Z(n1881) );
  XNOR U1671 ( .A(n1880), .B(n1877), .Z(n1879) );
  XOR U1672 ( .A(n1882), .B(n1883), .Z(n1877) );
  AND U1673 ( .A(n250), .B(n1884), .Z(n1883) );
  XOR U1674 ( .A(p_input[550]), .B(n1882), .Z(n1884) );
  XOR U1675 ( .A(n1885), .B(n1886), .Z(n1882) );
  AND U1676 ( .A(n254), .B(n1887), .Z(n1886) );
  XOR U1677 ( .A(n1888), .B(n1889), .Z(n1880) );
  AND U1678 ( .A(n258), .B(n1887), .Z(n1889) );
  XNOR U1679 ( .A(n1888), .B(n1885), .Z(n1887) );
  XOR U1680 ( .A(n1890), .B(n1891), .Z(n1885) );
  AND U1681 ( .A(n261), .B(n1892), .Z(n1891) );
  XOR U1682 ( .A(p_input[582]), .B(n1890), .Z(n1892) );
  XOR U1683 ( .A(n1893), .B(n1894), .Z(n1890) );
  AND U1684 ( .A(n265), .B(n1895), .Z(n1894) );
  XOR U1685 ( .A(n1896), .B(n1897), .Z(n1888) );
  AND U1686 ( .A(n269), .B(n1895), .Z(n1897) );
  XNOR U1687 ( .A(n1896), .B(n1893), .Z(n1895) );
  XOR U1688 ( .A(n1898), .B(n1899), .Z(n1893) );
  AND U1689 ( .A(n272), .B(n1900), .Z(n1899) );
  XOR U1690 ( .A(p_input[614]), .B(n1898), .Z(n1900) );
  XOR U1691 ( .A(n1901), .B(n1902), .Z(n1898) );
  AND U1692 ( .A(n276), .B(n1903), .Z(n1902) );
  XOR U1693 ( .A(n1904), .B(n1905), .Z(n1896) );
  AND U1694 ( .A(n280), .B(n1903), .Z(n1905) );
  XNOR U1695 ( .A(n1904), .B(n1901), .Z(n1903) );
  XOR U1696 ( .A(n1906), .B(n1907), .Z(n1901) );
  AND U1697 ( .A(n283), .B(n1908), .Z(n1907) );
  XOR U1698 ( .A(p_input[646]), .B(n1906), .Z(n1908) );
  XOR U1699 ( .A(n1909), .B(n1910), .Z(n1906) );
  AND U1700 ( .A(n287), .B(n1911), .Z(n1910) );
  XOR U1701 ( .A(n1912), .B(n1913), .Z(n1904) );
  AND U1702 ( .A(n291), .B(n1911), .Z(n1913) );
  XNOR U1703 ( .A(n1912), .B(n1909), .Z(n1911) );
  XOR U1704 ( .A(n1914), .B(n1915), .Z(n1909) );
  AND U1705 ( .A(n294), .B(n1916), .Z(n1915) );
  XOR U1706 ( .A(p_input[678]), .B(n1914), .Z(n1916) );
  XOR U1707 ( .A(n1917), .B(n1918), .Z(n1914) );
  AND U1708 ( .A(n298), .B(n1919), .Z(n1918) );
  XOR U1709 ( .A(n1920), .B(n1921), .Z(n1912) );
  AND U1710 ( .A(n302), .B(n1919), .Z(n1921) );
  XNOR U1711 ( .A(n1920), .B(n1917), .Z(n1919) );
  XOR U1712 ( .A(n1922), .B(n1923), .Z(n1917) );
  AND U1713 ( .A(n305), .B(n1924), .Z(n1923) );
  XOR U1714 ( .A(p_input[710]), .B(n1922), .Z(n1924) );
  XOR U1715 ( .A(n1925), .B(n1926), .Z(n1922) );
  AND U1716 ( .A(n309), .B(n1927), .Z(n1926) );
  XOR U1717 ( .A(n1928), .B(n1929), .Z(n1920) );
  AND U1718 ( .A(n313), .B(n1927), .Z(n1929) );
  XNOR U1719 ( .A(n1928), .B(n1925), .Z(n1927) );
  XOR U1720 ( .A(n1930), .B(n1931), .Z(n1925) );
  AND U1721 ( .A(n316), .B(n1932), .Z(n1931) );
  XOR U1722 ( .A(p_input[742]), .B(n1930), .Z(n1932) );
  XOR U1723 ( .A(n1933), .B(n1934), .Z(n1930) );
  AND U1724 ( .A(n320), .B(n1935), .Z(n1934) );
  XOR U1725 ( .A(n1936), .B(n1937), .Z(n1928) );
  AND U1726 ( .A(n324), .B(n1935), .Z(n1937) );
  XNOR U1727 ( .A(n1936), .B(n1933), .Z(n1935) );
  XOR U1728 ( .A(n1938), .B(n1939), .Z(n1933) );
  AND U1729 ( .A(n327), .B(n1940), .Z(n1939) );
  XOR U1730 ( .A(p_input[774]), .B(n1938), .Z(n1940) );
  XOR U1731 ( .A(n1941), .B(n1942), .Z(n1938) );
  AND U1732 ( .A(n331), .B(n1943), .Z(n1942) );
  XOR U1733 ( .A(n1944), .B(n1945), .Z(n1936) );
  AND U1734 ( .A(n335), .B(n1943), .Z(n1945) );
  XNOR U1735 ( .A(n1944), .B(n1941), .Z(n1943) );
  XOR U1736 ( .A(n1946), .B(n1947), .Z(n1941) );
  AND U1737 ( .A(n338), .B(n1948), .Z(n1947) );
  XOR U1738 ( .A(p_input[806]), .B(n1946), .Z(n1948) );
  XOR U1739 ( .A(n1949), .B(n1950), .Z(n1946) );
  AND U1740 ( .A(n342), .B(n1951), .Z(n1950) );
  XOR U1741 ( .A(n1952), .B(n1953), .Z(n1944) );
  AND U1742 ( .A(n346), .B(n1951), .Z(n1953) );
  XNOR U1743 ( .A(n1952), .B(n1949), .Z(n1951) );
  XOR U1744 ( .A(n1954), .B(n1955), .Z(n1949) );
  AND U1745 ( .A(n349), .B(n1956), .Z(n1955) );
  XOR U1746 ( .A(p_input[838]), .B(n1954), .Z(n1956) );
  XOR U1747 ( .A(n1957), .B(n1958), .Z(n1954) );
  AND U1748 ( .A(n353), .B(n1959), .Z(n1958) );
  XOR U1749 ( .A(n1960), .B(n1961), .Z(n1952) );
  AND U1750 ( .A(n357), .B(n1959), .Z(n1961) );
  XNOR U1751 ( .A(n1960), .B(n1957), .Z(n1959) );
  XOR U1752 ( .A(n1962), .B(n1963), .Z(n1957) );
  AND U1753 ( .A(n360), .B(n1964), .Z(n1963) );
  XOR U1754 ( .A(p_input[870]), .B(n1962), .Z(n1964) );
  XOR U1755 ( .A(n1965), .B(n1966), .Z(n1962) );
  AND U1756 ( .A(n364), .B(n1967), .Z(n1966) );
  XOR U1757 ( .A(n1968), .B(n1969), .Z(n1960) );
  AND U1758 ( .A(n368), .B(n1967), .Z(n1969) );
  XNOR U1759 ( .A(n1968), .B(n1965), .Z(n1967) );
  XOR U1760 ( .A(n1970), .B(n1971), .Z(n1965) );
  AND U1761 ( .A(n371), .B(n1972), .Z(n1971) );
  XOR U1762 ( .A(p_input[902]), .B(n1970), .Z(n1972) );
  XOR U1763 ( .A(n1973), .B(n1974), .Z(n1970) );
  AND U1764 ( .A(n375), .B(n1975), .Z(n1974) );
  XOR U1765 ( .A(n1976), .B(n1977), .Z(n1968) );
  AND U1766 ( .A(n379), .B(n1975), .Z(n1977) );
  XNOR U1767 ( .A(n1976), .B(n1973), .Z(n1975) );
  XOR U1768 ( .A(n1978), .B(n1979), .Z(n1973) );
  AND U1769 ( .A(n382), .B(n1980), .Z(n1979) );
  XOR U1770 ( .A(p_input[934]), .B(n1978), .Z(n1980) );
  XOR U1771 ( .A(n1981), .B(n1982), .Z(n1978) );
  AND U1772 ( .A(n386), .B(n1983), .Z(n1982) );
  XOR U1773 ( .A(n1984), .B(n1985), .Z(n1976) );
  AND U1774 ( .A(n390), .B(n1983), .Z(n1985) );
  XNOR U1775 ( .A(n1984), .B(n1981), .Z(n1983) );
  XOR U1776 ( .A(n1986), .B(n1987), .Z(n1981) );
  AND U1777 ( .A(n393), .B(n1988), .Z(n1987) );
  XOR U1778 ( .A(p_input[966]), .B(n1986), .Z(n1988) );
  XOR U1779 ( .A(n1989), .B(n1990), .Z(n1986) );
  AND U1780 ( .A(n397), .B(n1991), .Z(n1990) );
  XOR U1781 ( .A(n1992), .B(n1993), .Z(n1984) );
  AND U1782 ( .A(n401), .B(n1991), .Z(n1993) );
  XNOR U1783 ( .A(n1992), .B(n1989), .Z(n1991) );
  XOR U1784 ( .A(n1994), .B(n1995), .Z(n1989) );
  AND U1785 ( .A(n404), .B(n1996), .Z(n1995) );
  XOR U1786 ( .A(p_input[998]), .B(n1994), .Z(n1996) );
  XOR U1787 ( .A(n1997), .B(n1998), .Z(n1994) );
  AND U1788 ( .A(n408), .B(n1999), .Z(n1998) );
  XOR U1789 ( .A(n2000), .B(n2001), .Z(n1992) );
  AND U1790 ( .A(n412), .B(n1999), .Z(n2001) );
  XNOR U1791 ( .A(n2000), .B(n1997), .Z(n1999) );
  XOR U1792 ( .A(n2002), .B(n2003), .Z(n1997) );
  AND U1793 ( .A(n415), .B(n2004), .Z(n2003) );
  XOR U1794 ( .A(p_input[1030]), .B(n2002), .Z(n2004) );
  XOR U1795 ( .A(n2005), .B(n2006), .Z(n2002) );
  AND U1796 ( .A(n419), .B(n2007), .Z(n2006) );
  XOR U1797 ( .A(n2008), .B(n2009), .Z(n2000) );
  AND U1798 ( .A(n423), .B(n2007), .Z(n2009) );
  XNOR U1799 ( .A(n2008), .B(n2005), .Z(n2007) );
  XOR U1800 ( .A(n2010), .B(n2011), .Z(n2005) );
  AND U1801 ( .A(n426), .B(n2012), .Z(n2011) );
  XOR U1802 ( .A(p_input[1062]), .B(n2010), .Z(n2012) );
  XOR U1803 ( .A(n2013), .B(n2014), .Z(n2010) );
  AND U1804 ( .A(n430), .B(n2015), .Z(n2014) );
  XOR U1805 ( .A(n2016), .B(n2017), .Z(n2008) );
  AND U1806 ( .A(n434), .B(n2015), .Z(n2017) );
  XNOR U1807 ( .A(n2016), .B(n2013), .Z(n2015) );
  XOR U1808 ( .A(n2018), .B(n2019), .Z(n2013) );
  AND U1809 ( .A(n437), .B(n2020), .Z(n2019) );
  XOR U1810 ( .A(p_input[1094]), .B(n2018), .Z(n2020) );
  XOR U1811 ( .A(n2021), .B(n2022), .Z(n2018) );
  AND U1812 ( .A(n441), .B(n2023), .Z(n2022) );
  XOR U1813 ( .A(n2024), .B(n2025), .Z(n2016) );
  AND U1814 ( .A(n445), .B(n2023), .Z(n2025) );
  XNOR U1815 ( .A(n2024), .B(n2021), .Z(n2023) );
  XOR U1816 ( .A(n2026), .B(n2027), .Z(n2021) );
  AND U1817 ( .A(n448), .B(n2028), .Z(n2027) );
  XOR U1818 ( .A(p_input[1126]), .B(n2026), .Z(n2028) );
  XOR U1819 ( .A(n2029), .B(n2030), .Z(n2026) );
  AND U1820 ( .A(n452), .B(n2031), .Z(n2030) );
  XOR U1821 ( .A(n2032), .B(n2033), .Z(n2024) );
  AND U1822 ( .A(n456), .B(n2031), .Z(n2033) );
  XNOR U1823 ( .A(n2032), .B(n2029), .Z(n2031) );
  XOR U1824 ( .A(n2034), .B(n2035), .Z(n2029) );
  AND U1825 ( .A(n459), .B(n2036), .Z(n2035) );
  XOR U1826 ( .A(p_input[1158]), .B(n2034), .Z(n2036) );
  XOR U1827 ( .A(n2037), .B(n2038), .Z(n2034) );
  AND U1828 ( .A(n463), .B(n2039), .Z(n2038) );
  XOR U1829 ( .A(n2040), .B(n2041), .Z(n2032) );
  AND U1830 ( .A(n467), .B(n2039), .Z(n2041) );
  XNOR U1831 ( .A(n2040), .B(n2037), .Z(n2039) );
  XOR U1832 ( .A(n2042), .B(n2043), .Z(n2037) );
  AND U1833 ( .A(n470), .B(n2044), .Z(n2043) );
  XOR U1834 ( .A(p_input[1190]), .B(n2042), .Z(n2044) );
  XOR U1835 ( .A(n2045), .B(n2046), .Z(n2042) );
  AND U1836 ( .A(n474), .B(n2047), .Z(n2046) );
  XOR U1837 ( .A(n2048), .B(n2049), .Z(n2040) );
  AND U1838 ( .A(n478), .B(n2047), .Z(n2049) );
  XNOR U1839 ( .A(n2048), .B(n2045), .Z(n2047) );
  XOR U1840 ( .A(n2050), .B(n2051), .Z(n2045) );
  AND U1841 ( .A(n481), .B(n2052), .Z(n2051) );
  XOR U1842 ( .A(p_input[1222]), .B(n2050), .Z(n2052) );
  XOR U1843 ( .A(n2053), .B(n2054), .Z(n2050) );
  AND U1844 ( .A(n485), .B(n2055), .Z(n2054) );
  XOR U1845 ( .A(n2056), .B(n2057), .Z(n2048) );
  AND U1846 ( .A(n489), .B(n2055), .Z(n2057) );
  XNOR U1847 ( .A(n2056), .B(n2053), .Z(n2055) );
  XOR U1848 ( .A(n2058), .B(n2059), .Z(n2053) );
  AND U1849 ( .A(n492), .B(n2060), .Z(n2059) );
  XOR U1850 ( .A(p_input[1254]), .B(n2058), .Z(n2060) );
  XOR U1851 ( .A(n2061), .B(n2062), .Z(n2058) );
  AND U1852 ( .A(n496), .B(n2063), .Z(n2062) );
  XOR U1853 ( .A(n2064), .B(n2065), .Z(n2056) );
  AND U1854 ( .A(n500), .B(n2063), .Z(n2065) );
  XNOR U1855 ( .A(n2064), .B(n2061), .Z(n2063) );
  XOR U1856 ( .A(n2066), .B(n2067), .Z(n2061) );
  AND U1857 ( .A(n503), .B(n2068), .Z(n2067) );
  XOR U1858 ( .A(p_input[1286]), .B(n2066), .Z(n2068) );
  XOR U1859 ( .A(n2069), .B(n2070), .Z(n2066) );
  AND U1860 ( .A(n507), .B(n2071), .Z(n2070) );
  XOR U1861 ( .A(n2072), .B(n2073), .Z(n2064) );
  AND U1862 ( .A(n511), .B(n2071), .Z(n2073) );
  XNOR U1863 ( .A(n2072), .B(n2069), .Z(n2071) );
  XOR U1864 ( .A(n2074), .B(n2075), .Z(n2069) );
  AND U1865 ( .A(n514), .B(n2076), .Z(n2075) );
  XOR U1866 ( .A(p_input[1318]), .B(n2074), .Z(n2076) );
  XOR U1867 ( .A(n2077), .B(n2078), .Z(n2074) );
  AND U1868 ( .A(n518), .B(n2079), .Z(n2078) );
  XOR U1869 ( .A(n2080), .B(n2081), .Z(n2072) );
  AND U1870 ( .A(n522), .B(n2079), .Z(n2081) );
  XNOR U1871 ( .A(n2080), .B(n2077), .Z(n2079) );
  XOR U1872 ( .A(n2082), .B(n2083), .Z(n2077) );
  AND U1873 ( .A(n525), .B(n2084), .Z(n2083) );
  XOR U1874 ( .A(p_input[1350]), .B(n2082), .Z(n2084) );
  XOR U1875 ( .A(n2085), .B(n2086), .Z(n2082) );
  AND U1876 ( .A(n529), .B(n2087), .Z(n2086) );
  XOR U1877 ( .A(n2088), .B(n2089), .Z(n2080) );
  AND U1878 ( .A(n533), .B(n2087), .Z(n2089) );
  XNOR U1879 ( .A(n2088), .B(n2085), .Z(n2087) );
  XOR U1880 ( .A(n2090), .B(n2091), .Z(n2085) );
  AND U1881 ( .A(n536), .B(n2092), .Z(n2091) );
  XOR U1882 ( .A(p_input[1382]), .B(n2090), .Z(n2092) );
  XOR U1883 ( .A(n2093), .B(n2094), .Z(n2090) );
  AND U1884 ( .A(n540), .B(n2095), .Z(n2094) );
  XOR U1885 ( .A(n2096), .B(n2097), .Z(n2088) );
  AND U1886 ( .A(n544), .B(n2095), .Z(n2097) );
  XNOR U1887 ( .A(n2096), .B(n2093), .Z(n2095) );
  XOR U1888 ( .A(n2098), .B(n2099), .Z(n2093) );
  AND U1889 ( .A(n547), .B(n2100), .Z(n2099) );
  XOR U1890 ( .A(p_input[1414]), .B(n2098), .Z(n2100) );
  XOR U1891 ( .A(n2101), .B(n2102), .Z(n2098) );
  AND U1892 ( .A(n551), .B(n2103), .Z(n2102) );
  XOR U1893 ( .A(n2104), .B(n2105), .Z(n2096) );
  AND U1894 ( .A(n555), .B(n2103), .Z(n2105) );
  XNOR U1895 ( .A(n2104), .B(n2101), .Z(n2103) );
  XOR U1896 ( .A(n2106), .B(n2107), .Z(n2101) );
  AND U1897 ( .A(n558), .B(n2108), .Z(n2107) );
  XOR U1898 ( .A(p_input[1446]), .B(n2106), .Z(n2108) );
  XOR U1899 ( .A(n2109), .B(n2110), .Z(n2106) );
  AND U1900 ( .A(n562), .B(n2111), .Z(n2110) );
  XOR U1901 ( .A(n2112), .B(n2113), .Z(n2104) );
  AND U1902 ( .A(n566), .B(n2111), .Z(n2113) );
  XNOR U1903 ( .A(n2112), .B(n2109), .Z(n2111) );
  XOR U1904 ( .A(n2114), .B(n2115), .Z(n2109) );
  AND U1905 ( .A(n569), .B(n2116), .Z(n2115) );
  XOR U1906 ( .A(p_input[1478]), .B(n2114), .Z(n2116) );
  XOR U1907 ( .A(n2117), .B(n2118), .Z(n2114) );
  AND U1908 ( .A(n573), .B(n2119), .Z(n2118) );
  XOR U1909 ( .A(n2120), .B(n2121), .Z(n2112) );
  AND U1910 ( .A(n577), .B(n2119), .Z(n2121) );
  XNOR U1911 ( .A(n2120), .B(n2117), .Z(n2119) );
  XOR U1912 ( .A(n2122), .B(n2123), .Z(n2117) );
  AND U1913 ( .A(n580), .B(n2124), .Z(n2123) );
  XOR U1914 ( .A(p_input[1510]), .B(n2122), .Z(n2124) );
  XOR U1915 ( .A(n2125), .B(n2126), .Z(n2122) );
  AND U1916 ( .A(n584), .B(n2127), .Z(n2126) );
  XOR U1917 ( .A(n2128), .B(n2129), .Z(n2120) );
  AND U1918 ( .A(n588), .B(n2127), .Z(n2129) );
  XNOR U1919 ( .A(n2128), .B(n2125), .Z(n2127) );
  XOR U1920 ( .A(n2130), .B(n2131), .Z(n2125) );
  AND U1921 ( .A(n591), .B(n2132), .Z(n2131) );
  XOR U1922 ( .A(p_input[1542]), .B(n2130), .Z(n2132) );
  XOR U1923 ( .A(n2133), .B(n2134), .Z(n2130) );
  AND U1924 ( .A(n595), .B(n2135), .Z(n2134) );
  XOR U1925 ( .A(n2136), .B(n2137), .Z(n2128) );
  AND U1926 ( .A(n599), .B(n2135), .Z(n2137) );
  XNOR U1927 ( .A(n2136), .B(n2133), .Z(n2135) );
  XOR U1928 ( .A(n2138), .B(n2139), .Z(n2133) );
  AND U1929 ( .A(n602), .B(n2140), .Z(n2139) );
  XOR U1930 ( .A(p_input[1574]), .B(n2138), .Z(n2140) );
  XOR U1931 ( .A(n2141), .B(n2142), .Z(n2138) );
  AND U1932 ( .A(n606), .B(n2143), .Z(n2142) );
  XOR U1933 ( .A(n2144), .B(n2145), .Z(n2136) );
  AND U1934 ( .A(n610), .B(n2143), .Z(n2145) );
  XNOR U1935 ( .A(n2144), .B(n2141), .Z(n2143) );
  XOR U1936 ( .A(n2146), .B(n2147), .Z(n2141) );
  AND U1937 ( .A(n613), .B(n2148), .Z(n2147) );
  XOR U1938 ( .A(p_input[1606]), .B(n2146), .Z(n2148) );
  XOR U1939 ( .A(n2149), .B(n2150), .Z(n2146) );
  AND U1940 ( .A(n617), .B(n2151), .Z(n2150) );
  XOR U1941 ( .A(n2152), .B(n2153), .Z(n2144) );
  AND U1942 ( .A(n621), .B(n2151), .Z(n2153) );
  XNOR U1943 ( .A(n2152), .B(n2149), .Z(n2151) );
  XOR U1944 ( .A(n2154), .B(n2155), .Z(n2149) );
  AND U1945 ( .A(n624), .B(n2156), .Z(n2155) );
  XOR U1946 ( .A(p_input[1638]), .B(n2154), .Z(n2156) );
  XOR U1947 ( .A(n2157), .B(n2158), .Z(n2154) );
  AND U1948 ( .A(n628), .B(n2159), .Z(n2158) );
  XOR U1949 ( .A(n2160), .B(n2161), .Z(n2152) );
  AND U1950 ( .A(n632), .B(n2159), .Z(n2161) );
  XNOR U1951 ( .A(n2160), .B(n2157), .Z(n2159) );
  XOR U1952 ( .A(n2162), .B(n2163), .Z(n2157) );
  AND U1953 ( .A(n635), .B(n2164), .Z(n2163) );
  XOR U1954 ( .A(p_input[1670]), .B(n2162), .Z(n2164) );
  XOR U1955 ( .A(n2165), .B(n2166), .Z(n2162) );
  AND U1956 ( .A(n639), .B(n2167), .Z(n2166) );
  XOR U1957 ( .A(n2168), .B(n2169), .Z(n2160) );
  AND U1958 ( .A(n643), .B(n2167), .Z(n2169) );
  XNOR U1959 ( .A(n2168), .B(n2165), .Z(n2167) );
  XOR U1960 ( .A(n2170), .B(n2171), .Z(n2165) );
  AND U1961 ( .A(n646), .B(n2172), .Z(n2171) );
  XOR U1962 ( .A(p_input[1702]), .B(n2170), .Z(n2172) );
  XOR U1963 ( .A(n2173), .B(n2174), .Z(n2170) );
  AND U1964 ( .A(n650), .B(n2175), .Z(n2174) );
  XOR U1965 ( .A(n2176), .B(n2177), .Z(n2168) );
  AND U1966 ( .A(n654), .B(n2175), .Z(n2177) );
  XNOR U1967 ( .A(n2176), .B(n2173), .Z(n2175) );
  XOR U1968 ( .A(n2178), .B(n2179), .Z(n2173) );
  AND U1969 ( .A(n657), .B(n2180), .Z(n2179) );
  XOR U1970 ( .A(p_input[1734]), .B(n2178), .Z(n2180) );
  XOR U1971 ( .A(n2181), .B(n2182), .Z(n2178) );
  AND U1972 ( .A(n661), .B(n2183), .Z(n2182) );
  XOR U1973 ( .A(n2184), .B(n2185), .Z(n2176) );
  AND U1974 ( .A(n665), .B(n2183), .Z(n2185) );
  XNOR U1975 ( .A(n2184), .B(n2181), .Z(n2183) );
  XOR U1976 ( .A(n2186), .B(n2187), .Z(n2181) );
  AND U1977 ( .A(n668), .B(n2188), .Z(n2187) );
  XOR U1978 ( .A(p_input[1766]), .B(n2186), .Z(n2188) );
  XOR U1979 ( .A(n2189), .B(n2190), .Z(n2186) );
  AND U1980 ( .A(n672), .B(n2191), .Z(n2190) );
  XOR U1981 ( .A(n2192), .B(n2193), .Z(n2184) );
  AND U1982 ( .A(n676), .B(n2191), .Z(n2193) );
  XNOR U1983 ( .A(n2192), .B(n2189), .Z(n2191) );
  XOR U1984 ( .A(n2194), .B(n2195), .Z(n2189) );
  AND U1985 ( .A(n679), .B(n2196), .Z(n2195) );
  XOR U1986 ( .A(p_input[1798]), .B(n2194), .Z(n2196) );
  XOR U1987 ( .A(n2197), .B(n2198), .Z(n2194) );
  AND U1988 ( .A(n683), .B(n2199), .Z(n2198) );
  XOR U1989 ( .A(n2200), .B(n2201), .Z(n2192) );
  AND U1990 ( .A(n687), .B(n2199), .Z(n2201) );
  XNOR U1991 ( .A(n2200), .B(n2197), .Z(n2199) );
  XOR U1992 ( .A(n2202), .B(n2203), .Z(n2197) );
  AND U1993 ( .A(n690), .B(n2204), .Z(n2203) );
  XOR U1994 ( .A(p_input[1830]), .B(n2202), .Z(n2204) );
  XOR U1995 ( .A(n2205), .B(n2206), .Z(n2202) );
  AND U1996 ( .A(n694), .B(n2207), .Z(n2206) );
  XOR U1997 ( .A(n2208), .B(n2209), .Z(n2200) );
  AND U1998 ( .A(n698), .B(n2207), .Z(n2209) );
  XNOR U1999 ( .A(n2208), .B(n2205), .Z(n2207) );
  XOR U2000 ( .A(n2210), .B(n2211), .Z(n2205) );
  AND U2001 ( .A(n701), .B(n2212), .Z(n2211) );
  XOR U2002 ( .A(p_input[1862]), .B(n2210), .Z(n2212) );
  XOR U2003 ( .A(n2213), .B(n2214), .Z(n2210) );
  AND U2004 ( .A(n705), .B(n2215), .Z(n2214) );
  XOR U2005 ( .A(n2216), .B(n2217), .Z(n2208) );
  AND U2006 ( .A(n709), .B(n2215), .Z(n2217) );
  XNOR U2007 ( .A(n2216), .B(n2213), .Z(n2215) );
  XOR U2008 ( .A(n2218), .B(n2219), .Z(n2213) );
  AND U2009 ( .A(n712), .B(n2220), .Z(n2219) );
  XOR U2010 ( .A(p_input[1894]), .B(n2218), .Z(n2220) );
  XOR U2011 ( .A(n2221), .B(n2222), .Z(n2218) );
  AND U2012 ( .A(n716), .B(n2223), .Z(n2222) );
  XOR U2013 ( .A(n2224), .B(n2225), .Z(n2216) );
  AND U2014 ( .A(n720), .B(n2223), .Z(n2225) );
  XNOR U2015 ( .A(n2224), .B(n2221), .Z(n2223) );
  XOR U2016 ( .A(n2226), .B(n2227), .Z(n2221) );
  AND U2017 ( .A(n723), .B(n2228), .Z(n2227) );
  XOR U2018 ( .A(p_input[1926]), .B(n2226), .Z(n2228) );
  XOR U2019 ( .A(n2229), .B(n2230), .Z(n2226) );
  AND U2020 ( .A(n727), .B(n2231), .Z(n2230) );
  XOR U2021 ( .A(n2232), .B(n2233), .Z(n2224) );
  AND U2022 ( .A(n731), .B(n2231), .Z(n2233) );
  XNOR U2023 ( .A(n2232), .B(n2229), .Z(n2231) );
  XOR U2024 ( .A(n2234), .B(n2235), .Z(n2229) );
  AND U2025 ( .A(n734), .B(n2236), .Z(n2235) );
  XOR U2026 ( .A(p_input[1958]), .B(n2234), .Z(n2236) );
  XNOR U2027 ( .A(n2237), .B(n2238), .Z(n2234) );
  AND U2028 ( .A(n738), .B(n2239), .Z(n2238) );
  XNOR U2029 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n2240), .Z(n2232) );
  AND U2030 ( .A(n741), .B(n2239), .Z(n2240) );
  XOR U2031 ( .A(n2241), .B(n2237), .Z(n2239) );
  XOR U2032 ( .A(n17), .B(n2242), .Z(o[37]) );
  AND U2033 ( .A(n58), .B(n2243), .Z(n17) );
  XOR U2034 ( .A(n18), .B(n2242), .Z(n2243) );
  XOR U2035 ( .A(n2244), .B(n2245), .Z(n2242) );
  AND U2036 ( .A(n62), .B(n2246), .Z(n2245) );
  XOR U2037 ( .A(p_input[5]), .B(n2244), .Z(n2246) );
  XOR U2038 ( .A(n2247), .B(n2248), .Z(n2244) );
  AND U2039 ( .A(n66), .B(n2249), .Z(n2248) );
  XOR U2040 ( .A(n2250), .B(n2251), .Z(n18) );
  AND U2041 ( .A(n70), .B(n2249), .Z(n2251) );
  XNOR U2042 ( .A(n2252), .B(n2247), .Z(n2249) );
  XOR U2043 ( .A(n2253), .B(n2254), .Z(n2247) );
  AND U2044 ( .A(n74), .B(n2255), .Z(n2254) );
  XOR U2045 ( .A(p_input[37]), .B(n2253), .Z(n2255) );
  XOR U2046 ( .A(n2256), .B(n2257), .Z(n2253) );
  AND U2047 ( .A(n78), .B(n2258), .Z(n2257) );
  IV U2048 ( .A(n2250), .Z(n2252) );
  XNOR U2049 ( .A(n2259), .B(n2260), .Z(n2250) );
  AND U2050 ( .A(n82), .B(n2258), .Z(n2260) );
  XNOR U2051 ( .A(n2259), .B(n2256), .Z(n2258) );
  XOR U2052 ( .A(n2261), .B(n2262), .Z(n2256) );
  AND U2053 ( .A(n85), .B(n2263), .Z(n2262) );
  XOR U2054 ( .A(p_input[69]), .B(n2261), .Z(n2263) );
  XOR U2055 ( .A(n2264), .B(n2265), .Z(n2261) );
  AND U2056 ( .A(n89), .B(n2266), .Z(n2265) );
  XOR U2057 ( .A(n2267), .B(n2268), .Z(n2259) );
  AND U2058 ( .A(n93), .B(n2266), .Z(n2268) );
  XNOR U2059 ( .A(n2267), .B(n2264), .Z(n2266) );
  XOR U2060 ( .A(n2269), .B(n2270), .Z(n2264) );
  AND U2061 ( .A(n96), .B(n2271), .Z(n2270) );
  XOR U2062 ( .A(p_input[101]), .B(n2269), .Z(n2271) );
  XOR U2063 ( .A(n2272), .B(n2273), .Z(n2269) );
  AND U2064 ( .A(n100), .B(n2274), .Z(n2273) );
  XOR U2065 ( .A(n2275), .B(n2276), .Z(n2267) );
  AND U2066 ( .A(n104), .B(n2274), .Z(n2276) );
  XNOR U2067 ( .A(n2275), .B(n2272), .Z(n2274) );
  XOR U2068 ( .A(n2277), .B(n2278), .Z(n2272) );
  AND U2069 ( .A(n107), .B(n2279), .Z(n2278) );
  XOR U2070 ( .A(p_input[133]), .B(n2277), .Z(n2279) );
  XOR U2071 ( .A(n2280), .B(n2281), .Z(n2277) );
  AND U2072 ( .A(n111), .B(n2282), .Z(n2281) );
  XOR U2073 ( .A(n2283), .B(n2284), .Z(n2275) );
  AND U2074 ( .A(n115), .B(n2282), .Z(n2284) );
  XNOR U2075 ( .A(n2283), .B(n2280), .Z(n2282) );
  XOR U2076 ( .A(n2285), .B(n2286), .Z(n2280) );
  AND U2077 ( .A(n118), .B(n2287), .Z(n2286) );
  XOR U2078 ( .A(p_input[165]), .B(n2285), .Z(n2287) );
  XOR U2079 ( .A(n2288), .B(n2289), .Z(n2285) );
  AND U2080 ( .A(n122), .B(n2290), .Z(n2289) );
  XOR U2081 ( .A(n2291), .B(n2292), .Z(n2283) );
  AND U2082 ( .A(n126), .B(n2290), .Z(n2292) );
  XNOR U2083 ( .A(n2291), .B(n2288), .Z(n2290) );
  XOR U2084 ( .A(n2293), .B(n2294), .Z(n2288) );
  AND U2085 ( .A(n129), .B(n2295), .Z(n2294) );
  XOR U2086 ( .A(p_input[197]), .B(n2293), .Z(n2295) );
  XOR U2087 ( .A(n2296), .B(n2297), .Z(n2293) );
  AND U2088 ( .A(n133), .B(n2298), .Z(n2297) );
  XOR U2089 ( .A(n2299), .B(n2300), .Z(n2291) );
  AND U2090 ( .A(n137), .B(n2298), .Z(n2300) );
  XNOR U2091 ( .A(n2299), .B(n2296), .Z(n2298) );
  XOR U2092 ( .A(n2301), .B(n2302), .Z(n2296) );
  AND U2093 ( .A(n140), .B(n2303), .Z(n2302) );
  XOR U2094 ( .A(p_input[229]), .B(n2301), .Z(n2303) );
  XOR U2095 ( .A(n2304), .B(n2305), .Z(n2301) );
  AND U2096 ( .A(n144), .B(n2306), .Z(n2305) );
  XOR U2097 ( .A(n2307), .B(n2308), .Z(n2299) );
  AND U2098 ( .A(n148), .B(n2306), .Z(n2308) );
  XNOR U2099 ( .A(n2307), .B(n2304), .Z(n2306) );
  XOR U2100 ( .A(n2309), .B(n2310), .Z(n2304) );
  AND U2101 ( .A(n151), .B(n2311), .Z(n2310) );
  XOR U2102 ( .A(p_input[261]), .B(n2309), .Z(n2311) );
  XOR U2103 ( .A(n2312), .B(n2313), .Z(n2309) );
  AND U2104 ( .A(n155), .B(n2314), .Z(n2313) );
  XOR U2105 ( .A(n2315), .B(n2316), .Z(n2307) );
  AND U2106 ( .A(n159), .B(n2314), .Z(n2316) );
  XNOR U2107 ( .A(n2315), .B(n2312), .Z(n2314) );
  XOR U2108 ( .A(n2317), .B(n2318), .Z(n2312) );
  AND U2109 ( .A(n162), .B(n2319), .Z(n2318) );
  XOR U2110 ( .A(p_input[293]), .B(n2317), .Z(n2319) );
  XOR U2111 ( .A(n2320), .B(n2321), .Z(n2317) );
  AND U2112 ( .A(n166), .B(n2322), .Z(n2321) );
  XOR U2113 ( .A(n2323), .B(n2324), .Z(n2315) );
  AND U2114 ( .A(n170), .B(n2322), .Z(n2324) );
  XNOR U2115 ( .A(n2323), .B(n2320), .Z(n2322) );
  XOR U2116 ( .A(n2325), .B(n2326), .Z(n2320) );
  AND U2117 ( .A(n173), .B(n2327), .Z(n2326) );
  XOR U2118 ( .A(p_input[325]), .B(n2325), .Z(n2327) );
  XOR U2119 ( .A(n2328), .B(n2329), .Z(n2325) );
  AND U2120 ( .A(n177), .B(n2330), .Z(n2329) );
  XOR U2121 ( .A(n2331), .B(n2332), .Z(n2323) );
  AND U2122 ( .A(n181), .B(n2330), .Z(n2332) );
  XNOR U2123 ( .A(n2331), .B(n2328), .Z(n2330) );
  XOR U2124 ( .A(n2333), .B(n2334), .Z(n2328) );
  AND U2125 ( .A(n184), .B(n2335), .Z(n2334) );
  XOR U2126 ( .A(p_input[357]), .B(n2333), .Z(n2335) );
  XOR U2127 ( .A(n2336), .B(n2337), .Z(n2333) );
  AND U2128 ( .A(n188), .B(n2338), .Z(n2337) );
  XOR U2129 ( .A(n2339), .B(n2340), .Z(n2331) );
  AND U2130 ( .A(n192), .B(n2338), .Z(n2340) );
  XNOR U2131 ( .A(n2339), .B(n2336), .Z(n2338) );
  XOR U2132 ( .A(n2341), .B(n2342), .Z(n2336) );
  AND U2133 ( .A(n195), .B(n2343), .Z(n2342) );
  XOR U2134 ( .A(p_input[389]), .B(n2341), .Z(n2343) );
  XOR U2135 ( .A(n2344), .B(n2345), .Z(n2341) );
  AND U2136 ( .A(n199), .B(n2346), .Z(n2345) );
  XOR U2137 ( .A(n2347), .B(n2348), .Z(n2339) );
  AND U2138 ( .A(n203), .B(n2346), .Z(n2348) );
  XNOR U2139 ( .A(n2347), .B(n2344), .Z(n2346) );
  XOR U2140 ( .A(n2349), .B(n2350), .Z(n2344) );
  AND U2141 ( .A(n206), .B(n2351), .Z(n2350) );
  XOR U2142 ( .A(p_input[421]), .B(n2349), .Z(n2351) );
  XOR U2143 ( .A(n2352), .B(n2353), .Z(n2349) );
  AND U2144 ( .A(n210), .B(n2354), .Z(n2353) );
  XOR U2145 ( .A(n2355), .B(n2356), .Z(n2347) );
  AND U2146 ( .A(n214), .B(n2354), .Z(n2356) );
  XNOR U2147 ( .A(n2355), .B(n2352), .Z(n2354) );
  XOR U2148 ( .A(n2357), .B(n2358), .Z(n2352) );
  AND U2149 ( .A(n217), .B(n2359), .Z(n2358) );
  XOR U2150 ( .A(p_input[453]), .B(n2357), .Z(n2359) );
  XOR U2151 ( .A(n2360), .B(n2361), .Z(n2357) );
  AND U2152 ( .A(n221), .B(n2362), .Z(n2361) );
  XOR U2153 ( .A(n2363), .B(n2364), .Z(n2355) );
  AND U2154 ( .A(n225), .B(n2362), .Z(n2364) );
  XNOR U2155 ( .A(n2363), .B(n2360), .Z(n2362) );
  XOR U2156 ( .A(n2365), .B(n2366), .Z(n2360) );
  AND U2157 ( .A(n228), .B(n2367), .Z(n2366) );
  XOR U2158 ( .A(p_input[485]), .B(n2365), .Z(n2367) );
  XOR U2159 ( .A(n2368), .B(n2369), .Z(n2365) );
  AND U2160 ( .A(n232), .B(n2370), .Z(n2369) );
  XOR U2161 ( .A(n2371), .B(n2372), .Z(n2363) );
  AND U2162 ( .A(n236), .B(n2370), .Z(n2372) );
  XNOR U2163 ( .A(n2371), .B(n2368), .Z(n2370) );
  XOR U2164 ( .A(n2373), .B(n2374), .Z(n2368) );
  AND U2165 ( .A(n239), .B(n2375), .Z(n2374) );
  XOR U2166 ( .A(p_input[517]), .B(n2373), .Z(n2375) );
  XOR U2167 ( .A(n2376), .B(n2377), .Z(n2373) );
  AND U2168 ( .A(n243), .B(n2378), .Z(n2377) );
  XOR U2169 ( .A(n2379), .B(n2380), .Z(n2371) );
  AND U2170 ( .A(n247), .B(n2378), .Z(n2380) );
  XNOR U2171 ( .A(n2379), .B(n2376), .Z(n2378) );
  XOR U2172 ( .A(n2381), .B(n2382), .Z(n2376) );
  AND U2173 ( .A(n250), .B(n2383), .Z(n2382) );
  XOR U2174 ( .A(p_input[549]), .B(n2381), .Z(n2383) );
  XOR U2175 ( .A(n2384), .B(n2385), .Z(n2381) );
  AND U2176 ( .A(n254), .B(n2386), .Z(n2385) );
  XOR U2177 ( .A(n2387), .B(n2388), .Z(n2379) );
  AND U2178 ( .A(n258), .B(n2386), .Z(n2388) );
  XNOR U2179 ( .A(n2387), .B(n2384), .Z(n2386) );
  XOR U2180 ( .A(n2389), .B(n2390), .Z(n2384) );
  AND U2181 ( .A(n261), .B(n2391), .Z(n2390) );
  XOR U2182 ( .A(p_input[581]), .B(n2389), .Z(n2391) );
  XOR U2183 ( .A(n2392), .B(n2393), .Z(n2389) );
  AND U2184 ( .A(n265), .B(n2394), .Z(n2393) );
  XOR U2185 ( .A(n2395), .B(n2396), .Z(n2387) );
  AND U2186 ( .A(n269), .B(n2394), .Z(n2396) );
  XNOR U2187 ( .A(n2395), .B(n2392), .Z(n2394) );
  XOR U2188 ( .A(n2397), .B(n2398), .Z(n2392) );
  AND U2189 ( .A(n272), .B(n2399), .Z(n2398) );
  XOR U2190 ( .A(p_input[613]), .B(n2397), .Z(n2399) );
  XOR U2191 ( .A(n2400), .B(n2401), .Z(n2397) );
  AND U2192 ( .A(n276), .B(n2402), .Z(n2401) );
  XOR U2193 ( .A(n2403), .B(n2404), .Z(n2395) );
  AND U2194 ( .A(n280), .B(n2402), .Z(n2404) );
  XNOR U2195 ( .A(n2403), .B(n2400), .Z(n2402) );
  XOR U2196 ( .A(n2405), .B(n2406), .Z(n2400) );
  AND U2197 ( .A(n283), .B(n2407), .Z(n2406) );
  XOR U2198 ( .A(p_input[645]), .B(n2405), .Z(n2407) );
  XOR U2199 ( .A(n2408), .B(n2409), .Z(n2405) );
  AND U2200 ( .A(n287), .B(n2410), .Z(n2409) );
  XOR U2201 ( .A(n2411), .B(n2412), .Z(n2403) );
  AND U2202 ( .A(n291), .B(n2410), .Z(n2412) );
  XNOR U2203 ( .A(n2411), .B(n2408), .Z(n2410) );
  XOR U2204 ( .A(n2413), .B(n2414), .Z(n2408) );
  AND U2205 ( .A(n294), .B(n2415), .Z(n2414) );
  XOR U2206 ( .A(p_input[677]), .B(n2413), .Z(n2415) );
  XOR U2207 ( .A(n2416), .B(n2417), .Z(n2413) );
  AND U2208 ( .A(n298), .B(n2418), .Z(n2417) );
  XOR U2209 ( .A(n2419), .B(n2420), .Z(n2411) );
  AND U2210 ( .A(n302), .B(n2418), .Z(n2420) );
  XNOR U2211 ( .A(n2419), .B(n2416), .Z(n2418) );
  XOR U2212 ( .A(n2421), .B(n2422), .Z(n2416) );
  AND U2213 ( .A(n305), .B(n2423), .Z(n2422) );
  XOR U2214 ( .A(p_input[709]), .B(n2421), .Z(n2423) );
  XOR U2215 ( .A(n2424), .B(n2425), .Z(n2421) );
  AND U2216 ( .A(n309), .B(n2426), .Z(n2425) );
  XOR U2217 ( .A(n2427), .B(n2428), .Z(n2419) );
  AND U2218 ( .A(n313), .B(n2426), .Z(n2428) );
  XNOR U2219 ( .A(n2427), .B(n2424), .Z(n2426) );
  XOR U2220 ( .A(n2429), .B(n2430), .Z(n2424) );
  AND U2221 ( .A(n316), .B(n2431), .Z(n2430) );
  XOR U2222 ( .A(p_input[741]), .B(n2429), .Z(n2431) );
  XOR U2223 ( .A(n2432), .B(n2433), .Z(n2429) );
  AND U2224 ( .A(n320), .B(n2434), .Z(n2433) );
  XOR U2225 ( .A(n2435), .B(n2436), .Z(n2427) );
  AND U2226 ( .A(n324), .B(n2434), .Z(n2436) );
  XNOR U2227 ( .A(n2435), .B(n2432), .Z(n2434) );
  XOR U2228 ( .A(n2437), .B(n2438), .Z(n2432) );
  AND U2229 ( .A(n327), .B(n2439), .Z(n2438) );
  XOR U2230 ( .A(p_input[773]), .B(n2437), .Z(n2439) );
  XOR U2231 ( .A(n2440), .B(n2441), .Z(n2437) );
  AND U2232 ( .A(n331), .B(n2442), .Z(n2441) );
  XOR U2233 ( .A(n2443), .B(n2444), .Z(n2435) );
  AND U2234 ( .A(n335), .B(n2442), .Z(n2444) );
  XNOR U2235 ( .A(n2443), .B(n2440), .Z(n2442) );
  XOR U2236 ( .A(n2445), .B(n2446), .Z(n2440) );
  AND U2237 ( .A(n338), .B(n2447), .Z(n2446) );
  XOR U2238 ( .A(p_input[805]), .B(n2445), .Z(n2447) );
  XOR U2239 ( .A(n2448), .B(n2449), .Z(n2445) );
  AND U2240 ( .A(n342), .B(n2450), .Z(n2449) );
  XOR U2241 ( .A(n2451), .B(n2452), .Z(n2443) );
  AND U2242 ( .A(n346), .B(n2450), .Z(n2452) );
  XNOR U2243 ( .A(n2451), .B(n2448), .Z(n2450) );
  XOR U2244 ( .A(n2453), .B(n2454), .Z(n2448) );
  AND U2245 ( .A(n349), .B(n2455), .Z(n2454) );
  XOR U2246 ( .A(p_input[837]), .B(n2453), .Z(n2455) );
  XOR U2247 ( .A(n2456), .B(n2457), .Z(n2453) );
  AND U2248 ( .A(n353), .B(n2458), .Z(n2457) );
  XOR U2249 ( .A(n2459), .B(n2460), .Z(n2451) );
  AND U2250 ( .A(n357), .B(n2458), .Z(n2460) );
  XNOR U2251 ( .A(n2459), .B(n2456), .Z(n2458) );
  XOR U2252 ( .A(n2461), .B(n2462), .Z(n2456) );
  AND U2253 ( .A(n360), .B(n2463), .Z(n2462) );
  XOR U2254 ( .A(p_input[869]), .B(n2461), .Z(n2463) );
  XOR U2255 ( .A(n2464), .B(n2465), .Z(n2461) );
  AND U2256 ( .A(n364), .B(n2466), .Z(n2465) );
  XOR U2257 ( .A(n2467), .B(n2468), .Z(n2459) );
  AND U2258 ( .A(n368), .B(n2466), .Z(n2468) );
  XNOR U2259 ( .A(n2467), .B(n2464), .Z(n2466) );
  XOR U2260 ( .A(n2469), .B(n2470), .Z(n2464) );
  AND U2261 ( .A(n371), .B(n2471), .Z(n2470) );
  XOR U2262 ( .A(p_input[901]), .B(n2469), .Z(n2471) );
  XOR U2263 ( .A(n2472), .B(n2473), .Z(n2469) );
  AND U2264 ( .A(n375), .B(n2474), .Z(n2473) );
  XOR U2265 ( .A(n2475), .B(n2476), .Z(n2467) );
  AND U2266 ( .A(n379), .B(n2474), .Z(n2476) );
  XNOR U2267 ( .A(n2475), .B(n2472), .Z(n2474) );
  XOR U2268 ( .A(n2477), .B(n2478), .Z(n2472) );
  AND U2269 ( .A(n382), .B(n2479), .Z(n2478) );
  XOR U2270 ( .A(p_input[933]), .B(n2477), .Z(n2479) );
  XOR U2271 ( .A(n2480), .B(n2481), .Z(n2477) );
  AND U2272 ( .A(n386), .B(n2482), .Z(n2481) );
  XOR U2273 ( .A(n2483), .B(n2484), .Z(n2475) );
  AND U2274 ( .A(n390), .B(n2482), .Z(n2484) );
  XNOR U2275 ( .A(n2483), .B(n2480), .Z(n2482) );
  XOR U2276 ( .A(n2485), .B(n2486), .Z(n2480) );
  AND U2277 ( .A(n393), .B(n2487), .Z(n2486) );
  XOR U2278 ( .A(p_input[965]), .B(n2485), .Z(n2487) );
  XOR U2279 ( .A(n2488), .B(n2489), .Z(n2485) );
  AND U2280 ( .A(n397), .B(n2490), .Z(n2489) );
  XOR U2281 ( .A(n2491), .B(n2492), .Z(n2483) );
  AND U2282 ( .A(n401), .B(n2490), .Z(n2492) );
  XNOR U2283 ( .A(n2491), .B(n2488), .Z(n2490) );
  XOR U2284 ( .A(n2493), .B(n2494), .Z(n2488) );
  AND U2285 ( .A(n404), .B(n2495), .Z(n2494) );
  XOR U2286 ( .A(p_input[997]), .B(n2493), .Z(n2495) );
  XOR U2287 ( .A(n2496), .B(n2497), .Z(n2493) );
  AND U2288 ( .A(n408), .B(n2498), .Z(n2497) );
  XOR U2289 ( .A(n2499), .B(n2500), .Z(n2491) );
  AND U2290 ( .A(n412), .B(n2498), .Z(n2500) );
  XNOR U2291 ( .A(n2499), .B(n2496), .Z(n2498) );
  XOR U2292 ( .A(n2501), .B(n2502), .Z(n2496) );
  AND U2293 ( .A(n415), .B(n2503), .Z(n2502) );
  XOR U2294 ( .A(p_input[1029]), .B(n2501), .Z(n2503) );
  XOR U2295 ( .A(n2504), .B(n2505), .Z(n2501) );
  AND U2296 ( .A(n419), .B(n2506), .Z(n2505) );
  XOR U2297 ( .A(n2507), .B(n2508), .Z(n2499) );
  AND U2298 ( .A(n423), .B(n2506), .Z(n2508) );
  XNOR U2299 ( .A(n2507), .B(n2504), .Z(n2506) );
  XOR U2300 ( .A(n2509), .B(n2510), .Z(n2504) );
  AND U2301 ( .A(n426), .B(n2511), .Z(n2510) );
  XOR U2302 ( .A(p_input[1061]), .B(n2509), .Z(n2511) );
  XOR U2303 ( .A(n2512), .B(n2513), .Z(n2509) );
  AND U2304 ( .A(n430), .B(n2514), .Z(n2513) );
  XOR U2305 ( .A(n2515), .B(n2516), .Z(n2507) );
  AND U2306 ( .A(n434), .B(n2514), .Z(n2516) );
  XNOR U2307 ( .A(n2515), .B(n2512), .Z(n2514) );
  XOR U2308 ( .A(n2517), .B(n2518), .Z(n2512) );
  AND U2309 ( .A(n437), .B(n2519), .Z(n2518) );
  XOR U2310 ( .A(p_input[1093]), .B(n2517), .Z(n2519) );
  XOR U2311 ( .A(n2520), .B(n2521), .Z(n2517) );
  AND U2312 ( .A(n441), .B(n2522), .Z(n2521) );
  XOR U2313 ( .A(n2523), .B(n2524), .Z(n2515) );
  AND U2314 ( .A(n445), .B(n2522), .Z(n2524) );
  XNOR U2315 ( .A(n2523), .B(n2520), .Z(n2522) );
  XOR U2316 ( .A(n2525), .B(n2526), .Z(n2520) );
  AND U2317 ( .A(n448), .B(n2527), .Z(n2526) );
  XOR U2318 ( .A(p_input[1125]), .B(n2525), .Z(n2527) );
  XOR U2319 ( .A(n2528), .B(n2529), .Z(n2525) );
  AND U2320 ( .A(n452), .B(n2530), .Z(n2529) );
  XOR U2321 ( .A(n2531), .B(n2532), .Z(n2523) );
  AND U2322 ( .A(n456), .B(n2530), .Z(n2532) );
  XNOR U2323 ( .A(n2531), .B(n2528), .Z(n2530) );
  XOR U2324 ( .A(n2533), .B(n2534), .Z(n2528) );
  AND U2325 ( .A(n459), .B(n2535), .Z(n2534) );
  XOR U2326 ( .A(p_input[1157]), .B(n2533), .Z(n2535) );
  XOR U2327 ( .A(n2536), .B(n2537), .Z(n2533) );
  AND U2328 ( .A(n463), .B(n2538), .Z(n2537) );
  XOR U2329 ( .A(n2539), .B(n2540), .Z(n2531) );
  AND U2330 ( .A(n467), .B(n2538), .Z(n2540) );
  XNOR U2331 ( .A(n2539), .B(n2536), .Z(n2538) );
  XOR U2332 ( .A(n2541), .B(n2542), .Z(n2536) );
  AND U2333 ( .A(n470), .B(n2543), .Z(n2542) );
  XOR U2334 ( .A(p_input[1189]), .B(n2541), .Z(n2543) );
  XOR U2335 ( .A(n2544), .B(n2545), .Z(n2541) );
  AND U2336 ( .A(n474), .B(n2546), .Z(n2545) );
  XOR U2337 ( .A(n2547), .B(n2548), .Z(n2539) );
  AND U2338 ( .A(n478), .B(n2546), .Z(n2548) );
  XNOR U2339 ( .A(n2547), .B(n2544), .Z(n2546) );
  XOR U2340 ( .A(n2549), .B(n2550), .Z(n2544) );
  AND U2341 ( .A(n481), .B(n2551), .Z(n2550) );
  XOR U2342 ( .A(p_input[1221]), .B(n2549), .Z(n2551) );
  XOR U2343 ( .A(n2552), .B(n2553), .Z(n2549) );
  AND U2344 ( .A(n485), .B(n2554), .Z(n2553) );
  XOR U2345 ( .A(n2555), .B(n2556), .Z(n2547) );
  AND U2346 ( .A(n489), .B(n2554), .Z(n2556) );
  XNOR U2347 ( .A(n2555), .B(n2552), .Z(n2554) );
  XOR U2348 ( .A(n2557), .B(n2558), .Z(n2552) );
  AND U2349 ( .A(n492), .B(n2559), .Z(n2558) );
  XOR U2350 ( .A(p_input[1253]), .B(n2557), .Z(n2559) );
  XOR U2351 ( .A(n2560), .B(n2561), .Z(n2557) );
  AND U2352 ( .A(n496), .B(n2562), .Z(n2561) );
  XOR U2353 ( .A(n2563), .B(n2564), .Z(n2555) );
  AND U2354 ( .A(n500), .B(n2562), .Z(n2564) );
  XNOR U2355 ( .A(n2563), .B(n2560), .Z(n2562) );
  XOR U2356 ( .A(n2565), .B(n2566), .Z(n2560) );
  AND U2357 ( .A(n503), .B(n2567), .Z(n2566) );
  XOR U2358 ( .A(p_input[1285]), .B(n2565), .Z(n2567) );
  XOR U2359 ( .A(n2568), .B(n2569), .Z(n2565) );
  AND U2360 ( .A(n507), .B(n2570), .Z(n2569) );
  XOR U2361 ( .A(n2571), .B(n2572), .Z(n2563) );
  AND U2362 ( .A(n511), .B(n2570), .Z(n2572) );
  XNOR U2363 ( .A(n2571), .B(n2568), .Z(n2570) );
  XOR U2364 ( .A(n2573), .B(n2574), .Z(n2568) );
  AND U2365 ( .A(n514), .B(n2575), .Z(n2574) );
  XOR U2366 ( .A(p_input[1317]), .B(n2573), .Z(n2575) );
  XOR U2367 ( .A(n2576), .B(n2577), .Z(n2573) );
  AND U2368 ( .A(n518), .B(n2578), .Z(n2577) );
  XOR U2369 ( .A(n2579), .B(n2580), .Z(n2571) );
  AND U2370 ( .A(n522), .B(n2578), .Z(n2580) );
  XNOR U2371 ( .A(n2579), .B(n2576), .Z(n2578) );
  XOR U2372 ( .A(n2581), .B(n2582), .Z(n2576) );
  AND U2373 ( .A(n525), .B(n2583), .Z(n2582) );
  XOR U2374 ( .A(p_input[1349]), .B(n2581), .Z(n2583) );
  XOR U2375 ( .A(n2584), .B(n2585), .Z(n2581) );
  AND U2376 ( .A(n529), .B(n2586), .Z(n2585) );
  XOR U2377 ( .A(n2587), .B(n2588), .Z(n2579) );
  AND U2378 ( .A(n533), .B(n2586), .Z(n2588) );
  XNOR U2379 ( .A(n2587), .B(n2584), .Z(n2586) );
  XOR U2380 ( .A(n2589), .B(n2590), .Z(n2584) );
  AND U2381 ( .A(n536), .B(n2591), .Z(n2590) );
  XOR U2382 ( .A(p_input[1381]), .B(n2589), .Z(n2591) );
  XOR U2383 ( .A(n2592), .B(n2593), .Z(n2589) );
  AND U2384 ( .A(n540), .B(n2594), .Z(n2593) );
  XOR U2385 ( .A(n2595), .B(n2596), .Z(n2587) );
  AND U2386 ( .A(n544), .B(n2594), .Z(n2596) );
  XNOR U2387 ( .A(n2595), .B(n2592), .Z(n2594) );
  XOR U2388 ( .A(n2597), .B(n2598), .Z(n2592) );
  AND U2389 ( .A(n547), .B(n2599), .Z(n2598) );
  XOR U2390 ( .A(p_input[1413]), .B(n2597), .Z(n2599) );
  XOR U2391 ( .A(n2600), .B(n2601), .Z(n2597) );
  AND U2392 ( .A(n551), .B(n2602), .Z(n2601) );
  XOR U2393 ( .A(n2603), .B(n2604), .Z(n2595) );
  AND U2394 ( .A(n555), .B(n2602), .Z(n2604) );
  XNOR U2395 ( .A(n2603), .B(n2600), .Z(n2602) );
  XOR U2396 ( .A(n2605), .B(n2606), .Z(n2600) );
  AND U2397 ( .A(n558), .B(n2607), .Z(n2606) );
  XOR U2398 ( .A(p_input[1445]), .B(n2605), .Z(n2607) );
  XOR U2399 ( .A(n2608), .B(n2609), .Z(n2605) );
  AND U2400 ( .A(n562), .B(n2610), .Z(n2609) );
  XOR U2401 ( .A(n2611), .B(n2612), .Z(n2603) );
  AND U2402 ( .A(n566), .B(n2610), .Z(n2612) );
  XNOR U2403 ( .A(n2611), .B(n2608), .Z(n2610) );
  XOR U2404 ( .A(n2613), .B(n2614), .Z(n2608) );
  AND U2405 ( .A(n569), .B(n2615), .Z(n2614) );
  XOR U2406 ( .A(p_input[1477]), .B(n2613), .Z(n2615) );
  XOR U2407 ( .A(n2616), .B(n2617), .Z(n2613) );
  AND U2408 ( .A(n573), .B(n2618), .Z(n2617) );
  XOR U2409 ( .A(n2619), .B(n2620), .Z(n2611) );
  AND U2410 ( .A(n577), .B(n2618), .Z(n2620) );
  XNOR U2411 ( .A(n2619), .B(n2616), .Z(n2618) );
  XOR U2412 ( .A(n2621), .B(n2622), .Z(n2616) );
  AND U2413 ( .A(n580), .B(n2623), .Z(n2622) );
  XOR U2414 ( .A(p_input[1509]), .B(n2621), .Z(n2623) );
  XOR U2415 ( .A(n2624), .B(n2625), .Z(n2621) );
  AND U2416 ( .A(n584), .B(n2626), .Z(n2625) );
  XOR U2417 ( .A(n2627), .B(n2628), .Z(n2619) );
  AND U2418 ( .A(n588), .B(n2626), .Z(n2628) );
  XNOR U2419 ( .A(n2627), .B(n2624), .Z(n2626) );
  XOR U2420 ( .A(n2629), .B(n2630), .Z(n2624) );
  AND U2421 ( .A(n591), .B(n2631), .Z(n2630) );
  XOR U2422 ( .A(p_input[1541]), .B(n2629), .Z(n2631) );
  XOR U2423 ( .A(n2632), .B(n2633), .Z(n2629) );
  AND U2424 ( .A(n595), .B(n2634), .Z(n2633) );
  XOR U2425 ( .A(n2635), .B(n2636), .Z(n2627) );
  AND U2426 ( .A(n599), .B(n2634), .Z(n2636) );
  XNOR U2427 ( .A(n2635), .B(n2632), .Z(n2634) );
  XOR U2428 ( .A(n2637), .B(n2638), .Z(n2632) );
  AND U2429 ( .A(n602), .B(n2639), .Z(n2638) );
  XOR U2430 ( .A(p_input[1573]), .B(n2637), .Z(n2639) );
  XOR U2431 ( .A(n2640), .B(n2641), .Z(n2637) );
  AND U2432 ( .A(n606), .B(n2642), .Z(n2641) );
  XOR U2433 ( .A(n2643), .B(n2644), .Z(n2635) );
  AND U2434 ( .A(n610), .B(n2642), .Z(n2644) );
  XNOR U2435 ( .A(n2643), .B(n2640), .Z(n2642) );
  XOR U2436 ( .A(n2645), .B(n2646), .Z(n2640) );
  AND U2437 ( .A(n613), .B(n2647), .Z(n2646) );
  XOR U2438 ( .A(p_input[1605]), .B(n2645), .Z(n2647) );
  XOR U2439 ( .A(n2648), .B(n2649), .Z(n2645) );
  AND U2440 ( .A(n617), .B(n2650), .Z(n2649) );
  XOR U2441 ( .A(n2651), .B(n2652), .Z(n2643) );
  AND U2442 ( .A(n621), .B(n2650), .Z(n2652) );
  XNOR U2443 ( .A(n2651), .B(n2648), .Z(n2650) );
  XOR U2444 ( .A(n2653), .B(n2654), .Z(n2648) );
  AND U2445 ( .A(n624), .B(n2655), .Z(n2654) );
  XOR U2446 ( .A(p_input[1637]), .B(n2653), .Z(n2655) );
  XOR U2447 ( .A(n2656), .B(n2657), .Z(n2653) );
  AND U2448 ( .A(n628), .B(n2658), .Z(n2657) );
  XOR U2449 ( .A(n2659), .B(n2660), .Z(n2651) );
  AND U2450 ( .A(n632), .B(n2658), .Z(n2660) );
  XNOR U2451 ( .A(n2659), .B(n2656), .Z(n2658) );
  XOR U2452 ( .A(n2661), .B(n2662), .Z(n2656) );
  AND U2453 ( .A(n635), .B(n2663), .Z(n2662) );
  XOR U2454 ( .A(p_input[1669]), .B(n2661), .Z(n2663) );
  XOR U2455 ( .A(n2664), .B(n2665), .Z(n2661) );
  AND U2456 ( .A(n639), .B(n2666), .Z(n2665) );
  XOR U2457 ( .A(n2667), .B(n2668), .Z(n2659) );
  AND U2458 ( .A(n643), .B(n2666), .Z(n2668) );
  XNOR U2459 ( .A(n2667), .B(n2664), .Z(n2666) );
  XOR U2460 ( .A(n2669), .B(n2670), .Z(n2664) );
  AND U2461 ( .A(n646), .B(n2671), .Z(n2670) );
  XOR U2462 ( .A(p_input[1701]), .B(n2669), .Z(n2671) );
  XOR U2463 ( .A(n2672), .B(n2673), .Z(n2669) );
  AND U2464 ( .A(n650), .B(n2674), .Z(n2673) );
  XOR U2465 ( .A(n2675), .B(n2676), .Z(n2667) );
  AND U2466 ( .A(n654), .B(n2674), .Z(n2676) );
  XNOR U2467 ( .A(n2675), .B(n2672), .Z(n2674) );
  XOR U2468 ( .A(n2677), .B(n2678), .Z(n2672) );
  AND U2469 ( .A(n657), .B(n2679), .Z(n2678) );
  XOR U2470 ( .A(p_input[1733]), .B(n2677), .Z(n2679) );
  XOR U2471 ( .A(n2680), .B(n2681), .Z(n2677) );
  AND U2472 ( .A(n661), .B(n2682), .Z(n2681) );
  XOR U2473 ( .A(n2683), .B(n2684), .Z(n2675) );
  AND U2474 ( .A(n665), .B(n2682), .Z(n2684) );
  XNOR U2475 ( .A(n2683), .B(n2680), .Z(n2682) );
  XOR U2476 ( .A(n2685), .B(n2686), .Z(n2680) );
  AND U2477 ( .A(n668), .B(n2687), .Z(n2686) );
  XOR U2478 ( .A(p_input[1765]), .B(n2685), .Z(n2687) );
  XOR U2479 ( .A(n2688), .B(n2689), .Z(n2685) );
  AND U2480 ( .A(n672), .B(n2690), .Z(n2689) );
  XOR U2481 ( .A(n2691), .B(n2692), .Z(n2683) );
  AND U2482 ( .A(n676), .B(n2690), .Z(n2692) );
  XNOR U2483 ( .A(n2691), .B(n2688), .Z(n2690) );
  XOR U2484 ( .A(n2693), .B(n2694), .Z(n2688) );
  AND U2485 ( .A(n679), .B(n2695), .Z(n2694) );
  XOR U2486 ( .A(p_input[1797]), .B(n2693), .Z(n2695) );
  XOR U2487 ( .A(n2696), .B(n2697), .Z(n2693) );
  AND U2488 ( .A(n683), .B(n2698), .Z(n2697) );
  XOR U2489 ( .A(n2699), .B(n2700), .Z(n2691) );
  AND U2490 ( .A(n687), .B(n2698), .Z(n2700) );
  XNOR U2491 ( .A(n2699), .B(n2696), .Z(n2698) );
  XOR U2492 ( .A(n2701), .B(n2702), .Z(n2696) );
  AND U2493 ( .A(n690), .B(n2703), .Z(n2702) );
  XOR U2494 ( .A(p_input[1829]), .B(n2701), .Z(n2703) );
  XOR U2495 ( .A(n2704), .B(n2705), .Z(n2701) );
  AND U2496 ( .A(n694), .B(n2706), .Z(n2705) );
  XOR U2497 ( .A(n2707), .B(n2708), .Z(n2699) );
  AND U2498 ( .A(n698), .B(n2706), .Z(n2708) );
  XNOR U2499 ( .A(n2707), .B(n2704), .Z(n2706) );
  XOR U2500 ( .A(n2709), .B(n2710), .Z(n2704) );
  AND U2501 ( .A(n701), .B(n2711), .Z(n2710) );
  XOR U2502 ( .A(p_input[1861]), .B(n2709), .Z(n2711) );
  XOR U2503 ( .A(n2712), .B(n2713), .Z(n2709) );
  AND U2504 ( .A(n705), .B(n2714), .Z(n2713) );
  XOR U2505 ( .A(n2715), .B(n2716), .Z(n2707) );
  AND U2506 ( .A(n709), .B(n2714), .Z(n2716) );
  XNOR U2507 ( .A(n2715), .B(n2712), .Z(n2714) );
  XOR U2508 ( .A(n2717), .B(n2718), .Z(n2712) );
  AND U2509 ( .A(n712), .B(n2719), .Z(n2718) );
  XOR U2510 ( .A(p_input[1893]), .B(n2717), .Z(n2719) );
  XOR U2511 ( .A(n2720), .B(n2721), .Z(n2717) );
  AND U2512 ( .A(n716), .B(n2722), .Z(n2721) );
  XOR U2513 ( .A(n2723), .B(n2724), .Z(n2715) );
  AND U2514 ( .A(n720), .B(n2722), .Z(n2724) );
  XNOR U2515 ( .A(n2723), .B(n2720), .Z(n2722) );
  XOR U2516 ( .A(n2725), .B(n2726), .Z(n2720) );
  AND U2517 ( .A(n723), .B(n2727), .Z(n2726) );
  XOR U2518 ( .A(p_input[1925]), .B(n2725), .Z(n2727) );
  XOR U2519 ( .A(n2728), .B(n2729), .Z(n2725) );
  AND U2520 ( .A(n727), .B(n2730), .Z(n2729) );
  XOR U2521 ( .A(n2731), .B(n2732), .Z(n2723) );
  AND U2522 ( .A(n731), .B(n2730), .Z(n2732) );
  XNOR U2523 ( .A(n2731), .B(n2728), .Z(n2730) );
  XOR U2524 ( .A(n2733), .B(n2734), .Z(n2728) );
  AND U2525 ( .A(n734), .B(n2735), .Z(n2734) );
  XOR U2526 ( .A(p_input[1957]), .B(n2733), .Z(n2735) );
  XNOR U2527 ( .A(n2736), .B(n2737), .Z(n2733) );
  AND U2528 ( .A(n738), .B(n2738), .Z(n2737) );
  XNOR U2529 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n2739), .Z(n2731) );
  AND U2530 ( .A(n741), .B(n2738), .Z(n2739) );
  XOR U2531 ( .A(n2740), .B(n2736), .Z(n2738) );
  IV U2532 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .Z(n2736) );
  IV U2533 ( .A(\knn_comb_/min_val_out[0][5] ), .Z(n2740) );
  XOR U2534 ( .A(n39), .B(n2741), .Z(o[36]) );
  AND U2535 ( .A(n58), .B(n2742), .Z(n39) );
  XOR U2536 ( .A(n40), .B(n2741), .Z(n2742) );
  XOR U2537 ( .A(n2743), .B(n2744), .Z(n2741) );
  AND U2538 ( .A(n62), .B(n2745), .Z(n2744) );
  XOR U2539 ( .A(p_input[4]), .B(n2743), .Z(n2745) );
  XOR U2540 ( .A(n2746), .B(n2747), .Z(n2743) );
  AND U2541 ( .A(n66), .B(n2748), .Z(n2747) );
  XOR U2542 ( .A(n2749), .B(n2750), .Z(n40) );
  AND U2543 ( .A(n70), .B(n2748), .Z(n2750) );
  XNOR U2544 ( .A(n2751), .B(n2746), .Z(n2748) );
  XOR U2545 ( .A(n2752), .B(n2753), .Z(n2746) );
  AND U2546 ( .A(n74), .B(n2754), .Z(n2753) );
  XOR U2547 ( .A(p_input[36]), .B(n2752), .Z(n2754) );
  XOR U2548 ( .A(n2755), .B(n2756), .Z(n2752) );
  AND U2549 ( .A(n78), .B(n2757), .Z(n2756) );
  IV U2550 ( .A(n2749), .Z(n2751) );
  XNOR U2551 ( .A(n2758), .B(n2759), .Z(n2749) );
  AND U2552 ( .A(n82), .B(n2757), .Z(n2759) );
  XNOR U2553 ( .A(n2758), .B(n2755), .Z(n2757) );
  XOR U2554 ( .A(n2760), .B(n2761), .Z(n2755) );
  AND U2555 ( .A(n85), .B(n2762), .Z(n2761) );
  XOR U2556 ( .A(p_input[68]), .B(n2760), .Z(n2762) );
  XOR U2557 ( .A(n2763), .B(n2764), .Z(n2760) );
  AND U2558 ( .A(n89), .B(n2765), .Z(n2764) );
  XOR U2559 ( .A(n2766), .B(n2767), .Z(n2758) );
  AND U2560 ( .A(n93), .B(n2765), .Z(n2767) );
  XNOR U2561 ( .A(n2766), .B(n2763), .Z(n2765) );
  XOR U2562 ( .A(n2768), .B(n2769), .Z(n2763) );
  AND U2563 ( .A(n96), .B(n2770), .Z(n2769) );
  XOR U2564 ( .A(p_input[100]), .B(n2768), .Z(n2770) );
  XOR U2565 ( .A(n2771), .B(n2772), .Z(n2768) );
  AND U2566 ( .A(n100), .B(n2773), .Z(n2772) );
  XOR U2567 ( .A(n2774), .B(n2775), .Z(n2766) );
  AND U2568 ( .A(n104), .B(n2773), .Z(n2775) );
  XNOR U2569 ( .A(n2774), .B(n2771), .Z(n2773) );
  XOR U2570 ( .A(n2776), .B(n2777), .Z(n2771) );
  AND U2571 ( .A(n107), .B(n2778), .Z(n2777) );
  XOR U2572 ( .A(p_input[132]), .B(n2776), .Z(n2778) );
  XOR U2573 ( .A(n2779), .B(n2780), .Z(n2776) );
  AND U2574 ( .A(n111), .B(n2781), .Z(n2780) );
  XOR U2575 ( .A(n2782), .B(n2783), .Z(n2774) );
  AND U2576 ( .A(n115), .B(n2781), .Z(n2783) );
  XNOR U2577 ( .A(n2782), .B(n2779), .Z(n2781) );
  XOR U2578 ( .A(n2784), .B(n2785), .Z(n2779) );
  AND U2579 ( .A(n118), .B(n2786), .Z(n2785) );
  XOR U2580 ( .A(p_input[164]), .B(n2784), .Z(n2786) );
  XOR U2581 ( .A(n2787), .B(n2788), .Z(n2784) );
  AND U2582 ( .A(n122), .B(n2789), .Z(n2788) );
  XOR U2583 ( .A(n2790), .B(n2791), .Z(n2782) );
  AND U2584 ( .A(n126), .B(n2789), .Z(n2791) );
  XNOR U2585 ( .A(n2790), .B(n2787), .Z(n2789) );
  XOR U2586 ( .A(n2792), .B(n2793), .Z(n2787) );
  AND U2587 ( .A(n129), .B(n2794), .Z(n2793) );
  XOR U2588 ( .A(p_input[196]), .B(n2792), .Z(n2794) );
  XOR U2589 ( .A(n2795), .B(n2796), .Z(n2792) );
  AND U2590 ( .A(n133), .B(n2797), .Z(n2796) );
  XOR U2591 ( .A(n2798), .B(n2799), .Z(n2790) );
  AND U2592 ( .A(n137), .B(n2797), .Z(n2799) );
  XNOR U2593 ( .A(n2798), .B(n2795), .Z(n2797) );
  XOR U2594 ( .A(n2800), .B(n2801), .Z(n2795) );
  AND U2595 ( .A(n140), .B(n2802), .Z(n2801) );
  XOR U2596 ( .A(p_input[228]), .B(n2800), .Z(n2802) );
  XOR U2597 ( .A(n2803), .B(n2804), .Z(n2800) );
  AND U2598 ( .A(n144), .B(n2805), .Z(n2804) );
  XOR U2599 ( .A(n2806), .B(n2807), .Z(n2798) );
  AND U2600 ( .A(n148), .B(n2805), .Z(n2807) );
  XNOR U2601 ( .A(n2806), .B(n2803), .Z(n2805) );
  XOR U2602 ( .A(n2808), .B(n2809), .Z(n2803) );
  AND U2603 ( .A(n151), .B(n2810), .Z(n2809) );
  XOR U2604 ( .A(p_input[260]), .B(n2808), .Z(n2810) );
  XOR U2605 ( .A(n2811), .B(n2812), .Z(n2808) );
  AND U2606 ( .A(n155), .B(n2813), .Z(n2812) );
  XOR U2607 ( .A(n2814), .B(n2815), .Z(n2806) );
  AND U2608 ( .A(n159), .B(n2813), .Z(n2815) );
  XNOR U2609 ( .A(n2814), .B(n2811), .Z(n2813) );
  XOR U2610 ( .A(n2816), .B(n2817), .Z(n2811) );
  AND U2611 ( .A(n162), .B(n2818), .Z(n2817) );
  XOR U2612 ( .A(p_input[292]), .B(n2816), .Z(n2818) );
  XOR U2613 ( .A(n2819), .B(n2820), .Z(n2816) );
  AND U2614 ( .A(n166), .B(n2821), .Z(n2820) );
  XOR U2615 ( .A(n2822), .B(n2823), .Z(n2814) );
  AND U2616 ( .A(n170), .B(n2821), .Z(n2823) );
  XNOR U2617 ( .A(n2822), .B(n2819), .Z(n2821) );
  XOR U2618 ( .A(n2824), .B(n2825), .Z(n2819) );
  AND U2619 ( .A(n173), .B(n2826), .Z(n2825) );
  XOR U2620 ( .A(p_input[324]), .B(n2824), .Z(n2826) );
  XOR U2621 ( .A(n2827), .B(n2828), .Z(n2824) );
  AND U2622 ( .A(n177), .B(n2829), .Z(n2828) );
  XOR U2623 ( .A(n2830), .B(n2831), .Z(n2822) );
  AND U2624 ( .A(n181), .B(n2829), .Z(n2831) );
  XNOR U2625 ( .A(n2830), .B(n2827), .Z(n2829) );
  XOR U2626 ( .A(n2832), .B(n2833), .Z(n2827) );
  AND U2627 ( .A(n184), .B(n2834), .Z(n2833) );
  XOR U2628 ( .A(p_input[356]), .B(n2832), .Z(n2834) );
  XOR U2629 ( .A(n2835), .B(n2836), .Z(n2832) );
  AND U2630 ( .A(n188), .B(n2837), .Z(n2836) );
  XOR U2631 ( .A(n2838), .B(n2839), .Z(n2830) );
  AND U2632 ( .A(n192), .B(n2837), .Z(n2839) );
  XNOR U2633 ( .A(n2838), .B(n2835), .Z(n2837) );
  XOR U2634 ( .A(n2840), .B(n2841), .Z(n2835) );
  AND U2635 ( .A(n195), .B(n2842), .Z(n2841) );
  XOR U2636 ( .A(p_input[388]), .B(n2840), .Z(n2842) );
  XOR U2637 ( .A(n2843), .B(n2844), .Z(n2840) );
  AND U2638 ( .A(n199), .B(n2845), .Z(n2844) );
  XOR U2639 ( .A(n2846), .B(n2847), .Z(n2838) );
  AND U2640 ( .A(n203), .B(n2845), .Z(n2847) );
  XNOR U2641 ( .A(n2846), .B(n2843), .Z(n2845) );
  XOR U2642 ( .A(n2848), .B(n2849), .Z(n2843) );
  AND U2643 ( .A(n206), .B(n2850), .Z(n2849) );
  XOR U2644 ( .A(p_input[420]), .B(n2848), .Z(n2850) );
  XOR U2645 ( .A(n2851), .B(n2852), .Z(n2848) );
  AND U2646 ( .A(n210), .B(n2853), .Z(n2852) );
  XOR U2647 ( .A(n2854), .B(n2855), .Z(n2846) );
  AND U2648 ( .A(n214), .B(n2853), .Z(n2855) );
  XNOR U2649 ( .A(n2854), .B(n2851), .Z(n2853) );
  XOR U2650 ( .A(n2856), .B(n2857), .Z(n2851) );
  AND U2651 ( .A(n217), .B(n2858), .Z(n2857) );
  XOR U2652 ( .A(p_input[452]), .B(n2856), .Z(n2858) );
  XOR U2653 ( .A(n2859), .B(n2860), .Z(n2856) );
  AND U2654 ( .A(n221), .B(n2861), .Z(n2860) );
  XOR U2655 ( .A(n2862), .B(n2863), .Z(n2854) );
  AND U2656 ( .A(n225), .B(n2861), .Z(n2863) );
  XNOR U2657 ( .A(n2862), .B(n2859), .Z(n2861) );
  XOR U2658 ( .A(n2864), .B(n2865), .Z(n2859) );
  AND U2659 ( .A(n228), .B(n2866), .Z(n2865) );
  XOR U2660 ( .A(p_input[484]), .B(n2864), .Z(n2866) );
  XOR U2661 ( .A(n2867), .B(n2868), .Z(n2864) );
  AND U2662 ( .A(n232), .B(n2869), .Z(n2868) );
  XOR U2663 ( .A(n2870), .B(n2871), .Z(n2862) );
  AND U2664 ( .A(n236), .B(n2869), .Z(n2871) );
  XNOR U2665 ( .A(n2870), .B(n2867), .Z(n2869) );
  XOR U2666 ( .A(n2872), .B(n2873), .Z(n2867) );
  AND U2667 ( .A(n239), .B(n2874), .Z(n2873) );
  XOR U2668 ( .A(p_input[516]), .B(n2872), .Z(n2874) );
  XOR U2669 ( .A(n2875), .B(n2876), .Z(n2872) );
  AND U2670 ( .A(n243), .B(n2877), .Z(n2876) );
  XOR U2671 ( .A(n2878), .B(n2879), .Z(n2870) );
  AND U2672 ( .A(n247), .B(n2877), .Z(n2879) );
  XNOR U2673 ( .A(n2878), .B(n2875), .Z(n2877) );
  XOR U2674 ( .A(n2880), .B(n2881), .Z(n2875) );
  AND U2675 ( .A(n250), .B(n2882), .Z(n2881) );
  XOR U2676 ( .A(p_input[548]), .B(n2880), .Z(n2882) );
  XOR U2677 ( .A(n2883), .B(n2884), .Z(n2880) );
  AND U2678 ( .A(n254), .B(n2885), .Z(n2884) );
  XOR U2679 ( .A(n2886), .B(n2887), .Z(n2878) );
  AND U2680 ( .A(n258), .B(n2885), .Z(n2887) );
  XNOR U2681 ( .A(n2886), .B(n2883), .Z(n2885) );
  XOR U2682 ( .A(n2888), .B(n2889), .Z(n2883) );
  AND U2683 ( .A(n261), .B(n2890), .Z(n2889) );
  XOR U2684 ( .A(p_input[580]), .B(n2888), .Z(n2890) );
  XOR U2685 ( .A(n2891), .B(n2892), .Z(n2888) );
  AND U2686 ( .A(n265), .B(n2893), .Z(n2892) );
  XOR U2687 ( .A(n2894), .B(n2895), .Z(n2886) );
  AND U2688 ( .A(n269), .B(n2893), .Z(n2895) );
  XNOR U2689 ( .A(n2894), .B(n2891), .Z(n2893) );
  XOR U2690 ( .A(n2896), .B(n2897), .Z(n2891) );
  AND U2691 ( .A(n272), .B(n2898), .Z(n2897) );
  XOR U2692 ( .A(p_input[612]), .B(n2896), .Z(n2898) );
  XOR U2693 ( .A(n2899), .B(n2900), .Z(n2896) );
  AND U2694 ( .A(n276), .B(n2901), .Z(n2900) );
  XOR U2695 ( .A(n2902), .B(n2903), .Z(n2894) );
  AND U2696 ( .A(n280), .B(n2901), .Z(n2903) );
  XNOR U2697 ( .A(n2902), .B(n2899), .Z(n2901) );
  XOR U2698 ( .A(n2904), .B(n2905), .Z(n2899) );
  AND U2699 ( .A(n283), .B(n2906), .Z(n2905) );
  XOR U2700 ( .A(p_input[644]), .B(n2904), .Z(n2906) );
  XOR U2701 ( .A(n2907), .B(n2908), .Z(n2904) );
  AND U2702 ( .A(n287), .B(n2909), .Z(n2908) );
  XOR U2703 ( .A(n2910), .B(n2911), .Z(n2902) );
  AND U2704 ( .A(n291), .B(n2909), .Z(n2911) );
  XNOR U2705 ( .A(n2910), .B(n2907), .Z(n2909) );
  XOR U2706 ( .A(n2912), .B(n2913), .Z(n2907) );
  AND U2707 ( .A(n294), .B(n2914), .Z(n2913) );
  XOR U2708 ( .A(p_input[676]), .B(n2912), .Z(n2914) );
  XOR U2709 ( .A(n2915), .B(n2916), .Z(n2912) );
  AND U2710 ( .A(n298), .B(n2917), .Z(n2916) );
  XOR U2711 ( .A(n2918), .B(n2919), .Z(n2910) );
  AND U2712 ( .A(n302), .B(n2917), .Z(n2919) );
  XNOR U2713 ( .A(n2918), .B(n2915), .Z(n2917) );
  XOR U2714 ( .A(n2920), .B(n2921), .Z(n2915) );
  AND U2715 ( .A(n305), .B(n2922), .Z(n2921) );
  XOR U2716 ( .A(p_input[708]), .B(n2920), .Z(n2922) );
  XOR U2717 ( .A(n2923), .B(n2924), .Z(n2920) );
  AND U2718 ( .A(n309), .B(n2925), .Z(n2924) );
  XOR U2719 ( .A(n2926), .B(n2927), .Z(n2918) );
  AND U2720 ( .A(n313), .B(n2925), .Z(n2927) );
  XNOR U2721 ( .A(n2926), .B(n2923), .Z(n2925) );
  XOR U2722 ( .A(n2928), .B(n2929), .Z(n2923) );
  AND U2723 ( .A(n316), .B(n2930), .Z(n2929) );
  XOR U2724 ( .A(p_input[740]), .B(n2928), .Z(n2930) );
  XOR U2725 ( .A(n2931), .B(n2932), .Z(n2928) );
  AND U2726 ( .A(n320), .B(n2933), .Z(n2932) );
  XOR U2727 ( .A(n2934), .B(n2935), .Z(n2926) );
  AND U2728 ( .A(n324), .B(n2933), .Z(n2935) );
  XNOR U2729 ( .A(n2934), .B(n2931), .Z(n2933) );
  XOR U2730 ( .A(n2936), .B(n2937), .Z(n2931) );
  AND U2731 ( .A(n327), .B(n2938), .Z(n2937) );
  XOR U2732 ( .A(p_input[772]), .B(n2936), .Z(n2938) );
  XOR U2733 ( .A(n2939), .B(n2940), .Z(n2936) );
  AND U2734 ( .A(n331), .B(n2941), .Z(n2940) );
  XOR U2735 ( .A(n2942), .B(n2943), .Z(n2934) );
  AND U2736 ( .A(n335), .B(n2941), .Z(n2943) );
  XNOR U2737 ( .A(n2942), .B(n2939), .Z(n2941) );
  XOR U2738 ( .A(n2944), .B(n2945), .Z(n2939) );
  AND U2739 ( .A(n338), .B(n2946), .Z(n2945) );
  XOR U2740 ( .A(p_input[804]), .B(n2944), .Z(n2946) );
  XOR U2741 ( .A(n2947), .B(n2948), .Z(n2944) );
  AND U2742 ( .A(n342), .B(n2949), .Z(n2948) );
  XOR U2743 ( .A(n2950), .B(n2951), .Z(n2942) );
  AND U2744 ( .A(n346), .B(n2949), .Z(n2951) );
  XNOR U2745 ( .A(n2950), .B(n2947), .Z(n2949) );
  XOR U2746 ( .A(n2952), .B(n2953), .Z(n2947) );
  AND U2747 ( .A(n349), .B(n2954), .Z(n2953) );
  XOR U2748 ( .A(p_input[836]), .B(n2952), .Z(n2954) );
  XOR U2749 ( .A(n2955), .B(n2956), .Z(n2952) );
  AND U2750 ( .A(n353), .B(n2957), .Z(n2956) );
  XOR U2751 ( .A(n2958), .B(n2959), .Z(n2950) );
  AND U2752 ( .A(n357), .B(n2957), .Z(n2959) );
  XNOR U2753 ( .A(n2958), .B(n2955), .Z(n2957) );
  XOR U2754 ( .A(n2960), .B(n2961), .Z(n2955) );
  AND U2755 ( .A(n360), .B(n2962), .Z(n2961) );
  XOR U2756 ( .A(p_input[868]), .B(n2960), .Z(n2962) );
  XOR U2757 ( .A(n2963), .B(n2964), .Z(n2960) );
  AND U2758 ( .A(n364), .B(n2965), .Z(n2964) );
  XOR U2759 ( .A(n2966), .B(n2967), .Z(n2958) );
  AND U2760 ( .A(n368), .B(n2965), .Z(n2967) );
  XNOR U2761 ( .A(n2966), .B(n2963), .Z(n2965) );
  XOR U2762 ( .A(n2968), .B(n2969), .Z(n2963) );
  AND U2763 ( .A(n371), .B(n2970), .Z(n2969) );
  XOR U2764 ( .A(p_input[900]), .B(n2968), .Z(n2970) );
  XOR U2765 ( .A(n2971), .B(n2972), .Z(n2968) );
  AND U2766 ( .A(n375), .B(n2973), .Z(n2972) );
  XOR U2767 ( .A(n2974), .B(n2975), .Z(n2966) );
  AND U2768 ( .A(n379), .B(n2973), .Z(n2975) );
  XNOR U2769 ( .A(n2974), .B(n2971), .Z(n2973) );
  XOR U2770 ( .A(n2976), .B(n2977), .Z(n2971) );
  AND U2771 ( .A(n382), .B(n2978), .Z(n2977) );
  XOR U2772 ( .A(p_input[932]), .B(n2976), .Z(n2978) );
  XOR U2773 ( .A(n2979), .B(n2980), .Z(n2976) );
  AND U2774 ( .A(n386), .B(n2981), .Z(n2980) );
  XOR U2775 ( .A(n2982), .B(n2983), .Z(n2974) );
  AND U2776 ( .A(n390), .B(n2981), .Z(n2983) );
  XNOR U2777 ( .A(n2982), .B(n2979), .Z(n2981) );
  XOR U2778 ( .A(n2984), .B(n2985), .Z(n2979) );
  AND U2779 ( .A(n393), .B(n2986), .Z(n2985) );
  XOR U2780 ( .A(p_input[964]), .B(n2984), .Z(n2986) );
  XOR U2781 ( .A(n2987), .B(n2988), .Z(n2984) );
  AND U2782 ( .A(n397), .B(n2989), .Z(n2988) );
  XOR U2783 ( .A(n2990), .B(n2991), .Z(n2982) );
  AND U2784 ( .A(n401), .B(n2989), .Z(n2991) );
  XNOR U2785 ( .A(n2990), .B(n2987), .Z(n2989) );
  XOR U2786 ( .A(n2992), .B(n2993), .Z(n2987) );
  AND U2787 ( .A(n404), .B(n2994), .Z(n2993) );
  XOR U2788 ( .A(p_input[996]), .B(n2992), .Z(n2994) );
  XOR U2789 ( .A(n2995), .B(n2996), .Z(n2992) );
  AND U2790 ( .A(n408), .B(n2997), .Z(n2996) );
  XOR U2791 ( .A(n2998), .B(n2999), .Z(n2990) );
  AND U2792 ( .A(n412), .B(n2997), .Z(n2999) );
  XNOR U2793 ( .A(n2998), .B(n2995), .Z(n2997) );
  XOR U2794 ( .A(n3000), .B(n3001), .Z(n2995) );
  AND U2795 ( .A(n415), .B(n3002), .Z(n3001) );
  XOR U2796 ( .A(p_input[1028]), .B(n3000), .Z(n3002) );
  XOR U2797 ( .A(n3003), .B(n3004), .Z(n3000) );
  AND U2798 ( .A(n419), .B(n3005), .Z(n3004) );
  XOR U2799 ( .A(n3006), .B(n3007), .Z(n2998) );
  AND U2800 ( .A(n423), .B(n3005), .Z(n3007) );
  XNOR U2801 ( .A(n3006), .B(n3003), .Z(n3005) );
  XOR U2802 ( .A(n3008), .B(n3009), .Z(n3003) );
  AND U2803 ( .A(n426), .B(n3010), .Z(n3009) );
  XOR U2804 ( .A(p_input[1060]), .B(n3008), .Z(n3010) );
  XOR U2805 ( .A(n3011), .B(n3012), .Z(n3008) );
  AND U2806 ( .A(n430), .B(n3013), .Z(n3012) );
  XOR U2807 ( .A(n3014), .B(n3015), .Z(n3006) );
  AND U2808 ( .A(n434), .B(n3013), .Z(n3015) );
  XNOR U2809 ( .A(n3014), .B(n3011), .Z(n3013) );
  XOR U2810 ( .A(n3016), .B(n3017), .Z(n3011) );
  AND U2811 ( .A(n437), .B(n3018), .Z(n3017) );
  XOR U2812 ( .A(p_input[1092]), .B(n3016), .Z(n3018) );
  XOR U2813 ( .A(n3019), .B(n3020), .Z(n3016) );
  AND U2814 ( .A(n441), .B(n3021), .Z(n3020) );
  XOR U2815 ( .A(n3022), .B(n3023), .Z(n3014) );
  AND U2816 ( .A(n445), .B(n3021), .Z(n3023) );
  XNOR U2817 ( .A(n3022), .B(n3019), .Z(n3021) );
  XOR U2818 ( .A(n3024), .B(n3025), .Z(n3019) );
  AND U2819 ( .A(n448), .B(n3026), .Z(n3025) );
  XOR U2820 ( .A(p_input[1124]), .B(n3024), .Z(n3026) );
  XOR U2821 ( .A(n3027), .B(n3028), .Z(n3024) );
  AND U2822 ( .A(n452), .B(n3029), .Z(n3028) );
  XOR U2823 ( .A(n3030), .B(n3031), .Z(n3022) );
  AND U2824 ( .A(n456), .B(n3029), .Z(n3031) );
  XNOR U2825 ( .A(n3030), .B(n3027), .Z(n3029) );
  XOR U2826 ( .A(n3032), .B(n3033), .Z(n3027) );
  AND U2827 ( .A(n459), .B(n3034), .Z(n3033) );
  XOR U2828 ( .A(p_input[1156]), .B(n3032), .Z(n3034) );
  XOR U2829 ( .A(n3035), .B(n3036), .Z(n3032) );
  AND U2830 ( .A(n463), .B(n3037), .Z(n3036) );
  XOR U2831 ( .A(n3038), .B(n3039), .Z(n3030) );
  AND U2832 ( .A(n467), .B(n3037), .Z(n3039) );
  XNOR U2833 ( .A(n3038), .B(n3035), .Z(n3037) );
  XOR U2834 ( .A(n3040), .B(n3041), .Z(n3035) );
  AND U2835 ( .A(n470), .B(n3042), .Z(n3041) );
  XOR U2836 ( .A(p_input[1188]), .B(n3040), .Z(n3042) );
  XOR U2837 ( .A(n3043), .B(n3044), .Z(n3040) );
  AND U2838 ( .A(n474), .B(n3045), .Z(n3044) );
  XOR U2839 ( .A(n3046), .B(n3047), .Z(n3038) );
  AND U2840 ( .A(n478), .B(n3045), .Z(n3047) );
  XNOR U2841 ( .A(n3046), .B(n3043), .Z(n3045) );
  XOR U2842 ( .A(n3048), .B(n3049), .Z(n3043) );
  AND U2843 ( .A(n481), .B(n3050), .Z(n3049) );
  XOR U2844 ( .A(p_input[1220]), .B(n3048), .Z(n3050) );
  XOR U2845 ( .A(n3051), .B(n3052), .Z(n3048) );
  AND U2846 ( .A(n485), .B(n3053), .Z(n3052) );
  XOR U2847 ( .A(n3054), .B(n3055), .Z(n3046) );
  AND U2848 ( .A(n489), .B(n3053), .Z(n3055) );
  XNOR U2849 ( .A(n3054), .B(n3051), .Z(n3053) );
  XOR U2850 ( .A(n3056), .B(n3057), .Z(n3051) );
  AND U2851 ( .A(n492), .B(n3058), .Z(n3057) );
  XOR U2852 ( .A(p_input[1252]), .B(n3056), .Z(n3058) );
  XOR U2853 ( .A(n3059), .B(n3060), .Z(n3056) );
  AND U2854 ( .A(n496), .B(n3061), .Z(n3060) );
  XOR U2855 ( .A(n3062), .B(n3063), .Z(n3054) );
  AND U2856 ( .A(n500), .B(n3061), .Z(n3063) );
  XNOR U2857 ( .A(n3062), .B(n3059), .Z(n3061) );
  XOR U2858 ( .A(n3064), .B(n3065), .Z(n3059) );
  AND U2859 ( .A(n503), .B(n3066), .Z(n3065) );
  XOR U2860 ( .A(p_input[1284]), .B(n3064), .Z(n3066) );
  XOR U2861 ( .A(n3067), .B(n3068), .Z(n3064) );
  AND U2862 ( .A(n507), .B(n3069), .Z(n3068) );
  XOR U2863 ( .A(n3070), .B(n3071), .Z(n3062) );
  AND U2864 ( .A(n511), .B(n3069), .Z(n3071) );
  XNOR U2865 ( .A(n3070), .B(n3067), .Z(n3069) );
  XOR U2866 ( .A(n3072), .B(n3073), .Z(n3067) );
  AND U2867 ( .A(n514), .B(n3074), .Z(n3073) );
  XOR U2868 ( .A(p_input[1316]), .B(n3072), .Z(n3074) );
  XOR U2869 ( .A(n3075), .B(n3076), .Z(n3072) );
  AND U2870 ( .A(n518), .B(n3077), .Z(n3076) );
  XOR U2871 ( .A(n3078), .B(n3079), .Z(n3070) );
  AND U2872 ( .A(n522), .B(n3077), .Z(n3079) );
  XNOR U2873 ( .A(n3078), .B(n3075), .Z(n3077) );
  XOR U2874 ( .A(n3080), .B(n3081), .Z(n3075) );
  AND U2875 ( .A(n525), .B(n3082), .Z(n3081) );
  XOR U2876 ( .A(p_input[1348]), .B(n3080), .Z(n3082) );
  XOR U2877 ( .A(n3083), .B(n3084), .Z(n3080) );
  AND U2878 ( .A(n529), .B(n3085), .Z(n3084) );
  XOR U2879 ( .A(n3086), .B(n3087), .Z(n3078) );
  AND U2880 ( .A(n533), .B(n3085), .Z(n3087) );
  XNOR U2881 ( .A(n3086), .B(n3083), .Z(n3085) );
  XOR U2882 ( .A(n3088), .B(n3089), .Z(n3083) );
  AND U2883 ( .A(n536), .B(n3090), .Z(n3089) );
  XOR U2884 ( .A(p_input[1380]), .B(n3088), .Z(n3090) );
  XOR U2885 ( .A(n3091), .B(n3092), .Z(n3088) );
  AND U2886 ( .A(n540), .B(n3093), .Z(n3092) );
  XOR U2887 ( .A(n3094), .B(n3095), .Z(n3086) );
  AND U2888 ( .A(n544), .B(n3093), .Z(n3095) );
  XNOR U2889 ( .A(n3094), .B(n3091), .Z(n3093) );
  XOR U2890 ( .A(n3096), .B(n3097), .Z(n3091) );
  AND U2891 ( .A(n547), .B(n3098), .Z(n3097) );
  XOR U2892 ( .A(p_input[1412]), .B(n3096), .Z(n3098) );
  XOR U2893 ( .A(n3099), .B(n3100), .Z(n3096) );
  AND U2894 ( .A(n551), .B(n3101), .Z(n3100) );
  XOR U2895 ( .A(n3102), .B(n3103), .Z(n3094) );
  AND U2896 ( .A(n555), .B(n3101), .Z(n3103) );
  XNOR U2897 ( .A(n3102), .B(n3099), .Z(n3101) );
  XOR U2898 ( .A(n3104), .B(n3105), .Z(n3099) );
  AND U2899 ( .A(n558), .B(n3106), .Z(n3105) );
  XOR U2900 ( .A(p_input[1444]), .B(n3104), .Z(n3106) );
  XOR U2901 ( .A(n3107), .B(n3108), .Z(n3104) );
  AND U2902 ( .A(n562), .B(n3109), .Z(n3108) );
  XOR U2903 ( .A(n3110), .B(n3111), .Z(n3102) );
  AND U2904 ( .A(n566), .B(n3109), .Z(n3111) );
  XNOR U2905 ( .A(n3110), .B(n3107), .Z(n3109) );
  XOR U2906 ( .A(n3112), .B(n3113), .Z(n3107) );
  AND U2907 ( .A(n569), .B(n3114), .Z(n3113) );
  XOR U2908 ( .A(p_input[1476]), .B(n3112), .Z(n3114) );
  XOR U2909 ( .A(n3115), .B(n3116), .Z(n3112) );
  AND U2910 ( .A(n573), .B(n3117), .Z(n3116) );
  XOR U2911 ( .A(n3118), .B(n3119), .Z(n3110) );
  AND U2912 ( .A(n577), .B(n3117), .Z(n3119) );
  XNOR U2913 ( .A(n3118), .B(n3115), .Z(n3117) );
  XOR U2914 ( .A(n3120), .B(n3121), .Z(n3115) );
  AND U2915 ( .A(n580), .B(n3122), .Z(n3121) );
  XOR U2916 ( .A(p_input[1508]), .B(n3120), .Z(n3122) );
  XOR U2917 ( .A(n3123), .B(n3124), .Z(n3120) );
  AND U2918 ( .A(n584), .B(n3125), .Z(n3124) );
  XOR U2919 ( .A(n3126), .B(n3127), .Z(n3118) );
  AND U2920 ( .A(n588), .B(n3125), .Z(n3127) );
  XNOR U2921 ( .A(n3126), .B(n3123), .Z(n3125) );
  XOR U2922 ( .A(n3128), .B(n3129), .Z(n3123) );
  AND U2923 ( .A(n591), .B(n3130), .Z(n3129) );
  XOR U2924 ( .A(p_input[1540]), .B(n3128), .Z(n3130) );
  XOR U2925 ( .A(n3131), .B(n3132), .Z(n3128) );
  AND U2926 ( .A(n595), .B(n3133), .Z(n3132) );
  XOR U2927 ( .A(n3134), .B(n3135), .Z(n3126) );
  AND U2928 ( .A(n599), .B(n3133), .Z(n3135) );
  XNOR U2929 ( .A(n3134), .B(n3131), .Z(n3133) );
  XOR U2930 ( .A(n3136), .B(n3137), .Z(n3131) );
  AND U2931 ( .A(n602), .B(n3138), .Z(n3137) );
  XOR U2932 ( .A(p_input[1572]), .B(n3136), .Z(n3138) );
  XOR U2933 ( .A(n3139), .B(n3140), .Z(n3136) );
  AND U2934 ( .A(n606), .B(n3141), .Z(n3140) );
  XOR U2935 ( .A(n3142), .B(n3143), .Z(n3134) );
  AND U2936 ( .A(n610), .B(n3141), .Z(n3143) );
  XNOR U2937 ( .A(n3142), .B(n3139), .Z(n3141) );
  XOR U2938 ( .A(n3144), .B(n3145), .Z(n3139) );
  AND U2939 ( .A(n613), .B(n3146), .Z(n3145) );
  XOR U2940 ( .A(p_input[1604]), .B(n3144), .Z(n3146) );
  XOR U2941 ( .A(n3147), .B(n3148), .Z(n3144) );
  AND U2942 ( .A(n617), .B(n3149), .Z(n3148) );
  XOR U2943 ( .A(n3150), .B(n3151), .Z(n3142) );
  AND U2944 ( .A(n621), .B(n3149), .Z(n3151) );
  XNOR U2945 ( .A(n3150), .B(n3147), .Z(n3149) );
  XOR U2946 ( .A(n3152), .B(n3153), .Z(n3147) );
  AND U2947 ( .A(n624), .B(n3154), .Z(n3153) );
  XOR U2948 ( .A(p_input[1636]), .B(n3152), .Z(n3154) );
  XOR U2949 ( .A(n3155), .B(n3156), .Z(n3152) );
  AND U2950 ( .A(n628), .B(n3157), .Z(n3156) );
  XOR U2951 ( .A(n3158), .B(n3159), .Z(n3150) );
  AND U2952 ( .A(n632), .B(n3157), .Z(n3159) );
  XNOR U2953 ( .A(n3158), .B(n3155), .Z(n3157) );
  XOR U2954 ( .A(n3160), .B(n3161), .Z(n3155) );
  AND U2955 ( .A(n635), .B(n3162), .Z(n3161) );
  XOR U2956 ( .A(p_input[1668]), .B(n3160), .Z(n3162) );
  XOR U2957 ( .A(n3163), .B(n3164), .Z(n3160) );
  AND U2958 ( .A(n639), .B(n3165), .Z(n3164) );
  XOR U2959 ( .A(n3166), .B(n3167), .Z(n3158) );
  AND U2960 ( .A(n643), .B(n3165), .Z(n3167) );
  XNOR U2961 ( .A(n3166), .B(n3163), .Z(n3165) );
  XOR U2962 ( .A(n3168), .B(n3169), .Z(n3163) );
  AND U2963 ( .A(n646), .B(n3170), .Z(n3169) );
  XOR U2964 ( .A(p_input[1700]), .B(n3168), .Z(n3170) );
  XOR U2965 ( .A(n3171), .B(n3172), .Z(n3168) );
  AND U2966 ( .A(n650), .B(n3173), .Z(n3172) );
  XOR U2967 ( .A(n3174), .B(n3175), .Z(n3166) );
  AND U2968 ( .A(n654), .B(n3173), .Z(n3175) );
  XNOR U2969 ( .A(n3174), .B(n3171), .Z(n3173) );
  XOR U2970 ( .A(n3176), .B(n3177), .Z(n3171) );
  AND U2971 ( .A(n657), .B(n3178), .Z(n3177) );
  XOR U2972 ( .A(p_input[1732]), .B(n3176), .Z(n3178) );
  XOR U2973 ( .A(n3179), .B(n3180), .Z(n3176) );
  AND U2974 ( .A(n661), .B(n3181), .Z(n3180) );
  XOR U2975 ( .A(n3182), .B(n3183), .Z(n3174) );
  AND U2976 ( .A(n665), .B(n3181), .Z(n3183) );
  XNOR U2977 ( .A(n3182), .B(n3179), .Z(n3181) );
  XOR U2978 ( .A(n3184), .B(n3185), .Z(n3179) );
  AND U2979 ( .A(n668), .B(n3186), .Z(n3185) );
  XOR U2980 ( .A(p_input[1764]), .B(n3184), .Z(n3186) );
  XOR U2981 ( .A(n3187), .B(n3188), .Z(n3184) );
  AND U2982 ( .A(n672), .B(n3189), .Z(n3188) );
  XOR U2983 ( .A(n3190), .B(n3191), .Z(n3182) );
  AND U2984 ( .A(n676), .B(n3189), .Z(n3191) );
  XNOR U2985 ( .A(n3190), .B(n3187), .Z(n3189) );
  XOR U2986 ( .A(n3192), .B(n3193), .Z(n3187) );
  AND U2987 ( .A(n679), .B(n3194), .Z(n3193) );
  XOR U2988 ( .A(p_input[1796]), .B(n3192), .Z(n3194) );
  XOR U2989 ( .A(n3195), .B(n3196), .Z(n3192) );
  AND U2990 ( .A(n683), .B(n3197), .Z(n3196) );
  XOR U2991 ( .A(n3198), .B(n3199), .Z(n3190) );
  AND U2992 ( .A(n687), .B(n3197), .Z(n3199) );
  XNOR U2993 ( .A(n3198), .B(n3195), .Z(n3197) );
  XOR U2994 ( .A(n3200), .B(n3201), .Z(n3195) );
  AND U2995 ( .A(n690), .B(n3202), .Z(n3201) );
  XOR U2996 ( .A(p_input[1828]), .B(n3200), .Z(n3202) );
  XOR U2997 ( .A(n3203), .B(n3204), .Z(n3200) );
  AND U2998 ( .A(n694), .B(n3205), .Z(n3204) );
  XOR U2999 ( .A(n3206), .B(n3207), .Z(n3198) );
  AND U3000 ( .A(n698), .B(n3205), .Z(n3207) );
  XNOR U3001 ( .A(n3206), .B(n3203), .Z(n3205) );
  XOR U3002 ( .A(n3208), .B(n3209), .Z(n3203) );
  AND U3003 ( .A(n701), .B(n3210), .Z(n3209) );
  XOR U3004 ( .A(p_input[1860]), .B(n3208), .Z(n3210) );
  XOR U3005 ( .A(n3211), .B(n3212), .Z(n3208) );
  AND U3006 ( .A(n705), .B(n3213), .Z(n3212) );
  XOR U3007 ( .A(n3214), .B(n3215), .Z(n3206) );
  AND U3008 ( .A(n709), .B(n3213), .Z(n3215) );
  XNOR U3009 ( .A(n3214), .B(n3211), .Z(n3213) );
  XOR U3010 ( .A(n3216), .B(n3217), .Z(n3211) );
  AND U3011 ( .A(n712), .B(n3218), .Z(n3217) );
  XOR U3012 ( .A(p_input[1892]), .B(n3216), .Z(n3218) );
  XOR U3013 ( .A(n3219), .B(n3220), .Z(n3216) );
  AND U3014 ( .A(n716), .B(n3221), .Z(n3220) );
  XOR U3015 ( .A(n3222), .B(n3223), .Z(n3214) );
  AND U3016 ( .A(n720), .B(n3221), .Z(n3223) );
  XNOR U3017 ( .A(n3222), .B(n3219), .Z(n3221) );
  XOR U3018 ( .A(n3224), .B(n3225), .Z(n3219) );
  AND U3019 ( .A(n723), .B(n3226), .Z(n3225) );
  XOR U3020 ( .A(p_input[1924]), .B(n3224), .Z(n3226) );
  XOR U3021 ( .A(n3227), .B(n3228), .Z(n3224) );
  AND U3022 ( .A(n727), .B(n3229), .Z(n3228) );
  XOR U3023 ( .A(n3230), .B(n3231), .Z(n3222) );
  AND U3024 ( .A(n731), .B(n3229), .Z(n3231) );
  XNOR U3025 ( .A(n3230), .B(n3227), .Z(n3229) );
  XOR U3026 ( .A(n3232), .B(n3233), .Z(n3227) );
  AND U3027 ( .A(n734), .B(n3234), .Z(n3233) );
  XOR U3028 ( .A(p_input[1956]), .B(n3232), .Z(n3234) );
  XNOR U3029 ( .A(n3235), .B(n3236), .Z(n3232) );
  AND U3030 ( .A(n738), .B(n3237), .Z(n3236) );
  XNOR U3031 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n3238), .Z(n3230) );
  AND U3032 ( .A(n741), .B(n3237), .Z(n3238) );
  XOR U3033 ( .A(n3239), .B(n3235), .Z(n3237) );
  XOR U3034 ( .A(n1242), .B(n3240), .Z(o[35]) );
  AND U3035 ( .A(n58), .B(n3241), .Z(n1242) );
  XOR U3036 ( .A(n1243), .B(n3240), .Z(n3241) );
  XOR U3037 ( .A(n3242), .B(n3243), .Z(n3240) );
  AND U3038 ( .A(n62), .B(n3244), .Z(n3243) );
  XOR U3039 ( .A(p_input[3]), .B(n3242), .Z(n3244) );
  XOR U3040 ( .A(n3245), .B(n3246), .Z(n3242) );
  AND U3041 ( .A(n66), .B(n3247), .Z(n3246) );
  XOR U3042 ( .A(n3248), .B(n3249), .Z(n1243) );
  AND U3043 ( .A(n70), .B(n3247), .Z(n3249) );
  XNOR U3044 ( .A(n3250), .B(n3245), .Z(n3247) );
  XOR U3045 ( .A(n3251), .B(n3252), .Z(n3245) );
  AND U3046 ( .A(n74), .B(n3253), .Z(n3252) );
  XOR U3047 ( .A(p_input[35]), .B(n3251), .Z(n3253) );
  XOR U3048 ( .A(n3254), .B(n3255), .Z(n3251) );
  AND U3049 ( .A(n78), .B(n3256), .Z(n3255) );
  IV U3050 ( .A(n3248), .Z(n3250) );
  XNOR U3051 ( .A(n3257), .B(n3258), .Z(n3248) );
  AND U3052 ( .A(n82), .B(n3256), .Z(n3258) );
  XNOR U3053 ( .A(n3257), .B(n3254), .Z(n3256) );
  XOR U3054 ( .A(n3259), .B(n3260), .Z(n3254) );
  AND U3055 ( .A(n85), .B(n3261), .Z(n3260) );
  XOR U3056 ( .A(p_input[67]), .B(n3259), .Z(n3261) );
  XOR U3057 ( .A(n3262), .B(n3263), .Z(n3259) );
  AND U3058 ( .A(n89), .B(n3264), .Z(n3263) );
  XOR U3059 ( .A(n3265), .B(n3266), .Z(n3257) );
  AND U3060 ( .A(n93), .B(n3264), .Z(n3266) );
  XNOR U3061 ( .A(n3265), .B(n3262), .Z(n3264) );
  XOR U3062 ( .A(n3267), .B(n3268), .Z(n3262) );
  AND U3063 ( .A(n96), .B(n3269), .Z(n3268) );
  XOR U3064 ( .A(p_input[99]), .B(n3267), .Z(n3269) );
  XOR U3065 ( .A(n3270), .B(n3271), .Z(n3267) );
  AND U3066 ( .A(n100), .B(n3272), .Z(n3271) );
  XOR U3067 ( .A(n3273), .B(n3274), .Z(n3265) );
  AND U3068 ( .A(n104), .B(n3272), .Z(n3274) );
  XNOR U3069 ( .A(n3273), .B(n3270), .Z(n3272) );
  XOR U3070 ( .A(n3275), .B(n3276), .Z(n3270) );
  AND U3071 ( .A(n107), .B(n3277), .Z(n3276) );
  XOR U3072 ( .A(p_input[131]), .B(n3275), .Z(n3277) );
  XOR U3073 ( .A(n3278), .B(n3279), .Z(n3275) );
  AND U3074 ( .A(n111), .B(n3280), .Z(n3279) );
  XOR U3075 ( .A(n3281), .B(n3282), .Z(n3273) );
  AND U3076 ( .A(n115), .B(n3280), .Z(n3282) );
  XNOR U3077 ( .A(n3281), .B(n3278), .Z(n3280) );
  XOR U3078 ( .A(n3283), .B(n3284), .Z(n3278) );
  AND U3079 ( .A(n118), .B(n3285), .Z(n3284) );
  XOR U3080 ( .A(p_input[163]), .B(n3283), .Z(n3285) );
  XOR U3081 ( .A(n3286), .B(n3287), .Z(n3283) );
  AND U3082 ( .A(n122), .B(n3288), .Z(n3287) );
  XOR U3083 ( .A(n3289), .B(n3290), .Z(n3281) );
  AND U3084 ( .A(n126), .B(n3288), .Z(n3290) );
  XNOR U3085 ( .A(n3289), .B(n3286), .Z(n3288) );
  XOR U3086 ( .A(n3291), .B(n3292), .Z(n3286) );
  AND U3087 ( .A(n129), .B(n3293), .Z(n3292) );
  XOR U3088 ( .A(p_input[195]), .B(n3291), .Z(n3293) );
  XOR U3089 ( .A(n3294), .B(n3295), .Z(n3291) );
  AND U3090 ( .A(n133), .B(n3296), .Z(n3295) );
  XOR U3091 ( .A(n3297), .B(n3298), .Z(n3289) );
  AND U3092 ( .A(n137), .B(n3296), .Z(n3298) );
  XNOR U3093 ( .A(n3297), .B(n3294), .Z(n3296) );
  XOR U3094 ( .A(n3299), .B(n3300), .Z(n3294) );
  AND U3095 ( .A(n140), .B(n3301), .Z(n3300) );
  XOR U3096 ( .A(p_input[227]), .B(n3299), .Z(n3301) );
  XOR U3097 ( .A(n3302), .B(n3303), .Z(n3299) );
  AND U3098 ( .A(n144), .B(n3304), .Z(n3303) );
  XOR U3099 ( .A(n3305), .B(n3306), .Z(n3297) );
  AND U3100 ( .A(n148), .B(n3304), .Z(n3306) );
  XNOR U3101 ( .A(n3305), .B(n3302), .Z(n3304) );
  XOR U3102 ( .A(n3307), .B(n3308), .Z(n3302) );
  AND U3103 ( .A(n151), .B(n3309), .Z(n3308) );
  XOR U3104 ( .A(p_input[259]), .B(n3307), .Z(n3309) );
  XOR U3105 ( .A(n3310), .B(n3311), .Z(n3307) );
  AND U3106 ( .A(n155), .B(n3312), .Z(n3311) );
  XOR U3107 ( .A(n3313), .B(n3314), .Z(n3305) );
  AND U3108 ( .A(n159), .B(n3312), .Z(n3314) );
  XNOR U3109 ( .A(n3313), .B(n3310), .Z(n3312) );
  XOR U3110 ( .A(n3315), .B(n3316), .Z(n3310) );
  AND U3111 ( .A(n162), .B(n3317), .Z(n3316) );
  XOR U3112 ( .A(p_input[291]), .B(n3315), .Z(n3317) );
  XOR U3113 ( .A(n3318), .B(n3319), .Z(n3315) );
  AND U3114 ( .A(n166), .B(n3320), .Z(n3319) );
  XOR U3115 ( .A(n3321), .B(n3322), .Z(n3313) );
  AND U3116 ( .A(n170), .B(n3320), .Z(n3322) );
  XNOR U3117 ( .A(n3321), .B(n3318), .Z(n3320) );
  XOR U3118 ( .A(n3323), .B(n3324), .Z(n3318) );
  AND U3119 ( .A(n173), .B(n3325), .Z(n3324) );
  XOR U3120 ( .A(p_input[323]), .B(n3323), .Z(n3325) );
  XOR U3121 ( .A(n3326), .B(n3327), .Z(n3323) );
  AND U3122 ( .A(n177), .B(n3328), .Z(n3327) );
  XOR U3123 ( .A(n3329), .B(n3330), .Z(n3321) );
  AND U3124 ( .A(n181), .B(n3328), .Z(n3330) );
  XNOR U3125 ( .A(n3329), .B(n3326), .Z(n3328) );
  XOR U3126 ( .A(n3331), .B(n3332), .Z(n3326) );
  AND U3127 ( .A(n184), .B(n3333), .Z(n3332) );
  XOR U3128 ( .A(p_input[355]), .B(n3331), .Z(n3333) );
  XOR U3129 ( .A(n3334), .B(n3335), .Z(n3331) );
  AND U3130 ( .A(n188), .B(n3336), .Z(n3335) );
  XOR U3131 ( .A(n3337), .B(n3338), .Z(n3329) );
  AND U3132 ( .A(n192), .B(n3336), .Z(n3338) );
  XNOR U3133 ( .A(n3337), .B(n3334), .Z(n3336) );
  XOR U3134 ( .A(n3339), .B(n3340), .Z(n3334) );
  AND U3135 ( .A(n195), .B(n3341), .Z(n3340) );
  XOR U3136 ( .A(p_input[387]), .B(n3339), .Z(n3341) );
  XOR U3137 ( .A(n3342), .B(n3343), .Z(n3339) );
  AND U3138 ( .A(n199), .B(n3344), .Z(n3343) );
  XOR U3139 ( .A(n3345), .B(n3346), .Z(n3337) );
  AND U3140 ( .A(n203), .B(n3344), .Z(n3346) );
  XNOR U3141 ( .A(n3345), .B(n3342), .Z(n3344) );
  XOR U3142 ( .A(n3347), .B(n3348), .Z(n3342) );
  AND U3143 ( .A(n206), .B(n3349), .Z(n3348) );
  XOR U3144 ( .A(p_input[419]), .B(n3347), .Z(n3349) );
  XOR U3145 ( .A(n3350), .B(n3351), .Z(n3347) );
  AND U3146 ( .A(n210), .B(n3352), .Z(n3351) );
  XOR U3147 ( .A(n3353), .B(n3354), .Z(n3345) );
  AND U3148 ( .A(n214), .B(n3352), .Z(n3354) );
  XNOR U3149 ( .A(n3353), .B(n3350), .Z(n3352) );
  XOR U3150 ( .A(n3355), .B(n3356), .Z(n3350) );
  AND U3151 ( .A(n217), .B(n3357), .Z(n3356) );
  XOR U3152 ( .A(p_input[451]), .B(n3355), .Z(n3357) );
  XOR U3153 ( .A(n3358), .B(n3359), .Z(n3355) );
  AND U3154 ( .A(n221), .B(n3360), .Z(n3359) );
  XOR U3155 ( .A(n3361), .B(n3362), .Z(n3353) );
  AND U3156 ( .A(n225), .B(n3360), .Z(n3362) );
  XNOR U3157 ( .A(n3361), .B(n3358), .Z(n3360) );
  XOR U3158 ( .A(n3363), .B(n3364), .Z(n3358) );
  AND U3159 ( .A(n228), .B(n3365), .Z(n3364) );
  XOR U3160 ( .A(p_input[483]), .B(n3363), .Z(n3365) );
  XOR U3161 ( .A(n3366), .B(n3367), .Z(n3363) );
  AND U3162 ( .A(n232), .B(n3368), .Z(n3367) );
  XOR U3163 ( .A(n3369), .B(n3370), .Z(n3361) );
  AND U3164 ( .A(n236), .B(n3368), .Z(n3370) );
  XNOR U3165 ( .A(n3369), .B(n3366), .Z(n3368) );
  XOR U3166 ( .A(n3371), .B(n3372), .Z(n3366) );
  AND U3167 ( .A(n239), .B(n3373), .Z(n3372) );
  XOR U3168 ( .A(p_input[515]), .B(n3371), .Z(n3373) );
  XOR U3169 ( .A(n3374), .B(n3375), .Z(n3371) );
  AND U3170 ( .A(n243), .B(n3376), .Z(n3375) );
  XOR U3171 ( .A(n3377), .B(n3378), .Z(n3369) );
  AND U3172 ( .A(n247), .B(n3376), .Z(n3378) );
  XNOR U3173 ( .A(n3377), .B(n3374), .Z(n3376) );
  XOR U3174 ( .A(n3379), .B(n3380), .Z(n3374) );
  AND U3175 ( .A(n250), .B(n3381), .Z(n3380) );
  XOR U3176 ( .A(p_input[547]), .B(n3379), .Z(n3381) );
  XOR U3177 ( .A(n3382), .B(n3383), .Z(n3379) );
  AND U3178 ( .A(n254), .B(n3384), .Z(n3383) );
  XOR U3179 ( .A(n3385), .B(n3386), .Z(n3377) );
  AND U3180 ( .A(n258), .B(n3384), .Z(n3386) );
  XNOR U3181 ( .A(n3385), .B(n3382), .Z(n3384) );
  XOR U3182 ( .A(n3387), .B(n3388), .Z(n3382) );
  AND U3183 ( .A(n261), .B(n3389), .Z(n3388) );
  XOR U3184 ( .A(p_input[579]), .B(n3387), .Z(n3389) );
  XOR U3185 ( .A(n3390), .B(n3391), .Z(n3387) );
  AND U3186 ( .A(n265), .B(n3392), .Z(n3391) );
  XOR U3187 ( .A(n3393), .B(n3394), .Z(n3385) );
  AND U3188 ( .A(n269), .B(n3392), .Z(n3394) );
  XNOR U3189 ( .A(n3393), .B(n3390), .Z(n3392) );
  XOR U3190 ( .A(n3395), .B(n3396), .Z(n3390) );
  AND U3191 ( .A(n272), .B(n3397), .Z(n3396) );
  XOR U3192 ( .A(p_input[611]), .B(n3395), .Z(n3397) );
  XOR U3193 ( .A(n3398), .B(n3399), .Z(n3395) );
  AND U3194 ( .A(n276), .B(n3400), .Z(n3399) );
  XOR U3195 ( .A(n3401), .B(n3402), .Z(n3393) );
  AND U3196 ( .A(n280), .B(n3400), .Z(n3402) );
  XNOR U3197 ( .A(n3401), .B(n3398), .Z(n3400) );
  XOR U3198 ( .A(n3403), .B(n3404), .Z(n3398) );
  AND U3199 ( .A(n283), .B(n3405), .Z(n3404) );
  XOR U3200 ( .A(p_input[643]), .B(n3403), .Z(n3405) );
  XOR U3201 ( .A(n3406), .B(n3407), .Z(n3403) );
  AND U3202 ( .A(n287), .B(n3408), .Z(n3407) );
  XOR U3203 ( .A(n3409), .B(n3410), .Z(n3401) );
  AND U3204 ( .A(n291), .B(n3408), .Z(n3410) );
  XNOR U3205 ( .A(n3409), .B(n3406), .Z(n3408) );
  XOR U3206 ( .A(n3411), .B(n3412), .Z(n3406) );
  AND U3207 ( .A(n294), .B(n3413), .Z(n3412) );
  XOR U3208 ( .A(p_input[675]), .B(n3411), .Z(n3413) );
  XOR U3209 ( .A(n3414), .B(n3415), .Z(n3411) );
  AND U3210 ( .A(n298), .B(n3416), .Z(n3415) );
  XOR U3211 ( .A(n3417), .B(n3418), .Z(n3409) );
  AND U3212 ( .A(n302), .B(n3416), .Z(n3418) );
  XNOR U3213 ( .A(n3417), .B(n3414), .Z(n3416) );
  XOR U3214 ( .A(n3419), .B(n3420), .Z(n3414) );
  AND U3215 ( .A(n305), .B(n3421), .Z(n3420) );
  XOR U3216 ( .A(p_input[707]), .B(n3419), .Z(n3421) );
  XOR U3217 ( .A(n3422), .B(n3423), .Z(n3419) );
  AND U3218 ( .A(n309), .B(n3424), .Z(n3423) );
  XOR U3219 ( .A(n3425), .B(n3426), .Z(n3417) );
  AND U3220 ( .A(n313), .B(n3424), .Z(n3426) );
  XNOR U3221 ( .A(n3425), .B(n3422), .Z(n3424) );
  XOR U3222 ( .A(n3427), .B(n3428), .Z(n3422) );
  AND U3223 ( .A(n316), .B(n3429), .Z(n3428) );
  XOR U3224 ( .A(p_input[739]), .B(n3427), .Z(n3429) );
  XOR U3225 ( .A(n3430), .B(n3431), .Z(n3427) );
  AND U3226 ( .A(n320), .B(n3432), .Z(n3431) );
  XOR U3227 ( .A(n3433), .B(n3434), .Z(n3425) );
  AND U3228 ( .A(n324), .B(n3432), .Z(n3434) );
  XNOR U3229 ( .A(n3433), .B(n3430), .Z(n3432) );
  XOR U3230 ( .A(n3435), .B(n3436), .Z(n3430) );
  AND U3231 ( .A(n327), .B(n3437), .Z(n3436) );
  XOR U3232 ( .A(p_input[771]), .B(n3435), .Z(n3437) );
  XOR U3233 ( .A(n3438), .B(n3439), .Z(n3435) );
  AND U3234 ( .A(n331), .B(n3440), .Z(n3439) );
  XOR U3235 ( .A(n3441), .B(n3442), .Z(n3433) );
  AND U3236 ( .A(n335), .B(n3440), .Z(n3442) );
  XNOR U3237 ( .A(n3441), .B(n3438), .Z(n3440) );
  XOR U3238 ( .A(n3443), .B(n3444), .Z(n3438) );
  AND U3239 ( .A(n338), .B(n3445), .Z(n3444) );
  XOR U3240 ( .A(p_input[803]), .B(n3443), .Z(n3445) );
  XOR U3241 ( .A(n3446), .B(n3447), .Z(n3443) );
  AND U3242 ( .A(n342), .B(n3448), .Z(n3447) );
  XOR U3243 ( .A(n3449), .B(n3450), .Z(n3441) );
  AND U3244 ( .A(n346), .B(n3448), .Z(n3450) );
  XNOR U3245 ( .A(n3449), .B(n3446), .Z(n3448) );
  XOR U3246 ( .A(n3451), .B(n3452), .Z(n3446) );
  AND U3247 ( .A(n349), .B(n3453), .Z(n3452) );
  XOR U3248 ( .A(p_input[835]), .B(n3451), .Z(n3453) );
  XOR U3249 ( .A(n3454), .B(n3455), .Z(n3451) );
  AND U3250 ( .A(n353), .B(n3456), .Z(n3455) );
  XOR U3251 ( .A(n3457), .B(n3458), .Z(n3449) );
  AND U3252 ( .A(n357), .B(n3456), .Z(n3458) );
  XNOR U3253 ( .A(n3457), .B(n3454), .Z(n3456) );
  XOR U3254 ( .A(n3459), .B(n3460), .Z(n3454) );
  AND U3255 ( .A(n360), .B(n3461), .Z(n3460) );
  XOR U3256 ( .A(p_input[867]), .B(n3459), .Z(n3461) );
  XOR U3257 ( .A(n3462), .B(n3463), .Z(n3459) );
  AND U3258 ( .A(n364), .B(n3464), .Z(n3463) );
  XOR U3259 ( .A(n3465), .B(n3466), .Z(n3457) );
  AND U3260 ( .A(n368), .B(n3464), .Z(n3466) );
  XNOR U3261 ( .A(n3465), .B(n3462), .Z(n3464) );
  XOR U3262 ( .A(n3467), .B(n3468), .Z(n3462) );
  AND U3263 ( .A(n371), .B(n3469), .Z(n3468) );
  XOR U3264 ( .A(p_input[899]), .B(n3467), .Z(n3469) );
  XOR U3265 ( .A(n3470), .B(n3471), .Z(n3467) );
  AND U3266 ( .A(n375), .B(n3472), .Z(n3471) );
  XOR U3267 ( .A(n3473), .B(n3474), .Z(n3465) );
  AND U3268 ( .A(n379), .B(n3472), .Z(n3474) );
  XNOR U3269 ( .A(n3473), .B(n3470), .Z(n3472) );
  XOR U3270 ( .A(n3475), .B(n3476), .Z(n3470) );
  AND U3271 ( .A(n382), .B(n3477), .Z(n3476) );
  XOR U3272 ( .A(p_input[931]), .B(n3475), .Z(n3477) );
  XOR U3273 ( .A(n3478), .B(n3479), .Z(n3475) );
  AND U3274 ( .A(n386), .B(n3480), .Z(n3479) );
  XOR U3275 ( .A(n3481), .B(n3482), .Z(n3473) );
  AND U3276 ( .A(n390), .B(n3480), .Z(n3482) );
  XNOR U3277 ( .A(n3481), .B(n3478), .Z(n3480) );
  XOR U3278 ( .A(n3483), .B(n3484), .Z(n3478) );
  AND U3279 ( .A(n393), .B(n3485), .Z(n3484) );
  XOR U3280 ( .A(p_input[963]), .B(n3483), .Z(n3485) );
  XOR U3281 ( .A(n3486), .B(n3487), .Z(n3483) );
  AND U3282 ( .A(n397), .B(n3488), .Z(n3487) );
  XOR U3283 ( .A(n3489), .B(n3490), .Z(n3481) );
  AND U3284 ( .A(n401), .B(n3488), .Z(n3490) );
  XNOR U3285 ( .A(n3489), .B(n3486), .Z(n3488) );
  XOR U3286 ( .A(n3491), .B(n3492), .Z(n3486) );
  AND U3287 ( .A(n404), .B(n3493), .Z(n3492) );
  XOR U3288 ( .A(p_input[995]), .B(n3491), .Z(n3493) );
  XOR U3289 ( .A(n3494), .B(n3495), .Z(n3491) );
  AND U3290 ( .A(n408), .B(n3496), .Z(n3495) );
  XOR U3291 ( .A(n3497), .B(n3498), .Z(n3489) );
  AND U3292 ( .A(n412), .B(n3496), .Z(n3498) );
  XNOR U3293 ( .A(n3497), .B(n3494), .Z(n3496) );
  XOR U3294 ( .A(n3499), .B(n3500), .Z(n3494) );
  AND U3295 ( .A(n415), .B(n3501), .Z(n3500) );
  XOR U3296 ( .A(p_input[1027]), .B(n3499), .Z(n3501) );
  XOR U3297 ( .A(n3502), .B(n3503), .Z(n3499) );
  AND U3298 ( .A(n419), .B(n3504), .Z(n3503) );
  XOR U3299 ( .A(n3505), .B(n3506), .Z(n3497) );
  AND U3300 ( .A(n423), .B(n3504), .Z(n3506) );
  XNOR U3301 ( .A(n3505), .B(n3502), .Z(n3504) );
  XOR U3302 ( .A(n3507), .B(n3508), .Z(n3502) );
  AND U3303 ( .A(n426), .B(n3509), .Z(n3508) );
  XOR U3304 ( .A(p_input[1059]), .B(n3507), .Z(n3509) );
  XOR U3305 ( .A(n3510), .B(n3511), .Z(n3507) );
  AND U3306 ( .A(n430), .B(n3512), .Z(n3511) );
  XOR U3307 ( .A(n3513), .B(n3514), .Z(n3505) );
  AND U3308 ( .A(n434), .B(n3512), .Z(n3514) );
  XNOR U3309 ( .A(n3513), .B(n3510), .Z(n3512) );
  XOR U3310 ( .A(n3515), .B(n3516), .Z(n3510) );
  AND U3311 ( .A(n437), .B(n3517), .Z(n3516) );
  XOR U3312 ( .A(p_input[1091]), .B(n3515), .Z(n3517) );
  XOR U3313 ( .A(n3518), .B(n3519), .Z(n3515) );
  AND U3314 ( .A(n441), .B(n3520), .Z(n3519) );
  XOR U3315 ( .A(n3521), .B(n3522), .Z(n3513) );
  AND U3316 ( .A(n445), .B(n3520), .Z(n3522) );
  XNOR U3317 ( .A(n3521), .B(n3518), .Z(n3520) );
  XOR U3318 ( .A(n3523), .B(n3524), .Z(n3518) );
  AND U3319 ( .A(n448), .B(n3525), .Z(n3524) );
  XOR U3320 ( .A(p_input[1123]), .B(n3523), .Z(n3525) );
  XOR U3321 ( .A(n3526), .B(n3527), .Z(n3523) );
  AND U3322 ( .A(n452), .B(n3528), .Z(n3527) );
  XOR U3323 ( .A(n3529), .B(n3530), .Z(n3521) );
  AND U3324 ( .A(n456), .B(n3528), .Z(n3530) );
  XNOR U3325 ( .A(n3529), .B(n3526), .Z(n3528) );
  XOR U3326 ( .A(n3531), .B(n3532), .Z(n3526) );
  AND U3327 ( .A(n459), .B(n3533), .Z(n3532) );
  XOR U3328 ( .A(p_input[1155]), .B(n3531), .Z(n3533) );
  XOR U3329 ( .A(n3534), .B(n3535), .Z(n3531) );
  AND U3330 ( .A(n463), .B(n3536), .Z(n3535) );
  XOR U3331 ( .A(n3537), .B(n3538), .Z(n3529) );
  AND U3332 ( .A(n467), .B(n3536), .Z(n3538) );
  XNOR U3333 ( .A(n3537), .B(n3534), .Z(n3536) );
  XOR U3334 ( .A(n3539), .B(n3540), .Z(n3534) );
  AND U3335 ( .A(n470), .B(n3541), .Z(n3540) );
  XOR U3336 ( .A(p_input[1187]), .B(n3539), .Z(n3541) );
  XOR U3337 ( .A(n3542), .B(n3543), .Z(n3539) );
  AND U3338 ( .A(n474), .B(n3544), .Z(n3543) );
  XOR U3339 ( .A(n3545), .B(n3546), .Z(n3537) );
  AND U3340 ( .A(n478), .B(n3544), .Z(n3546) );
  XNOR U3341 ( .A(n3545), .B(n3542), .Z(n3544) );
  XOR U3342 ( .A(n3547), .B(n3548), .Z(n3542) );
  AND U3343 ( .A(n481), .B(n3549), .Z(n3548) );
  XOR U3344 ( .A(p_input[1219]), .B(n3547), .Z(n3549) );
  XOR U3345 ( .A(n3550), .B(n3551), .Z(n3547) );
  AND U3346 ( .A(n485), .B(n3552), .Z(n3551) );
  XOR U3347 ( .A(n3553), .B(n3554), .Z(n3545) );
  AND U3348 ( .A(n489), .B(n3552), .Z(n3554) );
  XNOR U3349 ( .A(n3553), .B(n3550), .Z(n3552) );
  XOR U3350 ( .A(n3555), .B(n3556), .Z(n3550) );
  AND U3351 ( .A(n492), .B(n3557), .Z(n3556) );
  XOR U3352 ( .A(p_input[1251]), .B(n3555), .Z(n3557) );
  XOR U3353 ( .A(n3558), .B(n3559), .Z(n3555) );
  AND U3354 ( .A(n496), .B(n3560), .Z(n3559) );
  XOR U3355 ( .A(n3561), .B(n3562), .Z(n3553) );
  AND U3356 ( .A(n500), .B(n3560), .Z(n3562) );
  XNOR U3357 ( .A(n3561), .B(n3558), .Z(n3560) );
  XOR U3358 ( .A(n3563), .B(n3564), .Z(n3558) );
  AND U3359 ( .A(n503), .B(n3565), .Z(n3564) );
  XOR U3360 ( .A(p_input[1283]), .B(n3563), .Z(n3565) );
  XOR U3361 ( .A(n3566), .B(n3567), .Z(n3563) );
  AND U3362 ( .A(n507), .B(n3568), .Z(n3567) );
  XOR U3363 ( .A(n3569), .B(n3570), .Z(n3561) );
  AND U3364 ( .A(n511), .B(n3568), .Z(n3570) );
  XNOR U3365 ( .A(n3569), .B(n3566), .Z(n3568) );
  XOR U3366 ( .A(n3571), .B(n3572), .Z(n3566) );
  AND U3367 ( .A(n514), .B(n3573), .Z(n3572) );
  XOR U3368 ( .A(p_input[1315]), .B(n3571), .Z(n3573) );
  XOR U3369 ( .A(n3574), .B(n3575), .Z(n3571) );
  AND U3370 ( .A(n518), .B(n3576), .Z(n3575) );
  XOR U3371 ( .A(n3577), .B(n3578), .Z(n3569) );
  AND U3372 ( .A(n522), .B(n3576), .Z(n3578) );
  XNOR U3373 ( .A(n3577), .B(n3574), .Z(n3576) );
  XOR U3374 ( .A(n3579), .B(n3580), .Z(n3574) );
  AND U3375 ( .A(n525), .B(n3581), .Z(n3580) );
  XOR U3376 ( .A(p_input[1347]), .B(n3579), .Z(n3581) );
  XOR U3377 ( .A(n3582), .B(n3583), .Z(n3579) );
  AND U3378 ( .A(n529), .B(n3584), .Z(n3583) );
  XOR U3379 ( .A(n3585), .B(n3586), .Z(n3577) );
  AND U3380 ( .A(n533), .B(n3584), .Z(n3586) );
  XNOR U3381 ( .A(n3585), .B(n3582), .Z(n3584) );
  XOR U3382 ( .A(n3587), .B(n3588), .Z(n3582) );
  AND U3383 ( .A(n536), .B(n3589), .Z(n3588) );
  XOR U3384 ( .A(p_input[1379]), .B(n3587), .Z(n3589) );
  XOR U3385 ( .A(n3590), .B(n3591), .Z(n3587) );
  AND U3386 ( .A(n540), .B(n3592), .Z(n3591) );
  XOR U3387 ( .A(n3593), .B(n3594), .Z(n3585) );
  AND U3388 ( .A(n544), .B(n3592), .Z(n3594) );
  XNOR U3389 ( .A(n3593), .B(n3590), .Z(n3592) );
  XOR U3390 ( .A(n3595), .B(n3596), .Z(n3590) );
  AND U3391 ( .A(n547), .B(n3597), .Z(n3596) );
  XOR U3392 ( .A(p_input[1411]), .B(n3595), .Z(n3597) );
  XOR U3393 ( .A(n3598), .B(n3599), .Z(n3595) );
  AND U3394 ( .A(n551), .B(n3600), .Z(n3599) );
  XOR U3395 ( .A(n3601), .B(n3602), .Z(n3593) );
  AND U3396 ( .A(n555), .B(n3600), .Z(n3602) );
  XNOR U3397 ( .A(n3601), .B(n3598), .Z(n3600) );
  XOR U3398 ( .A(n3603), .B(n3604), .Z(n3598) );
  AND U3399 ( .A(n558), .B(n3605), .Z(n3604) );
  XOR U3400 ( .A(p_input[1443]), .B(n3603), .Z(n3605) );
  XOR U3401 ( .A(n3606), .B(n3607), .Z(n3603) );
  AND U3402 ( .A(n562), .B(n3608), .Z(n3607) );
  XOR U3403 ( .A(n3609), .B(n3610), .Z(n3601) );
  AND U3404 ( .A(n566), .B(n3608), .Z(n3610) );
  XNOR U3405 ( .A(n3609), .B(n3606), .Z(n3608) );
  XOR U3406 ( .A(n3611), .B(n3612), .Z(n3606) );
  AND U3407 ( .A(n569), .B(n3613), .Z(n3612) );
  XOR U3408 ( .A(p_input[1475]), .B(n3611), .Z(n3613) );
  XOR U3409 ( .A(n3614), .B(n3615), .Z(n3611) );
  AND U3410 ( .A(n573), .B(n3616), .Z(n3615) );
  XOR U3411 ( .A(n3617), .B(n3618), .Z(n3609) );
  AND U3412 ( .A(n577), .B(n3616), .Z(n3618) );
  XNOR U3413 ( .A(n3617), .B(n3614), .Z(n3616) );
  XOR U3414 ( .A(n3619), .B(n3620), .Z(n3614) );
  AND U3415 ( .A(n580), .B(n3621), .Z(n3620) );
  XOR U3416 ( .A(p_input[1507]), .B(n3619), .Z(n3621) );
  XOR U3417 ( .A(n3622), .B(n3623), .Z(n3619) );
  AND U3418 ( .A(n584), .B(n3624), .Z(n3623) );
  XOR U3419 ( .A(n3625), .B(n3626), .Z(n3617) );
  AND U3420 ( .A(n588), .B(n3624), .Z(n3626) );
  XNOR U3421 ( .A(n3625), .B(n3622), .Z(n3624) );
  XOR U3422 ( .A(n3627), .B(n3628), .Z(n3622) );
  AND U3423 ( .A(n591), .B(n3629), .Z(n3628) );
  XOR U3424 ( .A(p_input[1539]), .B(n3627), .Z(n3629) );
  XOR U3425 ( .A(n3630), .B(n3631), .Z(n3627) );
  AND U3426 ( .A(n595), .B(n3632), .Z(n3631) );
  XOR U3427 ( .A(n3633), .B(n3634), .Z(n3625) );
  AND U3428 ( .A(n599), .B(n3632), .Z(n3634) );
  XNOR U3429 ( .A(n3633), .B(n3630), .Z(n3632) );
  XOR U3430 ( .A(n3635), .B(n3636), .Z(n3630) );
  AND U3431 ( .A(n602), .B(n3637), .Z(n3636) );
  XOR U3432 ( .A(p_input[1571]), .B(n3635), .Z(n3637) );
  XOR U3433 ( .A(n3638), .B(n3639), .Z(n3635) );
  AND U3434 ( .A(n606), .B(n3640), .Z(n3639) );
  XOR U3435 ( .A(n3641), .B(n3642), .Z(n3633) );
  AND U3436 ( .A(n610), .B(n3640), .Z(n3642) );
  XNOR U3437 ( .A(n3641), .B(n3638), .Z(n3640) );
  XOR U3438 ( .A(n3643), .B(n3644), .Z(n3638) );
  AND U3439 ( .A(n613), .B(n3645), .Z(n3644) );
  XOR U3440 ( .A(p_input[1603]), .B(n3643), .Z(n3645) );
  XOR U3441 ( .A(n3646), .B(n3647), .Z(n3643) );
  AND U3442 ( .A(n617), .B(n3648), .Z(n3647) );
  XOR U3443 ( .A(n3649), .B(n3650), .Z(n3641) );
  AND U3444 ( .A(n621), .B(n3648), .Z(n3650) );
  XNOR U3445 ( .A(n3649), .B(n3646), .Z(n3648) );
  XOR U3446 ( .A(n3651), .B(n3652), .Z(n3646) );
  AND U3447 ( .A(n624), .B(n3653), .Z(n3652) );
  XOR U3448 ( .A(p_input[1635]), .B(n3651), .Z(n3653) );
  XOR U3449 ( .A(n3654), .B(n3655), .Z(n3651) );
  AND U3450 ( .A(n628), .B(n3656), .Z(n3655) );
  XOR U3451 ( .A(n3657), .B(n3658), .Z(n3649) );
  AND U3452 ( .A(n632), .B(n3656), .Z(n3658) );
  XNOR U3453 ( .A(n3657), .B(n3654), .Z(n3656) );
  XOR U3454 ( .A(n3659), .B(n3660), .Z(n3654) );
  AND U3455 ( .A(n635), .B(n3661), .Z(n3660) );
  XOR U3456 ( .A(p_input[1667]), .B(n3659), .Z(n3661) );
  XOR U3457 ( .A(n3662), .B(n3663), .Z(n3659) );
  AND U3458 ( .A(n639), .B(n3664), .Z(n3663) );
  XOR U3459 ( .A(n3665), .B(n3666), .Z(n3657) );
  AND U3460 ( .A(n643), .B(n3664), .Z(n3666) );
  XNOR U3461 ( .A(n3665), .B(n3662), .Z(n3664) );
  XOR U3462 ( .A(n3667), .B(n3668), .Z(n3662) );
  AND U3463 ( .A(n646), .B(n3669), .Z(n3668) );
  XOR U3464 ( .A(p_input[1699]), .B(n3667), .Z(n3669) );
  XOR U3465 ( .A(n3670), .B(n3671), .Z(n3667) );
  AND U3466 ( .A(n650), .B(n3672), .Z(n3671) );
  XOR U3467 ( .A(n3673), .B(n3674), .Z(n3665) );
  AND U3468 ( .A(n654), .B(n3672), .Z(n3674) );
  XNOR U3469 ( .A(n3673), .B(n3670), .Z(n3672) );
  XOR U3470 ( .A(n3675), .B(n3676), .Z(n3670) );
  AND U3471 ( .A(n657), .B(n3677), .Z(n3676) );
  XOR U3472 ( .A(p_input[1731]), .B(n3675), .Z(n3677) );
  XOR U3473 ( .A(n3678), .B(n3679), .Z(n3675) );
  AND U3474 ( .A(n661), .B(n3680), .Z(n3679) );
  XOR U3475 ( .A(n3681), .B(n3682), .Z(n3673) );
  AND U3476 ( .A(n665), .B(n3680), .Z(n3682) );
  XNOR U3477 ( .A(n3681), .B(n3678), .Z(n3680) );
  XOR U3478 ( .A(n3683), .B(n3684), .Z(n3678) );
  AND U3479 ( .A(n668), .B(n3685), .Z(n3684) );
  XOR U3480 ( .A(p_input[1763]), .B(n3683), .Z(n3685) );
  XOR U3481 ( .A(n3686), .B(n3687), .Z(n3683) );
  AND U3482 ( .A(n672), .B(n3688), .Z(n3687) );
  XOR U3483 ( .A(n3689), .B(n3690), .Z(n3681) );
  AND U3484 ( .A(n676), .B(n3688), .Z(n3690) );
  XNOR U3485 ( .A(n3689), .B(n3686), .Z(n3688) );
  XOR U3486 ( .A(n3691), .B(n3692), .Z(n3686) );
  AND U3487 ( .A(n679), .B(n3693), .Z(n3692) );
  XOR U3488 ( .A(p_input[1795]), .B(n3691), .Z(n3693) );
  XOR U3489 ( .A(n3694), .B(n3695), .Z(n3691) );
  AND U3490 ( .A(n683), .B(n3696), .Z(n3695) );
  XOR U3491 ( .A(n3697), .B(n3698), .Z(n3689) );
  AND U3492 ( .A(n687), .B(n3696), .Z(n3698) );
  XNOR U3493 ( .A(n3697), .B(n3694), .Z(n3696) );
  XOR U3494 ( .A(n3699), .B(n3700), .Z(n3694) );
  AND U3495 ( .A(n690), .B(n3701), .Z(n3700) );
  XOR U3496 ( .A(p_input[1827]), .B(n3699), .Z(n3701) );
  XOR U3497 ( .A(n3702), .B(n3703), .Z(n3699) );
  AND U3498 ( .A(n694), .B(n3704), .Z(n3703) );
  XOR U3499 ( .A(n3705), .B(n3706), .Z(n3697) );
  AND U3500 ( .A(n698), .B(n3704), .Z(n3706) );
  XNOR U3501 ( .A(n3705), .B(n3702), .Z(n3704) );
  XOR U3502 ( .A(n3707), .B(n3708), .Z(n3702) );
  AND U3503 ( .A(n701), .B(n3709), .Z(n3708) );
  XOR U3504 ( .A(p_input[1859]), .B(n3707), .Z(n3709) );
  XOR U3505 ( .A(n3710), .B(n3711), .Z(n3707) );
  AND U3506 ( .A(n705), .B(n3712), .Z(n3711) );
  XOR U3507 ( .A(n3713), .B(n3714), .Z(n3705) );
  AND U3508 ( .A(n709), .B(n3712), .Z(n3714) );
  XNOR U3509 ( .A(n3713), .B(n3710), .Z(n3712) );
  XOR U3510 ( .A(n3715), .B(n3716), .Z(n3710) );
  AND U3511 ( .A(n712), .B(n3717), .Z(n3716) );
  XOR U3512 ( .A(p_input[1891]), .B(n3715), .Z(n3717) );
  XOR U3513 ( .A(n3718), .B(n3719), .Z(n3715) );
  AND U3514 ( .A(n716), .B(n3720), .Z(n3719) );
  XOR U3515 ( .A(n3721), .B(n3722), .Z(n3713) );
  AND U3516 ( .A(n720), .B(n3720), .Z(n3722) );
  XNOR U3517 ( .A(n3721), .B(n3718), .Z(n3720) );
  XOR U3518 ( .A(n3723), .B(n3724), .Z(n3718) );
  AND U3519 ( .A(n723), .B(n3725), .Z(n3724) );
  XOR U3520 ( .A(p_input[1923]), .B(n3723), .Z(n3725) );
  XOR U3521 ( .A(n3726), .B(n3727), .Z(n3723) );
  AND U3522 ( .A(n727), .B(n3728), .Z(n3727) );
  XOR U3523 ( .A(n3729), .B(n3730), .Z(n3721) );
  AND U3524 ( .A(n731), .B(n3728), .Z(n3730) );
  XNOR U3525 ( .A(n3729), .B(n3726), .Z(n3728) );
  XOR U3526 ( .A(n3731), .B(n3732), .Z(n3726) );
  AND U3527 ( .A(n734), .B(n3733), .Z(n3732) );
  XOR U3528 ( .A(p_input[1955]), .B(n3731), .Z(n3733) );
  XNOR U3529 ( .A(n3734), .B(n3735), .Z(n3731) );
  AND U3530 ( .A(n738), .B(n3736), .Z(n3735) );
  XNOR U3531 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n3737), .Z(n3729) );
  AND U3532 ( .A(n741), .B(n3736), .Z(n3737) );
  XOR U3533 ( .A(n3738), .B(n3734), .Z(n3736) );
  XOR U3534 ( .A(n3739), .B(n3740), .Z(o[34]) );
  XOR U3535 ( .A(n3741), .B(n3742), .Z(o[33]) );
  XOR U3536 ( .A(n3743), .B(n3744), .Z(o[32]) );
  XOR U3537 ( .A(n9), .B(n3745), .Z(o[31]) );
  AND U3538 ( .A(n58), .B(n3746), .Z(n9) );
  XOR U3539 ( .A(n10), .B(n3745), .Z(n3746) );
  XOR U3540 ( .A(n3747), .B(n3748), .Z(n3745) );
  AND U3541 ( .A(n70), .B(n3749), .Z(n3748) );
  XOR U3542 ( .A(n3750), .B(n3751), .Z(n10) );
  AND U3543 ( .A(n62), .B(n3752), .Z(n3751) );
  XOR U3544 ( .A(p_input[31]), .B(n3750), .Z(n3752) );
  XNOR U3545 ( .A(n3753), .B(n3754), .Z(n3750) );
  AND U3546 ( .A(n66), .B(n3749), .Z(n3754) );
  XNOR U3547 ( .A(n3753), .B(n3747), .Z(n3749) );
  XOR U3548 ( .A(n3755), .B(n3756), .Z(n3747) );
  AND U3549 ( .A(n82), .B(n3757), .Z(n3756) );
  XNOR U3550 ( .A(n3758), .B(n3759), .Z(n3753) );
  AND U3551 ( .A(n74), .B(n3760), .Z(n3759) );
  XOR U3552 ( .A(p_input[63]), .B(n3758), .Z(n3760) );
  XNOR U3553 ( .A(n3761), .B(n3762), .Z(n3758) );
  AND U3554 ( .A(n78), .B(n3757), .Z(n3762) );
  XNOR U3555 ( .A(n3761), .B(n3755), .Z(n3757) );
  XOR U3556 ( .A(n3763), .B(n3764), .Z(n3755) );
  AND U3557 ( .A(n93), .B(n3765), .Z(n3764) );
  XNOR U3558 ( .A(n3766), .B(n3767), .Z(n3761) );
  AND U3559 ( .A(n85), .B(n3768), .Z(n3767) );
  XOR U3560 ( .A(p_input[95]), .B(n3766), .Z(n3768) );
  XNOR U3561 ( .A(n3769), .B(n3770), .Z(n3766) );
  AND U3562 ( .A(n89), .B(n3765), .Z(n3770) );
  XNOR U3563 ( .A(n3769), .B(n3763), .Z(n3765) );
  XOR U3564 ( .A(n3771), .B(n3772), .Z(n3763) );
  AND U3565 ( .A(n104), .B(n3773), .Z(n3772) );
  XNOR U3566 ( .A(n3774), .B(n3775), .Z(n3769) );
  AND U3567 ( .A(n96), .B(n3776), .Z(n3775) );
  XOR U3568 ( .A(p_input[127]), .B(n3774), .Z(n3776) );
  XNOR U3569 ( .A(n3777), .B(n3778), .Z(n3774) );
  AND U3570 ( .A(n100), .B(n3773), .Z(n3778) );
  XNOR U3571 ( .A(n3777), .B(n3771), .Z(n3773) );
  XOR U3572 ( .A(n3779), .B(n3780), .Z(n3771) );
  AND U3573 ( .A(n115), .B(n3781), .Z(n3780) );
  XNOR U3574 ( .A(n3782), .B(n3783), .Z(n3777) );
  AND U3575 ( .A(n107), .B(n3784), .Z(n3783) );
  XOR U3576 ( .A(p_input[159]), .B(n3782), .Z(n3784) );
  XNOR U3577 ( .A(n3785), .B(n3786), .Z(n3782) );
  AND U3578 ( .A(n111), .B(n3781), .Z(n3786) );
  XNOR U3579 ( .A(n3785), .B(n3779), .Z(n3781) );
  XOR U3580 ( .A(n3787), .B(n3788), .Z(n3779) );
  AND U3581 ( .A(n126), .B(n3789), .Z(n3788) );
  XNOR U3582 ( .A(n3790), .B(n3791), .Z(n3785) );
  AND U3583 ( .A(n118), .B(n3792), .Z(n3791) );
  XOR U3584 ( .A(p_input[191]), .B(n3790), .Z(n3792) );
  XNOR U3585 ( .A(n3793), .B(n3794), .Z(n3790) );
  AND U3586 ( .A(n122), .B(n3789), .Z(n3794) );
  XNOR U3587 ( .A(n3793), .B(n3787), .Z(n3789) );
  XOR U3588 ( .A(n3795), .B(n3796), .Z(n3787) );
  AND U3589 ( .A(n137), .B(n3797), .Z(n3796) );
  XNOR U3590 ( .A(n3798), .B(n3799), .Z(n3793) );
  AND U3591 ( .A(n129), .B(n3800), .Z(n3799) );
  XOR U3592 ( .A(p_input[223]), .B(n3798), .Z(n3800) );
  XNOR U3593 ( .A(n3801), .B(n3802), .Z(n3798) );
  AND U3594 ( .A(n133), .B(n3797), .Z(n3802) );
  XNOR U3595 ( .A(n3801), .B(n3795), .Z(n3797) );
  XOR U3596 ( .A(n3803), .B(n3804), .Z(n3795) );
  AND U3597 ( .A(n148), .B(n3805), .Z(n3804) );
  XNOR U3598 ( .A(n3806), .B(n3807), .Z(n3801) );
  AND U3599 ( .A(n140), .B(n3808), .Z(n3807) );
  XOR U3600 ( .A(p_input[255]), .B(n3806), .Z(n3808) );
  XNOR U3601 ( .A(n3809), .B(n3810), .Z(n3806) );
  AND U3602 ( .A(n144), .B(n3805), .Z(n3810) );
  XNOR U3603 ( .A(n3809), .B(n3803), .Z(n3805) );
  XOR U3604 ( .A(n3811), .B(n3812), .Z(n3803) );
  AND U3605 ( .A(n159), .B(n3813), .Z(n3812) );
  XNOR U3606 ( .A(n3814), .B(n3815), .Z(n3809) );
  AND U3607 ( .A(n151), .B(n3816), .Z(n3815) );
  XOR U3608 ( .A(p_input[287]), .B(n3814), .Z(n3816) );
  XNOR U3609 ( .A(n3817), .B(n3818), .Z(n3814) );
  AND U3610 ( .A(n155), .B(n3813), .Z(n3818) );
  XNOR U3611 ( .A(n3817), .B(n3811), .Z(n3813) );
  XOR U3612 ( .A(n3819), .B(n3820), .Z(n3811) );
  AND U3613 ( .A(n170), .B(n3821), .Z(n3820) );
  XNOR U3614 ( .A(n3822), .B(n3823), .Z(n3817) );
  AND U3615 ( .A(n162), .B(n3824), .Z(n3823) );
  XOR U3616 ( .A(p_input[319]), .B(n3822), .Z(n3824) );
  XNOR U3617 ( .A(n3825), .B(n3826), .Z(n3822) );
  AND U3618 ( .A(n166), .B(n3821), .Z(n3826) );
  XNOR U3619 ( .A(n3825), .B(n3819), .Z(n3821) );
  XOR U3620 ( .A(n3827), .B(n3828), .Z(n3819) );
  AND U3621 ( .A(n181), .B(n3829), .Z(n3828) );
  XNOR U3622 ( .A(n3830), .B(n3831), .Z(n3825) );
  AND U3623 ( .A(n173), .B(n3832), .Z(n3831) );
  XOR U3624 ( .A(p_input[351]), .B(n3830), .Z(n3832) );
  XNOR U3625 ( .A(n3833), .B(n3834), .Z(n3830) );
  AND U3626 ( .A(n177), .B(n3829), .Z(n3834) );
  XNOR U3627 ( .A(n3833), .B(n3827), .Z(n3829) );
  XOR U3628 ( .A(n3835), .B(n3836), .Z(n3827) );
  AND U3629 ( .A(n192), .B(n3837), .Z(n3836) );
  XNOR U3630 ( .A(n3838), .B(n3839), .Z(n3833) );
  AND U3631 ( .A(n184), .B(n3840), .Z(n3839) );
  XOR U3632 ( .A(p_input[383]), .B(n3838), .Z(n3840) );
  XNOR U3633 ( .A(n3841), .B(n3842), .Z(n3838) );
  AND U3634 ( .A(n188), .B(n3837), .Z(n3842) );
  XNOR U3635 ( .A(n3841), .B(n3835), .Z(n3837) );
  XOR U3636 ( .A(n3843), .B(n3844), .Z(n3835) );
  AND U3637 ( .A(n203), .B(n3845), .Z(n3844) );
  XNOR U3638 ( .A(n3846), .B(n3847), .Z(n3841) );
  AND U3639 ( .A(n195), .B(n3848), .Z(n3847) );
  XOR U3640 ( .A(p_input[415]), .B(n3846), .Z(n3848) );
  XNOR U3641 ( .A(n3849), .B(n3850), .Z(n3846) );
  AND U3642 ( .A(n199), .B(n3845), .Z(n3850) );
  XNOR U3643 ( .A(n3849), .B(n3843), .Z(n3845) );
  XOR U3644 ( .A(n3851), .B(n3852), .Z(n3843) );
  AND U3645 ( .A(n214), .B(n3853), .Z(n3852) );
  XNOR U3646 ( .A(n3854), .B(n3855), .Z(n3849) );
  AND U3647 ( .A(n206), .B(n3856), .Z(n3855) );
  XOR U3648 ( .A(p_input[447]), .B(n3854), .Z(n3856) );
  XNOR U3649 ( .A(n3857), .B(n3858), .Z(n3854) );
  AND U3650 ( .A(n210), .B(n3853), .Z(n3858) );
  XNOR U3651 ( .A(n3857), .B(n3851), .Z(n3853) );
  XOR U3652 ( .A(n3859), .B(n3860), .Z(n3851) );
  AND U3653 ( .A(n225), .B(n3861), .Z(n3860) );
  XNOR U3654 ( .A(n3862), .B(n3863), .Z(n3857) );
  AND U3655 ( .A(n217), .B(n3864), .Z(n3863) );
  XOR U3656 ( .A(p_input[479]), .B(n3862), .Z(n3864) );
  XNOR U3657 ( .A(n3865), .B(n3866), .Z(n3862) );
  AND U3658 ( .A(n221), .B(n3861), .Z(n3866) );
  XNOR U3659 ( .A(n3865), .B(n3859), .Z(n3861) );
  XOR U3660 ( .A(n3867), .B(n3868), .Z(n3859) );
  AND U3661 ( .A(n236), .B(n3869), .Z(n3868) );
  XNOR U3662 ( .A(n3870), .B(n3871), .Z(n3865) );
  AND U3663 ( .A(n228), .B(n3872), .Z(n3871) );
  XOR U3664 ( .A(p_input[511]), .B(n3870), .Z(n3872) );
  XNOR U3665 ( .A(n3873), .B(n3874), .Z(n3870) );
  AND U3666 ( .A(n232), .B(n3869), .Z(n3874) );
  XNOR U3667 ( .A(n3873), .B(n3867), .Z(n3869) );
  XOR U3668 ( .A(n3875), .B(n3876), .Z(n3867) );
  AND U3669 ( .A(n247), .B(n3877), .Z(n3876) );
  XNOR U3670 ( .A(n3878), .B(n3879), .Z(n3873) );
  AND U3671 ( .A(n239), .B(n3880), .Z(n3879) );
  XOR U3672 ( .A(p_input[543]), .B(n3878), .Z(n3880) );
  XNOR U3673 ( .A(n3881), .B(n3882), .Z(n3878) );
  AND U3674 ( .A(n243), .B(n3877), .Z(n3882) );
  XNOR U3675 ( .A(n3881), .B(n3875), .Z(n3877) );
  XOR U3676 ( .A(n3883), .B(n3884), .Z(n3875) );
  AND U3677 ( .A(n258), .B(n3885), .Z(n3884) );
  XNOR U3678 ( .A(n3886), .B(n3887), .Z(n3881) );
  AND U3679 ( .A(n250), .B(n3888), .Z(n3887) );
  XOR U3680 ( .A(p_input[575]), .B(n3886), .Z(n3888) );
  XNOR U3681 ( .A(n3889), .B(n3890), .Z(n3886) );
  AND U3682 ( .A(n254), .B(n3885), .Z(n3890) );
  XNOR U3683 ( .A(n3889), .B(n3883), .Z(n3885) );
  XOR U3684 ( .A(n3891), .B(n3892), .Z(n3883) );
  AND U3685 ( .A(n269), .B(n3893), .Z(n3892) );
  XNOR U3686 ( .A(n3894), .B(n3895), .Z(n3889) );
  AND U3687 ( .A(n261), .B(n3896), .Z(n3895) );
  XOR U3688 ( .A(p_input[607]), .B(n3894), .Z(n3896) );
  XNOR U3689 ( .A(n3897), .B(n3898), .Z(n3894) );
  AND U3690 ( .A(n265), .B(n3893), .Z(n3898) );
  XNOR U3691 ( .A(n3897), .B(n3891), .Z(n3893) );
  XOR U3692 ( .A(n3899), .B(n3900), .Z(n3891) );
  AND U3693 ( .A(n280), .B(n3901), .Z(n3900) );
  XNOR U3694 ( .A(n3902), .B(n3903), .Z(n3897) );
  AND U3695 ( .A(n272), .B(n3904), .Z(n3903) );
  XOR U3696 ( .A(p_input[639]), .B(n3902), .Z(n3904) );
  XNOR U3697 ( .A(n3905), .B(n3906), .Z(n3902) );
  AND U3698 ( .A(n276), .B(n3901), .Z(n3906) );
  XNOR U3699 ( .A(n3905), .B(n3899), .Z(n3901) );
  XOR U3700 ( .A(n3907), .B(n3908), .Z(n3899) );
  AND U3701 ( .A(n291), .B(n3909), .Z(n3908) );
  XNOR U3702 ( .A(n3910), .B(n3911), .Z(n3905) );
  AND U3703 ( .A(n283), .B(n3912), .Z(n3911) );
  XOR U3704 ( .A(p_input[671]), .B(n3910), .Z(n3912) );
  XNOR U3705 ( .A(n3913), .B(n3914), .Z(n3910) );
  AND U3706 ( .A(n287), .B(n3909), .Z(n3914) );
  XNOR U3707 ( .A(n3913), .B(n3907), .Z(n3909) );
  XOR U3708 ( .A(n3915), .B(n3916), .Z(n3907) );
  AND U3709 ( .A(n302), .B(n3917), .Z(n3916) );
  XNOR U3710 ( .A(n3918), .B(n3919), .Z(n3913) );
  AND U3711 ( .A(n294), .B(n3920), .Z(n3919) );
  XOR U3712 ( .A(p_input[703]), .B(n3918), .Z(n3920) );
  XNOR U3713 ( .A(n3921), .B(n3922), .Z(n3918) );
  AND U3714 ( .A(n298), .B(n3917), .Z(n3922) );
  XNOR U3715 ( .A(n3921), .B(n3915), .Z(n3917) );
  XOR U3716 ( .A(n3923), .B(n3924), .Z(n3915) );
  AND U3717 ( .A(n313), .B(n3925), .Z(n3924) );
  XNOR U3718 ( .A(n3926), .B(n3927), .Z(n3921) );
  AND U3719 ( .A(n305), .B(n3928), .Z(n3927) );
  XOR U3720 ( .A(p_input[735]), .B(n3926), .Z(n3928) );
  XNOR U3721 ( .A(n3929), .B(n3930), .Z(n3926) );
  AND U3722 ( .A(n309), .B(n3925), .Z(n3930) );
  XNOR U3723 ( .A(n3929), .B(n3923), .Z(n3925) );
  XOR U3724 ( .A(n3931), .B(n3932), .Z(n3923) );
  AND U3725 ( .A(n324), .B(n3933), .Z(n3932) );
  XNOR U3726 ( .A(n3934), .B(n3935), .Z(n3929) );
  AND U3727 ( .A(n316), .B(n3936), .Z(n3935) );
  XOR U3728 ( .A(p_input[767]), .B(n3934), .Z(n3936) );
  XNOR U3729 ( .A(n3937), .B(n3938), .Z(n3934) );
  AND U3730 ( .A(n320), .B(n3933), .Z(n3938) );
  XNOR U3731 ( .A(n3937), .B(n3931), .Z(n3933) );
  XOR U3732 ( .A(n3939), .B(n3940), .Z(n3931) );
  AND U3733 ( .A(n335), .B(n3941), .Z(n3940) );
  XNOR U3734 ( .A(n3942), .B(n3943), .Z(n3937) );
  AND U3735 ( .A(n327), .B(n3944), .Z(n3943) );
  XOR U3736 ( .A(p_input[799]), .B(n3942), .Z(n3944) );
  XNOR U3737 ( .A(n3945), .B(n3946), .Z(n3942) );
  AND U3738 ( .A(n331), .B(n3941), .Z(n3946) );
  XNOR U3739 ( .A(n3945), .B(n3939), .Z(n3941) );
  XOR U3740 ( .A(n3947), .B(n3948), .Z(n3939) );
  AND U3741 ( .A(n346), .B(n3949), .Z(n3948) );
  XNOR U3742 ( .A(n3950), .B(n3951), .Z(n3945) );
  AND U3743 ( .A(n338), .B(n3952), .Z(n3951) );
  XOR U3744 ( .A(p_input[831]), .B(n3950), .Z(n3952) );
  XNOR U3745 ( .A(n3953), .B(n3954), .Z(n3950) );
  AND U3746 ( .A(n342), .B(n3949), .Z(n3954) );
  XNOR U3747 ( .A(n3953), .B(n3947), .Z(n3949) );
  XOR U3748 ( .A(n3955), .B(n3956), .Z(n3947) );
  AND U3749 ( .A(n357), .B(n3957), .Z(n3956) );
  XNOR U3750 ( .A(n3958), .B(n3959), .Z(n3953) );
  AND U3751 ( .A(n349), .B(n3960), .Z(n3959) );
  XOR U3752 ( .A(p_input[863]), .B(n3958), .Z(n3960) );
  XNOR U3753 ( .A(n3961), .B(n3962), .Z(n3958) );
  AND U3754 ( .A(n353), .B(n3957), .Z(n3962) );
  XNOR U3755 ( .A(n3961), .B(n3955), .Z(n3957) );
  XOR U3756 ( .A(n3963), .B(n3964), .Z(n3955) );
  AND U3757 ( .A(n368), .B(n3965), .Z(n3964) );
  XNOR U3758 ( .A(n3966), .B(n3967), .Z(n3961) );
  AND U3759 ( .A(n360), .B(n3968), .Z(n3967) );
  XOR U3760 ( .A(p_input[895]), .B(n3966), .Z(n3968) );
  XNOR U3761 ( .A(n3969), .B(n3970), .Z(n3966) );
  AND U3762 ( .A(n364), .B(n3965), .Z(n3970) );
  XNOR U3763 ( .A(n3969), .B(n3963), .Z(n3965) );
  XOR U3764 ( .A(n3971), .B(n3972), .Z(n3963) );
  AND U3765 ( .A(n379), .B(n3973), .Z(n3972) );
  XNOR U3766 ( .A(n3974), .B(n3975), .Z(n3969) );
  AND U3767 ( .A(n371), .B(n3976), .Z(n3975) );
  XOR U3768 ( .A(p_input[927]), .B(n3974), .Z(n3976) );
  XNOR U3769 ( .A(n3977), .B(n3978), .Z(n3974) );
  AND U3770 ( .A(n375), .B(n3973), .Z(n3978) );
  XNOR U3771 ( .A(n3977), .B(n3971), .Z(n3973) );
  XOR U3772 ( .A(n3979), .B(n3980), .Z(n3971) );
  AND U3773 ( .A(n390), .B(n3981), .Z(n3980) );
  XNOR U3774 ( .A(n3982), .B(n3983), .Z(n3977) );
  AND U3775 ( .A(n382), .B(n3984), .Z(n3983) );
  XOR U3776 ( .A(p_input[959]), .B(n3982), .Z(n3984) );
  XNOR U3777 ( .A(n3985), .B(n3986), .Z(n3982) );
  AND U3778 ( .A(n386), .B(n3981), .Z(n3986) );
  XNOR U3779 ( .A(n3985), .B(n3979), .Z(n3981) );
  XOR U3780 ( .A(n3987), .B(n3988), .Z(n3979) );
  AND U3781 ( .A(n401), .B(n3989), .Z(n3988) );
  XNOR U3782 ( .A(n3990), .B(n3991), .Z(n3985) );
  AND U3783 ( .A(n393), .B(n3992), .Z(n3991) );
  XOR U3784 ( .A(p_input[991]), .B(n3990), .Z(n3992) );
  XNOR U3785 ( .A(n3993), .B(n3994), .Z(n3990) );
  AND U3786 ( .A(n397), .B(n3989), .Z(n3994) );
  XNOR U3787 ( .A(n3993), .B(n3987), .Z(n3989) );
  XOR U3788 ( .A(n3995), .B(n3996), .Z(n3987) );
  AND U3789 ( .A(n412), .B(n3997), .Z(n3996) );
  XNOR U3790 ( .A(n3998), .B(n3999), .Z(n3993) );
  AND U3791 ( .A(n404), .B(n4000), .Z(n3999) );
  XOR U3792 ( .A(p_input[1023]), .B(n3998), .Z(n4000) );
  XNOR U3793 ( .A(n4001), .B(n4002), .Z(n3998) );
  AND U3794 ( .A(n408), .B(n3997), .Z(n4002) );
  XNOR U3795 ( .A(n4001), .B(n3995), .Z(n3997) );
  XOR U3796 ( .A(n4003), .B(n4004), .Z(n3995) );
  AND U3797 ( .A(n423), .B(n4005), .Z(n4004) );
  XNOR U3798 ( .A(n4006), .B(n4007), .Z(n4001) );
  AND U3799 ( .A(n415), .B(n4008), .Z(n4007) );
  XOR U3800 ( .A(p_input[1055]), .B(n4006), .Z(n4008) );
  XNOR U3801 ( .A(n4009), .B(n4010), .Z(n4006) );
  AND U3802 ( .A(n419), .B(n4005), .Z(n4010) );
  XNOR U3803 ( .A(n4009), .B(n4003), .Z(n4005) );
  XOR U3804 ( .A(n4011), .B(n4012), .Z(n4003) );
  AND U3805 ( .A(n434), .B(n4013), .Z(n4012) );
  XNOR U3806 ( .A(n4014), .B(n4015), .Z(n4009) );
  AND U3807 ( .A(n426), .B(n4016), .Z(n4015) );
  XOR U3808 ( .A(p_input[1087]), .B(n4014), .Z(n4016) );
  XNOR U3809 ( .A(n4017), .B(n4018), .Z(n4014) );
  AND U3810 ( .A(n430), .B(n4013), .Z(n4018) );
  XNOR U3811 ( .A(n4017), .B(n4011), .Z(n4013) );
  XOR U3812 ( .A(n4019), .B(n4020), .Z(n4011) );
  AND U3813 ( .A(n445), .B(n4021), .Z(n4020) );
  XNOR U3814 ( .A(n4022), .B(n4023), .Z(n4017) );
  AND U3815 ( .A(n437), .B(n4024), .Z(n4023) );
  XOR U3816 ( .A(p_input[1119]), .B(n4022), .Z(n4024) );
  XNOR U3817 ( .A(n4025), .B(n4026), .Z(n4022) );
  AND U3818 ( .A(n441), .B(n4021), .Z(n4026) );
  XNOR U3819 ( .A(n4025), .B(n4019), .Z(n4021) );
  XOR U3820 ( .A(n4027), .B(n4028), .Z(n4019) );
  AND U3821 ( .A(n456), .B(n4029), .Z(n4028) );
  XNOR U3822 ( .A(n4030), .B(n4031), .Z(n4025) );
  AND U3823 ( .A(n448), .B(n4032), .Z(n4031) );
  XOR U3824 ( .A(p_input[1151]), .B(n4030), .Z(n4032) );
  XNOR U3825 ( .A(n4033), .B(n4034), .Z(n4030) );
  AND U3826 ( .A(n452), .B(n4029), .Z(n4034) );
  XNOR U3827 ( .A(n4033), .B(n4027), .Z(n4029) );
  XOR U3828 ( .A(n4035), .B(n4036), .Z(n4027) );
  AND U3829 ( .A(n467), .B(n4037), .Z(n4036) );
  XNOR U3830 ( .A(n4038), .B(n4039), .Z(n4033) );
  AND U3831 ( .A(n459), .B(n4040), .Z(n4039) );
  XOR U3832 ( .A(p_input[1183]), .B(n4038), .Z(n4040) );
  XNOR U3833 ( .A(n4041), .B(n4042), .Z(n4038) );
  AND U3834 ( .A(n463), .B(n4037), .Z(n4042) );
  XNOR U3835 ( .A(n4041), .B(n4035), .Z(n4037) );
  XOR U3836 ( .A(n4043), .B(n4044), .Z(n4035) );
  AND U3837 ( .A(n478), .B(n4045), .Z(n4044) );
  XNOR U3838 ( .A(n4046), .B(n4047), .Z(n4041) );
  AND U3839 ( .A(n470), .B(n4048), .Z(n4047) );
  XOR U3840 ( .A(p_input[1215]), .B(n4046), .Z(n4048) );
  XNOR U3841 ( .A(n4049), .B(n4050), .Z(n4046) );
  AND U3842 ( .A(n474), .B(n4045), .Z(n4050) );
  XNOR U3843 ( .A(n4049), .B(n4043), .Z(n4045) );
  XOR U3844 ( .A(n4051), .B(n4052), .Z(n4043) );
  AND U3845 ( .A(n489), .B(n4053), .Z(n4052) );
  XNOR U3846 ( .A(n4054), .B(n4055), .Z(n4049) );
  AND U3847 ( .A(n481), .B(n4056), .Z(n4055) );
  XOR U3848 ( .A(p_input[1247]), .B(n4054), .Z(n4056) );
  XNOR U3849 ( .A(n4057), .B(n4058), .Z(n4054) );
  AND U3850 ( .A(n485), .B(n4053), .Z(n4058) );
  XNOR U3851 ( .A(n4057), .B(n4051), .Z(n4053) );
  XOR U3852 ( .A(n4059), .B(n4060), .Z(n4051) );
  AND U3853 ( .A(n500), .B(n4061), .Z(n4060) );
  XNOR U3854 ( .A(n4062), .B(n4063), .Z(n4057) );
  AND U3855 ( .A(n492), .B(n4064), .Z(n4063) );
  XOR U3856 ( .A(p_input[1279]), .B(n4062), .Z(n4064) );
  XNOR U3857 ( .A(n4065), .B(n4066), .Z(n4062) );
  AND U3858 ( .A(n496), .B(n4061), .Z(n4066) );
  XNOR U3859 ( .A(n4065), .B(n4059), .Z(n4061) );
  XOR U3860 ( .A(n4067), .B(n4068), .Z(n4059) );
  AND U3861 ( .A(n511), .B(n4069), .Z(n4068) );
  XNOR U3862 ( .A(n4070), .B(n4071), .Z(n4065) );
  AND U3863 ( .A(n503), .B(n4072), .Z(n4071) );
  XOR U3864 ( .A(p_input[1311]), .B(n4070), .Z(n4072) );
  XNOR U3865 ( .A(n4073), .B(n4074), .Z(n4070) );
  AND U3866 ( .A(n507), .B(n4069), .Z(n4074) );
  XNOR U3867 ( .A(n4073), .B(n4067), .Z(n4069) );
  XOR U3868 ( .A(n4075), .B(n4076), .Z(n4067) );
  AND U3869 ( .A(n522), .B(n4077), .Z(n4076) );
  XNOR U3870 ( .A(n4078), .B(n4079), .Z(n4073) );
  AND U3871 ( .A(n514), .B(n4080), .Z(n4079) );
  XOR U3872 ( .A(p_input[1343]), .B(n4078), .Z(n4080) );
  XNOR U3873 ( .A(n4081), .B(n4082), .Z(n4078) );
  AND U3874 ( .A(n518), .B(n4077), .Z(n4082) );
  XNOR U3875 ( .A(n4081), .B(n4075), .Z(n4077) );
  XOR U3876 ( .A(n4083), .B(n4084), .Z(n4075) );
  AND U3877 ( .A(n533), .B(n4085), .Z(n4084) );
  XNOR U3878 ( .A(n4086), .B(n4087), .Z(n4081) );
  AND U3879 ( .A(n525), .B(n4088), .Z(n4087) );
  XOR U3880 ( .A(p_input[1375]), .B(n4086), .Z(n4088) );
  XNOR U3881 ( .A(n4089), .B(n4090), .Z(n4086) );
  AND U3882 ( .A(n529), .B(n4085), .Z(n4090) );
  XNOR U3883 ( .A(n4089), .B(n4083), .Z(n4085) );
  XOR U3884 ( .A(n4091), .B(n4092), .Z(n4083) );
  AND U3885 ( .A(n544), .B(n4093), .Z(n4092) );
  XNOR U3886 ( .A(n4094), .B(n4095), .Z(n4089) );
  AND U3887 ( .A(n536), .B(n4096), .Z(n4095) );
  XOR U3888 ( .A(p_input[1407]), .B(n4094), .Z(n4096) );
  XNOR U3889 ( .A(n4097), .B(n4098), .Z(n4094) );
  AND U3890 ( .A(n540), .B(n4093), .Z(n4098) );
  XNOR U3891 ( .A(n4097), .B(n4091), .Z(n4093) );
  XOR U3892 ( .A(n4099), .B(n4100), .Z(n4091) );
  AND U3893 ( .A(n555), .B(n4101), .Z(n4100) );
  XNOR U3894 ( .A(n4102), .B(n4103), .Z(n4097) );
  AND U3895 ( .A(n547), .B(n4104), .Z(n4103) );
  XOR U3896 ( .A(p_input[1439]), .B(n4102), .Z(n4104) );
  XNOR U3897 ( .A(n4105), .B(n4106), .Z(n4102) );
  AND U3898 ( .A(n551), .B(n4101), .Z(n4106) );
  XNOR U3899 ( .A(n4105), .B(n4099), .Z(n4101) );
  XOR U3900 ( .A(n4107), .B(n4108), .Z(n4099) );
  AND U3901 ( .A(n566), .B(n4109), .Z(n4108) );
  XNOR U3902 ( .A(n4110), .B(n4111), .Z(n4105) );
  AND U3903 ( .A(n558), .B(n4112), .Z(n4111) );
  XOR U3904 ( .A(p_input[1471]), .B(n4110), .Z(n4112) );
  XNOR U3905 ( .A(n4113), .B(n4114), .Z(n4110) );
  AND U3906 ( .A(n562), .B(n4109), .Z(n4114) );
  XNOR U3907 ( .A(n4113), .B(n4107), .Z(n4109) );
  XOR U3908 ( .A(n4115), .B(n4116), .Z(n4107) );
  AND U3909 ( .A(n577), .B(n4117), .Z(n4116) );
  XNOR U3910 ( .A(n4118), .B(n4119), .Z(n4113) );
  AND U3911 ( .A(n569), .B(n4120), .Z(n4119) );
  XOR U3912 ( .A(p_input[1503]), .B(n4118), .Z(n4120) );
  XNOR U3913 ( .A(n4121), .B(n4122), .Z(n4118) );
  AND U3914 ( .A(n573), .B(n4117), .Z(n4122) );
  XNOR U3915 ( .A(n4121), .B(n4115), .Z(n4117) );
  XOR U3916 ( .A(n4123), .B(n4124), .Z(n4115) );
  AND U3917 ( .A(n588), .B(n4125), .Z(n4124) );
  XNOR U3918 ( .A(n4126), .B(n4127), .Z(n4121) );
  AND U3919 ( .A(n580), .B(n4128), .Z(n4127) );
  XOR U3920 ( .A(p_input[1535]), .B(n4126), .Z(n4128) );
  XNOR U3921 ( .A(n4129), .B(n4130), .Z(n4126) );
  AND U3922 ( .A(n584), .B(n4125), .Z(n4130) );
  XNOR U3923 ( .A(n4129), .B(n4123), .Z(n4125) );
  XOR U3924 ( .A(n4131), .B(n4132), .Z(n4123) );
  AND U3925 ( .A(n599), .B(n4133), .Z(n4132) );
  XNOR U3926 ( .A(n4134), .B(n4135), .Z(n4129) );
  AND U3927 ( .A(n591), .B(n4136), .Z(n4135) );
  XOR U3928 ( .A(p_input[1567]), .B(n4134), .Z(n4136) );
  XNOR U3929 ( .A(n4137), .B(n4138), .Z(n4134) );
  AND U3930 ( .A(n595), .B(n4133), .Z(n4138) );
  XNOR U3931 ( .A(n4137), .B(n4131), .Z(n4133) );
  XOR U3932 ( .A(n4139), .B(n4140), .Z(n4131) );
  AND U3933 ( .A(n610), .B(n4141), .Z(n4140) );
  XNOR U3934 ( .A(n4142), .B(n4143), .Z(n4137) );
  AND U3935 ( .A(n602), .B(n4144), .Z(n4143) );
  XOR U3936 ( .A(p_input[1599]), .B(n4142), .Z(n4144) );
  XNOR U3937 ( .A(n4145), .B(n4146), .Z(n4142) );
  AND U3938 ( .A(n606), .B(n4141), .Z(n4146) );
  XNOR U3939 ( .A(n4145), .B(n4139), .Z(n4141) );
  XOR U3940 ( .A(n4147), .B(n4148), .Z(n4139) );
  AND U3941 ( .A(n621), .B(n4149), .Z(n4148) );
  XNOR U3942 ( .A(n4150), .B(n4151), .Z(n4145) );
  AND U3943 ( .A(n613), .B(n4152), .Z(n4151) );
  XOR U3944 ( .A(p_input[1631]), .B(n4150), .Z(n4152) );
  XNOR U3945 ( .A(n4153), .B(n4154), .Z(n4150) );
  AND U3946 ( .A(n617), .B(n4149), .Z(n4154) );
  XNOR U3947 ( .A(n4153), .B(n4147), .Z(n4149) );
  XOR U3948 ( .A(n4155), .B(n4156), .Z(n4147) );
  AND U3949 ( .A(n632), .B(n4157), .Z(n4156) );
  XNOR U3950 ( .A(n4158), .B(n4159), .Z(n4153) );
  AND U3951 ( .A(n624), .B(n4160), .Z(n4159) );
  XOR U3952 ( .A(p_input[1663]), .B(n4158), .Z(n4160) );
  XNOR U3953 ( .A(n4161), .B(n4162), .Z(n4158) );
  AND U3954 ( .A(n628), .B(n4157), .Z(n4162) );
  XNOR U3955 ( .A(n4161), .B(n4155), .Z(n4157) );
  XOR U3956 ( .A(n4163), .B(n4164), .Z(n4155) );
  AND U3957 ( .A(n643), .B(n4165), .Z(n4164) );
  XNOR U3958 ( .A(n4166), .B(n4167), .Z(n4161) );
  AND U3959 ( .A(n635), .B(n4168), .Z(n4167) );
  XOR U3960 ( .A(p_input[1695]), .B(n4166), .Z(n4168) );
  XNOR U3961 ( .A(n4169), .B(n4170), .Z(n4166) );
  AND U3962 ( .A(n639), .B(n4165), .Z(n4170) );
  XNOR U3963 ( .A(n4169), .B(n4163), .Z(n4165) );
  XOR U3964 ( .A(n4171), .B(n4172), .Z(n4163) );
  AND U3965 ( .A(n654), .B(n4173), .Z(n4172) );
  XNOR U3966 ( .A(n4174), .B(n4175), .Z(n4169) );
  AND U3967 ( .A(n646), .B(n4176), .Z(n4175) );
  XOR U3968 ( .A(p_input[1727]), .B(n4174), .Z(n4176) );
  XNOR U3969 ( .A(n4177), .B(n4178), .Z(n4174) );
  AND U3970 ( .A(n650), .B(n4173), .Z(n4178) );
  XNOR U3971 ( .A(n4177), .B(n4171), .Z(n4173) );
  XOR U3972 ( .A(n4179), .B(n4180), .Z(n4171) );
  AND U3973 ( .A(n665), .B(n4181), .Z(n4180) );
  XNOR U3974 ( .A(n4182), .B(n4183), .Z(n4177) );
  AND U3975 ( .A(n657), .B(n4184), .Z(n4183) );
  XOR U3976 ( .A(p_input[1759]), .B(n4182), .Z(n4184) );
  XNOR U3977 ( .A(n4185), .B(n4186), .Z(n4182) );
  AND U3978 ( .A(n661), .B(n4181), .Z(n4186) );
  XNOR U3979 ( .A(n4185), .B(n4179), .Z(n4181) );
  XOR U3980 ( .A(n4187), .B(n4188), .Z(n4179) );
  AND U3981 ( .A(n676), .B(n4189), .Z(n4188) );
  XNOR U3982 ( .A(n4190), .B(n4191), .Z(n4185) );
  AND U3983 ( .A(n668), .B(n4192), .Z(n4191) );
  XOR U3984 ( .A(p_input[1791]), .B(n4190), .Z(n4192) );
  XNOR U3985 ( .A(n4193), .B(n4194), .Z(n4190) );
  AND U3986 ( .A(n672), .B(n4189), .Z(n4194) );
  XNOR U3987 ( .A(n4193), .B(n4187), .Z(n4189) );
  XOR U3988 ( .A(n4195), .B(n4196), .Z(n4187) );
  AND U3989 ( .A(n687), .B(n4197), .Z(n4196) );
  XNOR U3990 ( .A(n4198), .B(n4199), .Z(n4193) );
  AND U3991 ( .A(n679), .B(n4200), .Z(n4199) );
  XOR U3992 ( .A(p_input[1823]), .B(n4198), .Z(n4200) );
  XNOR U3993 ( .A(n4201), .B(n4202), .Z(n4198) );
  AND U3994 ( .A(n683), .B(n4197), .Z(n4202) );
  XNOR U3995 ( .A(n4201), .B(n4195), .Z(n4197) );
  XOR U3996 ( .A(n4203), .B(n4204), .Z(n4195) );
  AND U3997 ( .A(n698), .B(n4205), .Z(n4204) );
  XNOR U3998 ( .A(n4206), .B(n4207), .Z(n4201) );
  AND U3999 ( .A(n690), .B(n4208), .Z(n4207) );
  XOR U4000 ( .A(p_input[1855]), .B(n4206), .Z(n4208) );
  XNOR U4001 ( .A(n4209), .B(n4210), .Z(n4206) );
  AND U4002 ( .A(n694), .B(n4205), .Z(n4210) );
  XNOR U4003 ( .A(n4209), .B(n4203), .Z(n4205) );
  XOR U4004 ( .A(n4211), .B(n4212), .Z(n4203) );
  AND U4005 ( .A(n709), .B(n4213), .Z(n4212) );
  XNOR U4006 ( .A(n4214), .B(n4215), .Z(n4209) );
  AND U4007 ( .A(n701), .B(n4216), .Z(n4215) );
  XOR U4008 ( .A(p_input[1887]), .B(n4214), .Z(n4216) );
  XNOR U4009 ( .A(n4217), .B(n4218), .Z(n4214) );
  AND U4010 ( .A(n705), .B(n4213), .Z(n4218) );
  XNOR U4011 ( .A(n4217), .B(n4211), .Z(n4213) );
  XOR U4012 ( .A(n4219), .B(n4220), .Z(n4211) );
  AND U4013 ( .A(n720), .B(n4221), .Z(n4220) );
  XNOR U4014 ( .A(n4222), .B(n4223), .Z(n4217) );
  AND U4015 ( .A(n712), .B(n4224), .Z(n4223) );
  XOR U4016 ( .A(p_input[1919]), .B(n4222), .Z(n4224) );
  XNOR U4017 ( .A(n4225), .B(n4226), .Z(n4222) );
  AND U4018 ( .A(n716), .B(n4221), .Z(n4226) );
  XNOR U4019 ( .A(n4225), .B(n4219), .Z(n4221) );
  XOR U4020 ( .A(n4227), .B(n4228), .Z(n4219) );
  AND U4021 ( .A(n731), .B(n4229), .Z(n4228) );
  XNOR U4022 ( .A(n4230), .B(n4231), .Z(n4225) );
  AND U4023 ( .A(n723), .B(n4232), .Z(n4231) );
  XOR U4024 ( .A(p_input[1951]), .B(n4230), .Z(n4232) );
  XNOR U4025 ( .A(n4233), .B(n4234), .Z(n4230) );
  AND U4026 ( .A(n727), .B(n4229), .Z(n4234) );
  XNOR U4027 ( .A(n4233), .B(n4227), .Z(n4229) );
  XOR U4028 ( .A(\knn_comb_/min_val_out[0][31] ), .B(n4235), .Z(n4227) );
  AND U4029 ( .A(n741), .B(n4236), .Z(n4235) );
  XNOR U4030 ( .A(n4237), .B(n4238), .Z(n4233) );
  AND U4031 ( .A(n734), .B(n4239), .Z(n4238) );
  XOR U4032 ( .A(p_input[1983]), .B(n4237), .Z(n4239) );
  XNOR U4033 ( .A(n4240), .B(n4241), .Z(n4237) );
  AND U4034 ( .A(n738), .B(n4236), .Z(n4241) );
  XOR U4035 ( .A(n4242), .B(n4240), .Z(n4236) );
  IV U4036 ( .A(\knn_comb_/min_val_out[0][31] ), .Z(n4242) );
  IV U4037 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .Z(n4240) );
  XOR U4038 ( .A(n11), .B(n4243), .Z(o[30]) );
  AND U4039 ( .A(n58), .B(n4244), .Z(n11) );
  XOR U4040 ( .A(n12), .B(n4243), .Z(n4244) );
  XOR U4041 ( .A(n4245), .B(n4246), .Z(n4243) );
  AND U4042 ( .A(n70), .B(n4247), .Z(n4246) );
  XOR U4043 ( .A(n4248), .B(n4249), .Z(n12) );
  AND U4044 ( .A(n62), .B(n4250), .Z(n4249) );
  XOR U4045 ( .A(p_input[30]), .B(n4248), .Z(n4250) );
  XNOR U4046 ( .A(n4251), .B(n4252), .Z(n4248) );
  AND U4047 ( .A(n66), .B(n4247), .Z(n4252) );
  XNOR U4048 ( .A(n4251), .B(n4245), .Z(n4247) );
  XOR U4049 ( .A(n4253), .B(n4254), .Z(n4245) );
  AND U4050 ( .A(n82), .B(n4255), .Z(n4254) );
  XNOR U4051 ( .A(n4256), .B(n4257), .Z(n4251) );
  AND U4052 ( .A(n74), .B(n4258), .Z(n4257) );
  XOR U4053 ( .A(p_input[62]), .B(n4256), .Z(n4258) );
  XNOR U4054 ( .A(n4259), .B(n4260), .Z(n4256) );
  AND U4055 ( .A(n78), .B(n4255), .Z(n4260) );
  XNOR U4056 ( .A(n4259), .B(n4253), .Z(n4255) );
  XOR U4057 ( .A(n4261), .B(n4262), .Z(n4253) );
  AND U4058 ( .A(n93), .B(n4263), .Z(n4262) );
  XNOR U4059 ( .A(n4264), .B(n4265), .Z(n4259) );
  AND U4060 ( .A(n85), .B(n4266), .Z(n4265) );
  XOR U4061 ( .A(p_input[94]), .B(n4264), .Z(n4266) );
  XNOR U4062 ( .A(n4267), .B(n4268), .Z(n4264) );
  AND U4063 ( .A(n89), .B(n4263), .Z(n4268) );
  XNOR U4064 ( .A(n4267), .B(n4261), .Z(n4263) );
  XOR U4065 ( .A(n4269), .B(n4270), .Z(n4261) );
  AND U4066 ( .A(n104), .B(n4271), .Z(n4270) );
  XNOR U4067 ( .A(n4272), .B(n4273), .Z(n4267) );
  AND U4068 ( .A(n96), .B(n4274), .Z(n4273) );
  XOR U4069 ( .A(p_input[126]), .B(n4272), .Z(n4274) );
  XNOR U4070 ( .A(n4275), .B(n4276), .Z(n4272) );
  AND U4071 ( .A(n100), .B(n4271), .Z(n4276) );
  XNOR U4072 ( .A(n4275), .B(n4269), .Z(n4271) );
  XOR U4073 ( .A(n4277), .B(n4278), .Z(n4269) );
  AND U4074 ( .A(n115), .B(n4279), .Z(n4278) );
  XNOR U4075 ( .A(n4280), .B(n4281), .Z(n4275) );
  AND U4076 ( .A(n107), .B(n4282), .Z(n4281) );
  XOR U4077 ( .A(p_input[158]), .B(n4280), .Z(n4282) );
  XNOR U4078 ( .A(n4283), .B(n4284), .Z(n4280) );
  AND U4079 ( .A(n111), .B(n4279), .Z(n4284) );
  XNOR U4080 ( .A(n4283), .B(n4277), .Z(n4279) );
  XOR U4081 ( .A(n4285), .B(n4286), .Z(n4277) );
  AND U4082 ( .A(n126), .B(n4287), .Z(n4286) );
  XNOR U4083 ( .A(n4288), .B(n4289), .Z(n4283) );
  AND U4084 ( .A(n118), .B(n4290), .Z(n4289) );
  XOR U4085 ( .A(p_input[190]), .B(n4288), .Z(n4290) );
  XNOR U4086 ( .A(n4291), .B(n4292), .Z(n4288) );
  AND U4087 ( .A(n122), .B(n4287), .Z(n4292) );
  XNOR U4088 ( .A(n4291), .B(n4285), .Z(n4287) );
  XOR U4089 ( .A(n4293), .B(n4294), .Z(n4285) );
  AND U4090 ( .A(n137), .B(n4295), .Z(n4294) );
  XNOR U4091 ( .A(n4296), .B(n4297), .Z(n4291) );
  AND U4092 ( .A(n129), .B(n4298), .Z(n4297) );
  XOR U4093 ( .A(p_input[222]), .B(n4296), .Z(n4298) );
  XNOR U4094 ( .A(n4299), .B(n4300), .Z(n4296) );
  AND U4095 ( .A(n133), .B(n4295), .Z(n4300) );
  XNOR U4096 ( .A(n4299), .B(n4293), .Z(n4295) );
  XOR U4097 ( .A(n4301), .B(n4302), .Z(n4293) );
  AND U4098 ( .A(n148), .B(n4303), .Z(n4302) );
  XNOR U4099 ( .A(n4304), .B(n4305), .Z(n4299) );
  AND U4100 ( .A(n140), .B(n4306), .Z(n4305) );
  XOR U4101 ( .A(p_input[254]), .B(n4304), .Z(n4306) );
  XNOR U4102 ( .A(n4307), .B(n4308), .Z(n4304) );
  AND U4103 ( .A(n144), .B(n4303), .Z(n4308) );
  XNOR U4104 ( .A(n4307), .B(n4301), .Z(n4303) );
  XOR U4105 ( .A(n4309), .B(n4310), .Z(n4301) );
  AND U4106 ( .A(n159), .B(n4311), .Z(n4310) );
  XNOR U4107 ( .A(n4312), .B(n4313), .Z(n4307) );
  AND U4108 ( .A(n151), .B(n4314), .Z(n4313) );
  XOR U4109 ( .A(p_input[286]), .B(n4312), .Z(n4314) );
  XNOR U4110 ( .A(n4315), .B(n4316), .Z(n4312) );
  AND U4111 ( .A(n155), .B(n4311), .Z(n4316) );
  XNOR U4112 ( .A(n4315), .B(n4309), .Z(n4311) );
  XOR U4113 ( .A(n4317), .B(n4318), .Z(n4309) );
  AND U4114 ( .A(n170), .B(n4319), .Z(n4318) );
  XNOR U4115 ( .A(n4320), .B(n4321), .Z(n4315) );
  AND U4116 ( .A(n162), .B(n4322), .Z(n4321) );
  XOR U4117 ( .A(p_input[318]), .B(n4320), .Z(n4322) );
  XNOR U4118 ( .A(n4323), .B(n4324), .Z(n4320) );
  AND U4119 ( .A(n166), .B(n4319), .Z(n4324) );
  XNOR U4120 ( .A(n4323), .B(n4317), .Z(n4319) );
  XOR U4121 ( .A(n4325), .B(n4326), .Z(n4317) );
  AND U4122 ( .A(n181), .B(n4327), .Z(n4326) );
  XNOR U4123 ( .A(n4328), .B(n4329), .Z(n4323) );
  AND U4124 ( .A(n173), .B(n4330), .Z(n4329) );
  XOR U4125 ( .A(p_input[350]), .B(n4328), .Z(n4330) );
  XNOR U4126 ( .A(n4331), .B(n4332), .Z(n4328) );
  AND U4127 ( .A(n177), .B(n4327), .Z(n4332) );
  XNOR U4128 ( .A(n4331), .B(n4325), .Z(n4327) );
  XOR U4129 ( .A(n4333), .B(n4334), .Z(n4325) );
  AND U4130 ( .A(n192), .B(n4335), .Z(n4334) );
  XNOR U4131 ( .A(n4336), .B(n4337), .Z(n4331) );
  AND U4132 ( .A(n184), .B(n4338), .Z(n4337) );
  XOR U4133 ( .A(p_input[382]), .B(n4336), .Z(n4338) );
  XNOR U4134 ( .A(n4339), .B(n4340), .Z(n4336) );
  AND U4135 ( .A(n188), .B(n4335), .Z(n4340) );
  XNOR U4136 ( .A(n4339), .B(n4333), .Z(n4335) );
  XOR U4137 ( .A(n4341), .B(n4342), .Z(n4333) );
  AND U4138 ( .A(n203), .B(n4343), .Z(n4342) );
  XNOR U4139 ( .A(n4344), .B(n4345), .Z(n4339) );
  AND U4140 ( .A(n195), .B(n4346), .Z(n4345) );
  XOR U4141 ( .A(p_input[414]), .B(n4344), .Z(n4346) );
  XNOR U4142 ( .A(n4347), .B(n4348), .Z(n4344) );
  AND U4143 ( .A(n199), .B(n4343), .Z(n4348) );
  XNOR U4144 ( .A(n4347), .B(n4341), .Z(n4343) );
  XOR U4145 ( .A(n4349), .B(n4350), .Z(n4341) );
  AND U4146 ( .A(n214), .B(n4351), .Z(n4350) );
  XNOR U4147 ( .A(n4352), .B(n4353), .Z(n4347) );
  AND U4148 ( .A(n206), .B(n4354), .Z(n4353) );
  XOR U4149 ( .A(p_input[446]), .B(n4352), .Z(n4354) );
  XNOR U4150 ( .A(n4355), .B(n4356), .Z(n4352) );
  AND U4151 ( .A(n210), .B(n4351), .Z(n4356) );
  XNOR U4152 ( .A(n4355), .B(n4349), .Z(n4351) );
  XOR U4153 ( .A(n4357), .B(n4358), .Z(n4349) );
  AND U4154 ( .A(n225), .B(n4359), .Z(n4358) );
  XNOR U4155 ( .A(n4360), .B(n4361), .Z(n4355) );
  AND U4156 ( .A(n217), .B(n4362), .Z(n4361) );
  XOR U4157 ( .A(p_input[478]), .B(n4360), .Z(n4362) );
  XNOR U4158 ( .A(n4363), .B(n4364), .Z(n4360) );
  AND U4159 ( .A(n221), .B(n4359), .Z(n4364) );
  XNOR U4160 ( .A(n4363), .B(n4357), .Z(n4359) );
  XOR U4161 ( .A(n4365), .B(n4366), .Z(n4357) );
  AND U4162 ( .A(n236), .B(n4367), .Z(n4366) );
  XNOR U4163 ( .A(n4368), .B(n4369), .Z(n4363) );
  AND U4164 ( .A(n228), .B(n4370), .Z(n4369) );
  XOR U4165 ( .A(p_input[510]), .B(n4368), .Z(n4370) );
  XNOR U4166 ( .A(n4371), .B(n4372), .Z(n4368) );
  AND U4167 ( .A(n232), .B(n4367), .Z(n4372) );
  XNOR U4168 ( .A(n4371), .B(n4365), .Z(n4367) );
  XOR U4169 ( .A(n4373), .B(n4374), .Z(n4365) );
  AND U4170 ( .A(n247), .B(n4375), .Z(n4374) );
  XNOR U4171 ( .A(n4376), .B(n4377), .Z(n4371) );
  AND U4172 ( .A(n239), .B(n4378), .Z(n4377) );
  XOR U4173 ( .A(p_input[542]), .B(n4376), .Z(n4378) );
  XNOR U4174 ( .A(n4379), .B(n4380), .Z(n4376) );
  AND U4175 ( .A(n243), .B(n4375), .Z(n4380) );
  XNOR U4176 ( .A(n4379), .B(n4373), .Z(n4375) );
  XOR U4177 ( .A(n4381), .B(n4382), .Z(n4373) );
  AND U4178 ( .A(n258), .B(n4383), .Z(n4382) );
  XNOR U4179 ( .A(n4384), .B(n4385), .Z(n4379) );
  AND U4180 ( .A(n250), .B(n4386), .Z(n4385) );
  XOR U4181 ( .A(p_input[574]), .B(n4384), .Z(n4386) );
  XNOR U4182 ( .A(n4387), .B(n4388), .Z(n4384) );
  AND U4183 ( .A(n254), .B(n4383), .Z(n4388) );
  XNOR U4184 ( .A(n4387), .B(n4381), .Z(n4383) );
  XOR U4185 ( .A(n4389), .B(n4390), .Z(n4381) );
  AND U4186 ( .A(n269), .B(n4391), .Z(n4390) );
  XNOR U4187 ( .A(n4392), .B(n4393), .Z(n4387) );
  AND U4188 ( .A(n261), .B(n4394), .Z(n4393) );
  XOR U4189 ( .A(p_input[606]), .B(n4392), .Z(n4394) );
  XNOR U4190 ( .A(n4395), .B(n4396), .Z(n4392) );
  AND U4191 ( .A(n265), .B(n4391), .Z(n4396) );
  XNOR U4192 ( .A(n4395), .B(n4389), .Z(n4391) );
  XOR U4193 ( .A(n4397), .B(n4398), .Z(n4389) );
  AND U4194 ( .A(n280), .B(n4399), .Z(n4398) );
  XNOR U4195 ( .A(n4400), .B(n4401), .Z(n4395) );
  AND U4196 ( .A(n272), .B(n4402), .Z(n4401) );
  XOR U4197 ( .A(p_input[638]), .B(n4400), .Z(n4402) );
  XNOR U4198 ( .A(n4403), .B(n4404), .Z(n4400) );
  AND U4199 ( .A(n276), .B(n4399), .Z(n4404) );
  XNOR U4200 ( .A(n4403), .B(n4397), .Z(n4399) );
  XOR U4201 ( .A(n4405), .B(n4406), .Z(n4397) );
  AND U4202 ( .A(n291), .B(n4407), .Z(n4406) );
  XNOR U4203 ( .A(n4408), .B(n4409), .Z(n4403) );
  AND U4204 ( .A(n283), .B(n4410), .Z(n4409) );
  XOR U4205 ( .A(p_input[670]), .B(n4408), .Z(n4410) );
  XNOR U4206 ( .A(n4411), .B(n4412), .Z(n4408) );
  AND U4207 ( .A(n287), .B(n4407), .Z(n4412) );
  XNOR U4208 ( .A(n4411), .B(n4405), .Z(n4407) );
  XOR U4209 ( .A(n4413), .B(n4414), .Z(n4405) );
  AND U4210 ( .A(n302), .B(n4415), .Z(n4414) );
  XNOR U4211 ( .A(n4416), .B(n4417), .Z(n4411) );
  AND U4212 ( .A(n294), .B(n4418), .Z(n4417) );
  XOR U4213 ( .A(p_input[702]), .B(n4416), .Z(n4418) );
  XNOR U4214 ( .A(n4419), .B(n4420), .Z(n4416) );
  AND U4215 ( .A(n298), .B(n4415), .Z(n4420) );
  XNOR U4216 ( .A(n4419), .B(n4413), .Z(n4415) );
  XOR U4217 ( .A(n4421), .B(n4422), .Z(n4413) );
  AND U4218 ( .A(n313), .B(n4423), .Z(n4422) );
  XNOR U4219 ( .A(n4424), .B(n4425), .Z(n4419) );
  AND U4220 ( .A(n305), .B(n4426), .Z(n4425) );
  XOR U4221 ( .A(p_input[734]), .B(n4424), .Z(n4426) );
  XNOR U4222 ( .A(n4427), .B(n4428), .Z(n4424) );
  AND U4223 ( .A(n309), .B(n4423), .Z(n4428) );
  XNOR U4224 ( .A(n4427), .B(n4421), .Z(n4423) );
  XOR U4225 ( .A(n4429), .B(n4430), .Z(n4421) );
  AND U4226 ( .A(n324), .B(n4431), .Z(n4430) );
  XNOR U4227 ( .A(n4432), .B(n4433), .Z(n4427) );
  AND U4228 ( .A(n316), .B(n4434), .Z(n4433) );
  XOR U4229 ( .A(p_input[766]), .B(n4432), .Z(n4434) );
  XNOR U4230 ( .A(n4435), .B(n4436), .Z(n4432) );
  AND U4231 ( .A(n320), .B(n4431), .Z(n4436) );
  XNOR U4232 ( .A(n4435), .B(n4429), .Z(n4431) );
  XOR U4233 ( .A(n4437), .B(n4438), .Z(n4429) );
  AND U4234 ( .A(n335), .B(n4439), .Z(n4438) );
  XNOR U4235 ( .A(n4440), .B(n4441), .Z(n4435) );
  AND U4236 ( .A(n327), .B(n4442), .Z(n4441) );
  XOR U4237 ( .A(p_input[798]), .B(n4440), .Z(n4442) );
  XNOR U4238 ( .A(n4443), .B(n4444), .Z(n4440) );
  AND U4239 ( .A(n331), .B(n4439), .Z(n4444) );
  XNOR U4240 ( .A(n4443), .B(n4437), .Z(n4439) );
  XOR U4241 ( .A(n4445), .B(n4446), .Z(n4437) );
  AND U4242 ( .A(n346), .B(n4447), .Z(n4446) );
  XNOR U4243 ( .A(n4448), .B(n4449), .Z(n4443) );
  AND U4244 ( .A(n338), .B(n4450), .Z(n4449) );
  XOR U4245 ( .A(p_input[830]), .B(n4448), .Z(n4450) );
  XNOR U4246 ( .A(n4451), .B(n4452), .Z(n4448) );
  AND U4247 ( .A(n342), .B(n4447), .Z(n4452) );
  XNOR U4248 ( .A(n4451), .B(n4445), .Z(n4447) );
  XOR U4249 ( .A(n4453), .B(n4454), .Z(n4445) );
  AND U4250 ( .A(n357), .B(n4455), .Z(n4454) );
  XNOR U4251 ( .A(n4456), .B(n4457), .Z(n4451) );
  AND U4252 ( .A(n349), .B(n4458), .Z(n4457) );
  XOR U4253 ( .A(p_input[862]), .B(n4456), .Z(n4458) );
  XNOR U4254 ( .A(n4459), .B(n4460), .Z(n4456) );
  AND U4255 ( .A(n353), .B(n4455), .Z(n4460) );
  XNOR U4256 ( .A(n4459), .B(n4453), .Z(n4455) );
  XOR U4257 ( .A(n4461), .B(n4462), .Z(n4453) );
  AND U4258 ( .A(n368), .B(n4463), .Z(n4462) );
  XNOR U4259 ( .A(n4464), .B(n4465), .Z(n4459) );
  AND U4260 ( .A(n360), .B(n4466), .Z(n4465) );
  XOR U4261 ( .A(p_input[894]), .B(n4464), .Z(n4466) );
  XNOR U4262 ( .A(n4467), .B(n4468), .Z(n4464) );
  AND U4263 ( .A(n364), .B(n4463), .Z(n4468) );
  XNOR U4264 ( .A(n4467), .B(n4461), .Z(n4463) );
  XOR U4265 ( .A(n4469), .B(n4470), .Z(n4461) );
  AND U4266 ( .A(n379), .B(n4471), .Z(n4470) );
  XNOR U4267 ( .A(n4472), .B(n4473), .Z(n4467) );
  AND U4268 ( .A(n371), .B(n4474), .Z(n4473) );
  XOR U4269 ( .A(p_input[926]), .B(n4472), .Z(n4474) );
  XNOR U4270 ( .A(n4475), .B(n4476), .Z(n4472) );
  AND U4271 ( .A(n375), .B(n4471), .Z(n4476) );
  XNOR U4272 ( .A(n4475), .B(n4469), .Z(n4471) );
  XOR U4273 ( .A(n4477), .B(n4478), .Z(n4469) );
  AND U4274 ( .A(n390), .B(n4479), .Z(n4478) );
  XNOR U4275 ( .A(n4480), .B(n4481), .Z(n4475) );
  AND U4276 ( .A(n382), .B(n4482), .Z(n4481) );
  XOR U4277 ( .A(p_input[958]), .B(n4480), .Z(n4482) );
  XNOR U4278 ( .A(n4483), .B(n4484), .Z(n4480) );
  AND U4279 ( .A(n386), .B(n4479), .Z(n4484) );
  XNOR U4280 ( .A(n4483), .B(n4477), .Z(n4479) );
  XOR U4281 ( .A(n4485), .B(n4486), .Z(n4477) );
  AND U4282 ( .A(n401), .B(n4487), .Z(n4486) );
  XNOR U4283 ( .A(n4488), .B(n4489), .Z(n4483) );
  AND U4284 ( .A(n393), .B(n4490), .Z(n4489) );
  XOR U4285 ( .A(p_input[990]), .B(n4488), .Z(n4490) );
  XNOR U4286 ( .A(n4491), .B(n4492), .Z(n4488) );
  AND U4287 ( .A(n397), .B(n4487), .Z(n4492) );
  XNOR U4288 ( .A(n4491), .B(n4485), .Z(n4487) );
  XOR U4289 ( .A(n4493), .B(n4494), .Z(n4485) );
  AND U4290 ( .A(n412), .B(n4495), .Z(n4494) );
  XNOR U4291 ( .A(n4496), .B(n4497), .Z(n4491) );
  AND U4292 ( .A(n404), .B(n4498), .Z(n4497) );
  XOR U4293 ( .A(p_input[1022]), .B(n4496), .Z(n4498) );
  XNOR U4294 ( .A(n4499), .B(n4500), .Z(n4496) );
  AND U4295 ( .A(n408), .B(n4495), .Z(n4500) );
  XNOR U4296 ( .A(n4499), .B(n4493), .Z(n4495) );
  XOR U4297 ( .A(n4501), .B(n4502), .Z(n4493) );
  AND U4298 ( .A(n423), .B(n4503), .Z(n4502) );
  XNOR U4299 ( .A(n4504), .B(n4505), .Z(n4499) );
  AND U4300 ( .A(n415), .B(n4506), .Z(n4505) );
  XOR U4301 ( .A(p_input[1054]), .B(n4504), .Z(n4506) );
  XNOR U4302 ( .A(n4507), .B(n4508), .Z(n4504) );
  AND U4303 ( .A(n419), .B(n4503), .Z(n4508) );
  XNOR U4304 ( .A(n4507), .B(n4501), .Z(n4503) );
  XOR U4305 ( .A(n4509), .B(n4510), .Z(n4501) );
  AND U4306 ( .A(n434), .B(n4511), .Z(n4510) );
  XNOR U4307 ( .A(n4512), .B(n4513), .Z(n4507) );
  AND U4308 ( .A(n426), .B(n4514), .Z(n4513) );
  XOR U4309 ( .A(p_input[1086]), .B(n4512), .Z(n4514) );
  XNOR U4310 ( .A(n4515), .B(n4516), .Z(n4512) );
  AND U4311 ( .A(n430), .B(n4511), .Z(n4516) );
  XNOR U4312 ( .A(n4515), .B(n4509), .Z(n4511) );
  XOR U4313 ( .A(n4517), .B(n4518), .Z(n4509) );
  AND U4314 ( .A(n445), .B(n4519), .Z(n4518) );
  XNOR U4315 ( .A(n4520), .B(n4521), .Z(n4515) );
  AND U4316 ( .A(n437), .B(n4522), .Z(n4521) );
  XOR U4317 ( .A(p_input[1118]), .B(n4520), .Z(n4522) );
  XNOR U4318 ( .A(n4523), .B(n4524), .Z(n4520) );
  AND U4319 ( .A(n441), .B(n4519), .Z(n4524) );
  XNOR U4320 ( .A(n4523), .B(n4517), .Z(n4519) );
  XOR U4321 ( .A(n4525), .B(n4526), .Z(n4517) );
  AND U4322 ( .A(n456), .B(n4527), .Z(n4526) );
  XNOR U4323 ( .A(n4528), .B(n4529), .Z(n4523) );
  AND U4324 ( .A(n448), .B(n4530), .Z(n4529) );
  XOR U4325 ( .A(p_input[1150]), .B(n4528), .Z(n4530) );
  XNOR U4326 ( .A(n4531), .B(n4532), .Z(n4528) );
  AND U4327 ( .A(n452), .B(n4527), .Z(n4532) );
  XNOR U4328 ( .A(n4531), .B(n4525), .Z(n4527) );
  XOR U4329 ( .A(n4533), .B(n4534), .Z(n4525) );
  AND U4330 ( .A(n467), .B(n4535), .Z(n4534) );
  XNOR U4331 ( .A(n4536), .B(n4537), .Z(n4531) );
  AND U4332 ( .A(n459), .B(n4538), .Z(n4537) );
  XOR U4333 ( .A(p_input[1182]), .B(n4536), .Z(n4538) );
  XNOR U4334 ( .A(n4539), .B(n4540), .Z(n4536) );
  AND U4335 ( .A(n463), .B(n4535), .Z(n4540) );
  XNOR U4336 ( .A(n4539), .B(n4533), .Z(n4535) );
  XOR U4337 ( .A(n4541), .B(n4542), .Z(n4533) );
  AND U4338 ( .A(n478), .B(n4543), .Z(n4542) );
  XNOR U4339 ( .A(n4544), .B(n4545), .Z(n4539) );
  AND U4340 ( .A(n470), .B(n4546), .Z(n4545) );
  XOR U4341 ( .A(p_input[1214]), .B(n4544), .Z(n4546) );
  XNOR U4342 ( .A(n4547), .B(n4548), .Z(n4544) );
  AND U4343 ( .A(n474), .B(n4543), .Z(n4548) );
  XNOR U4344 ( .A(n4547), .B(n4541), .Z(n4543) );
  XOR U4345 ( .A(n4549), .B(n4550), .Z(n4541) );
  AND U4346 ( .A(n489), .B(n4551), .Z(n4550) );
  XNOR U4347 ( .A(n4552), .B(n4553), .Z(n4547) );
  AND U4348 ( .A(n481), .B(n4554), .Z(n4553) );
  XOR U4349 ( .A(p_input[1246]), .B(n4552), .Z(n4554) );
  XNOR U4350 ( .A(n4555), .B(n4556), .Z(n4552) );
  AND U4351 ( .A(n485), .B(n4551), .Z(n4556) );
  XNOR U4352 ( .A(n4555), .B(n4549), .Z(n4551) );
  XOR U4353 ( .A(n4557), .B(n4558), .Z(n4549) );
  AND U4354 ( .A(n500), .B(n4559), .Z(n4558) );
  XNOR U4355 ( .A(n4560), .B(n4561), .Z(n4555) );
  AND U4356 ( .A(n492), .B(n4562), .Z(n4561) );
  XOR U4357 ( .A(p_input[1278]), .B(n4560), .Z(n4562) );
  XNOR U4358 ( .A(n4563), .B(n4564), .Z(n4560) );
  AND U4359 ( .A(n496), .B(n4559), .Z(n4564) );
  XNOR U4360 ( .A(n4563), .B(n4557), .Z(n4559) );
  XOR U4361 ( .A(n4565), .B(n4566), .Z(n4557) );
  AND U4362 ( .A(n511), .B(n4567), .Z(n4566) );
  XNOR U4363 ( .A(n4568), .B(n4569), .Z(n4563) );
  AND U4364 ( .A(n503), .B(n4570), .Z(n4569) );
  XOR U4365 ( .A(p_input[1310]), .B(n4568), .Z(n4570) );
  XNOR U4366 ( .A(n4571), .B(n4572), .Z(n4568) );
  AND U4367 ( .A(n507), .B(n4567), .Z(n4572) );
  XNOR U4368 ( .A(n4571), .B(n4565), .Z(n4567) );
  XOR U4369 ( .A(n4573), .B(n4574), .Z(n4565) );
  AND U4370 ( .A(n522), .B(n4575), .Z(n4574) );
  XNOR U4371 ( .A(n4576), .B(n4577), .Z(n4571) );
  AND U4372 ( .A(n514), .B(n4578), .Z(n4577) );
  XOR U4373 ( .A(p_input[1342]), .B(n4576), .Z(n4578) );
  XNOR U4374 ( .A(n4579), .B(n4580), .Z(n4576) );
  AND U4375 ( .A(n518), .B(n4575), .Z(n4580) );
  XNOR U4376 ( .A(n4579), .B(n4573), .Z(n4575) );
  XOR U4377 ( .A(n4581), .B(n4582), .Z(n4573) );
  AND U4378 ( .A(n533), .B(n4583), .Z(n4582) );
  XNOR U4379 ( .A(n4584), .B(n4585), .Z(n4579) );
  AND U4380 ( .A(n525), .B(n4586), .Z(n4585) );
  XOR U4381 ( .A(p_input[1374]), .B(n4584), .Z(n4586) );
  XNOR U4382 ( .A(n4587), .B(n4588), .Z(n4584) );
  AND U4383 ( .A(n529), .B(n4583), .Z(n4588) );
  XNOR U4384 ( .A(n4587), .B(n4581), .Z(n4583) );
  XOR U4385 ( .A(n4589), .B(n4590), .Z(n4581) );
  AND U4386 ( .A(n544), .B(n4591), .Z(n4590) );
  XNOR U4387 ( .A(n4592), .B(n4593), .Z(n4587) );
  AND U4388 ( .A(n536), .B(n4594), .Z(n4593) );
  XOR U4389 ( .A(p_input[1406]), .B(n4592), .Z(n4594) );
  XNOR U4390 ( .A(n4595), .B(n4596), .Z(n4592) );
  AND U4391 ( .A(n540), .B(n4591), .Z(n4596) );
  XNOR U4392 ( .A(n4595), .B(n4589), .Z(n4591) );
  XOR U4393 ( .A(n4597), .B(n4598), .Z(n4589) );
  AND U4394 ( .A(n555), .B(n4599), .Z(n4598) );
  XNOR U4395 ( .A(n4600), .B(n4601), .Z(n4595) );
  AND U4396 ( .A(n547), .B(n4602), .Z(n4601) );
  XOR U4397 ( .A(p_input[1438]), .B(n4600), .Z(n4602) );
  XNOR U4398 ( .A(n4603), .B(n4604), .Z(n4600) );
  AND U4399 ( .A(n551), .B(n4599), .Z(n4604) );
  XNOR U4400 ( .A(n4603), .B(n4597), .Z(n4599) );
  XOR U4401 ( .A(n4605), .B(n4606), .Z(n4597) );
  AND U4402 ( .A(n566), .B(n4607), .Z(n4606) );
  XNOR U4403 ( .A(n4608), .B(n4609), .Z(n4603) );
  AND U4404 ( .A(n558), .B(n4610), .Z(n4609) );
  XOR U4405 ( .A(p_input[1470]), .B(n4608), .Z(n4610) );
  XNOR U4406 ( .A(n4611), .B(n4612), .Z(n4608) );
  AND U4407 ( .A(n562), .B(n4607), .Z(n4612) );
  XNOR U4408 ( .A(n4611), .B(n4605), .Z(n4607) );
  XOR U4409 ( .A(n4613), .B(n4614), .Z(n4605) );
  AND U4410 ( .A(n577), .B(n4615), .Z(n4614) );
  XNOR U4411 ( .A(n4616), .B(n4617), .Z(n4611) );
  AND U4412 ( .A(n569), .B(n4618), .Z(n4617) );
  XOR U4413 ( .A(p_input[1502]), .B(n4616), .Z(n4618) );
  XNOR U4414 ( .A(n4619), .B(n4620), .Z(n4616) );
  AND U4415 ( .A(n573), .B(n4615), .Z(n4620) );
  XNOR U4416 ( .A(n4619), .B(n4613), .Z(n4615) );
  XOR U4417 ( .A(n4621), .B(n4622), .Z(n4613) );
  AND U4418 ( .A(n588), .B(n4623), .Z(n4622) );
  XNOR U4419 ( .A(n4624), .B(n4625), .Z(n4619) );
  AND U4420 ( .A(n580), .B(n4626), .Z(n4625) );
  XOR U4421 ( .A(p_input[1534]), .B(n4624), .Z(n4626) );
  XNOR U4422 ( .A(n4627), .B(n4628), .Z(n4624) );
  AND U4423 ( .A(n584), .B(n4623), .Z(n4628) );
  XNOR U4424 ( .A(n4627), .B(n4621), .Z(n4623) );
  XOR U4425 ( .A(n4629), .B(n4630), .Z(n4621) );
  AND U4426 ( .A(n599), .B(n4631), .Z(n4630) );
  XNOR U4427 ( .A(n4632), .B(n4633), .Z(n4627) );
  AND U4428 ( .A(n591), .B(n4634), .Z(n4633) );
  XOR U4429 ( .A(p_input[1566]), .B(n4632), .Z(n4634) );
  XNOR U4430 ( .A(n4635), .B(n4636), .Z(n4632) );
  AND U4431 ( .A(n595), .B(n4631), .Z(n4636) );
  XNOR U4432 ( .A(n4635), .B(n4629), .Z(n4631) );
  XOR U4433 ( .A(n4637), .B(n4638), .Z(n4629) );
  AND U4434 ( .A(n610), .B(n4639), .Z(n4638) );
  XNOR U4435 ( .A(n4640), .B(n4641), .Z(n4635) );
  AND U4436 ( .A(n602), .B(n4642), .Z(n4641) );
  XOR U4437 ( .A(p_input[1598]), .B(n4640), .Z(n4642) );
  XNOR U4438 ( .A(n4643), .B(n4644), .Z(n4640) );
  AND U4439 ( .A(n606), .B(n4639), .Z(n4644) );
  XNOR U4440 ( .A(n4643), .B(n4637), .Z(n4639) );
  XOR U4441 ( .A(n4645), .B(n4646), .Z(n4637) );
  AND U4442 ( .A(n621), .B(n4647), .Z(n4646) );
  XNOR U4443 ( .A(n4648), .B(n4649), .Z(n4643) );
  AND U4444 ( .A(n613), .B(n4650), .Z(n4649) );
  XOR U4445 ( .A(p_input[1630]), .B(n4648), .Z(n4650) );
  XNOR U4446 ( .A(n4651), .B(n4652), .Z(n4648) );
  AND U4447 ( .A(n617), .B(n4647), .Z(n4652) );
  XNOR U4448 ( .A(n4651), .B(n4645), .Z(n4647) );
  XOR U4449 ( .A(n4653), .B(n4654), .Z(n4645) );
  AND U4450 ( .A(n632), .B(n4655), .Z(n4654) );
  XNOR U4451 ( .A(n4656), .B(n4657), .Z(n4651) );
  AND U4452 ( .A(n624), .B(n4658), .Z(n4657) );
  XOR U4453 ( .A(p_input[1662]), .B(n4656), .Z(n4658) );
  XNOR U4454 ( .A(n4659), .B(n4660), .Z(n4656) );
  AND U4455 ( .A(n628), .B(n4655), .Z(n4660) );
  XNOR U4456 ( .A(n4659), .B(n4653), .Z(n4655) );
  XOR U4457 ( .A(n4661), .B(n4662), .Z(n4653) );
  AND U4458 ( .A(n643), .B(n4663), .Z(n4662) );
  XNOR U4459 ( .A(n4664), .B(n4665), .Z(n4659) );
  AND U4460 ( .A(n635), .B(n4666), .Z(n4665) );
  XOR U4461 ( .A(p_input[1694]), .B(n4664), .Z(n4666) );
  XNOR U4462 ( .A(n4667), .B(n4668), .Z(n4664) );
  AND U4463 ( .A(n639), .B(n4663), .Z(n4668) );
  XNOR U4464 ( .A(n4667), .B(n4661), .Z(n4663) );
  XOR U4465 ( .A(n4669), .B(n4670), .Z(n4661) );
  AND U4466 ( .A(n654), .B(n4671), .Z(n4670) );
  XNOR U4467 ( .A(n4672), .B(n4673), .Z(n4667) );
  AND U4468 ( .A(n646), .B(n4674), .Z(n4673) );
  XOR U4469 ( .A(p_input[1726]), .B(n4672), .Z(n4674) );
  XNOR U4470 ( .A(n4675), .B(n4676), .Z(n4672) );
  AND U4471 ( .A(n650), .B(n4671), .Z(n4676) );
  XNOR U4472 ( .A(n4675), .B(n4669), .Z(n4671) );
  XOR U4473 ( .A(n4677), .B(n4678), .Z(n4669) );
  AND U4474 ( .A(n665), .B(n4679), .Z(n4678) );
  XNOR U4475 ( .A(n4680), .B(n4681), .Z(n4675) );
  AND U4476 ( .A(n657), .B(n4682), .Z(n4681) );
  XOR U4477 ( .A(p_input[1758]), .B(n4680), .Z(n4682) );
  XNOR U4478 ( .A(n4683), .B(n4684), .Z(n4680) );
  AND U4479 ( .A(n661), .B(n4679), .Z(n4684) );
  XNOR U4480 ( .A(n4683), .B(n4677), .Z(n4679) );
  XOR U4481 ( .A(n4685), .B(n4686), .Z(n4677) );
  AND U4482 ( .A(n676), .B(n4687), .Z(n4686) );
  XNOR U4483 ( .A(n4688), .B(n4689), .Z(n4683) );
  AND U4484 ( .A(n668), .B(n4690), .Z(n4689) );
  XOR U4485 ( .A(p_input[1790]), .B(n4688), .Z(n4690) );
  XNOR U4486 ( .A(n4691), .B(n4692), .Z(n4688) );
  AND U4487 ( .A(n672), .B(n4687), .Z(n4692) );
  XNOR U4488 ( .A(n4691), .B(n4685), .Z(n4687) );
  XOR U4489 ( .A(n4693), .B(n4694), .Z(n4685) );
  AND U4490 ( .A(n687), .B(n4695), .Z(n4694) );
  XNOR U4491 ( .A(n4696), .B(n4697), .Z(n4691) );
  AND U4492 ( .A(n679), .B(n4698), .Z(n4697) );
  XOR U4493 ( .A(p_input[1822]), .B(n4696), .Z(n4698) );
  XNOR U4494 ( .A(n4699), .B(n4700), .Z(n4696) );
  AND U4495 ( .A(n683), .B(n4695), .Z(n4700) );
  XNOR U4496 ( .A(n4699), .B(n4693), .Z(n4695) );
  XOR U4497 ( .A(n4701), .B(n4702), .Z(n4693) );
  AND U4498 ( .A(n698), .B(n4703), .Z(n4702) );
  XNOR U4499 ( .A(n4704), .B(n4705), .Z(n4699) );
  AND U4500 ( .A(n690), .B(n4706), .Z(n4705) );
  XOR U4501 ( .A(p_input[1854]), .B(n4704), .Z(n4706) );
  XNOR U4502 ( .A(n4707), .B(n4708), .Z(n4704) );
  AND U4503 ( .A(n694), .B(n4703), .Z(n4708) );
  XNOR U4504 ( .A(n4707), .B(n4701), .Z(n4703) );
  XOR U4505 ( .A(n4709), .B(n4710), .Z(n4701) );
  AND U4506 ( .A(n709), .B(n4711), .Z(n4710) );
  XNOR U4507 ( .A(n4712), .B(n4713), .Z(n4707) );
  AND U4508 ( .A(n701), .B(n4714), .Z(n4713) );
  XOR U4509 ( .A(p_input[1886]), .B(n4712), .Z(n4714) );
  XNOR U4510 ( .A(n4715), .B(n4716), .Z(n4712) );
  AND U4511 ( .A(n705), .B(n4711), .Z(n4716) );
  XNOR U4512 ( .A(n4715), .B(n4709), .Z(n4711) );
  XOR U4513 ( .A(n4717), .B(n4718), .Z(n4709) );
  AND U4514 ( .A(n720), .B(n4719), .Z(n4718) );
  XNOR U4515 ( .A(n4720), .B(n4721), .Z(n4715) );
  AND U4516 ( .A(n712), .B(n4722), .Z(n4721) );
  XOR U4517 ( .A(p_input[1918]), .B(n4720), .Z(n4722) );
  XNOR U4518 ( .A(n4723), .B(n4724), .Z(n4720) );
  AND U4519 ( .A(n716), .B(n4719), .Z(n4724) );
  XNOR U4520 ( .A(n4723), .B(n4717), .Z(n4719) );
  XOR U4521 ( .A(n4725), .B(n4726), .Z(n4717) );
  AND U4522 ( .A(n731), .B(n4727), .Z(n4726) );
  XNOR U4523 ( .A(n4728), .B(n4729), .Z(n4723) );
  AND U4524 ( .A(n723), .B(n4730), .Z(n4729) );
  XOR U4525 ( .A(p_input[1950]), .B(n4728), .Z(n4730) );
  XNOR U4526 ( .A(n4731), .B(n4732), .Z(n4728) );
  AND U4527 ( .A(n727), .B(n4727), .Z(n4732) );
  XNOR U4528 ( .A(n4731), .B(n4725), .Z(n4727) );
  XOR U4529 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n4733), .Z(n4725) );
  AND U4530 ( .A(n741), .B(n4734), .Z(n4733) );
  XNOR U4531 ( .A(n4735), .B(n4736), .Z(n4731) );
  AND U4532 ( .A(n734), .B(n4737), .Z(n4736) );
  XOR U4533 ( .A(p_input[1982]), .B(n4735), .Z(n4737) );
  XNOR U4534 ( .A(n4738), .B(n4739), .Z(n4735) );
  AND U4535 ( .A(n738), .B(n4734), .Z(n4739) );
  XOR U4536 ( .A(n4740), .B(n4738), .Z(n4734) );
  IV U4537 ( .A(\knn_comb_/min_val_out[0][30] ), .Z(n4740) );
  IV U4538 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .Z(n4738) );
  XOR U4539 ( .A(n3739), .B(n4741), .Z(o[2]) );
  AND U4540 ( .A(n58), .B(n4742), .Z(n3739) );
  XOR U4541 ( .A(n3740), .B(n4741), .Z(n4742) );
  XOR U4542 ( .A(n4743), .B(n4744), .Z(n4741) );
  AND U4543 ( .A(n70), .B(n4745), .Z(n4744) );
  XOR U4544 ( .A(n4746), .B(n4747), .Z(n3740) );
  AND U4545 ( .A(n62), .B(n4748), .Z(n4747) );
  XOR U4546 ( .A(p_input[2]), .B(n4746), .Z(n4748) );
  XNOR U4547 ( .A(n4749), .B(n4750), .Z(n4746) );
  AND U4548 ( .A(n66), .B(n4745), .Z(n4750) );
  XNOR U4549 ( .A(n4749), .B(n4743), .Z(n4745) );
  XOR U4550 ( .A(n4751), .B(n4752), .Z(n4743) );
  AND U4551 ( .A(n82), .B(n4753), .Z(n4752) );
  XNOR U4552 ( .A(n4754), .B(n4755), .Z(n4749) );
  AND U4553 ( .A(n74), .B(n4756), .Z(n4755) );
  XOR U4554 ( .A(p_input[34]), .B(n4754), .Z(n4756) );
  XNOR U4555 ( .A(n4757), .B(n4758), .Z(n4754) );
  AND U4556 ( .A(n78), .B(n4753), .Z(n4758) );
  XNOR U4557 ( .A(n4757), .B(n4751), .Z(n4753) );
  XOR U4558 ( .A(n4759), .B(n4760), .Z(n4751) );
  AND U4559 ( .A(n93), .B(n4761), .Z(n4760) );
  XNOR U4560 ( .A(n4762), .B(n4763), .Z(n4757) );
  AND U4561 ( .A(n85), .B(n4764), .Z(n4763) );
  XOR U4562 ( .A(p_input[66]), .B(n4762), .Z(n4764) );
  XNOR U4563 ( .A(n4765), .B(n4766), .Z(n4762) );
  AND U4564 ( .A(n89), .B(n4761), .Z(n4766) );
  XNOR U4565 ( .A(n4765), .B(n4759), .Z(n4761) );
  XOR U4566 ( .A(n4767), .B(n4768), .Z(n4759) );
  AND U4567 ( .A(n104), .B(n4769), .Z(n4768) );
  XNOR U4568 ( .A(n4770), .B(n4771), .Z(n4765) );
  AND U4569 ( .A(n96), .B(n4772), .Z(n4771) );
  XOR U4570 ( .A(p_input[98]), .B(n4770), .Z(n4772) );
  XNOR U4571 ( .A(n4773), .B(n4774), .Z(n4770) );
  AND U4572 ( .A(n100), .B(n4769), .Z(n4774) );
  XNOR U4573 ( .A(n4773), .B(n4767), .Z(n4769) );
  XOR U4574 ( .A(n4775), .B(n4776), .Z(n4767) );
  AND U4575 ( .A(n115), .B(n4777), .Z(n4776) );
  XNOR U4576 ( .A(n4778), .B(n4779), .Z(n4773) );
  AND U4577 ( .A(n107), .B(n4780), .Z(n4779) );
  XOR U4578 ( .A(p_input[130]), .B(n4778), .Z(n4780) );
  XNOR U4579 ( .A(n4781), .B(n4782), .Z(n4778) );
  AND U4580 ( .A(n111), .B(n4777), .Z(n4782) );
  XNOR U4581 ( .A(n4781), .B(n4775), .Z(n4777) );
  XOR U4582 ( .A(n4783), .B(n4784), .Z(n4775) );
  AND U4583 ( .A(n126), .B(n4785), .Z(n4784) );
  XNOR U4584 ( .A(n4786), .B(n4787), .Z(n4781) );
  AND U4585 ( .A(n118), .B(n4788), .Z(n4787) );
  XOR U4586 ( .A(p_input[162]), .B(n4786), .Z(n4788) );
  XNOR U4587 ( .A(n4789), .B(n4790), .Z(n4786) );
  AND U4588 ( .A(n122), .B(n4785), .Z(n4790) );
  XNOR U4589 ( .A(n4789), .B(n4783), .Z(n4785) );
  XOR U4590 ( .A(n4791), .B(n4792), .Z(n4783) );
  AND U4591 ( .A(n137), .B(n4793), .Z(n4792) );
  XNOR U4592 ( .A(n4794), .B(n4795), .Z(n4789) );
  AND U4593 ( .A(n129), .B(n4796), .Z(n4795) );
  XOR U4594 ( .A(p_input[194]), .B(n4794), .Z(n4796) );
  XNOR U4595 ( .A(n4797), .B(n4798), .Z(n4794) );
  AND U4596 ( .A(n133), .B(n4793), .Z(n4798) );
  XNOR U4597 ( .A(n4797), .B(n4791), .Z(n4793) );
  XOR U4598 ( .A(n4799), .B(n4800), .Z(n4791) );
  AND U4599 ( .A(n148), .B(n4801), .Z(n4800) );
  XNOR U4600 ( .A(n4802), .B(n4803), .Z(n4797) );
  AND U4601 ( .A(n140), .B(n4804), .Z(n4803) );
  XOR U4602 ( .A(p_input[226]), .B(n4802), .Z(n4804) );
  XNOR U4603 ( .A(n4805), .B(n4806), .Z(n4802) );
  AND U4604 ( .A(n144), .B(n4801), .Z(n4806) );
  XNOR U4605 ( .A(n4805), .B(n4799), .Z(n4801) );
  XOR U4606 ( .A(n4807), .B(n4808), .Z(n4799) );
  AND U4607 ( .A(n159), .B(n4809), .Z(n4808) );
  XNOR U4608 ( .A(n4810), .B(n4811), .Z(n4805) );
  AND U4609 ( .A(n151), .B(n4812), .Z(n4811) );
  XOR U4610 ( .A(p_input[258]), .B(n4810), .Z(n4812) );
  XNOR U4611 ( .A(n4813), .B(n4814), .Z(n4810) );
  AND U4612 ( .A(n155), .B(n4809), .Z(n4814) );
  XNOR U4613 ( .A(n4813), .B(n4807), .Z(n4809) );
  XOR U4614 ( .A(n4815), .B(n4816), .Z(n4807) );
  AND U4615 ( .A(n170), .B(n4817), .Z(n4816) );
  XNOR U4616 ( .A(n4818), .B(n4819), .Z(n4813) );
  AND U4617 ( .A(n162), .B(n4820), .Z(n4819) );
  XOR U4618 ( .A(p_input[290]), .B(n4818), .Z(n4820) );
  XNOR U4619 ( .A(n4821), .B(n4822), .Z(n4818) );
  AND U4620 ( .A(n166), .B(n4817), .Z(n4822) );
  XNOR U4621 ( .A(n4821), .B(n4815), .Z(n4817) );
  XOR U4622 ( .A(n4823), .B(n4824), .Z(n4815) );
  AND U4623 ( .A(n181), .B(n4825), .Z(n4824) );
  XNOR U4624 ( .A(n4826), .B(n4827), .Z(n4821) );
  AND U4625 ( .A(n173), .B(n4828), .Z(n4827) );
  XOR U4626 ( .A(p_input[322]), .B(n4826), .Z(n4828) );
  XNOR U4627 ( .A(n4829), .B(n4830), .Z(n4826) );
  AND U4628 ( .A(n177), .B(n4825), .Z(n4830) );
  XNOR U4629 ( .A(n4829), .B(n4823), .Z(n4825) );
  XOR U4630 ( .A(n4831), .B(n4832), .Z(n4823) );
  AND U4631 ( .A(n192), .B(n4833), .Z(n4832) );
  XNOR U4632 ( .A(n4834), .B(n4835), .Z(n4829) );
  AND U4633 ( .A(n184), .B(n4836), .Z(n4835) );
  XOR U4634 ( .A(p_input[354]), .B(n4834), .Z(n4836) );
  XNOR U4635 ( .A(n4837), .B(n4838), .Z(n4834) );
  AND U4636 ( .A(n188), .B(n4833), .Z(n4838) );
  XNOR U4637 ( .A(n4837), .B(n4831), .Z(n4833) );
  XOR U4638 ( .A(n4839), .B(n4840), .Z(n4831) );
  AND U4639 ( .A(n203), .B(n4841), .Z(n4840) );
  XNOR U4640 ( .A(n4842), .B(n4843), .Z(n4837) );
  AND U4641 ( .A(n195), .B(n4844), .Z(n4843) );
  XOR U4642 ( .A(p_input[386]), .B(n4842), .Z(n4844) );
  XNOR U4643 ( .A(n4845), .B(n4846), .Z(n4842) );
  AND U4644 ( .A(n199), .B(n4841), .Z(n4846) );
  XNOR U4645 ( .A(n4845), .B(n4839), .Z(n4841) );
  XOR U4646 ( .A(n4847), .B(n4848), .Z(n4839) );
  AND U4647 ( .A(n214), .B(n4849), .Z(n4848) );
  XNOR U4648 ( .A(n4850), .B(n4851), .Z(n4845) );
  AND U4649 ( .A(n206), .B(n4852), .Z(n4851) );
  XOR U4650 ( .A(p_input[418]), .B(n4850), .Z(n4852) );
  XNOR U4651 ( .A(n4853), .B(n4854), .Z(n4850) );
  AND U4652 ( .A(n210), .B(n4849), .Z(n4854) );
  XNOR U4653 ( .A(n4853), .B(n4847), .Z(n4849) );
  XOR U4654 ( .A(n4855), .B(n4856), .Z(n4847) );
  AND U4655 ( .A(n225), .B(n4857), .Z(n4856) );
  XNOR U4656 ( .A(n4858), .B(n4859), .Z(n4853) );
  AND U4657 ( .A(n217), .B(n4860), .Z(n4859) );
  XOR U4658 ( .A(p_input[450]), .B(n4858), .Z(n4860) );
  XNOR U4659 ( .A(n4861), .B(n4862), .Z(n4858) );
  AND U4660 ( .A(n221), .B(n4857), .Z(n4862) );
  XNOR U4661 ( .A(n4861), .B(n4855), .Z(n4857) );
  XOR U4662 ( .A(n4863), .B(n4864), .Z(n4855) );
  AND U4663 ( .A(n236), .B(n4865), .Z(n4864) );
  XNOR U4664 ( .A(n4866), .B(n4867), .Z(n4861) );
  AND U4665 ( .A(n228), .B(n4868), .Z(n4867) );
  XOR U4666 ( .A(p_input[482]), .B(n4866), .Z(n4868) );
  XNOR U4667 ( .A(n4869), .B(n4870), .Z(n4866) );
  AND U4668 ( .A(n232), .B(n4865), .Z(n4870) );
  XNOR U4669 ( .A(n4869), .B(n4863), .Z(n4865) );
  XOR U4670 ( .A(n4871), .B(n4872), .Z(n4863) );
  AND U4671 ( .A(n247), .B(n4873), .Z(n4872) );
  XNOR U4672 ( .A(n4874), .B(n4875), .Z(n4869) );
  AND U4673 ( .A(n239), .B(n4876), .Z(n4875) );
  XOR U4674 ( .A(p_input[514]), .B(n4874), .Z(n4876) );
  XNOR U4675 ( .A(n4877), .B(n4878), .Z(n4874) );
  AND U4676 ( .A(n243), .B(n4873), .Z(n4878) );
  XNOR U4677 ( .A(n4877), .B(n4871), .Z(n4873) );
  XOR U4678 ( .A(n4879), .B(n4880), .Z(n4871) );
  AND U4679 ( .A(n258), .B(n4881), .Z(n4880) );
  XNOR U4680 ( .A(n4882), .B(n4883), .Z(n4877) );
  AND U4681 ( .A(n250), .B(n4884), .Z(n4883) );
  XOR U4682 ( .A(p_input[546]), .B(n4882), .Z(n4884) );
  XNOR U4683 ( .A(n4885), .B(n4886), .Z(n4882) );
  AND U4684 ( .A(n254), .B(n4881), .Z(n4886) );
  XNOR U4685 ( .A(n4885), .B(n4879), .Z(n4881) );
  XOR U4686 ( .A(n4887), .B(n4888), .Z(n4879) );
  AND U4687 ( .A(n269), .B(n4889), .Z(n4888) );
  XNOR U4688 ( .A(n4890), .B(n4891), .Z(n4885) );
  AND U4689 ( .A(n261), .B(n4892), .Z(n4891) );
  XOR U4690 ( .A(p_input[578]), .B(n4890), .Z(n4892) );
  XNOR U4691 ( .A(n4893), .B(n4894), .Z(n4890) );
  AND U4692 ( .A(n265), .B(n4889), .Z(n4894) );
  XNOR U4693 ( .A(n4893), .B(n4887), .Z(n4889) );
  XOR U4694 ( .A(n4895), .B(n4896), .Z(n4887) );
  AND U4695 ( .A(n280), .B(n4897), .Z(n4896) );
  XNOR U4696 ( .A(n4898), .B(n4899), .Z(n4893) );
  AND U4697 ( .A(n272), .B(n4900), .Z(n4899) );
  XOR U4698 ( .A(p_input[610]), .B(n4898), .Z(n4900) );
  XNOR U4699 ( .A(n4901), .B(n4902), .Z(n4898) );
  AND U4700 ( .A(n276), .B(n4897), .Z(n4902) );
  XNOR U4701 ( .A(n4901), .B(n4895), .Z(n4897) );
  XOR U4702 ( .A(n4903), .B(n4904), .Z(n4895) );
  AND U4703 ( .A(n291), .B(n4905), .Z(n4904) );
  XNOR U4704 ( .A(n4906), .B(n4907), .Z(n4901) );
  AND U4705 ( .A(n283), .B(n4908), .Z(n4907) );
  XOR U4706 ( .A(p_input[642]), .B(n4906), .Z(n4908) );
  XNOR U4707 ( .A(n4909), .B(n4910), .Z(n4906) );
  AND U4708 ( .A(n287), .B(n4905), .Z(n4910) );
  XNOR U4709 ( .A(n4909), .B(n4903), .Z(n4905) );
  XOR U4710 ( .A(n4911), .B(n4912), .Z(n4903) );
  AND U4711 ( .A(n302), .B(n4913), .Z(n4912) );
  XNOR U4712 ( .A(n4914), .B(n4915), .Z(n4909) );
  AND U4713 ( .A(n294), .B(n4916), .Z(n4915) );
  XOR U4714 ( .A(p_input[674]), .B(n4914), .Z(n4916) );
  XNOR U4715 ( .A(n4917), .B(n4918), .Z(n4914) );
  AND U4716 ( .A(n298), .B(n4913), .Z(n4918) );
  XNOR U4717 ( .A(n4917), .B(n4911), .Z(n4913) );
  XOR U4718 ( .A(n4919), .B(n4920), .Z(n4911) );
  AND U4719 ( .A(n313), .B(n4921), .Z(n4920) );
  XNOR U4720 ( .A(n4922), .B(n4923), .Z(n4917) );
  AND U4721 ( .A(n305), .B(n4924), .Z(n4923) );
  XOR U4722 ( .A(p_input[706]), .B(n4922), .Z(n4924) );
  XNOR U4723 ( .A(n4925), .B(n4926), .Z(n4922) );
  AND U4724 ( .A(n309), .B(n4921), .Z(n4926) );
  XNOR U4725 ( .A(n4925), .B(n4919), .Z(n4921) );
  XOR U4726 ( .A(n4927), .B(n4928), .Z(n4919) );
  AND U4727 ( .A(n324), .B(n4929), .Z(n4928) );
  XNOR U4728 ( .A(n4930), .B(n4931), .Z(n4925) );
  AND U4729 ( .A(n316), .B(n4932), .Z(n4931) );
  XOR U4730 ( .A(p_input[738]), .B(n4930), .Z(n4932) );
  XNOR U4731 ( .A(n4933), .B(n4934), .Z(n4930) );
  AND U4732 ( .A(n320), .B(n4929), .Z(n4934) );
  XNOR U4733 ( .A(n4933), .B(n4927), .Z(n4929) );
  XOR U4734 ( .A(n4935), .B(n4936), .Z(n4927) );
  AND U4735 ( .A(n335), .B(n4937), .Z(n4936) );
  XNOR U4736 ( .A(n4938), .B(n4939), .Z(n4933) );
  AND U4737 ( .A(n327), .B(n4940), .Z(n4939) );
  XOR U4738 ( .A(p_input[770]), .B(n4938), .Z(n4940) );
  XNOR U4739 ( .A(n4941), .B(n4942), .Z(n4938) );
  AND U4740 ( .A(n331), .B(n4937), .Z(n4942) );
  XNOR U4741 ( .A(n4941), .B(n4935), .Z(n4937) );
  XOR U4742 ( .A(n4943), .B(n4944), .Z(n4935) );
  AND U4743 ( .A(n346), .B(n4945), .Z(n4944) );
  XNOR U4744 ( .A(n4946), .B(n4947), .Z(n4941) );
  AND U4745 ( .A(n338), .B(n4948), .Z(n4947) );
  XOR U4746 ( .A(p_input[802]), .B(n4946), .Z(n4948) );
  XNOR U4747 ( .A(n4949), .B(n4950), .Z(n4946) );
  AND U4748 ( .A(n342), .B(n4945), .Z(n4950) );
  XNOR U4749 ( .A(n4949), .B(n4943), .Z(n4945) );
  XOR U4750 ( .A(n4951), .B(n4952), .Z(n4943) );
  AND U4751 ( .A(n357), .B(n4953), .Z(n4952) );
  XNOR U4752 ( .A(n4954), .B(n4955), .Z(n4949) );
  AND U4753 ( .A(n349), .B(n4956), .Z(n4955) );
  XOR U4754 ( .A(p_input[834]), .B(n4954), .Z(n4956) );
  XNOR U4755 ( .A(n4957), .B(n4958), .Z(n4954) );
  AND U4756 ( .A(n353), .B(n4953), .Z(n4958) );
  XNOR U4757 ( .A(n4957), .B(n4951), .Z(n4953) );
  XOR U4758 ( .A(n4959), .B(n4960), .Z(n4951) );
  AND U4759 ( .A(n368), .B(n4961), .Z(n4960) );
  XNOR U4760 ( .A(n4962), .B(n4963), .Z(n4957) );
  AND U4761 ( .A(n360), .B(n4964), .Z(n4963) );
  XOR U4762 ( .A(p_input[866]), .B(n4962), .Z(n4964) );
  XNOR U4763 ( .A(n4965), .B(n4966), .Z(n4962) );
  AND U4764 ( .A(n364), .B(n4961), .Z(n4966) );
  XNOR U4765 ( .A(n4965), .B(n4959), .Z(n4961) );
  XOR U4766 ( .A(n4967), .B(n4968), .Z(n4959) );
  AND U4767 ( .A(n379), .B(n4969), .Z(n4968) );
  XNOR U4768 ( .A(n4970), .B(n4971), .Z(n4965) );
  AND U4769 ( .A(n371), .B(n4972), .Z(n4971) );
  XOR U4770 ( .A(p_input[898]), .B(n4970), .Z(n4972) );
  XNOR U4771 ( .A(n4973), .B(n4974), .Z(n4970) );
  AND U4772 ( .A(n375), .B(n4969), .Z(n4974) );
  XNOR U4773 ( .A(n4973), .B(n4967), .Z(n4969) );
  XOR U4774 ( .A(n4975), .B(n4976), .Z(n4967) );
  AND U4775 ( .A(n390), .B(n4977), .Z(n4976) );
  XNOR U4776 ( .A(n4978), .B(n4979), .Z(n4973) );
  AND U4777 ( .A(n382), .B(n4980), .Z(n4979) );
  XOR U4778 ( .A(p_input[930]), .B(n4978), .Z(n4980) );
  XNOR U4779 ( .A(n4981), .B(n4982), .Z(n4978) );
  AND U4780 ( .A(n386), .B(n4977), .Z(n4982) );
  XNOR U4781 ( .A(n4981), .B(n4975), .Z(n4977) );
  XOR U4782 ( .A(n4983), .B(n4984), .Z(n4975) );
  AND U4783 ( .A(n401), .B(n4985), .Z(n4984) );
  XNOR U4784 ( .A(n4986), .B(n4987), .Z(n4981) );
  AND U4785 ( .A(n393), .B(n4988), .Z(n4987) );
  XOR U4786 ( .A(p_input[962]), .B(n4986), .Z(n4988) );
  XNOR U4787 ( .A(n4989), .B(n4990), .Z(n4986) );
  AND U4788 ( .A(n397), .B(n4985), .Z(n4990) );
  XNOR U4789 ( .A(n4989), .B(n4983), .Z(n4985) );
  XOR U4790 ( .A(n4991), .B(n4992), .Z(n4983) );
  AND U4791 ( .A(n412), .B(n4993), .Z(n4992) );
  XNOR U4792 ( .A(n4994), .B(n4995), .Z(n4989) );
  AND U4793 ( .A(n404), .B(n4996), .Z(n4995) );
  XOR U4794 ( .A(p_input[994]), .B(n4994), .Z(n4996) );
  XNOR U4795 ( .A(n4997), .B(n4998), .Z(n4994) );
  AND U4796 ( .A(n408), .B(n4993), .Z(n4998) );
  XNOR U4797 ( .A(n4997), .B(n4991), .Z(n4993) );
  XOR U4798 ( .A(n4999), .B(n5000), .Z(n4991) );
  AND U4799 ( .A(n423), .B(n5001), .Z(n5000) );
  XNOR U4800 ( .A(n5002), .B(n5003), .Z(n4997) );
  AND U4801 ( .A(n415), .B(n5004), .Z(n5003) );
  XOR U4802 ( .A(p_input[1026]), .B(n5002), .Z(n5004) );
  XNOR U4803 ( .A(n5005), .B(n5006), .Z(n5002) );
  AND U4804 ( .A(n419), .B(n5001), .Z(n5006) );
  XNOR U4805 ( .A(n5005), .B(n4999), .Z(n5001) );
  XOR U4806 ( .A(n5007), .B(n5008), .Z(n4999) );
  AND U4807 ( .A(n434), .B(n5009), .Z(n5008) );
  XNOR U4808 ( .A(n5010), .B(n5011), .Z(n5005) );
  AND U4809 ( .A(n426), .B(n5012), .Z(n5011) );
  XOR U4810 ( .A(p_input[1058]), .B(n5010), .Z(n5012) );
  XNOR U4811 ( .A(n5013), .B(n5014), .Z(n5010) );
  AND U4812 ( .A(n430), .B(n5009), .Z(n5014) );
  XNOR U4813 ( .A(n5013), .B(n5007), .Z(n5009) );
  XOR U4814 ( .A(n5015), .B(n5016), .Z(n5007) );
  AND U4815 ( .A(n445), .B(n5017), .Z(n5016) );
  XNOR U4816 ( .A(n5018), .B(n5019), .Z(n5013) );
  AND U4817 ( .A(n437), .B(n5020), .Z(n5019) );
  XOR U4818 ( .A(p_input[1090]), .B(n5018), .Z(n5020) );
  XNOR U4819 ( .A(n5021), .B(n5022), .Z(n5018) );
  AND U4820 ( .A(n441), .B(n5017), .Z(n5022) );
  XNOR U4821 ( .A(n5021), .B(n5015), .Z(n5017) );
  XOR U4822 ( .A(n5023), .B(n5024), .Z(n5015) );
  AND U4823 ( .A(n456), .B(n5025), .Z(n5024) );
  XNOR U4824 ( .A(n5026), .B(n5027), .Z(n5021) );
  AND U4825 ( .A(n448), .B(n5028), .Z(n5027) );
  XOR U4826 ( .A(p_input[1122]), .B(n5026), .Z(n5028) );
  XNOR U4827 ( .A(n5029), .B(n5030), .Z(n5026) );
  AND U4828 ( .A(n452), .B(n5025), .Z(n5030) );
  XNOR U4829 ( .A(n5029), .B(n5023), .Z(n5025) );
  XOR U4830 ( .A(n5031), .B(n5032), .Z(n5023) );
  AND U4831 ( .A(n467), .B(n5033), .Z(n5032) );
  XNOR U4832 ( .A(n5034), .B(n5035), .Z(n5029) );
  AND U4833 ( .A(n459), .B(n5036), .Z(n5035) );
  XOR U4834 ( .A(p_input[1154]), .B(n5034), .Z(n5036) );
  XNOR U4835 ( .A(n5037), .B(n5038), .Z(n5034) );
  AND U4836 ( .A(n463), .B(n5033), .Z(n5038) );
  XNOR U4837 ( .A(n5037), .B(n5031), .Z(n5033) );
  XOR U4838 ( .A(n5039), .B(n5040), .Z(n5031) );
  AND U4839 ( .A(n478), .B(n5041), .Z(n5040) );
  XNOR U4840 ( .A(n5042), .B(n5043), .Z(n5037) );
  AND U4841 ( .A(n470), .B(n5044), .Z(n5043) );
  XOR U4842 ( .A(p_input[1186]), .B(n5042), .Z(n5044) );
  XNOR U4843 ( .A(n5045), .B(n5046), .Z(n5042) );
  AND U4844 ( .A(n474), .B(n5041), .Z(n5046) );
  XNOR U4845 ( .A(n5045), .B(n5039), .Z(n5041) );
  XOR U4846 ( .A(n5047), .B(n5048), .Z(n5039) );
  AND U4847 ( .A(n489), .B(n5049), .Z(n5048) );
  XNOR U4848 ( .A(n5050), .B(n5051), .Z(n5045) );
  AND U4849 ( .A(n481), .B(n5052), .Z(n5051) );
  XOR U4850 ( .A(p_input[1218]), .B(n5050), .Z(n5052) );
  XNOR U4851 ( .A(n5053), .B(n5054), .Z(n5050) );
  AND U4852 ( .A(n485), .B(n5049), .Z(n5054) );
  XNOR U4853 ( .A(n5053), .B(n5047), .Z(n5049) );
  XOR U4854 ( .A(n5055), .B(n5056), .Z(n5047) );
  AND U4855 ( .A(n500), .B(n5057), .Z(n5056) );
  XNOR U4856 ( .A(n5058), .B(n5059), .Z(n5053) );
  AND U4857 ( .A(n492), .B(n5060), .Z(n5059) );
  XOR U4858 ( .A(p_input[1250]), .B(n5058), .Z(n5060) );
  XNOR U4859 ( .A(n5061), .B(n5062), .Z(n5058) );
  AND U4860 ( .A(n496), .B(n5057), .Z(n5062) );
  XNOR U4861 ( .A(n5061), .B(n5055), .Z(n5057) );
  XOR U4862 ( .A(n5063), .B(n5064), .Z(n5055) );
  AND U4863 ( .A(n511), .B(n5065), .Z(n5064) );
  XNOR U4864 ( .A(n5066), .B(n5067), .Z(n5061) );
  AND U4865 ( .A(n503), .B(n5068), .Z(n5067) );
  XOR U4866 ( .A(p_input[1282]), .B(n5066), .Z(n5068) );
  XNOR U4867 ( .A(n5069), .B(n5070), .Z(n5066) );
  AND U4868 ( .A(n507), .B(n5065), .Z(n5070) );
  XNOR U4869 ( .A(n5069), .B(n5063), .Z(n5065) );
  XOR U4870 ( .A(n5071), .B(n5072), .Z(n5063) );
  AND U4871 ( .A(n522), .B(n5073), .Z(n5072) );
  XNOR U4872 ( .A(n5074), .B(n5075), .Z(n5069) );
  AND U4873 ( .A(n514), .B(n5076), .Z(n5075) );
  XOR U4874 ( .A(p_input[1314]), .B(n5074), .Z(n5076) );
  XNOR U4875 ( .A(n5077), .B(n5078), .Z(n5074) );
  AND U4876 ( .A(n518), .B(n5073), .Z(n5078) );
  XNOR U4877 ( .A(n5077), .B(n5071), .Z(n5073) );
  XOR U4878 ( .A(n5079), .B(n5080), .Z(n5071) );
  AND U4879 ( .A(n533), .B(n5081), .Z(n5080) );
  XNOR U4880 ( .A(n5082), .B(n5083), .Z(n5077) );
  AND U4881 ( .A(n525), .B(n5084), .Z(n5083) );
  XOR U4882 ( .A(p_input[1346]), .B(n5082), .Z(n5084) );
  XNOR U4883 ( .A(n5085), .B(n5086), .Z(n5082) );
  AND U4884 ( .A(n529), .B(n5081), .Z(n5086) );
  XNOR U4885 ( .A(n5085), .B(n5079), .Z(n5081) );
  XOR U4886 ( .A(n5087), .B(n5088), .Z(n5079) );
  AND U4887 ( .A(n544), .B(n5089), .Z(n5088) );
  XNOR U4888 ( .A(n5090), .B(n5091), .Z(n5085) );
  AND U4889 ( .A(n536), .B(n5092), .Z(n5091) );
  XOR U4890 ( .A(p_input[1378]), .B(n5090), .Z(n5092) );
  XNOR U4891 ( .A(n5093), .B(n5094), .Z(n5090) );
  AND U4892 ( .A(n540), .B(n5089), .Z(n5094) );
  XNOR U4893 ( .A(n5093), .B(n5087), .Z(n5089) );
  XOR U4894 ( .A(n5095), .B(n5096), .Z(n5087) );
  AND U4895 ( .A(n555), .B(n5097), .Z(n5096) );
  XNOR U4896 ( .A(n5098), .B(n5099), .Z(n5093) );
  AND U4897 ( .A(n547), .B(n5100), .Z(n5099) );
  XOR U4898 ( .A(p_input[1410]), .B(n5098), .Z(n5100) );
  XNOR U4899 ( .A(n5101), .B(n5102), .Z(n5098) );
  AND U4900 ( .A(n551), .B(n5097), .Z(n5102) );
  XNOR U4901 ( .A(n5101), .B(n5095), .Z(n5097) );
  XOR U4902 ( .A(n5103), .B(n5104), .Z(n5095) );
  AND U4903 ( .A(n566), .B(n5105), .Z(n5104) );
  XNOR U4904 ( .A(n5106), .B(n5107), .Z(n5101) );
  AND U4905 ( .A(n558), .B(n5108), .Z(n5107) );
  XOR U4906 ( .A(p_input[1442]), .B(n5106), .Z(n5108) );
  XNOR U4907 ( .A(n5109), .B(n5110), .Z(n5106) );
  AND U4908 ( .A(n562), .B(n5105), .Z(n5110) );
  XNOR U4909 ( .A(n5109), .B(n5103), .Z(n5105) );
  XOR U4910 ( .A(n5111), .B(n5112), .Z(n5103) );
  AND U4911 ( .A(n577), .B(n5113), .Z(n5112) );
  XNOR U4912 ( .A(n5114), .B(n5115), .Z(n5109) );
  AND U4913 ( .A(n569), .B(n5116), .Z(n5115) );
  XOR U4914 ( .A(p_input[1474]), .B(n5114), .Z(n5116) );
  XNOR U4915 ( .A(n5117), .B(n5118), .Z(n5114) );
  AND U4916 ( .A(n573), .B(n5113), .Z(n5118) );
  XNOR U4917 ( .A(n5117), .B(n5111), .Z(n5113) );
  XOR U4918 ( .A(n5119), .B(n5120), .Z(n5111) );
  AND U4919 ( .A(n588), .B(n5121), .Z(n5120) );
  XNOR U4920 ( .A(n5122), .B(n5123), .Z(n5117) );
  AND U4921 ( .A(n580), .B(n5124), .Z(n5123) );
  XOR U4922 ( .A(p_input[1506]), .B(n5122), .Z(n5124) );
  XNOR U4923 ( .A(n5125), .B(n5126), .Z(n5122) );
  AND U4924 ( .A(n584), .B(n5121), .Z(n5126) );
  XNOR U4925 ( .A(n5125), .B(n5119), .Z(n5121) );
  XOR U4926 ( .A(n5127), .B(n5128), .Z(n5119) );
  AND U4927 ( .A(n599), .B(n5129), .Z(n5128) );
  XNOR U4928 ( .A(n5130), .B(n5131), .Z(n5125) );
  AND U4929 ( .A(n591), .B(n5132), .Z(n5131) );
  XOR U4930 ( .A(p_input[1538]), .B(n5130), .Z(n5132) );
  XNOR U4931 ( .A(n5133), .B(n5134), .Z(n5130) );
  AND U4932 ( .A(n595), .B(n5129), .Z(n5134) );
  XNOR U4933 ( .A(n5133), .B(n5127), .Z(n5129) );
  XOR U4934 ( .A(n5135), .B(n5136), .Z(n5127) );
  AND U4935 ( .A(n610), .B(n5137), .Z(n5136) );
  XNOR U4936 ( .A(n5138), .B(n5139), .Z(n5133) );
  AND U4937 ( .A(n602), .B(n5140), .Z(n5139) );
  XOR U4938 ( .A(p_input[1570]), .B(n5138), .Z(n5140) );
  XNOR U4939 ( .A(n5141), .B(n5142), .Z(n5138) );
  AND U4940 ( .A(n606), .B(n5137), .Z(n5142) );
  XNOR U4941 ( .A(n5141), .B(n5135), .Z(n5137) );
  XOR U4942 ( .A(n5143), .B(n5144), .Z(n5135) );
  AND U4943 ( .A(n621), .B(n5145), .Z(n5144) );
  XNOR U4944 ( .A(n5146), .B(n5147), .Z(n5141) );
  AND U4945 ( .A(n613), .B(n5148), .Z(n5147) );
  XOR U4946 ( .A(p_input[1602]), .B(n5146), .Z(n5148) );
  XNOR U4947 ( .A(n5149), .B(n5150), .Z(n5146) );
  AND U4948 ( .A(n617), .B(n5145), .Z(n5150) );
  XNOR U4949 ( .A(n5149), .B(n5143), .Z(n5145) );
  XOR U4950 ( .A(n5151), .B(n5152), .Z(n5143) );
  AND U4951 ( .A(n632), .B(n5153), .Z(n5152) );
  XNOR U4952 ( .A(n5154), .B(n5155), .Z(n5149) );
  AND U4953 ( .A(n624), .B(n5156), .Z(n5155) );
  XOR U4954 ( .A(p_input[1634]), .B(n5154), .Z(n5156) );
  XNOR U4955 ( .A(n5157), .B(n5158), .Z(n5154) );
  AND U4956 ( .A(n628), .B(n5153), .Z(n5158) );
  XNOR U4957 ( .A(n5157), .B(n5151), .Z(n5153) );
  XOR U4958 ( .A(n5159), .B(n5160), .Z(n5151) );
  AND U4959 ( .A(n643), .B(n5161), .Z(n5160) );
  XNOR U4960 ( .A(n5162), .B(n5163), .Z(n5157) );
  AND U4961 ( .A(n635), .B(n5164), .Z(n5163) );
  XOR U4962 ( .A(p_input[1666]), .B(n5162), .Z(n5164) );
  XNOR U4963 ( .A(n5165), .B(n5166), .Z(n5162) );
  AND U4964 ( .A(n639), .B(n5161), .Z(n5166) );
  XNOR U4965 ( .A(n5165), .B(n5159), .Z(n5161) );
  XOR U4966 ( .A(n5167), .B(n5168), .Z(n5159) );
  AND U4967 ( .A(n654), .B(n5169), .Z(n5168) );
  XNOR U4968 ( .A(n5170), .B(n5171), .Z(n5165) );
  AND U4969 ( .A(n646), .B(n5172), .Z(n5171) );
  XOR U4970 ( .A(p_input[1698]), .B(n5170), .Z(n5172) );
  XNOR U4971 ( .A(n5173), .B(n5174), .Z(n5170) );
  AND U4972 ( .A(n650), .B(n5169), .Z(n5174) );
  XNOR U4973 ( .A(n5173), .B(n5167), .Z(n5169) );
  XOR U4974 ( .A(n5175), .B(n5176), .Z(n5167) );
  AND U4975 ( .A(n665), .B(n5177), .Z(n5176) );
  XNOR U4976 ( .A(n5178), .B(n5179), .Z(n5173) );
  AND U4977 ( .A(n657), .B(n5180), .Z(n5179) );
  XOR U4978 ( .A(p_input[1730]), .B(n5178), .Z(n5180) );
  XNOR U4979 ( .A(n5181), .B(n5182), .Z(n5178) );
  AND U4980 ( .A(n661), .B(n5177), .Z(n5182) );
  XNOR U4981 ( .A(n5181), .B(n5175), .Z(n5177) );
  XOR U4982 ( .A(n5183), .B(n5184), .Z(n5175) );
  AND U4983 ( .A(n676), .B(n5185), .Z(n5184) );
  XNOR U4984 ( .A(n5186), .B(n5187), .Z(n5181) );
  AND U4985 ( .A(n668), .B(n5188), .Z(n5187) );
  XOR U4986 ( .A(p_input[1762]), .B(n5186), .Z(n5188) );
  XNOR U4987 ( .A(n5189), .B(n5190), .Z(n5186) );
  AND U4988 ( .A(n672), .B(n5185), .Z(n5190) );
  XNOR U4989 ( .A(n5189), .B(n5183), .Z(n5185) );
  XOR U4990 ( .A(n5191), .B(n5192), .Z(n5183) );
  AND U4991 ( .A(n687), .B(n5193), .Z(n5192) );
  XNOR U4992 ( .A(n5194), .B(n5195), .Z(n5189) );
  AND U4993 ( .A(n679), .B(n5196), .Z(n5195) );
  XOR U4994 ( .A(p_input[1794]), .B(n5194), .Z(n5196) );
  XNOR U4995 ( .A(n5197), .B(n5198), .Z(n5194) );
  AND U4996 ( .A(n683), .B(n5193), .Z(n5198) );
  XNOR U4997 ( .A(n5197), .B(n5191), .Z(n5193) );
  XOR U4998 ( .A(n5199), .B(n5200), .Z(n5191) );
  AND U4999 ( .A(n698), .B(n5201), .Z(n5200) );
  XNOR U5000 ( .A(n5202), .B(n5203), .Z(n5197) );
  AND U5001 ( .A(n690), .B(n5204), .Z(n5203) );
  XOR U5002 ( .A(p_input[1826]), .B(n5202), .Z(n5204) );
  XNOR U5003 ( .A(n5205), .B(n5206), .Z(n5202) );
  AND U5004 ( .A(n694), .B(n5201), .Z(n5206) );
  XNOR U5005 ( .A(n5205), .B(n5199), .Z(n5201) );
  XOR U5006 ( .A(n5207), .B(n5208), .Z(n5199) );
  AND U5007 ( .A(n709), .B(n5209), .Z(n5208) );
  XNOR U5008 ( .A(n5210), .B(n5211), .Z(n5205) );
  AND U5009 ( .A(n701), .B(n5212), .Z(n5211) );
  XOR U5010 ( .A(p_input[1858]), .B(n5210), .Z(n5212) );
  XNOR U5011 ( .A(n5213), .B(n5214), .Z(n5210) );
  AND U5012 ( .A(n705), .B(n5209), .Z(n5214) );
  XNOR U5013 ( .A(n5213), .B(n5207), .Z(n5209) );
  XOR U5014 ( .A(n5215), .B(n5216), .Z(n5207) );
  AND U5015 ( .A(n720), .B(n5217), .Z(n5216) );
  XNOR U5016 ( .A(n5218), .B(n5219), .Z(n5213) );
  AND U5017 ( .A(n712), .B(n5220), .Z(n5219) );
  XOR U5018 ( .A(p_input[1890]), .B(n5218), .Z(n5220) );
  XNOR U5019 ( .A(n5221), .B(n5222), .Z(n5218) );
  AND U5020 ( .A(n716), .B(n5217), .Z(n5222) );
  XNOR U5021 ( .A(n5221), .B(n5215), .Z(n5217) );
  XOR U5022 ( .A(n5223), .B(n5224), .Z(n5215) );
  AND U5023 ( .A(n731), .B(n5225), .Z(n5224) );
  XNOR U5024 ( .A(n5226), .B(n5227), .Z(n5221) );
  AND U5025 ( .A(n723), .B(n5228), .Z(n5227) );
  XOR U5026 ( .A(p_input[1922]), .B(n5226), .Z(n5228) );
  XNOR U5027 ( .A(n5229), .B(n5230), .Z(n5226) );
  AND U5028 ( .A(n727), .B(n5225), .Z(n5230) );
  XNOR U5029 ( .A(n5229), .B(n5223), .Z(n5225) );
  XOR U5030 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n5231), .Z(n5223) );
  AND U5031 ( .A(n741), .B(n5232), .Z(n5231) );
  XNOR U5032 ( .A(n5233), .B(n5234), .Z(n5229) );
  AND U5033 ( .A(n734), .B(n5235), .Z(n5234) );
  XOR U5034 ( .A(p_input[1954]), .B(n5233), .Z(n5235) );
  XNOR U5035 ( .A(n5236), .B(n5237), .Z(n5233) );
  AND U5036 ( .A(n738), .B(n5232), .Z(n5237) );
  XOR U5037 ( .A(\knn_comb_/min_val_out[0][2] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n5232) );
  XOR U5038 ( .A(n13), .B(n5238), .Z(o[29]) );
  AND U5039 ( .A(n58), .B(n5239), .Z(n13) );
  XOR U5040 ( .A(n14), .B(n5238), .Z(n5239) );
  XOR U5041 ( .A(n5240), .B(n5241), .Z(n5238) );
  AND U5042 ( .A(n70), .B(n5242), .Z(n5241) );
  XOR U5043 ( .A(n5243), .B(n5244), .Z(n14) );
  AND U5044 ( .A(n62), .B(n5245), .Z(n5244) );
  XOR U5045 ( .A(p_input[29]), .B(n5243), .Z(n5245) );
  XNOR U5046 ( .A(n5246), .B(n5247), .Z(n5243) );
  AND U5047 ( .A(n66), .B(n5242), .Z(n5247) );
  XNOR U5048 ( .A(n5246), .B(n5240), .Z(n5242) );
  XOR U5049 ( .A(n5248), .B(n5249), .Z(n5240) );
  AND U5050 ( .A(n82), .B(n5250), .Z(n5249) );
  XNOR U5051 ( .A(n5251), .B(n5252), .Z(n5246) );
  AND U5052 ( .A(n74), .B(n5253), .Z(n5252) );
  XOR U5053 ( .A(p_input[61]), .B(n5251), .Z(n5253) );
  XNOR U5054 ( .A(n5254), .B(n5255), .Z(n5251) );
  AND U5055 ( .A(n78), .B(n5250), .Z(n5255) );
  XNOR U5056 ( .A(n5254), .B(n5248), .Z(n5250) );
  XOR U5057 ( .A(n5256), .B(n5257), .Z(n5248) );
  AND U5058 ( .A(n93), .B(n5258), .Z(n5257) );
  XNOR U5059 ( .A(n5259), .B(n5260), .Z(n5254) );
  AND U5060 ( .A(n85), .B(n5261), .Z(n5260) );
  XOR U5061 ( .A(p_input[93]), .B(n5259), .Z(n5261) );
  XNOR U5062 ( .A(n5262), .B(n5263), .Z(n5259) );
  AND U5063 ( .A(n89), .B(n5258), .Z(n5263) );
  XNOR U5064 ( .A(n5262), .B(n5256), .Z(n5258) );
  XOR U5065 ( .A(n5264), .B(n5265), .Z(n5256) );
  AND U5066 ( .A(n104), .B(n5266), .Z(n5265) );
  XNOR U5067 ( .A(n5267), .B(n5268), .Z(n5262) );
  AND U5068 ( .A(n96), .B(n5269), .Z(n5268) );
  XOR U5069 ( .A(p_input[125]), .B(n5267), .Z(n5269) );
  XNOR U5070 ( .A(n5270), .B(n5271), .Z(n5267) );
  AND U5071 ( .A(n100), .B(n5266), .Z(n5271) );
  XNOR U5072 ( .A(n5270), .B(n5264), .Z(n5266) );
  XOR U5073 ( .A(n5272), .B(n5273), .Z(n5264) );
  AND U5074 ( .A(n115), .B(n5274), .Z(n5273) );
  XNOR U5075 ( .A(n5275), .B(n5276), .Z(n5270) );
  AND U5076 ( .A(n107), .B(n5277), .Z(n5276) );
  XOR U5077 ( .A(p_input[157]), .B(n5275), .Z(n5277) );
  XNOR U5078 ( .A(n5278), .B(n5279), .Z(n5275) );
  AND U5079 ( .A(n111), .B(n5274), .Z(n5279) );
  XNOR U5080 ( .A(n5278), .B(n5272), .Z(n5274) );
  XOR U5081 ( .A(n5280), .B(n5281), .Z(n5272) );
  AND U5082 ( .A(n126), .B(n5282), .Z(n5281) );
  XNOR U5083 ( .A(n5283), .B(n5284), .Z(n5278) );
  AND U5084 ( .A(n118), .B(n5285), .Z(n5284) );
  XOR U5085 ( .A(p_input[189]), .B(n5283), .Z(n5285) );
  XNOR U5086 ( .A(n5286), .B(n5287), .Z(n5283) );
  AND U5087 ( .A(n122), .B(n5282), .Z(n5287) );
  XNOR U5088 ( .A(n5286), .B(n5280), .Z(n5282) );
  XOR U5089 ( .A(n5288), .B(n5289), .Z(n5280) );
  AND U5090 ( .A(n137), .B(n5290), .Z(n5289) );
  XNOR U5091 ( .A(n5291), .B(n5292), .Z(n5286) );
  AND U5092 ( .A(n129), .B(n5293), .Z(n5292) );
  XOR U5093 ( .A(p_input[221]), .B(n5291), .Z(n5293) );
  XNOR U5094 ( .A(n5294), .B(n5295), .Z(n5291) );
  AND U5095 ( .A(n133), .B(n5290), .Z(n5295) );
  XNOR U5096 ( .A(n5294), .B(n5288), .Z(n5290) );
  XOR U5097 ( .A(n5296), .B(n5297), .Z(n5288) );
  AND U5098 ( .A(n148), .B(n5298), .Z(n5297) );
  XNOR U5099 ( .A(n5299), .B(n5300), .Z(n5294) );
  AND U5100 ( .A(n140), .B(n5301), .Z(n5300) );
  XOR U5101 ( .A(p_input[253]), .B(n5299), .Z(n5301) );
  XNOR U5102 ( .A(n5302), .B(n5303), .Z(n5299) );
  AND U5103 ( .A(n144), .B(n5298), .Z(n5303) );
  XNOR U5104 ( .A(n5302), .B(n5296), .Z(n5298) );
  XOR U5105 ( .A(n5304), .B(n5305), .Z(n5296) );
  AND U5106 ( .A(n159), .B(n5306), .Z(n5305) );
  XNOR U5107 ( .A(n5307), .B(n5308), .Z(n5302) );
  AND U5108 ( .A(n151), .B(n5309), .Z(n5308) );
  XOR U5109 ( .A(p_input[285]), .B(n5307), .Z(n5309) );
  XNOR U5110 ( .A(n5310), .B(n5311), .Z(n5307) );
  AND U5111 ( .A(n155), .B(n5306), .Z(n5311) );
  XNOR U5112 ( .A(n5310), .B(n5304), .Z(n5306) );
  XOR U5113 ( .A(n5312), .B(n5313), .Z(n5304) );
  AND U5114 ( .A(n170), .B(n5314), .Z(n5313) );
  XNOR U5115 ( .A(n5315), .B(n5316), .Z(n5310) );
  AND U5116 ( .A(n162), .B(n5317), .Z(n5316) );
  XOR U5117 ( .A(p_input[317]), .B(n5315), .Z(n5317) );
  XNOR U5118 ( .A(n5318), .B(n5319), .Z(n5315) );
  AND U5119 ( .A(n166), .B(n5314), .Z(n5319) );
  XNOR U5120 ( .A(n5318), .B(n5312), .Z(n5314) );
  XOR U5121 ( .A(n5320), .B(n5321), .Z(n5312) );
  AND U5122 ( .A(n181), .B(n5322), .Z(n5321) );
  XNOR U5123 ( .A(n5323), .B(n5324), .Z(n5318) );
  AND U5124 ( .A(n173), .B(n5325), .Z(n5324) );
  XOR U5125 ( .A(p_input[349]), .B(n5323), .Z(n5325) );
  XNOR U5126 ( .A(n5326), .B(n5327), .Z(n5323) );
  AND U5127 ( .A(n177), .B(n5322), .Z(n5327) );
  XNOR U5128 ( .A(n5326), .B(n5320), .Z(n5322) );
  XOR U5129 ( .A(n5328), .B(n5329), .Z(n5320) );
  AND U5130 ( .A(n192), .B(n5330), .Z(n5329) );
  XNOR U5131 ( .A(n5331), .B(n5332), .Z(n5326) );
  AND U5132 ( .A(n184), .B(n5333), .Z(n5332) );
  XOR U5133 ( .A(p_input[381]), .B(n5331), .Z(n5333) );
  XNOR U5134 ( .A(n5334), .B(n5335), .Z(n5331) );
  AND U5135 ( .A(n188), .B(n5330), .Z(n5335) );
  XNOR U5136 ( .A(n5334), .B(n5328), .Z(n5330) );
  XOR U5137 ( .A(n5336), .B(n5337), .Z(n5328) );
  AND U5138 ( .A(n203), .B(n5338), .Z(n5337) );
  XNOR U5139 ( .A(n5339), .B(n5340), .Z(n5334) );
  AND U5140 ( .A(n195), .B(n5341), .Z(n5340) );
  XOR U5141 ( .A(p_input[413]), .B(n5339), .Z(n5341) );
  XNOR U5142 ( .A(n5342), .B(n5343), .Z(n5339) );
  AND U5143 ( .A(n199), .B(n5338), .Z(n5343) );
  XNOR U5144 ( .A(n5342), .B(n5336), .Z(n5338) );
  XOR U5145 ( .A(n5344), .B(n5345), .Z(n5336) );
  AND U5146 ( .A(n214), .B(n5346), .Z(n5345) );
  XNOR U5147 ( .A(n5347), .B(n5348), .Z(n5342) );
  AND U5148 ( .A(n206), .B(n5349), .Z(n5348) );
  XOR U5149 ( .A(p_input[445]), .B(n5347), .Z(n5349) );
  XNOR U5150 ( .A(n5350), .B(n5351), .Z(n5347) );
  AND U5151 ( .A(n210), .B(n5346), .Z(n5351) );
  XNOR U5152 ( .A(n5350), .B(n5344), .Z(n5346) );
  XOR U5153 ( .A(n5352), .B(n5353), .Z(n5344) );
  AND U5154 ( .A(n225), .B(n5354), .Z(n5353) );
  XNOR U5155 ( .A(n5355), .B(n5356), .Z(n5350) );
  AND U5156 ( .A(n217), .B(n5357), .Z(n5356) );
  XOR U5157 ( .A(p_input[477]), .B(n5355), .Z(n5357) );
  XNOR U5158 ( .A(n5358), .B(n5359), .Z(n5355) );
  AND U5159 ( .A(n221), .B(n5354), .Z(n5359) );
  XNOR U5160 ( .A(n5358), .B(n5352), .Z(n5354) );
  XOR U5161 ( .A(n5360), .B(n5361), .Z(n5352) );
  AND U5162 ( .A(n236), .B(n5362), .Z(n5361) );
  XNOR U5163 ( .A(n5363), .B(n5364), .Z(n5358) );
  AND U5164 ( .A(n228), .B(n5365), .Z(n5364) );
  XOR U5165 ( .A(p_input[509]), .B(n5363), .Z(n5365) );
  XNOR U5166 ( .A(n5366), .B(n5367), .Z(n5363) );
  AND U5167 ( .A(n232), .B(n5362), .Z(n5367) );
  XNOR U5168 ( .A(n5366), .B(n5360), .Z(n5362) );
  XOR U5169 ( .A(n5368), .B(n5369), .Z(n5360) );
  AND U5170 ( .A(n247), .B(n5370), .Z(n5369) );
  XNOR U5171 ( .A(n5371), .B(n5372), .Z(n5366) );
  AND U5172 ( .A(n239), .B(n5373), .Z(n5372) );
  XOR U5173 ( .A(p_input[541]), .B(n5371), .Z(n5373) );
  XNOR U5174 ( .A(n5374), .B(n5375), .Z(n5371) );
  AND U5175 ( .A(n243), .B(n5370), .Z(n5375) );
  XNOR U5176 ( .A(n5374), .B(n5368), .Z(n5370) );
  XOR U5177 ( .A(n5376), .B(n5377), .Z(n5368) );
  AND U5178 ( .A(n258), .B(n5378), .Z(n5377) );
  XNOR U5179 ( .A(n5379), .B(n5380), .Z(n5374) );
  AND U5180 ( .A(n250), .B(n5381), .Z(n5380) );
  XOR U5181 ( .A(p_input[573]), .B(n5379), .Z(n5381) );
  XNOR U5182 ( .A(n5382), .B(n5383), .Z(n5379) );
  AND U5183 ( .A(n254), .B(n5378), .Z(n5383) );
  XNOR U5184 ( .A(n5382), .B(n5376), .Z(n5378) );
  XOR U5185 ( .A(n5384), .B(n5385), .Z(n5376) );
  AND U5186 ( .A(n269), .B(n5386), .Z(n5385) );
  XNOR U5187 ( .A(n5387), .B(n5388), .Z(n5382) );
  AND U5188 ( .A(n261), .B(n5389), .Z(n5388) );
  XOR U5189 ( .A(p_input[605]), .B(n5387), .Z(n5389) );
  XNOR U5190 ( .A(n5390), .B(n5391), .Z(n5387) );
  AND U5191 ( .A(n265), .B(n5386), .Z(n5391) );
  XNOR U5192 ( .A(n5390), .B(n5384), .Z(n5386) );
  XOR U5193 ( .A(n5392), .B(n5393), .Z(n5384) );
  AND U5194 ( .A(n280), .B(n5394), .Z(n5393) );
  XNOR U5195 ( .A(n5395), .B(n5396), .Z(n5390) );
  AND U5196 ( .A(n272), .B(n5397), .Z(n5396) );
  XOR U5197 ( .A(p_input[637]), .B(n5395), .Z(n5397) );
  XNOR U5198 ( .A(n5398), .B(n5399), .Z(n5395) );
  AND U5199 ( .A(n276), .B(n5394), .Z(n5399) );
  XNOR U5200 ( .A(n5398), .B(n5392), .Z(n5394) );
  XOR U5201 ( .A(n5400), .B(n5401), .Z(n5392) );
  AND U5202 ( .A(n291), .B(n5402), .Z(n5401) );
  XNOR U5203 ( .A(n5403), .B(n5404), .Z(n5398) );
  AND U5204 ( .A(n283), .B(n5405), .Z(n5404) );
  XOR U5205 ( .A(p_input[669]), .B(n5403), .Z(n5405) );
  XNOR U5206 ( .A(n5406), .B(n5407), .Z(n5403) );
  AND U5207 ( .A(n287), .B(n5402), .Z(n5407) );
  XNOR U5208 ( .A(n5406), .B(n5400), .Z(n5402) );
  XOR U5209 ( .A(n5408), .B(n5409), .Z(n5400) );
  AND U5210 ( .A(n302), .B(n5410), .Z(n5409) );
  XNOR U5211 ( .A(n5411), .B(n5412), .Z(n5406) );
  AND U5212 ( .A(n294), .B(n5413), .Z(n5412) );
  XOR U5213 ( .A(p_input[701]), .B(n5411), .Z(n5413) );
  XNOR U5214 ( .A(n5414), .B(n5415), .Z(n5411) );
  AND U5215 ( .A(n298), .B(n5410), .Z(n5415) );
  XNOR U5216 ( .A(n5414), .B(n5408), .Z(n5410) );
  XOR U5217 ( .A(n5416), .B(n5417), .Z(n5408) );
  AND U5218 ( .A(n313), .B(n5418), .Z(n5417) );
  XNOR U5219 ( .A(n5419), .B(n5420), .Z(n5414) );
  AND U5220 ( .A(n305), .B(n5421), .Z(n5420) );
  XOR U5221 ( .A(p_input[733]), .B(n5419), .Z(n5421) );
  XNOR U5222 ( .A(n5422), .B(n5423), .Z(n5419) );
  AND U5223 ( .A(n309), .B(n5418), .Z(n5423) );
  XNOR U5224 ( .A(n5422), .B(n5416), .Z(n5418) );
  XOR U5225 ( .A(n5424), .B(n5425), .Z(n5416) );
  AND U5226 ( .A(n324), .B(n5426), .Z(n5425) );
  XNOR U5227 ( .A(n5427), .B(n5428), .Z(n5422) );
  AND U5228 ( .A(n316), .B(n5429), .Z(n5428) );
  XOR U5229 ( .A(p_input[765]), .B(n5427), .Z(n5429) );
  XNOR U5230 ( .A(n5430), .B(n5431), .Z(n5427) );
  AND U5231 ( .A(n320), .B(n5426), .Z(n5431) );
  XNOR U5232 ( .A(n5430), .B(n5424), .Z(n5426) );
  XOR U5233 ( .A(n5432), .B(n5433), .Z(n5424) );
  AND U5234 ( .A(n335), .B(n5434), .Z(n5433) );
  XNOR U5235 ( .A(n5435), .B(n5436), .Z(n5430) );
  AND U5236 ( .A(n327), .B(n5437), .Z(n5436) );
  XOR U5237 ( .A(p_input[797]), .B(n5435), .Z(n5437) );
  XNOR U5238 ( .A(n5438), .B(n5439), .Z(n5435) );
  AND U5239 ( .A(n331), .B(n5434), .Z(n5439) );
  XNOR U5240 ( .A(n5438), .B(n5432), .Z(n5434) );
  XOR U5241 ( .A(n5440), .B(n5441), .Z(n5432) );
  AND U5242 ( .A(n346), .B(n5442), .Z(n5441) );
  XNOR U5243 ( .A(n5443), .B(n5444), .Z(n5438) );
  AND U5244 ( .A(n338), .B(n5445), .Z(n5444) );
  XOR U5245 ( .A(p_input[829]), .B(n5443), .Z(n5445) );
  XNOR U5246 ( .A(n5446), .B(n5447), .Z(n5443) );
  AND U5247 ( .A(n342), .B(n5442), .Z(n5447) );
  XNOR U5248 ( .A(n5446), .B(n5440), .Z(n5442) );
  XOR U5249 ( .A(n5448), .B(n5449), .Z(n5440) );
  AND U5250 ( .A(n357), .B(n5450), .Z(n5449) );
  XNOR U5251 ( .A(n5451), .B(n5452), .Z(n5446) );
  AND U5252 ( .A(n349), .B(n5453), .Z(n5452) );
  XOR U5253 ( .A(p_input[861]), .B(n5451), .Z(n5453) );
  XNOR U5254 ( .A(n5454), .B(n5455), .Z(n5451) );
  AND U5255 ( .A(n353), .B(n5450), .Z(n5455) );
  XNOR U5256 ( .A(n5454), .B(n5448), .Z(n5450) );
  XOR U5257 ( .A(n5456), .B(n5457), .Z(n5448) );
  AND U5258 ( .A(n368), .B(n5458), .Z(n5457) );
  XNOR U5259 ( .A(n5459), .B(n5460), .Z(n5454) );
  AND U5260 ( .A(n360), .B(n5461), .Z(n5460) );
  XOR U5261 ( .A(p_input[893]), .B(n5459), .Z(n5461) );
  XNOR U5262 ( .A(n5462), .B(n5463), .Z(n5459) );
  AND U5263 ( .A(n364), .B(n5458), .Z(n5463) );
  XNOR U5264 ( .A(n5462), .B(n5456), .Z(n5458) );
  XOR U5265 ( .A(n5464), .B(n5465), .Z(n5456) );
  AND U5266 ( .A(n379), .B(n5466), .Z(n5465) );
  XNOR U5267 ( .A(n5467), .B(n5468), .Z(n5462) );
  AND U5268 ( .A(n371), .B(n5469), .Z(n5468) );
  XOR U5269 ( .A(p_input[925]), .B(n5467), .Z(n5469) );
  XNOR U5270 ( .A(n5470), .B(n5471), .Z(n5467) );
  AND U5271 ( .A(n375), .B(n5466), .Z(n5471) );
  XNOR U5272 ( .A(n5470), .B(n5464), .Z(n5466) );
  XOR U5273 ( .A(n5472), .B(n5473), .Z(n5464) );
  AND U5274 ( .A(n390), .B(n5474), .Z(n5473) );
  XNOR U5275 ( .A(n5475), .B(n5476), .Z(n5470) );
  AND U5276 ( .A(n382), .B(n5477), .Z(n5476) );
  XOR U5277 ( .A(p_input[957]), .B(n5475), .Z(n5477) );
  XNOR U5278 ( .A(n5478), .B(n5479), .Z(n5475) );
  AND U5279 ( .A(n386), .B(n5474), .Z(n5479) );
  XNOR U5280 ( .A(n5478), .B(n5472), .Z(n5474) );
  XOR U5281 ( .A(n5480), .B(n5481), .Z(n5472) );
  AND U5282 ( .A(n401), .B(n5482), .Z(n5481) );
  XNOR U5283 ( .A(n5483), .B(n5484), .Z(n5478) );
  AND U5284 ( .A(n393), .B(n5485), .Z(n5484) );
  XOR U5285 ( .A(p_input[989]), .B(n5483), .Z(n5485) );
  XNOR U5286 ( .A(n5486), .B(n5487), .Z(n5483) );
  AND U5287 ( .A(n397), .B(n5482), .Z(n5487) );
  XNOR U5288 ( .A(n5486), .B(n5480), .Z(n5482) );
  XOR U5289 ( .A(n5488), .B(n5489), .Z(n5480) );
  AND U5290 ( .A(n412), .B(n5490), .Z(n5489) );
  XNOR U5291 ( .A(n5491), .B(n5492), .Z(n5486) );
  AND U5292 ( .A(n404), .B(n5493), .Z(n5492) );
  XOR U5293 ( .A(p_input[1021]), .B(n5491), .Z(n5493) );
  XNOR U5294 ( .A(n5494), .B(n5495), .Z(n5491) );
  AND U5295 ( .A(n408), .B(n5490), .Z(n5495) );
  XNOR U5296 ( .A(n5494), .B(n5488), .Z(n5490) );
  XOR U5297 ( .A(n5496), .B(n5497), .Z(n5488) );
  AND U5298 ( .A(n423), .B(n5498), .Z(n5497) );
  XNOR U5299 ( .A(n5499), .B(n5500), .Z(n5494) );
  AND U5300 ( .A(n415), .B(n5501), .Z(n5500) );
  XOR U5301 ( .A(p_input[1053]), .B(n5499), .Z(n5501) );
  XNOR U5302 ( .A(n5502), .B(n5503), .Z(n5499) );
  AND U5303 ( .A(n419), .B(n5498), .Z(n5503) );
  XNOR U5304 ( .A(n5502), .B(n5496), .Z(n5498) );
  XOR U5305 ( .A(n5504), .B(n5505), .Z(n5496) );
  AND U5306 ( .A(n434), .B(n5506), .Z(n5505) );
  XNOR U5307 ( .A(n5507), .B(n5508), .Z(n5502) );
  AND U5308 ( .A(n426), .B(n5509), .Z(n5508) );
  XOR U5309 ( .A(p_input[1085]), .B(n5507), .Z(n5509) );
  XNOR U5310 ( .A(n5510), .B(n5511), .Z(n5507) );
  AND U5311 ( .A(n430), .B(n5506), .Z(n5511) );
  XNOR U5312 ( .A(n5510), .B(n5504), .Z(n5506) );
  XOR U5313 ( .A(n5512), .B(n5513), .Z(n5504) );
  AND U5314 ( .A(n445), .B(n5514), .Z(n5513) );
  XNOR U5315 ( .A(n5515), .B(n5516), .Z(n5510) );
  AND U5316 ( .A(n437), .B(n5517), .Z(n5516) );
  XOR U5317 ( .A(p_input[1117]), .B(n5515), .Z(n5517) );
  XNOR U5318 ( .A(n5518), .B(n5519), .Z(n5515) );
  AND U5319 ( .A(n441), .B(n5514), .Z(n5519) );
  XNOR U5320 ( .A(n5518), .B(n5512), .Z(n5514) );
  XOR U5321 ( .A(n5520), .B(n5521), .Z(n5512) );
  AND U5322 ( .A(n456), .B(n5522), .Z(n5521) );
  XNOR U5323 ( .A(n5523), .B(n5524), .Z(n5518) );
  AND U5324 ( .A(n448), .B(n5525), .Z(n5524) );
  XOR U5325 ( .A(p_input[1149]), .B(n5523), .Z(n5525) );
  XNOR U5326 ( .A(n5526), .B(n5527), .Z(n5523) );
  AND U5327 ( .A(n452), .B(n5522), .Z(n5527) );
  XNOR U5328 ( .A(n5526), .B(n5520), .Z(n5522) );
  XOR U5329 ( .A(n5528), .B(n5529), .Z(n5520) );
  AND U5330 ( .A(n467), .B(n5530), .Z(n5529) );
  XNOR U5331 ( .A(n5531), .B(n5532), .Z(n5526) );
  AND U5332 ( .A(n459), .B(n5533), .Z(n5532) );
  XOR U5333 ( .A(p_input[1181]), .B(n5531), .Z(n5533) );
  XNOR U5334 ( .A(n5534), .B(n5535), .Z(n5531) );
  AND U5335 ( .A(n463), .B(n5530), .Z(n5535) );
  XNOR U5336 ( .A(n5534), .B(n5528), .Z(n5530) );
  XOR U5337 ( .A(n5536), .B(n5537), .Z(n5528) );
  AND U5338 ( .A(n478), .B(n5538), .Z(n5537) );
  XNOR U5339 ( .A(n5539), .B(n5540), .Z(n5534) );
  AND U5340 ( .A(n470), .B(n5541), .Z(n5540) );
  XOR U5341 ( .A(p_input[1213]), .B(n5539), .Z(n5541) );
  XNOR U5342 ( .A(n5542), .B(n5543), .Z(n5539) );
  AND U5343 ( .A(n474), .B(n5538), .Z(n5543) );
  XNOR U5344 ( .A(n5542), .B(n5536), .Z(n5538) );
  XOR U5345 ( .A(n5544), .B(n5545), .Z(n5536) );
  AND U5346 ( .A(n489), .B(n5546), .Z(n5545) );
  XNOR U5347 ( .A(n5547), .B(n5548), .Z(n5542) );
  AND U5348 ( .A(n481), .B(n5549), .Z(n5548) );
  XOR U5349 ( .A(p_input[1245]), .B(n5547), .Z(n5549) );
  XNOR U5350 ( .A(n5550), .B(n5551), .Z(n5547) );
  AND U5351 ( .A(n485), .B(n5546), .Z(n5551) );
  XNOR U5352 ( .A(n5550), .B(n5544), .Z(n5546) );
  XOR U5353 ( .A(n5552), .B(n5553), .Z(n5544) );
  AND U5354 ( .A(n500), .B(n5554), .Z(n5553) );
  XNOR U5355 ( .A(n5555), .B(n5556), .Z(n5550) );
  AND U5356 ( .A(n492), .B(n5557), .Z(n5556) );
  XOR U5357 ( .A(p_input[1277]), .B(n5555), .Z(n5557) );
  XNOR U5358 ( .A(n5558), .B(n5559), .Z(n5555) );
  AND U5359 ( .A(n496), .B(n5554), .Z(n5559) );
  XNOR U5360 ( .A(n5558), .B(n5552), .Z(n5554) );
  XOR U5361 ( .A(n5560), .B(n5561), .Z(n5552) );
  AND U5362 ( .A(n511), .B(n5562), .Z(n5561) );
  XNOR U5363 ( .A(n5563), .B(n5564), .Z(n5558) );
  AND U5364 ( .A(n503), .B(n5565), .Z(n5564) );
  XOR U5365 ( .A(p_input[1309]), .B(n5563), .Z(n5565) );
  XNOR U5366 ( .A(n5566), .B(n5567), .Z(n5563) );
  AND U5367 ( .A(n507), .B(n5562), .Z(n5567) );
  XNOR U5368 ( .A(n5566), .B(n5560), .Z(n5562) );
  XOR U5369 ( .A(n5568), .B(n5569), .Z(n5560) );
  AND U5370 ( .A(n522), .B(n5570), .Z(n5569) );
  XNOR U5371 ( .A(n5571), .B(n5572), .Z(n5566) );
  AND U5372 ( .A(n514), .B(n5573), .Z(n5572) );
  XOR U5373 ( .A(p_input[1341]), .B(n5571), .Z(n5573) );
  XNOR U5374 ( .A(n5574), .B(n5575), .Z(n5571) );
  AND U5375 ( .A(n518), .B(n5570), .Z(n5575) );
  XNOR U5376 ( .A(n5574), .B(n5568), .Z(n5570) );
  XOR U5377 ( .A(n5576), .B(n5577), .Z(n5568) );
  AND U5378 ( .A(n533), .B(n5578), .Z(n5577) );
  XNOR U5379 ( .A(n5579), .B(n5580), .Z(n5574) );
  AND U5380 ( .A(n525), .B(n5581), .Z(n5580) );
  XOR U5381 ( .A(p_input[1373]), .B(n5579), .Z(n5581) );
  XNOR U5382 ( .A(n5582), .B(n5583), .Z(n5579) );
  AND U5383 ( .A(n529), .B(n5578), .Z(n5583) );
  XNOR U5384 ( .A(n5582), .B(n5576), .Z(n5578) );
  XOR U5385 ( .A(n5584), .B(n5585), .Z(n5576) );
  AND U5386 ( .A(n544), .B(n5586), .Z(n5585) );
  XNOR U5387 ( .A(n5587), .B(n5588), .Z(n5582) );
  AND U5388 ( .A(n536), .B(n5589), .Z(n5588) );
  XOR U5389 ( .A(p_input[1405]), .B(n5587), .Z(n5589) );
  XNOR U5390 ( .A(n5590), .B(n5591), .Z(n5587) );
  AND U5391 ( .A(n540), .B(n5586), .Z(n5591) );
  XNOR U5392 ( .A(n5590), .B(n5584), .Z(n5586) );
  XOR U5393 ( .A(n5592), .B(n5593), .Z(n5584) );
  AND U5394 ( .A(n555), .B(n5594), .Z(n5593) );
  XNOR U5395 ( .A(n5595), .B(n5596), .Z(n5590) );
  AND U5396 ( .A(n547), .B(n5597), .Z(n5596) );
  XOR U5397 ( .A(p_input[1437]), .B(n5595), .Z(n5597) );
  XNOR U5398 ( .A(n5598), .B(n5599), .Z(n5595) );
  AND U5399 ( .A(n551), .B(n5594), .Z(n5599) );
  XNOR U5400 ( .A(n5598), .B(n5592), .Z(n5594) );
  XOR U5401 ( .A(n5600), .B(n5601), .Z(n5592) );
  AND U5402 ( .A(n566), .B(n5602), .Z(n5601) );
  XNOR U5403 ( .A(n5603), .B(n5604), .Z(n5598) );
  AND U5404 ( .A(n558), .B(n5605), .Z(n5604) );
  XOR U5405 ( .A(p_input[1469]), .B(n5603), .Z(n5605) );
  XNOR U5406 ( .A(n5606), .B(n5607), .Z(n5603) );
  AND U5407 ( .A(n562), .B(n5602), .Z(n5607) );
  XNOR U5408 ( .A(n5606), .B(n5600), .Z(n5602) );
  XOR U5409 ( .A(n5608), .B(n5609), .Z(n5600) );
  AND U5410 ( .A(n577), .B(n5610), .Z(n5609) );
  XNOR U5411 ( .A(n5611), .B(n5612), .Z(n5606) );
  AND U5412 ( .A(n569), .B(n5613), .Z(n5612) );
  XOR U5413 ( .A(p_input[1501]), .B(n5611), .Z(n5613) );
  XNOR U5414 ( .A(n5614), .B(n5615), .Z(n5611) );
  AND U5415 ( .A(n573), .B(n5610), .Z(n5615) );
  XNOR U5416 ( .A(n5614), .B(n5608), .Z(n5610) );
  XOR U5417 ( .A(n5616), .B(n5617), .Z(n5608) );
  AND U5418 ( .A(n588), .B(n5618), .Z(n5617) );
  XNOR U5419 ( .A(n5619), .B(n5620), .Z(n5614) );
  AND U5420 ( .A(n580), .B(n5621), .Z(n5620) );
  XOR U5421 ( .A(p_input[1533]), .B(n5619), .Z(n5621) );
  XNOR U5422 ( .A(n5622), .B(n5623), .Z(n5619) );
  AND U5423 ( .A(n584), .B(n5618), .Z(n5623) );
  XNOR U5424 ( .A(n5622), .B(n5616), .Z(n5618) );
  XOR U5425 ( .A(n5624), .B(n5625), .Z(n5616) );
  AND U5426 ( .A(n599), .B(n5626), .Z(n5625) );
  XNOR U5427 ( .A(n5627), .B(n5628), .Z(n5622) );
  AND U5428 ( .A(n591), .B(n5629), .Z(n5628) );
  XOR U5429 ( .A(p_input[1565]), .B(n5627), .Z(n5629) );
  XNOR U5430 ( .A(n5630), .B(n5631), .Z(n5627) );
  AND U5431 ( .A(n595), .B(n5626), .Z(n5631) );
  XNOR U5432 ( .A(n5630), .B(n5624), .Z(n5626) );
  XOR U5433 ( .A(n5632), .B(n5633), .Z(n5624) );
  AND U5434 ( .A(n610), .B(n5634), .Z(n5633) );
  XNOR U5435 ( .A(n5635), .B(n5636), .Z(n5630) );
  AND U5436 ( .A(n602), .B(n5637), .Z(n5636) );
  XOR U5437 ( .A(p_input[1597]), .B(n5635), .Z(n5637) );
  XNOR U5438 ( .A(n5638), .B(n5639), .Z(n5635) );
  AND U5439 ( .A(n606), .B(n5634), .Z(n5639) );
  XNOR U5440 ( .A(n5638), .B(n5632), .Z(n5634) );
  XOR U5441 ( .A(n5640), .B(n5641), .Z(n5632) );
  AND U5442 ( .A(n621), .B(n5642), .Z(n5641) );
  XNOR U5443 ( .A(n5643), .B(n5644), .Z(n5638) );
  AND U5444 ( .A(n613), .B(n5645), .Z(n5644) );
  XOR U5445 ( .A(p_input[1629]), .B(n5643), .Z(n5645) );
  XNOR U5446 ( .A(n5646), .B(n5647), .Z(n5643) );
  AND U5447 ( .A(n617), .B(n5642), .Z(n5647) );
  XNOR U5448 ( .A(n5646), .B(n5640), .Z(n5642) );
  XOR U5449 ( .A(n5648), .B(n5649), .Z(n5640) );
  AND U5450 ( .A(n632), .B(n5650), .Z(n5649) );
  XNOR U5451 ( .A(n5651), .B(n5652), .Z(n5646) );
  AND U5452 ( .A(n624), .B(n5653), .Z(n5652) );
  XOR U5453 ( .A(p_input[1661]), .B(n5651), .Z(n5653) );
  XNOR U5454 ( .A(n5654), .B(n5655), .Z(n5651) );
  AND U5455 ( .A(n628), .B(n5650), .Z(n5655) );
  XNOR U5456 ( .A(n5654), .B(n5648), .Z(n5650) );
  XOR U5457 ( .A(n5656), .B(n5657), .Z(n5648) );
  AND U5458 ( .A(n643), .B(n5658), .Z(n5657) );
  XNOR U5459 ( .A(n5659), .B(n5660), .Z(n5654) );
  AND U5460 ( .A(n635), .B(n5661), .Z(n5660) );
  XOR U5461 ( .A(p_input[1693]), .B(n5659), .Z(n5661) );
  XNOR U5462 ( .A(n5662), .B(n5663), .Z(n5659) );
  AND U5463 ( .A(n639), .B(n5658), .Z(n5663) );
  XNOR U5464 ( .A(n5662), .B(n5656), .Z(n5658) );
  XOR U5465 ( .A(n5664), .B(n5665), .Z(n5656) );
  AND U5466 ( .A(n654), .B(n5666), .Z(n5665) );
  XNOR U5467 ( .A(n5667), .B(n5668), .Z(n5662) );
  AND U5468 ( .A(n646), .B(n5669), .Z(n5668) );
  XOR U5469 ( .A(p_input[1725]), .B(n5667), .Z(n5669) );
  XNOR U5470 ( .A(n5670), .B(n5671), .Z(n5667) );
  AND U5471 ( .A(n650), .B(n5666), .Z(n5671) );
  XNOR U5472 ( .A(n5670), .B(n5664), .Z(n5666) );
  XOR U5473 ( .A(n5672), .B(n5673), .Z(n5664) );
  AND U5474 ( .A(n665), .B(n5674), .Z(n5673) );
  XNOR U5475 ( .A(n5675), .B(n5676), .Z(n5670) );
  AND U5476 ( .A(n657), .B(n5677), .Z(n5676) );
  XOR U5477 ( .A(p_input[1757]), .B(n5675), .Z(n5677) );
  XNOR U5478 ( .A(n5678), .B(n5679), .Z(n5675) );
  AND U5479 ( .A(n661), .B(n5674), .Z(n5679) );
  XNOR U5480 ( .A(n5678), .B(n5672), .Z(n5674) );
  XOR U5481 ( .A(n5680), .B(n5681), .Z(n5672) );
  AND U5482 ( .A(n676), .B(n5682), .Z(n5681) );
  XNOR U5483 ( .A(n5683), .B(n5684), .Z(n5678) );
  AND U5484 ( .A(n668), .B(n5685), .Z(n5684) );
  XOR U5485 ( .A(p_input[1789]), .B(n5683), .Z(n5685) );
  XNOR U5486 ( .A(n5686), .B(n5687), .Z(n5683) );
  AND U5487 ( .A(n672), .B(n5682), .Z(n5687) );
  XNOR U5488 ( .A(n5686), .B(n5680), .Z(n5682) );
  XOR U5489 ( .A(n5688), .B(n5689), .Z(n5680) );
  AND U5490 ( .A(n687), .B(n5690), .Z(n5689) );
  XNOR U5491 ( .A(n5691), .B(n5692), .Z(n5686) );
  AND U5492 ( .A(n679), .B(n5693), .Z(n5692) );
  XOR U5493 ( .A(p_input[1821]), .B(n5691), .Z(n5693) );
  XNOR U5494 ( .A(n5694), .B(n5695), .Z(n5691) );
  AND U5495 ( .A(n683), .B(n5690), .Z(n5695) );
  XNOR U5496 ( .A(n5694), .B(n5688), .Z(n5690) );
  XOR U5497 ( .A(n5696), .B(n5697), .Z(n5688) );
  AND U5498 ( .A(n698), .B(n5698), .Z(n5697) );
  XNOR U5499 ( .A(n5699), .B(n5700), .Z(n5694) );
  AND U5500 ( .A(n690), .B(n5701), .Z(n5700) );
  XOR U5501 ( .A(p_input[1853]), .B(n5699), .Z(n5701) );
  XNOR U5502 ( .A(n5702), .B(n5703), .Z(n5699) );
  AND U5503 ( .A(n694), .B(n5698), .Z(n5703) );
  XNOR U5504 ( .A(n5702), .B(n5696), .Z(n5698) );
  XOR U5505 ( .A(n5704), .B(n5705), .Z(n5696) );
  AND U5506 ( .A(n709), .B(n5706), .Z(n5705) );
  XNOR U5507 ( .A(n5707), .B(n5708), .Z(n5702) );
  AND U5508 ( .A(n701), .B(n5709), .Z(n5708) );
  XOR U5509 ( .A(p_input[1885]), .B(n5707), .Z(n5709) );
  XNOR U5510 ( .A(n5710), .B(n5711), .Z(n5707) );
  AND U5511 ( .A(n705), .B(n5706), .Z(n5711) );
  XNOR U5512 ( .A(n5710), .B(n5704), .Z(n5706) );
  XOR U5513 ( .A(n5712), .B(n5713), .Z(n5704) );
  AND U5514 ( .A(n720), .B(n5714), .Z(n5713) );
  XNOR U5515 ( .A(n5715), .B(n5716), .Z(n5710) );
  AND U5516 ( .A(n712), .B(n5717), .Z(n5716) );
  XOR U5517 ( .A(p_input[1917]), .B(n5715), .Z(n5717) );
  XNOR U5518 ( .A(n5718), .B(n5719), .Z(n5715) );
  AND U5519 ( .A(n716), .B(n5714), .Z(n5719) );
  XNOR U5520 ( .A(n5718), .B(n5712), .Z(n5714) );
  XOR U5521 ( .A(n5720), .B(n5721), .Z(n5712) );
  AND U5522 ( .A(n731), .B(n5722), .Z(n5721) );
  XNOR U5523 ( .A(n5723), .B(n5724), .Z(n5718) );
  AND U5524 ( .A(n723), .B(n5725), .Z(n5724) );
  XOR U5525 ( .A(p_input[1949]), .B(n5723), .Z(n5725) );
  XNOR U5526 ( .A(n5726), .B(n5727), .Z(n5723) );
  AND U5527 ( .A(n727), .B(n5722), .Z(n5727) );
  XNOR U5528 ( .A(n5726), .B(n5720), .Z(n5722) );
  XOR U5529 ( .A(\knn_comb_/min_val_out[0][29] ), .B(n5728), .Z(n5720) );
  AND U5530 ( .A(n741), .B(n5729), .Z(n5728) );
  XNOR U5531 ( .A(n5730), .B(n5731), .Z(n5726) );
  AND U5532 ( .A(n734), .B(n5732), .Z(n5731) );
  XOR U5533 ( .A(p_input[1981]), .B(n5730), .Z(n5732) );
  XNOR U5534 ( .A(n5733), .B(n5734), .Z(n5730) );
  AND U5535 ( .A(n738), .B(n5729), .Z(n5734) );
  XOR U5536 ( .A(\knn_comb_/min_val_out[0][29] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .Z(n5729) );
  XOR U5537 ( .A(n15), .B(n5735), .Z(o[28]) );
  AND U5538 ( .A(n58), .B(n5736), .Z(n15) );
  XOR U5539 ( .A(n16), .B(n5735), .Z(n5736) );
  XOR U5540 ( .A(n5737), .B(n5738), .Z(n5735) );
  AND U5541 ( .A(n70), .B(n5739), .Z(n5738) );
  XOR U5542 ( .A(n5740), .B(n5741), .Z(n16) );
  AND U5543 ( .A(n62), .B(n5742), .Z(n5741) );
  XOR U5544 ( .A(p_input[28]), .B(n5740), .Z(n5742) );
  XNOR U5545 ( .A(n5743), .B(n5744), .Z(n5740) );
  AND U5546 ( .A(n66), .B(n5739), .Z(n5744) );
  XNOR U5547 ( .A(n5743), .B(n5737), .Z(n5739) );
  XOR U5548 ( .A(n5745), .B(n5746), .Z(n5737) );
  AND U5549 ( .A(n82), .B(n5747), .Z(n5746) );
  XNOR U5550 ( .A(n5748), .B(n5749), .Z(n5743) );
  AND U5551 ( .A(n74), .B(n5750), .Z(n5749) );
  XOR U5552 ( .A(p_input[60]), .B(n5748), .Z(n5750) );
  XNOR U5553 ( .A(n5751), .B(n5752), .Z(n5748) );
  AND U5554 ( .A(n78), .B(n5747), .Z(n5752) );
  XNOR U5555 ( .A(n5751), .B(n5745), .Z(n5747) );
  XOR U5556 ( .A(n5753), .B(n5754), .Z(n5745) );
  AND U5557 ( .A(n93), .B(n5755), .Z(n5754) );
  XNOR U5558 ( .A(n5756), .B(n5757), .Z(n5751) );
  AND U5559 ( .A(n85), .B(n5758), .Z(n5757) );
  XOR U5560 ( .A(p_input[92]), .B(n5756), .Z(n5758) );
  XNOR U5561 ( .A(n5759), .B(n5760), .Z(n5756) );
  AND U5562 ( .A(n89), .B(n5755), .Z(n5760) );
  XNOR U5563 ( .A(n5759), .B(n5753), .Z(n5755) );
  XOR U5564 ( .A(n5761), .B(n5762), .Z(n5753) );
  AND U5565 ( .A(n104), .B(n5763), .Z(n5762) );
  XNOR U5566 ( .A(n5764), .B(n5765), .Z(n5759) );
  AND U5567 ( .A(n96), .B(n5766), .Z(n5765) );
  XOR U5568 ( .A(p_input[124]), .B(n5764), .Z(n5766) );
  XNOR U5569 ( .A(n5767), .B(n5768), .Z(n5764) );
  AND U5570 ( .A(n100), .B(n5763), .Z(n5768) );
  XNOR U5571 ( .A(n5767), .B(n5761), .Z(n5763) );
  XOR U5572 ( .A(n5769), .B(n5770), .Z(n5761) );
  AND U5573 ( .A(n115), .B(n5771), .Z(n5770) );
  XNOR U5574 ( .A(n5772), .B(n5773), .Z(n5767) );
  AND U5575 ( .A(n107), .B(n5774), .Z(n5773) );
  XOR U5576 ( .A(p_input[156]), .B(n5772), .Z(n5774) );
  XNOR U5577 ( .A(n5775), .B(n5776), .Z(n5772) );
  AND U5578 ( .A(n111), .B(n5771), .Z(n5776) );
  XNOR U5579 ( .A(n5775), .B(n5769), .Z(n5771) );
  XOR U5580 ( .A(n5777), .B(n5778), .Z(n5769) );
  AND U5581 ( .A(n126), .B(n5779), .Z(n5778) );
  XNOR U5582 ( .A(n5780), .B(n5781), .Z(n5775) );
  AND U5583 ( .A(n118), .B(n5782), .Z(n5781) );
  XOR U5584 ( .A(p_input[188]), .B(n5780), .Z(n5782) );
  XNOR U5585 ( .A(n5783), .B(n5784), .Z(n5780) );
  AND U5586 ( .A(n122), .B(n5779), .Z(n5784) );
  XNOR U5587 ( .A(n5783), .B(n5777), .Z(n5779) );
  XOR U5588 ( .A(n5785), .B(n5786), .Z(n5777) );
  AND U5589 ( .A(n137), .B(n5787), .Z(n5786) );
  XNOR U5590 ( .A(n5788), .B(n5789), .Z(n5783) );
  AND U5591 ( .A(n129), .B(n5790), .Z(n5789) );
  XOR U5592 ( .A(p_input[220]), .B(n5788), .Z(n5790) );
  XNOR U5593 ( .A(n5791), .B(n5792), .Z(n5788) );
  AND U5594 ( .A(n133), .B(n5787), .Z(n5792) );
  XNOR U5595 ( .A(n5791), .B(n5785), .Z(n5787) );
  XOR U5596 ( .A(n5793), .B(n5794), .Z(n5785) );
  AND U5597 ( .A(n148), .B(n5795), .Z(n5794) );
  XNOR U5598 ( .A(n5796), .B(n5797), .Z(n5791) );
  AND U5599 ( .A(n140), .B(n5798), .Z(n5797) );
  XOR U5600 ( .A(p_input[252]), .B(n5796), .Z(n5798) );
  XNOR U5601 ( .A(n5799), .B(n5800), .Z(n5796) );
  AND U5602 ( .A(n144), .B(n5795), .Z(n5800) );
  XNOR U5603 ( .A(n5799), .B(n5793), .Z(n5795) );
  XOR U5604 ( .A(n5801), .B(n5802), .Z(n5793) );
  AND U5605 ( .A(n159), .B(n5803), .Z(n5802) );
  XNOR U5606 ( .A(n5804), .B(n5805), .Z(n5799) );
  AND U5607 ( .A(n151), .B(n5806), .Z(n5805) );
  XOR U5608 ( .A(p_input[284]), .B(n5804), .Z(n5806) );
  XNOR U5609 ( .A(n5807), .B(n5808), .Z(n5804) );
  AND U5610 ( .A(n155), .B(n5803), .Z(n5808) );
  XNOR U5611 ( .A(n5807), .B(n5801), .Z(n5803) );
  XOR U5612 ( .A(n5809), .B(n5810), .Z(n5801) );
  AND U5613 ( .A(n170), .B(n5811), .Z(n5810) );
  XNOR U5614 ( .A(n5812), .B(n5813), .Z(n5807) );
  AND U5615 ( .A(n162), .B(n5814), .Z(n5813) );
  XOR U5616 ( .A(p_input[316]), .B(n5812), .Z(n5814) );
  XNOR U5617 ( .A(n5815), .B(n5816), .Z(n5812) );
  AND U5618 ( .A(n166), .B(n5811), .Z(n5816) );
  XNOR U5619 ( .A(n5815), .B(n5809), .Z(n5811) );
  XOR U5620 ( .A(n5817), .B(n5818), .Z(n5809) );
  AND U5621 ( .A(n181), .B(n5819), .Z(n5818) );
  XNOR U5622 ( .A(n5820), .B(n5821), .Z(n5815) );
  AND U5623 ( .A(n173), .B(n5822), .Z(n5821) );
  XOR U5624 ( .A(p_input[348]), .B(n5820), .Z(n5822) );
  XNOR U5625 ( .A(n5823), .B(n5824), .Z(n5820) );
  AND U5626 ( .A(n177), .B(n5819), .Z(n5824) );
  XNOR U5627 ( .A(n5823), .B(n5817), .Z(n5819) );
  XOR U5628 ( .A(n5825), .B(n5826), .Z(n5817) );
  AND U5629 ( .A(n192), .B(n5827), .Z(n5826) );
  XNOR U5630 ( .A(n5828), .B(n5829), .Z(n5823) );
  AND U5631 ( .A(n184), .B(n5830), .Z(n5829) );
  XOR U5632 ( .A(p_input[380]), .B(n5828), .Z(n5830) );
  XNOR U5633 ( .A(n5831), .B(n5832), .Z(n5828) );
  AND U5634 ( .A(n188), .B(n5827), .Z(n5832) );
  XNOR U5635 ( .A(n5831), .B(n5825), .Z(n5827) );
  XOR U5636 ( .A(n5833), .B(n5834), .Z(n5825) );
  AND U5637 ( .A(n203), .B(n5835), .Z(n5834) );
  XNOR U5638 ( .A(n5836), .B(n5837), .Z(n5831) );
  AND U5639 ( .A(n195), .B(n5838), .Z(n5837) );
  XOR U5640 ( .A(p_input[412]), .B(n5836), .Z(n5838) );
  XNOR U5641 ( .A(n5839), .B(n5840), .Z(n5836) );
  AND U5642 ( .A(n199), .B(n5835), .Z(n5840) );
  XNOR U5643 ( .A(n5839), .B(n5833), .Z(n5835) );
  XOR U5644 ( .A(n5841), .B(n5842), .Z(n5833) );
  AND U5645 ( .A(n214), .B(n5843), .Z(n5842) );
  XNOR U5646 ( .A(n5844), .B(n5845), .Z(n5839) );
  AND U5647 ( .A(n206), .B(n5846), .Z(n5845) );
  XOR U5648 ( .A(p_input[444]), .B(n5844), .Z(n5846) );
  XNOR U5649 ( .A(n5847), .B(n5848), .Z(n5844) );
  AND U5650 ( .A(n210), .B(n5843), .Z(n5848) );
  XNOR U5651 ( .A(n5847), .B(n5841), .Z(n5843) );
  XOR U5652 ( .A(n5849), .B(n5850), .Z(n5841) );
  AND U5653 ( .A(n225), .B(n5851), .Z(n5850) );
  XNOR U5654 ( .A(n5852), .B(n5853), .Z(n5847) );
  AND U5655 ( .A(n217), .B(n5854), .Z(n5853) );
  XOR U5656 ( .A(p_input[476]), .B(n5852), .Z(n5854) );
  XNOR U5657 ( .A(n5855), .B(n5856), .Z(n5852) );
  AND U5658 ( .A(n221), .B(n5851), .Z(n5856) );
  XNOR U5659 ( .A(n5855), .B(n5849), .Z(n5851) );
  XOR U5660 ( .A(n5857), .B(n5858), .Z(n5849) );
  AND U5661 ( .A(n236), .B(n5859), .Z(n5858) );
  XNOR U5662 ( .A(n5860), .B(n5861), .Z(n5855) );
  AND U5663 ( .A(n228), .B(n5862), .Z(n5861) );
  XOR U5664 ( .A(p_input[508]), .B(n5860), .Z(n5862) );
  XNOR U5665 ( .A(n5863), .B(n5864), .Z(n5860) );
  AND U5666 ( .A(n232), .B(n5859), .Z(n5864) );
  XNOR U5667 ( .A(n5863), .B(n5857), .Z(n5859) );
  XOR U5668 ( .A(n5865), .B(n5866), .Z(n5857) );
  AND U5669 ( .A(n247), .B(n5867), .Z(n5866) );
  XNOR U5670 ( .A(n5868), .B(n5869), .Z(n5863) );
  AND U5671 ( .A(n239), .B(n5870), .Z(n5869) );
  XOR U5672 ( .A(p_input[540]), .B(n5868), .Z(n5870) );
  XNOR U5673 ( .A(n5871), .B(n5872), .Z(n5868) );
  AND U5674 ( .A(n243), .B(n5867), .Z(n5872) );
  XNOR U5675 ( .A(n5871), .B(n5865), .Z(n5867) );
  XOR U5676 ( .A(n5873), .B(n5874), .Z(n5865) );
  AND U5677 ( .A(n258), .B(n5875), .Z(n5874) );
  XNOR U5678 ( .A(n5876), .B(n5877), .Z(n5871) );
  AND U5679 ( .A(n250), .B(n5878), .Z(n5877) );
  XOR U5680 ( .A(p_input[572]), .B(n5876), .Z(n5878) );
  XNOR U5681 ( .A(n5879), .B(n5880), .Z(n5876) );
  AND U5682 ( .A(n254), .B(n5875), .Z(n5880) );
  XNOR U5683 ( .A(n5879), .B(n5873), .Z(n5875) );
  XOR U5684 ( .A(n5881), .B(n5882), .Z(n5873) );
  AND U5685 ( .A(n269), .B(n5883), .Z(n5882) );
  XNOR U5686 ( .A(n5884), .B(n5885), .Z(n5879) );
  AND U5687 ( .A(n261), .B(n5886), .Z(n5885) );
  XOR U5688 ( .A(p_input[604]), .B(n5884), .Z(n5886) );
  XNOR U5689 ( .A(n5887), .B(n5888), .Z(n5884) );
  AND U5690 ( .A(n265), .B(n5883), .Z(n5888) );
  XNOR U5691 ( .A(n5887), .B(n5881), .Z(n5883) );
  XOR U5692 ( .A(n5889), .B(n5890), .Z(n5881) );
  AND U5693 ( .A(n280), .B(n5891), .Z(n5890) );
  XNOR U5694 ( .A(n5892), .B(n5893), .Z(n5887) );
  AND U5695 ( .A(n272), .B(n5894), .Z(n5893) );
  XOR U5696 ( .A(p_input[636]), .B(n5892), .Z(n5894) );
  XNOR U5697 ( .A(n5895), .B(n5896), .Z(n5892) );
  AND U5698 ( .A(n276), .B(n5891), .Z(n5896) );
  XNOR U5699 ( .A(n5895), .B(n5889), .Z(n5891) );
  XOR U5700 ( .A(n5897), .B(n5898), .Z(n5889) );
  AND U5701 ( .A(n291), .B(n5899), .Z(n5898) );
  XNOR U5702 ( .A(n5900), .B(n5901), .Z(n5895) );
  AND U5703 ( .A(n283), .B(n5902), .Z(n5901) );
  XOR U5704 ( .A(p_input[668]), .B(n5900), .Z(n5902) );
  XNOR U5705 ( .A(n5903), .B(n5904), .Z(n5900) );
  AND U5706 ( .A(n287), .B(n5899), .Z(n5904) );
  XNOR U5707 ( .A(n5903), .B(n5897), .Z(n5899) );
  XOR U5708 ( .A(n5905), .B(n5906), .Z(n5897) );
  AND U5709 ( .A(n302), .B(n5907), .Z(n5906) );
  XNOR U5710 ( .A(n5908), .B(n5909), .Z(n5903) );
  AND U5711 ( .A(n294), .B(n5910), .Z(n5909) );
  XOR U5712 ( .A(p_input[700]), .B(n5908), .Z(n5910) );
  XNOR U5713 ( .A(n5911), .B(n5912), .Z(n5908) );
  AND U5714 ( .A(n298), .B(n5907), .Z(n5912) );
  XNOR U5715 ( .A(n5911), .B(n5905), .Z(n5907) );
  XOR U5716 ( .A(n5913), .B(n5914), .Z(n5905) );
  AND U5717 ( .A(n313), .B(n5915), .Z(n5914) );
  XNOR U5718 ( .A(n5916), .B(n5917), .Z(n5911) );
  AND U5719 ( .A(n305), .B(n5918), .Z(n5917) );
  XOR U5720 ( .A(p_input[732]), .B(n5916), .Z(n5918) );
  XNOR U5721 ( .A(n5919), .B(n5920), .Z(n5916) );
  AND U5722 ( .A(n309), .B(n5915), .Z(n5920) );
  XNOR U5723 ( .A(n5919), .B(n5913), .Z(n5915) );
  XOR U5724 ( .A(n5921), .B(n5922), .Z(n5913) );
  AND U5725 ( .A(n324), .B(n5923), .Z(n5922) );
  XNOR U5726 ( .A(n5924), .B(n5925), .Z(n5919) );
  AND U5727 ( .A(n316), .B(n5926), .Z(n5925) );
  XOR U5728 ( .A(p_input[764]), .B(n5924), .Z(n5926) );
  XNOR U5729 ( .A(n5927), .B(n5928), .Z(n5924) );
  AND U5730 ( .A(n320), .B(n5923), .Z(n5928) );
  XNOR U5731 ( .A(n5927), .B(n5921), .Z(n5923) );
  XOR U5732 ( .A(n5929), .B(n5930), .Z(n5921) );
  AND U5733 ( .A(n335), .B(n5931), .Z(n5930) );
  XNOR U5734 ( .A(n5932), .B(n5933), .Z(n5927) );
  AND U5735 ( .A(n327), .B(n5934), .Z(n5933) );
  XOR U5736 ( .A(p_input[796]), .B(n5932), .Z(n5934) );
  XNOR U5737 ( .A(n5935), .B(n5936), .Z(n5932) );
  AND U5738 ( .A(n331), .B(n5931), .Z(n5936) );
  XNOR U5739 ( .A(n5935), .B(n5929), .Z(n5931) );
  XOR U5740 ( .A(n5937), .B(n5938), .Z(n5929) );
  AND U5741 ( .A(n346), .B(n5939), .Z(n5938) );
  XNOR U5742 ( .A(n5940), .B(n5941), .Z(n5935) );
  AND U5743 ( .A(n338), .B(n5942), .Z(n5941) );
  XOR U5744 ( .A(p_input[828]), .B(n5940), .Z(n5942) );
  XNOR U5745 ( .A(n5943), .B(n5944), .Z(n5940) );
  AND U5746 ( .A(n342), .B(n5939), .Z(n5944) );
  XNOR U5747 ( .A(n5943), .B(n5937), .Z(n5939) );
  XOR U5748 ( .A(n5945), .B(n5946), .Z(n5937) );
  AND U5749 ( .A(n357), .B(n5947), .Z(n5946) );
  XNOR U5750 ( .A(n5948), .B(n5949), .Z(n5943) );
  AND U5751 ( .A(n349), .B(n5950), .Z(n5949) );
  XOR U5752 ( .A(p_input[860]), .B(n5948), .Z(n5950) );
  XNOR U5753 ( .A(n5951), .B(n5952), .Z(n5948) );
  AND U5754 ( .A(n353), .B(n5947), .Z(n5952) );
  XNOR U5755 ( .A(n5951), .B(n5945), .Z(n5947) );
  XOR U5756 ( .A(n5953), .B(n5954), .Z(n5945) );
  AND U5757 ( .A(n368), .B(n5955), .Z(n5954) );
  XNOR U5758 ( .A(n5956), .B(n5957), .Z(n5951) );
  AND U5759 ( .A(n360), .B(n5958), .Z(n5957) );
  XOR U5760 ( .A(p_input[892]), .B(n5956), .Z(n5958) );
  XNOR U5761 ( .A(n5959), .B(n5960), .Z(n5956) );
  AND U5762 ( .A(n364), .B(n5955), .Z(n5960) );
  XNOR U5763 ( .A(n5959), .B(n5953), .Z(n5955) );
  XOR U5764 ( .A(n5961), .B(n5962), .Z(n5953) );
  AND U5765 ( .A(n379), .B(n5963), .Z(n5962) );
  XNOR U5766 ( .A(n5964), .B(n5965), .Z(n5959) );
  AND U5767 ( .A(n371), .B(n5966), .Z(n5965) );
  XOR U5768 ( .A(p_input[924]), .B(n5964), .Z(n5966) );
  XNOR U5769 ( .A(n5967), .B(n5968), .Z(n5964) );
  AND U5770 ( .A(n375), .B(n5963), .Z(n5968) );
  XNOR U5771 ( .A(n5967), .B(n5961), .Z(n5963) );
  XOR U5772 ( .A(n5969), .B(n5970), .Z(n5961) );
  AND U5773 ( .A(n390), .B(n5971), .Z(n5970) );
  XNOR U5774 ( .A(n5972), .B(n5973), .Z(n5967) );
  AND U5775 ( .A(n382), .B(n5974), .Z(n5973) );
  XOR U5776 ( .A(p_input[956]), .B(n5972), .Z(n5974) );
  XNOR U5777 ( .A(n5975), .B(n5976), .Z(n5972) );
  AND U5778 ( .A(n386), .B(n5971), .Z(n5976) );
  XNOR U5779 ( .A(n5975), .B(n5969), .Z(n5971) );
  XOR U5780 ( .A(n5977), .B(n5978), .Z(n5969) );
  AND U5781 ( .A(n401), .B(n5979), .Z(n5978) );
  XNOR U5782 ( .A(n5980), .B(n5981), .Z(n5975) );
  AND U5783 ( .A(n393), .B(n5982), .Z(n5981) );
  XOR U5784 ( .A(p_input[988]), .B(n5980), .Z(n5982) );
  XNOR U5785 ( .A(n5983), .B(n5984), .Z(n5980) );
  AND U5786 ( .A(n397), .B(n5979), .Z(n5984) );
  XNOR U5787 ( .A(n5983), .B(n5977), .Z(n5979) );
  XOR U5788 ( .A(n5985), .B(n5986), .Z(n5977) );
  AND U5789 ( .A(n412), .B(n5987), .Z(n5986) );
  XNOR U5790 ( .A(n5988), .B(n5989), .Z(n5983) );
  AND U5791 ( .A(n404), .B(n5990), .Z(n5989) );
  XOR U5792 ( .A(p_input[1020]), .B(n5988), .Z(n5990) );
  XNOR U5793 ( .A(n5991), .B(n5992), .Z(n5988) );
  AND U5794 ( .A(n408), .B(n5987), .Z(n5992) );
  XNOR U5795 ( .A(n5991), .B(n5985), .Z(n5987) );
  XOR U5796 ( .A(n5993), .B(n5994), .Z(n5985) );
  AND U5797 ( .A(n423), .B(n5995), .Z(n5994) );
  XNOR U5798 ( .A(n5996), .B(n5997), .Z(n5991) );
  AND U5799 ( .A(n415), .B(n5998), .Z(n5997) );
  XOR U5800 ( .A(p_input[1052]), .B(n5996), .Z(n5998) );
  XNOR U5801 ( .A(n5999), .B(n6000), .Z(n5996) );
  AND U5802 ( .A(n419), .B(n5995), .Z(n6000) );
  XNOR U5803 ( .A(n5999), .B(n5993), .Z(n5995) );
  XOR U5804 ( .A(n6001), .B(n6002), .Z(n5993) );
  AND U5805 ( .A(n434), .B(n6003), .Z(n6002) );
  XNOR U5806 ( .A(n6004), .B(n6005), .Z(n5999) );
  AND U5807 ( .A(n426), .B(n6006), .Z(n6005) );
  XOR U5808 ( .A(p_input[1084]), .B(n6004), .Z(n6006) );
  XNOR U5809 ( .A(n6007), .B(n6008), .Z(n6004) );
  AND U5810 ( .A(n430), .B(n6003), .Z(n6008) );
  XNOR U5811 ( .A(n6007), .B(n6001), .Z(n6003) );
  XOR U5812 ( .A(n6009), .B(n6010), .Z(n6001) );
  AND U5813 ( .A(n445), .B(n6011), .Z(n6010) );
  XNOR U5814 ( .A(n6012), .B(n6013), .Z(n6007) );
  AND U5815 ( .A(n437), .B(n6014), .Z(n6013) );
  XOR U5816 ( .A(p_input[1116]), .B(n6012), .Z(n6014) );
  XNOR U5817 ( .A(n6015), .B(n6016), .Z(n6012) );
  AND U5818 ( .A(n441), .B(n6011), .Z(n6016) );
  XNOR U5819 ( .A(n6015), .B(n6009), .Z(n6011) );
  XOR U5820 ( .A(n6017), .B(n6018), .Z(n6009) );
  AND U5821 ( .A(n456), .B(n6019), .Z(n6018) );
  XNOR U5822 ( .A(n6020), .B(n6021), .Z(n6015) );
  AND U5823 ( .A(n448), .B(n6022), .Z(n6021) );
  XOR U5824 ( .A(p_input[1148]), .B(n6020), .Z(n6022) );
  XNOR U5825 ( .A(n6023), .B(n6024), .Z(n6020) );
  AND U5826 ( .A(n452), .B(n6019), .Z(n6024) );
  XNOR U5827 ( .A(n6023), .B(n6017), .Z(n6019) );
  XOR U5828 ( .A(n6025), .B(n6026), .Z(n6017) );
  AND U5829 ( .A(n467), .B(n6027), .Z(n6026) );
  XNOR U5830 ( .A(n6028), .B(n6029), .Z(n6023) );
  AND U5831 ( .A(n459), .B(n6030), .Z(n6029) );
  XOR U5832 ( .A(p_input[1180]), .B(n6028), .Z(n6030) );
  XNOR U5833 ( .A(n6031), .B(n6032), .Z(n6028) );
  AND U5834 ( .A(n463), .B(n6027), .Z(n6032) );
  XNOR U5835 ( .A(n6031), .B(n6025), .Z(n6027) );
  XOR U5836 ( .A(n6033), .B(n6034), .Z(n6025) );
  AND U5837 ( .A(n478), .B(n6035), .Z(n6034) );
  XNOR U5838 ( .A(n6036), .B(n6037), .Z(n6031) );
  AND U5839 ( .A(n470), .B(n6038), .Z(n6037) );
  XOR U5840 ( .A(p_input[1212]), .B(n6036), .Z(n6038) );
  XNOR U5841 ( .A(n6039), .B(n6040), .Z(n6036) );
  AND U5842 ( .A(n474), .B(n6035), .Z(n6040) );
  XNOR U5843 ( .A(n6039), .B(n6033), .Z(n6035) );
  XOR U5844 ( .A(n6041), .B(n6042), .Z(n6033) );
  AND U5845 ( .A(n489), .B(n6043), .Z(n6042) );
  XNOR U5846 ( .A(n6044), .B(n6045), .Z(n6039) );
  AND U5847 ( .A(n481), .B(n6046), .Z(n6045) );
  XOR U5848 ( .A(p_input[1244]), .B(n6044), .Z(n6046) );
  XNOR U5849 ( .A(n6047), .B(n6048), .Z(n6044) );
  AND U5850 ( .A(n485), .B(n6043), .Z(n6048) );
  XNOR U5851 ( .A(n6047), .B(n6041), .Z(n6043) );
  XOR U5852 ( .A(n6049), .B(n6050), .Z(n6041) );
  AND U5853 ( .A(n500), .B(n6051), .Z(n6050) );
  XNOR U5854 ( .A(n6052), .B(n6053), .Z(n6047) );
  AND U5855 ( .A(n492), .B(n6054), .Z(n6053) );
  XOR U5856 ( .A(p_input[1276]), .B(n6052), .Z(n6054) );
  XNOR U5857 ( .A(n6055), .B(n6056), .Z(n6052) );
  AND U5858 ( .A(n496), .B(n6051), .Z(n6056) );
  XNOR U5859 ( .A(n6055), .B(n6049), .Z(n6051) );
  XOR U5860 ( .A(n6057), .B(n6058), .Z(n6049) );
  AND U5861 ( .A(n511), .B(n6059), .Z(n6058) );
  XNOR U5862 ( .A(n6060), .B(n6061), .Z(n6055) );
  AND U5863 ( .A(n503), .B(n6062), .Z(n6061) );
  XOR U5864 ( .A(p_input[1308]), .B(n6060), .Z(n6062) );
  XNOR U5865 ( .A(n6063), .B(n6064), .Z(n6060) );
  AND U5866 ( .A(n507), .B(n6059), .Z(n6064) );
  XNOR U5867 ( .A(n6063), .B(n6057), .Z(n6059) );
  XOR U5868 ( .A(n6065), .B(n6066), .Z(n6057) );
  AND U5869 ( .A(n522), .B(n6067), .Z(n6066) );
  XNOR U5870 ( .A(n6068), .B(n6069), .Z(n6063) );
  AND U5871 ( .A(n514), .B(n6070), .Z(n6069) );
  XOR U5872 ( .A(p_input[1340]), .B(n6068), .Z(n6070) );
  XNOR U5873 ( .A(n6071), .B(n6072), .Z(n6068) );
  AND U5874 ( .A(n518), .B(n6067), .Z(n6072) );
  XNOR U5875 ( .A(n6071), .B(n6065), .Z(n6067) );
  XOR U5876 ( .A(n6073), .B(n6074), .Z(n6065) );
  AND U5877 ( .A(n533), .B(n6075), .Z(n6074) );
  XNOR U5878 ( .A(n6076), .B(n6077), .Z(n6071) );
  AND U5879 ( .A(n525), .B(n6078), .Z(n6077) );
  XOR U5880 ( .A(p_input[1372]), .B(n6076), .Z(n6078) );
  XNOR U5881 ( .A(n6079), .B(n6080), .Z(n6076) );
  AND U5882 ( .A(n529), .B(n6075), .Z(n6080) );
  XNOR U5883 ( .A(n6079), .B(n6073), .Z(n6075) );
  XOR U5884 ( .A(n6081), .B(n6082), .Z(n6073) );
  AND U5885 ( .A(n544), .B(n6083), .Z(n6082) );
  XNOR U5886 ( .A(n6084), .B(n6085), .Z(n6079) );
  AND U5887 ( .A(n536), .B(n6086), .Z(n6085) );
  XOR U5888 ( .A(p_input[1404]), .B(n6084), .Z(n6086) );
  XNOR U5889 ( .A(n6087), .B(n6088), .Z(n6084) );
  AND U5890 ( .A(n540), .B(n6083), .Z(n6088) );
  XNOR U5891 ( .A(n6087), .B(n6081), .Z(n6083) );
  XOR U5892 ( .A(n6089), .B(n6090), .Z(n6081) );
  AND U5893 ( .A(n555), .B(n6091), .Z(n6090) );
  XNOR U5894 ( .A(n6092), .B(n6093), .Z(n6087) );
  AND U5895 ( .A(n547), .B(n6094), .Z(n6093) );
  XOR U5896 ( .A(p_input[1436]), .B(n6092), .Z(n6094) );
  XNOR U5897 ( .A(n6095), .B(n6096), .Z(n6092) );
  AND U5898 ( .A(n551), .B(n6091), .Z(n6096) );
  XNOR U5899 ( .A(n6095), .B(n6089), .Z(n6091) );
  XOR U5900 ( .A(n6097), .B(n6098), .Z(n6089) );
  AND U5901 ( .A(n566), .B(n6099), .Z(n6098) );
  XNOR U5902 ( .A(n6100), .B(n6101), .Z(n6095) );
  AND U5903 ( .A(n558), .B(n6102), .Z(n6101) );
  XOR U5904 ( .A(p_input[1468]), .B(n6100), .Z(n6102) );
  XNOR U5905 ( .A(n6103), .B(n6104), .Z(n6100) );
  AND U5906 ( .A(n562), .B(n6099), .Z(n6104) );
  XNOR U5907 ( .A(n6103), .B(n6097), .Z(n6099) );
  XOR U5908 ( .A(n6105), .B(n6106), .Z(n6097) );
  AND U5909 ( .A(n577), .B(n6107), .Z(n6106) );
  XNOR U5910 ( .A(n6108), .B(n6109), .Z(n6103) );
  AND U5911 ( .A(n569), .B(n6110), .Z(n6109) );
  XOR U5912 ( .A(p_input[1500]), .B(n6108), .Z(n6110) );
  XNOR U5913 ( .A(n6111), .B(n6112), .Z(n6108) );
  AND U5914 ( .A(n573), .B(n6107), .Z(n6112) );
  XNOR U5915 ( .A(n6111), .B(n6105), .Z(n6107) );
  XOR U5916 ( .A(n6113), .B(n6114), .Z(n6105) );
  AND U5917 ( .A(n588), .B(n6115), .Z(n6114) );
  XNOR U5918 ( .A(n6116), .B(n6117), .Z(n6111) );
  AND U5919 ( .A(n580), .B(n6118), .Z(n6117) );
  XOR U5920 ( .A(p_input[1532]), .B(n6116), .Z(n6118) );
  XNOR U5921 ( .A(n6119), .B(n6120), .Z(n6116) );
  AND U5922 ( .A(n584), .B(n6115), .Z(n6120) );
  XNOR U5923 ( .A(n6119), .B(n6113), .Z(n6115) );
  XOR U5924 ( .A(n6121), .B(n6122), .Z(n6113) );
  AND U5925 ( .A(n599), .B(n6123), .Z(n6122) );
  XNOR U5926 ( .A(n6124), .B(n6125), .Z(n6119) );
  AND U5927 ( .A(n591), .B(n6126), .Z(n6125) );
  XOR U5928 ( .A(p_input[1564]), .B(n6124), .Z(n6126) );
  XNOR U5929 ( .A(n6127), .B(n6128), .Z(n6124) );
  AND U5930 ( .A(n595), .B(n6123), .Z(n6128) );
  XNOR U5931 ( .A(n6127), .B(n6121), .Z(n6123) );
  XOR U5932 ( .A(n6129), .B(n6130), .Z(n6121) );
  AND U5933 ( .A(n610), .B(n6131), .Z(n6130) );
  XNOR U5934 ( .A(n6132), .B(n6133), .Z(n6127) );
  AND U5935 ( .A(n602), .B(n6134), .Z(n6133) );
  XOR U5936 ( .A(p_input[1596]), .B(n6132), .Z(n6134) );
  XNOR U5937 ( .A(n6135), .B(n6136), .Z(n6132) );
  AND U5938 ( .A(n606), .B(n6131), .Z(n6136) );
  XNOR U5939 ( .A(n6135), .B(n6129), .Z(n6131) );
  XOR U5940 ( .A(n6137), .B(n6138), .Z(n6129) );
  AND U5941 ( .A(n621), .B(n6139), .Z(n6138) );
  XNOR U5942 ( .A(n6140), .B(n6141), .Z(n6135) );
  AND U5943 ( .A(n613), .B(n6142), .Z(n6141) );
  XOR U5944 ( .A(p_input[1628]), .B(n6140), .Z(n6142) );
  XNOR U5945 ( .A(n6143), .B(n6144), .Z(n6140) );
  AND U5946 ( .A(n617), .B(n6139), .Z(n6144) );
  XNOR U5947 ( .A(n6143), .B(n6137), .Z(n6139) );
  XOR U5948 ( .A(n6145), .B(n6146), .Z(n6137) );
  AND U5949 ( .A(n632), .B(n6147), .Z(n6146) );
  XNOR U5950 ( .A(n6148), .B(n6149), .Z(n6143) );
  AND U5951 ( .A(n624), .B(n6150), .Z(n6149) );
  XOR U5952 ( .A(p_input[1660]), .B(n6148), .Z(n6150) );
  XNOR U5953 ( .A(n6151), .B(n6152), .Z(n6148) );
  AND U5954 ( .A(n628), .B(n6147), .Z(n6152) );
  XNOR U5955 ( .A(n6151), .B(n6145), .Z(n6147) );
  XOR U5956 ( .A(n6153), .B(n6154), .Z(n6145) );
  AND U5957 ( .A(n643), .B(n6155), .Z(n6154) );
  XNOR U5958 ( .A(n6156), .B(n6157), .Z(n6151) );
  AND U5959 ( .A(n635), .B(n6158), .Z(n6157) );
  XOR U5960 ( .A(p_input[1692]), .B(n6156), .Z(n6158) );
  XNOR U5961 ( .A(n6159), .B(n6160), .Z(n6156) );
  AND U5962 ( .A(n639), .B(n6155), .Z(n6160) );
  XNOR U5963 ( .A(n6159), .B(n6153), .Z(n6155) );
  XOR U5964 ( .A(n6161), .B(n6162), .Z(n6153) );
  AND U5965 ( .A(n654), .B(n6163), .Z(n6162) );
  XNOR U5966 ( .A(n6164), .B(n6165), .Z(n6159) );
  AND U5967 ( .A(n646), .B(n6166), .Z(n6165) );
  XOR U5968 ( .A(p_input[1724]), .B(n6164), .Z(n6166) );
  XNOR U5969 ( .A(n6167), .B(n6168), .Z(n6164) );
  AND U5970 ( .A(n650), .B(n6163), .Z(n6168) );
  XNOR U5971 ( .A(n6167), .B(n6161), .Z(n6163) );
  XOR U5972 ( .A(n6169), .B(n6170), .Z(n6161) );
  AND U5973 ( .A(n665), .B(n6171), .Z(n6170) );
  XNOR U5974 ( .A(n6172), .B(n6173), .Z(n6167) );
  AND U5975 ( .A(n657), .B(n6174), .Z(n6173) );
  XOR U5976 ( .A(p_input[1756]), .B(n6172), .Z(n6174) );
  XNOR U5977 ( .A(n6175), .B(n6176), .Z(n6172) );
  AND U5978 ( .A(n661), .B(n6171), .Z(n6176) );
  XNOR U5979 ( .A(n6175), .B(n6169), .Z(n6171) );
  XOR U5980 ( .A(n6177), .B(n6178), .Z(n6169) );
  AND U5981 ( .A(n676), .B(n6179), .Z(n6178) );
  XNOR U5982 ( .A(n6180), .B(n6181), .Z(n6175) );
  AND U5983 ( .A(n668), .B(n6182), .Z(n6181) );
  XOR U5984 ( .A(p_input[1788]), .B(n6180), .Z(n6182) );
  XNOR U5985 ( .A(n6183), .B(n6184), .Z(n6180) );
  AND U5986 ( .A(n672), .B(n6179), .Z(n6184) );
  XNOR U5987 ( .A(n6183), .B(n6177), .Z(n6179) );
  XOR U5988 ( .A(n6185), .B(n6186), .Z(n6177) );
  AND U5989 ( .A(n687), .B(n6187), .Z(n6186) );
  XNOR U5990 ( .A(n6188), .B(n6189), .Z(n6183) );
  AND U5991 ( .A(n679), .B(n6190), .Z(n6189) );
  XOR U5992 ( .A(p_input[1820]), .B(n6188), .Z(n6190) );
  XNOR U5993 ( .A(n6191), .B(n6192), .Z(n6188) );
  AND U5994 ( .A(n683), .B(n6187), .Z(n6192) );
  XNOR U5995 ( .A(n6191), .B(n6185), .Z(n6187) );
  XOR U5996 ( .A(n6193), .B(n6194), .Z(n6185) );
  AND U5997 ( .A(n698), .B(n6195), .Z(n6194) );
  XNOR U5998 ( .A(n6196), .B(n6197), .Z(n6191) );
  AND U5999 ( .A(n690), .B(n6198), .Z(n6197) );
  XOR U6000 ( .A(p_input[1852]), .B(n6196), .Z(n6198) );
  XNOR U6001 ( .A(n6199), .B(n6200), .Z(n6196) );
  AND U6002 ( .A(n694), .B(n6195), .Z(n6200) );
  XNOR U6003 ( .A(n6199), .B(n6193), .Z(n6195) );
  XOR U6004 ( .A(n6201), .B(n6202), .Z(n6193) );
  AND U6005 ( .A(n709), .B(n6203), .Z(n6202) );
  XNOR U6006 ( .A(n6204), .B(n6205), .Z(n6199) );
  AND U6007 ( .A(n701), .B(n6206), .Z(n6205) );
  XOR U6008 ( .A(p_input[1884]), .B(n6204), .Z(n6206) );
  XNOR U6009 ( .A(n6207), .B(n6208), .Z(n6204) );
  AND U6010 ( .A(n705), .B(n6203), .Z(n6208) );
  XNOR U6011 ( .A(n6207), .B(n6201), .Z(n6203) );
  XOR U6012 ( .A(n6209), .B(n6210), .Z(n6201) );
  AND U6013 ( .A(n720), .B(n6211), .Z(n6210) );
  XNOR U6014 ( .A(n6212), .B(n6213), .Z(n6207) );
  AND U6015 ( .A(n712), .B(n6214), .Z(n6213) );
  XOR U6016 ( .A(p_input[1916]), .B(n6212), .Z(n6214) );
  XNOR U6017 ( .A(n6215), .B(n6216), .Z(n6212) );
  AND U6018 ( .A(n716), .B(n6211), .Z(n6216) );
  XNOR U6019 ( .A(n6215), .B(n6209), .Z(n6211) );
  XOR U6020 ( .A(n6217), .B(n6218), .Z(n6209) );
  AND U6021 ( .A(n731), .B(n6219), .Z(n6218) );
  XNOR U6022 ( .A(n6220), .B(n6221), .Z(n6215) );
  AND U6023 ( .A(n723), .B(n6222), .Z(n6221) );
  XOR U6024 ( .A(p_input[1948]), .B(n6220), .Z(n6222) );
  XNOR U6025 ( .A(n6223), .B(n6224), .Z(n6220) );
  AND U6026 ( .A(n727), .B(n6219), .Z(n6224) );
  XNOR U6027 ( .A(n6223), .B(n6217), .Z(n6219) );
  XOR U6028 ( .A(\knn_comb_/min_val_out[0][28] ), .B(n6225), .Z(n6217) );
  AND U6029 ( .A(n741), .B(n6226), .Z(n6225) );
  XNOR U6030 ( .A(n6227), .B(n6228), .Z(n6223) );
  AND U6031 ( .A(n734), .B(n6229), .Z(n6228) );
  XOR U6032 ( .A(p_input[1980]), .B(n6227), .Z(n6229) );
  XNOR U6033 ( .A(n6230), .B(n6231), .Z(n6227) );
  AND U6034 ( .A(n738), .B(n6226), .Z(n6231) );
  XOR U6035 ( .A(\knn_comb_/min_val_out[0][28] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .Z(n6226) );
  XOR U6036 ( .A(n19), .B(n6232), .Z(o[27]) );
  AND U6037 ( .A(n58), .B(n6233), .Z(n19) );
  XOR U6038 ( .A(n20), .B(n6232), .Z(n6233) );
  XOR U6039 ( .A(n6234), .B(n6235), .Z(n6232) );
  AND U6040 ( .A(n70), .B(n6236), .Z(n6235) );
  XOR U6041 ( .A(n6237), .B(n6238), .Z(n20) );
  AND U6042 ( .A(n62), .B(n6239), .Z(n6238) );
  XOR U6043 ( .A(p_input[27]), .B(n6237), .Z(n6239) );
  XNOR U6044 ( .A(n6240), .B(n6241), .Z(n6237) );
  AND U6045 ( .A(n66), .B(n6236), .Z(n6241) );
  XNOR U6046 ( .A(n6240), .B(n6234), .Z(n6236) );
  XOR U6047 ( .A(n6242), .B(n6243), .Z(n6234) );
  AND U6048 ( .A(n82), .B(n6244), .Z(n6243) );
  XNOR U6049 ( .A(n6245), .B(n6246), .Z(n6240) );
  AND U6050 ( .A(n74), .B(n6247), .Z(n6246) );
  XOR U6051 ( .A(p_input[59]), .B(n6245), .Z(n6247) );
  XNOR U6052 ( .A(n6248), .B(n6249), .Z(n6245) );
  AND U6053 ( .A(n78), .B(n6244), .Z(n6249) );
  XNOR U6054 ( .A(n6248), .B(n6242), .Z(n6244) );
  XOR U6055 ( .A(n6250), .B(n6251), .Z(n6242) );
  AND U6056 ( .A(n93), .B(n6252), .Z(n6251) );
  XNOR U6057 ( .A(n6253), .B(n6254), .Z(n6248) );
  AND U6058 ( .A(n85), .B(n6255), .Z(n6254) );
  XOR U6059 ( .A(p_input[91]), .B(n6253), .Z(n6255) );
  XNOR U6060 ( .A(n6256), .B(n6257), .Z(n6253) );
  AND U6061 ( .A(n89), .B(n6252), .Z(n6257) );
  XNOR U6062 ( .A(n6256), .B(n6250), .Z(n6252) );
  XOR U6063 ( .A(n6258), .B(n6259), .Z(n6250) );
  AND U6064 ( .A(n104), .B(n6260), .Z(n6259) );
  XNOR U6065 ( .A(n6261), .B(n6262), .Z(n6256) );
  AND U6066 ( .A(n96), .B(n6263), .Z(n6262) );
  XOR U6067 ( .A(p_input[123]), .B(n6261), .Z(n6263) );
  XNOR U6068 ( .A(n6264), .B(n6265), .Z(n6261) );
  AND U6069 ( .A(n100), .B(n6260), .Z(n6265) );
  XNOR U6070 ( .A(n6264), .B(n6258), .Z(n6260) );
  XOR U6071 ( .A(n6266), .B(n6267), .Z(n6258) );
  AND U6072 ( .A(n115), .B(n6268), .Z(n6267) );
  XNOR U6073 ( .A(n6269), .B(n6270), .Z(n6264) );
  AND U6074 ( .A(n107), .B(n6271), .Z(n6270) );
  XOR U6075 ( .A(p_input[155]), .B(n6269), .Z(n6271) );
  XNOR U6076 ( .A(n6272), .B(n6273), .Z(n6269) );
  AND U6077 ( .A(n111), .B(n6268), .Z(n6273) );
  XNOR U6078 ( .A(n6272), .B(n6266), .Z(n6268) );
  XOR U6079 ( .A(n6274), .B(n6275), .Z(n6266) );
  AND U6080 ( .A(n126), .B(n6276), .Z(n6275) );
  XNOR U6081 ( .A(n6277), .B(n6278), .Z(n6272) );
  AND U6082 ( .A(n118), .B(n6279), .Z(n6278) );
  XOR U6083 ( .A(p_input[187]), .B(n6277), .Z(n6279) );
  XNOR U6084 ( .A(n6280), .B(n6281), .Z(n6277) );
  AND U6085 ( .A(n122), .B(n6276), .Z(n6281) );
  XNOR U6086 ( .A(n6280), .B(n6274), .Z(n6276) );
  XOR U6087 ( .A(n6282), .B(n6283), .Z(n6274) );
  AND U6088 ( .A(n137), .B(n6284), .Z(n6283) );
  XNOR U6089 ( .A(n6285), .B(n6286), .Z(n6280) );
  AND U6090 ( .A(n129), .B(n6287), .Z(n6286) );
  XOR U6091 ( .A(p_input[219]), .B(n6285), .Z(n6287) );
  XNOR U6092 ( .A(n6288), .B(n6289), .Z(n6285) );
  AND U6093 ( .A(n133), .B(n6284), .Z(n6289) );
  XNOR U6094 ( .A(n6288), .B(n6282), .Z(n6284) );
  XOR U6095 ( .A(n6290), .B(n6291), .Z(n6282) );
  AND U6096 ( .A(n148), .B(n6292), .Z(n6291) );
  XNOR U6097 ( .A(n6293), .B(n6294), .Z(n6288) );
  AND U6098 ( .A(n140), .B(n6295), .Z(n6294) );
  XOR U6099 ( .A(p_input[251]), .B(n6293), .Z(n6295) );
  XNOR U6100 ( .A(n6296), .B(n6297), .Z(n6293) );
  AND U6101 ( .A(n144), .B(n6292), .Z(n6297) );
  XNOR U6102 ( .A(n6296), .B(n6290), .Z(n6292) );
  XOR U6103 ( .A(n6298), .B(n6299), .Z(n6290) );
  AND U6104 ( .A(n159), .B(n6300), .Z(n6299) );
  XNOR U6105 ( .A(n6301), .B(n6302), .Z(n6296) );
  AND U6106 ( .A(n151), .B(n6303), .Z(n6302) );
  XOR U6107 ( .A(p_input[283]), .B(n6301), .Z(n6303) );
  XNOR U6108 ( .A(n6304), .B(n6305), .Z(n6301) );
  AND U6109 ( .A(n155), .B(n6300), .Z(n6305) );
  XNOR U6110 ( .A(n6304), .B(n6298), .Z(n6300) );
  XOR U6111 ( .A(n6306), .B(n6307), .Z(n6298) );
  AND U6112 ( .A(n170), .B(n6308), .Z(n6307) );
  XNOR U6113 ( .A(n6309), .B(n6310), .Z(n6304) );
  AND U6114 ( .A(n162), .B(n6311), .Z(n6310) );
  XOR U6115 ( .A(p_input[315]), .B(n6309), .Z(n6311) );
  XNOR U6116 ( .A(n6312), .B(n6313), .Z(n6309) );
  AND U6117 ( .A(n166), .B(n6308), .Z(n6313) );
  XNOR U6118 ( .A(n6312), .B(n6306), .Z(n6308) );
  XOR U6119 ( .A(n6314), .B(n6315), .Z(n6306) );
  AND U6120 ( .A(n181), .B(n6316), .Z(n6315) );
  XNOR U6121 ( .A(n6317), .B(n6318), .Z(n6312) );
  AND U6122 ( .A(n173), .B(n6319), .Z(n6318) );
  XOR U6123 ( .A(p_input[347]), .B(n6317), .Z(n6319) );
  XNOR U6124 ( .A(n6320), .B(n6321), .Z(n6317) );
  AND U6125 ( .A(n177), .B(n6316), .Z(n6321) );
  XNOR U6126 ( .A(n6320), .B(n6314), .Z(n6316) );
  XOR U6127 ( .A(n6322), .B(n6323), .Z(n6314) );
  AND U6128 ( .A(n192), .B(n6324), .Z(n6323) );
  XNOR U6129 ( .A(n6325), .B(n6326), .Z(n6320) );
  AND U6130 ( .A(n184), .B(n6327), .Z(n6326) );
  XOR U6131 ( .A(p_input[379]), .B(n6325), .Z(n6327) );
  XNOR U6132 ( .A(n6328), .B(n6329), .Z(n6325) );
  AND U6133 ( .A(n188), .B(n6324), .Z(n6329) );
  XNOR U6134 ( .A(n6328), .B(n6322), .Z(n6324) );
  XOR U6135 ( .A(n6330), .B(n6331), .Z(n6322) );
  AND U6136 ( .A(n203), .B(n6332), .Z(n6331) );
  XNOR U6137 ( .A(n6333), .B(n6334), .Z(n6328) );
  AND U6138 ( .A(n195), .B(n6335), .Z(n6334) );
  XOR U6139 ( .A(p_input[411]), .B(n6333), .Z(n6335) );
  XNOR U6140 ( .A(n6336), .B(n6337), .Z(n6333) );
  AND U6141 ( .A(n199), .B(n6332), .Z(n6337) );
  XNOR U6142 ( .A(n6336), .B(n6330), .Z(n6332) );
  XOR U6143 ( .A(n6338), .B(n6339), .Z(n6330) );
  AND U6144 ( .A(n214), .B(n6340), .Z(n6339) );
  XNOR U6145 ( .A(n6341), .B(n6342), .Z(n6336) );
  AND U6146 ( .A(n206), .B(n6343), .Z(n6342) );
  XOR U6147 ( .A(p_input[443]), .B(n6341), .Z(n6343) );
  XNOR U6148 ( .A(n6344), .B(n6345), .Z(n6341) );
  AND U6149 ( .A(n210), .B(n6340), .Z(n6345) );
  XNOR U6150 ( .A(n6344), .B(n6338), .Z(n6340) );
  XOR U6151 ( .A(n6346), .B(n6347), .Z(n6338) );
  AND U6152 ( .A(n225), .B(n6348), .Z(n6347) );
  XNOR U6153 ( .A(n6349), .B(n6350), .Z(n6344) );
  AND U6154 ( .A(n217), .B(n6351), .Z(n6350) );
  XOR U6155 ( .A(p_input[475]), .B(n6349), .Z(n6351) );
  XNOR U6156 ( .A(n6352), .B(n6353), .Z(n6349) );
  AND U6157 ( .A(n221), .B(n6348), .Z(n6353) );
  XNOR U6158 ( .A(n6352), .B(n6346), .Z(n6348) );
  XOR U6159 ( .A(n6354), .B(n6355), .Z(n6346) );
  AND U6160 ( .A(n236), .B(n6356), .Z(n6355) );
  XNOR U6161 ( .A(n6357), .B(n6358), .Z(n6352) );
  AND U6162 ( .A(n228), .B(n6359), .Z(n6358) );
  XOR U6163 ( .A(p_input[507]), .B(n6357), .Z(n6359) );
  XNOR U6164 ( .A(n6360), .B(n6361), .Z(n6357) );
  AND U6165 ( .A(n232), .B(n6356), .Z(n6361) );
  XNOR U6166 ( .A(n6360), .B(n6354), .Z(n6356) );
  XOR U6167 ( .A(n6362), .B(n6363), .Z(n6354) );
  AND U6168 ( .A(n247), .B(n6364), .Z(n6363) );
  XNOR U6169 ( .A(n6365), .B(n6366), .Z(n6360) );
  AND U6170 ( .A(n239), .B(n6367), .Z(n6366) );
  XOR U6171 ( .A(p_input[539]), .B(n6365), .Z(n6367) );
  XNOR U6172 ( .A(n6368), .B(n6369), .Z(n6365) );
  AND U6173 ( .A(n243), .B(n6364), .Z(n6369) );
  XNOR U6174 ( .A(n6368), .B(n6362), .Z(n6364) );
  XOR U6175 ( .A(n6370), .B(n6371), .Z(n6362) );
  AND U6176 ( .A(n258), .B(n6372), .Z(n6371) );
  XNOR U6177 ( .A(n6373), .B(n6374), .Z(n6368) );
  AND U6178 ( .A(n250), .B(n6375), .Z(n6374) );
  XOR U6179 ( .A(p_input[571]), .B(n6373), .Z(n6375) );
  XNOR U6180 ( .A(n6376), .B(n6377), .Z(n6373) );
  AND U6181 ( .A(n254), .B(n6372), .Z(n6377) );
  XNOR U6182 ( .A(n6376), .B(n6370), .Z(n6372) );
  XOR U6183 ( .A(n6378), .B(n6379), .Z(n6370) );
  AND U6184 ( .A(n269), .B(n6380), .Z(n6379) );
  XNOR U6185 ( .A(n6381), .B(n6382), .Z(n6376) );
  AND U6186 ( .A(n261), .B(n6383), .Z(n6382) );
  XOR U6187 ( .A(p_input[603]), .B(n6381), .Z(n6383) );
  XNOR U6188 ( .A(n6384), .B(n6385), .Z(n6381) );
  AND U6189 ( .A(n265), .B(n6380), .Z(n6385) );
  XNOR U6190 ( .A(n6384), .B(n6378), .Z(n6380) );
  XOR U6191 ( .A(n6386), .B(n6387), .Z(n6378) );
  AND U6192 ( .A(n280), .B(n6388), .Z(n6387) );
  XNOR U6193 ( .A(n6389), .B(n6390), .Z(n6384) );
  AND U6194 ( .A(n272), .B(n6391), .Z(n6390) );
  XOR U6195 ( .A(p_input[635]), .B(n6389), .Z(n6391) );
  XNOR U6196 ( .A(n6392), .B(n6393), .Z(n6389) );
  AND U6197 ( .A(n276), .B(n6388), .Z(n6393) );
  XNOR U6198 ( .A(n6392), .B(n6386), .Z(n6388) );
  XOR U6199 ( .A(n6394), .B(n6395), .Z(n6386) );
  AND U6200 ( .A(n291), .B(n6396), .Z(n6395) );
  XNOR U6201 ( .A(n6397), .B(n6398), .Z(n6392) );
  AND U6202 ( .A(n283), .B(n6399), .Z(n6398) );
  XOR U6203 ( .A(p_input[667]), .B(n6397), .Z(n6399) );
  XNOR U6204 ( .A(n6400), .B(n6401), .Z(n6397) );
  AND U6205 ( .A(n287), .B(n6396), .Z(n6401) );
  XNOR U6206 ( .A(n6400), .B(n6394), .Z(n6396) );
  XOR U6207 ( .A(n6402), .B(n6403), .Z(n6394) );
  AND U6208 ( .A(n302), .B(n6404), .Z(n6403) );
  XNOR U6209 ( .A(n6405), .B(n6406), .Z(n6400) );
  AND U6210 ( .A(n294), .B(n6407), .Z(n6406) );
  XOR U6211 ( .A(p_input[699]), .B(n6405), .Z(n6407) );
  XNOR U6212 ( .A(n6408), .B(n6409), .Z(n6405) );
  AND U6213 ( .A(n298), .B(n6404), .Z(n6409) );
  XNOR U6214 ( .A(n6408), .B(n6402), .Z(n6404) );
  XOR U6215 ( .A(n6410), .B(n6411), .Z(n6402) );
  AND U6216 ( .A(n313), .B(n6412), .Z(n6411) );
  XNOR U6217 ( .A(n6413), .B(n6414), .Z(n6408) );
  AND U6218 ( .A(n305), .B(n6415), .Z(n6414) );
  XOR U6219 ( .A(p_input[731]), .B(n6413), .Z(n6415) );
  XNOR U6220 ( .A(n6416), .B(n6417), .Z(n6413) );
  AND U6221 ( .A(n309), .B(n6412), .Z(n6417) );
  XNOR U6222 ( .A(n6416), .B(n6410), .Z(n6412) );
  XOR U6223 ( .A(n6418), .B(n6419), .Z(n6410) );
  AND U6224 ( .A(n324), .B(n6420), .Z(n6419) );
  XNOR U6225 ( .A(n6421), .B(n6422), .Z(n6416) );
  AND U6226 ( .A(n316), .B(n6423), .Z(n6422) );
  XOR U6227 ( .A(p_input[763]), .B(n6421), .Z(n6423) );
  XNOR U6228 ( .A(n6424), .B(n6425), .Z(n6421) );
  AND U6229 ( .A(n320), .B(n6420), .Z(n6425) );
  XNOR U6230 ( .A(n6424), .B(n6418), .Z(n6420) );
  XOR U6231 ( .A(n6426), .B(n6427), .Z(n6418) );
  AND U6232 ( .A(n335), .B(n6428), .Z(n6427) );
  XNOR U6233 ( .A(n6429), .B(n6430), .Z(n6424) );
  AND U6234 ( .A(n327), .B(n6431), .Z(n6430) );
  XOR U6235 ( .A(p_input[795]), .B(n6429), .Z(n6431) );
  XNOR U6236 ( .A(n6432), .B(n6433), .Z(n6429) );
  AND U6237 ( .A(n331), .B(n6428), .Z(n6433) );
  XNOR U6238 ( .A(n6432), .B(n6426), .Z(n6428) );
  XOR U6239 ( .A(n6434), .B(n6435), .Z(n6426) );
  AND U6240 ( .A(n346), .B(n6436), .Z(n6435) );
  XNOR U6241 ( .A(n6437), .B(n6438), .Z(n6432) );
  AND U6242 ( .A(n338), .B(n6439), .Z(n6438) );
  XOR U6243 ( .A(p_input[827]), .B(n6437), .Z(n6439) );
  XNOR U6244 ( .A(n6440), .B(n6441), .Z(n6437) );
  AND U6245 ( .A(n342), .B(n6436), .Z(n6441) );
  XNOR U6246 ( .A(n6440), .B(n6434), .Z(n6436) );
  XOR U6247 ( .A(n6442), .B(n6443), .Z(n6434) );
  AND U6248 ( .A(n357), .B(n6444), .Z(n6443) );
  XNOR U6249 ( .A(n6445), .B(n6446), .Z(n6440) );
  AND U6250 ( .A(n349), .B(n6447), .Z(n6446) );
  XOR U6251 ( .A(p_input[859]), .B(n6445), .Z(n6447) );
  XNOR U6252 ( .A(n6448), .B(n6449), .Z(n6445) );
  AND U6253 ( .A(n353), .B(n6444), .Z(n6449) );
  XNOR U6254 ( .A(n6448), .B(n6442), .Z(n6444) );
  XOR U6255 ( .A(n6450), .B(n6451), .Z(n6442) );
  AND U6256 ( .A(n368), .B(n6452), .Z(n6451) );
  XNOR U6257 ( .A(n6453), .B(n6454), .Z(n6448) );
  AND U6258 ( .A(n360), .B(n6455), .Z(n6454) );
  XOR U6259 ( .A(p_input[891]), .B(n6453), .Z(n6455) );
  XNOR U6260 ( .A(n6456), .B(n6457), .Z(n6453) );
  AND U6261 ( .A(n364), .B(n6452), .Z(n6457) );
  XNOR U6262 ( .A(n6456), .B(n6450), .Z(n6452) );
  XOR U6263 ( .A(n6458), .B(n6459), .Z(n6450) );
  AND U6264 ( .A(n379), .B(n6460), .Z(n6459) );
  XNOR U6265 ( .A(n6461), .B(n6462), .Z(n6456) );
  AND U6266 ( .A(n371), .B(n6463), .Z(n6462) );
  XOR U6267 ( .A(p_input[923]), .B(n6461), .Z(n6463) );
  XNOR U6268 ( .A(n6464), .B(n6465), .Z(n6461) );
  AND U6269 ( .A(n375), .B(n6460), .Z(n6465) );
  XNOR U6270 ( .A(n6464), .B(n6458), .Z(n6460) );
  XOR U6271 ( .A(n6466), .B(n6467), .Z(n6458) );
  AND U6272 ( .A(n390), .B(n6468), .Z(n6467) );
  XNOR U6273 ( .A(n6469), .B(n6470), .Z(n6464) );
  AND U6274 ( .A(n382), .B(n6471), .Z(n6470) );
  XOR U6275 ( .A(p_input[955]), .B(n6469), .Z(n6471) );
  XNOR U6276 ( .A(n6472), .B(n6473), .Z(n6469) );
  AND U6277 ( .A(n386), .B(n6468), .Z(n6473) );
  XNOR U6278 ( .A(n6472), .B(n6466), .Z(n6468) );
  XOR U6279 ( .A(n6474), .B(n6475), .Z(n6466) );
  AND U6280 ( .A(n401), .B(n6476), .Z(n6475) );
  XNOR U6281 ( .A(n6477), .B(n6478), .Z(n6472) );
  AND U6282 ( .A(n393), .B(n6479), .Z(n6478) );
  XOR U6283 ( .A(p_input[987]), .B(n6477), .Z(n6479) );
  XNOR U6284 ( .A(n6480), .B(n6481), .Z(n6477) );
  AND U6285 ( .A(n397), .B(n6476), .Z(n6481) );
  XNOR U6286 ( .A(n6480), .B(n6474), .Z(n6476) );
  XOR U6287 ( .A(n6482), .B(n6483), .Z(n6474) );
  AND U6288 ( .A(n412), .B(n6484), .Z(n6483) );
  XNOR U6289 ( .A(n6485), .B(n6486), .Z(n6480) );
  AND U6290 ( .A(n404), .B(n6487), .Z(n6486) );
  XOR U6291 ( .A(p_input[1019]), .B(n6485), .Z(n6487) );
  XNOR U6292 ( .A(n6488), .B(n6489), .Z(n6485) );
  AND U6293 ( .A(n408), .B(n6484), .Z(n6489) );
  XNOR U6294 ( .A(n6488), .B(n6482), .Z(n6484) );
  XOR U6295 ( .A(n6490), .B(n6491), .Z(n6482) );
  AND U6296 ( .A(n423), .B(n6492), .Z(n6491) );
  XNOR U6297 ( .A(n6493), .B(n6494), .Z(n6488) );
  AND U6298 ( .A(n415), .B(n6495), .Z(n6494) );
  XOR U6299 ( .A(p_input[1051]), .B(n6493), .Z(n6495) );
  XNOR U6300 ( .A(n6496), .B(n6497), .Z(n6493) );
  AND U6301 ( .A(n419), .B(n6492), .Z(n6497) );
  XNOR U6302 ( .A(n6496), .B(n6490), .Z(n6492) );
  XOR U6303 ( .A(n6498), .B(n6499), .Z(n6490) );
  AND U6304 ( .A(n434), .B(n6500), .Z(n6499) );
  XNOR U6305 ( .A(n6501), .B(n6502), .Z(n6496) );
  AND U6306 ( .A(n426), .B(n6503), .Z(n6502) );
  XOR U6307 ( .A(p_input[1083]), .B(n6501), .Z(n6503) );
  XNOR U6308 ( .A(n6504), .B(n6505), .Z(n6501) );
  AND U6309 ( .A(n430), .B(n6500), .Z(n6505) );
  XNOR U6310 ( .A(n6504), .B(n6498), .Z(n6500) );
  XOR U6311 ( .A(n6506), .B(n6507), .Z(n6498) );
  AND U6312 ( .A(n445), .B(n6508), .Z(n6507) );
  XNOR U6313 ( .A(n6509), .B(n6510), .Z(n6504) );
  AND U6314 ( .A(n437), .B(n6511), .Z(n6510) );
  XOR U6315 ( .A(p_input[1115]), .B(n6509), .Z(n6511) );
  XNOR U6316 ( .A(n6512), .B(n6513), .Z(n6509) );
  AND U6317 ( .A(n441), .B(n6508), .Z(n6513) );
  XNOR U6318 ( .A(n6512), .B(n6506), .Z(n6508) );
  XOR U6319 ( .A(n6514), .B(n6515), .Z(n6506) );
  AND U6320 ( .A(n456), .B(n6516), .Z(n6515) );
  XNOR U6321 ( .A(n6517), .B(n6518), .Z(n6512) );
  AND U6322 ( .A(n448), .B(n6519), .Z(n6518) );
  XOR U6323 ( .A(p_input[1147]), .B(n6517), .Z(n6519) );
  XNOR U6324 ( .A(n6520), .B(n6521), .Z(n6517) );
  AND U6325 ( .A(n452), .B(n6516), .Z(n6521) );
  XNOR U6326 ( .A(n6520), .B(n6514), .Z(n6516) );
  XOR U6327 ( .A(n6522), .B(n6523), .Z(n6514) );
  AND U6328 ( .A(n467), .B(n6524), .Z(n6523) );
  XNOR U6329 ( .A(n6525), .B(n6526), .Z(n6520) );
  AND U6330 ( .A(n459), .B(n6527), .Z(n6526) );
  XOR U6331 ( .A(p_input[1179]), .B(n6525), .Z(n6527) );
  XNOR U6332 ( .A(n6528), .B(n6529), .Z(n6525) );
  AND U6333 ( .A(n463), .B(n6524), .Z(n6529) );
  XNOR U6334 ( .A(n6528), .B(n6522), .Z(n6524) );
  XOR U6335 ( .A(n6530), .B(n6531), .Z(n6522) );
  AND U6336 ( .A(n478), .B(n6532), .Z(n6531) );
  XNOR U6337 ( .A(n6533), .B(n6534), .Z(n6528) );
  AND U6338 ( .A(n470), .B(n6535), .Z(n6534) );
  XOR U6339 ( .A(p_input[1211]), .B(n6533), .Z(n6535) );
  XNOR U6340 ( .A(n6536), .B(n6537), .Z(n6533) );
  AND U6341 ( .A(n474), .B(n6532), .Z(n6537) );
  XNOR U6342 ( .A(n6536), .B(n6530), .Z(n6532) );
  XOR U6343 ( .A(n6538), .B(n6539), .Z(n6530) );
  AND U6344 ( .A(n489), .B(n6540), .Z(n6539) );
  XNOR U6345 ( .A(n6541), .B(n6542), .Z(n6536) );
  AND U6346 ( .A(n481), .B(n6543), .Z(n6542) );
  XOR U6347 ( .A(p_input[1243]), .B(n6541), .Z(n6543) );
  XNOR U6348 ( .A(n6544), .B(n6545), .Z(n6541) );
  AND U6349 ( .A(n485), .B(n6540), .Z(n6545) );
  XNOR U6350 ( .A(n6544), .B(n6538), .Z(n6540) );
  XOR U6351 ( .A(n6546), .B(n6547), .Z(n6538) );
  AND U6352 ( .A(n500), .B(n6548), .Z(n6547) );
  XNOR U6353 ( .A(n6549), .B(n6550), .Z(n6544) );
  AND U6354 ( .A(n492), .B(n6551), .Z(n6550) );
  XOR U6355 ( .A(p_input[1275]), .B(n6549), .Z(n6551) );
  XNOR U6356 ( .A(n6552), .B(n6553), .Z(n6549) );
  AND U6357 ( .A(n496), .B(n6548), .Z(n6553) );
  XNOR U6358 ( .A(n6552), .B(n6546), .Z(n6548) );
  XOR U6359 ( .A(n6554), .B(n6555), .Z(n6546) );
  AND U6360 ( .A(n511), .B(n6556), .Z(n6555) );
  XNOR U6361 ( .A(n6557), .B(n6558), .Z(n6552) );
  AND U6362 ( .A(n503), .B(n6559), .Z(n6558) );
  XOR U6363 ( .A(p_input[1307]), .B(n6557), .Z(n6559) );
  XNOR U6364 ( .A(n6560), .B(n6561), .Z(n6557) );
  AND U6365 ( .A(n507), .B(n6556), .Z(n6561) );
  XNOR U6366 ( .A(n6560), .B(n6554), .Z(n6556) );
  XOR U6367 ( .A(n6562), .B(n6563), .Z(n6554) );
  AND U6368 ( .A(n522), .B(n6564), .Z(n6563) );
  XNOR U6369 ( .A(n6565), .B(n6566), .Z(n6560) );
  AND U6370 ( .A(n514), .B(n6567), .Z(n6566) );
  XOR U6371 ( .A(p_input[1339]), .B(n6565), .Z(n6567) );
  XNOR U6372 ( .A(n6568), .B(n6569), .Z(n6565) );
  AND U6373 ( .A(n518), .B(n6564), .Z(n6569) );
  XNOR U6374 ( .A(n6568), .B(n6562), .Z(n6564) );
  XOR U6375 ( .A(n6570), .B(n6571), .Z(n6562) );
  AND U6376 ( .A(n533), .B(n6572), .Z(n6571) );
  XNOR U6377 ( .A(n6573), .B(n6574), .Z(n6568) );
  AND U6378 ( .A(n525), .B(n6575), .Z(n6574) );
  XOR U6379 ( .A(p_input[1371]), .B(n6573), .Z(n6575) );
  XNOR U6380 ( .A(n6576), .B(n6577), .Z(n6573) );
  AND U6381 ( .A(n529), .B(n6572), .Z(n6577) );
  XNOR U6382 ( .A(n6576), .B(n6570), .Z(n6572) );
  XOR U6383 ( .A(n6578), .B(n6579), .Z(n6570) );
  AND U6384 ( .A(n544), .B(n6580), .Z(n6579) );
  XNOR U6385 ( .A(n6581), .B(n6582), .Z(n6576) );
  AND U6386 ( .A(n536), .B(n6583), .Z(n6582) );
  XOR U6387 ( .A(p_input[1403]), .B(n6581), .Z(n6583) );
  XNOR U6388 ( .A(n6584), .B(n6585), .Z(n6581) );
  AND U6389 ( .A(n540), .B(n6580), .Z(n6585) );
  XNOR U6390 ( .A(n6584), .B(n6578), .Z(n6580) );
  XOR U6391 ( .A(n6586), .B(n6587), .Z(n6578) );
  AND U6392 ( .A(n555), .B(n6588), .Z(n6587) );
  XNOR U6393 ( .A(n6589), .B(n6590), .Z(n6584) );
  AND U6394 ( .A(n547), .B(n6591), .Z(n6590) );
  XOR U6395 ( .A(p_input[1435]), .B(n6589), .Z(n6591) );
  XNOR U6396 ( .A(n6592), .B(n6593), .Z(n6589) );
  AND U6397 ( .A(n551), .B(n6588), .Z(n6593) );
  XNOR U6398 ( .A(n6592), .B(n6586), .Z(n6588) );
  XOR U6399 ( .A(n6594), .B(n6595), .Z(n6586) );
  AND U6400 ( .A(n566), .B(n6596), .Z(n6595) );
  XNOR U6401 ( .A(n6597), .B(n6598), .Z(n6592) );
  AND U6402 ( .A(n558), .B(n6599), .Z(n6598) );
  XOR U6403 ( .A(p_input[1467]), .B(n6597), .Z(n6599) );
  XNOR U6404 ( .A(n6600), .B(n6601), .Z(n6597) );
  AND U6405 ( .A(n562), .B(n6596), .Z(n6601) );
  XNOR U6406 ( .A(n6600), .B(n6594), .Z(n6596) );
  XOR U6407 ( .A(n6602), .B(n6603), .Z(n6594) );
  AND U6408 ( .A(n577), .B(n6604), .Z(n6603) );
  XNOR U6409 ( .A(n6605), .B(n6606), .Z(n6600) );
  AND U6410 ( .A(n569), .B(n6607), .Z(n6606) );
  XOR U6411 ( .A(p_input[1499]), .B(n6605), .Z(n6607) );
  XNOR U6412 ( .A(n6608), .B(n6609), .Z(n6605) );
  AND U6413 ( .A(n573), .B(n6604), .Z(n6609) );
  XNOR U6414 ( .A(n6608), .B(n6602), .Z(n6604) );
  XOR U6415 ( .A(n6610), .B(n6611), .Z(n6602) );
  AND U6416 ( .A(n588), .B(n6612), .Z(n6611) );
  XNOR U6417 ( .A(n6613), .B(n6614), .Z(n6608) );
  AND U6418 ( .A(n580), .B(n6615), .Z(n6614) );
  XOR U6419 ( .A(p_input[1531]), .B(n6613), .Z(n6615) );
  XNOR U6420 ( .A(n6616), .B(n6617), .Z(n6613) );
  AND U6421 ( .A(n584), .B(n6612), .Z(n6617) );
  XNOR U6422 ( .A(n6616), .B(n6610), .Z(n6612) );
  XOR U6423 ( .A(n6618), .B(n6619), .Z(n6610) );
  AND U6424 ( .A(n599), .B(n6620), .Z(n6619) );
  XNOR U6425 ( .A(n6621), .B(n6622), .Z(n6616) );
  AND U6426 ( .A(n591), .B(n6623), .Z(n6622) );
  XOR U6427 ( .A(p_input[1563]), .B(n6621), .Z(n6623) );
  XNOR U6428 ( .A(n6624), .B(n6625), .Z(n6621) );
  AND U6429 ( .A(n595), .B(n6620), .Z(n6625) );
  XNOR U6430 ( .A(n6624), .B(n6618), .Z(n6620) );
  XOR U6431 ( .A(n6626), .B(n6627), .Z(n6618) );
  AND U6432 ( .A(n610), .B(n6628), .Z(n6627) );
  XNOR U6433 ( .A(n6629), .B(n6630), .Z(n6624) );
  AND U6434 ( .A(n602), .B(n6631), .Z(n6630) );
  XOR U6435 ( .A(p_input[1595]), .B(n6629), .Z(n6631) );
  XNOR U6436 ( .A(n6632), .B(n6633), .Z(n6629) );
  AND U6437 ( .A(n606), .B(n6628), .Z(n6633) );
  XNOR U6438 ( .A(n6632), .B(n6626), .Z(n6628) );
  XOR U6439 ( .A(n6634), .B(n6635), .Z(n6626) );
  AND U6440 ( .A(n621), .B(n6636), .Z(n6635) );
  XNOR U6441 ( .A(n6637), .B(n6638), .Z(n6632) );
  AND U6442 ( .A(n613), .B(n6639), .Z(n6638) );
  XOR U6443 ( .A(p_input[1627]), .B(n6637), .Z(n6639) );
  XNOR U6444 ( .A(n6640), .B(n6641), .Z(n6637) );
  AND U6445 ( .A(n617), .B(n6636), .Z(n6641) );
  XNOR U6446 ( .A(n6640), .B(n6634), .Z(n6636) );
  XOR U6447 ( .A(n6642), .B(n6643), .Z(n6634) );
  AND U6448 ( .A(n632), .B(n6644), .Z(n6643) );
  XNOR U6449 ( .A(n6645), .B(n6646), .Z(n6640) );
  AND U6450 ( .A(n624), .B(n6647), .Z(n6646) );
  XOR U6451 ( .A(p_input[1659]), .B(n6645), .Z(n6647) );
  XNOR U6452 ( .A(n6648), .B(n6649), .Z(n6645) );
  AND U6453 ( .A(n628), .B(n6644), .Z(n6649) );
  XNOR U6454 ( .A(n6648), .B(n6642), .Z(n6644) );
  XOR U6455 ( .A(n6650), .B(n6651), .Z(n6642) );
  AND U6456 ( .A(n643), .B(n6652), .Z(n6651) );
  XNOR U6457 ( .A(n6653), .B(n6654), .Z(n6648) );
  AND U6458 ( .A(n635), .B(n6655), .Z(n6654) );
  XOR U6459 ( .A(p_input[1691]), .B(n6653), .Z(n6655) );
  XNOR U6460 ( .A(n6656), .B(n6657), .Z(n6653) );
  AND U6461 ( .A(n639), .B(n6652), .Z(n6657) );
  XNOR U6462 ( .A(n6656), .B(n6650), .Z(n6652) );
  XOR U6463 ( .A(n6658), .B(n6659), .Z(n6650) );
  AND U6464 ( .A(n654), .B(n6660), .Z(n6659) );
  XNOR U6465 ( .A(n6661), .B(n6662), .Z(n6656) );
  AND U6466 ( .A(n646), .B(n6663), .Z(n6662) );
  XOR U6467 ( .A(p_input[1723]), .B(n6661), .Z(n6663) );
  XNOR U6468 ( .A(n6664), .B(n6665), .Z(n6661) );
  AND U6469 ( .A(n650), .B(n6660), .Z(n6665) );
  XNOR U6470 ( .A(n6664), .B(n6658), .Z(n6660) );
  XOR U6471 ( .A(n6666), .B(n6667), .Z(n6658) );
  AND U6472 ( .A(n665), .B(n6668), .Z(n6667) );
  XNOR U6473 ( .A(n6669), .B(n6670), .Z(n6664) );
  AND U6474 ( .A(n657), .B(n6671), .Z(n6670) );
  XOR U6475 ( .A(p_input[1755]), .B(n6669), .Z(n6671) );
  XNOR U6476 ( .A(n6672), .B(n6673), .Z(n6669) );
  AND U6477 ( .A(n661), .B(n6668), .Z(n6673) );
  XNOR U6478 ( .A(n6672), .B(n6666), .Z(n6668) );
  XOR U6479 ( .A(n6674), .B(n6675), .Z(n6666) );
  AND U6480 ( .A(n676), .B(n6676), .Z(n6675) );
  XNOR U6481 ( .A(n6677), .B(n6678), .Z(n6672) );
  AND U6482 ( .A(n668), .B(n6679), .Z(n6678) );
  XOR U6483 ( .A(p_input[1787]), .B(n6677), .Z(n6679) );
  XNOR U6484 ( .A(n6680), .B(n6681), .Z(n6677) );
  AND U6485 ( .A(n672), .B(n6676), .Z(n6681) );
  XNOR U6486 ( .A(n6680), .B(n6674), .Z(n6676) );
  XOR U6487 ( .A(n6682), .B(n6683), .Z(n6674) );
  AND U6488 ( .A(n687), .B(n6684), .Z(n6683) );
  XNOR U6489 ( .A(n6685), .B(n6686), .Z(n6680) );
  AND U6490 ( .A(n679), .B(n6687), .Z(n6686) );
  XOR U6491 ( .A(p_input[1819]), .B(n6685), .Z(n6687) );
  XNOR U6492 ( .A(n6688), .B(n6689), .Z(n6685) );
  AND U6493 ( .A(n683), .B(n6684), .Z(n6689) );
  XNOR U6494 ( .A(n6688), .B(n6682), .Z(n6684) );
  XOR U6495 ( .A(n6690), .B(n6691), .Z(n6682) );
  AND U6496 ( .A(n698), .B(n6692), .Z(n6691) );
  XNOR U6497 ( .A(n6693), .B(n6694), .Z(n6688) );
  AND U6498 ( .A(n690), .B(n6695), .Z(n6694) );
  XOR U6499 ( .A(p_input[1851]), .B(n6693), .Z(n6695) );
  XNOR U6500 ( .A(n6696), .B(n6697), .Z(n6693) );
  AND U6501 ( .A(n694), .B(n6692), .Z(n6697) );
  XNOR U6502 ( .A(n6696), .B(n6690), .Z(n6692) );
  XOR U6503 ( .A(n6698), .B(n6699), .Z(n6690) );
  AND U6504 ( .A(n709), .B(n6700), .Z(n6699) );
  XNOR U6505 ( .A(n6701), .B(n6702), .Z(n6696) );
  AND U6506 ( .A(n701), .B(n6703), .Z(n6702) );
  XOR U6507 ( .A(p_input[1883]), .B(n6701), .Z(n6703) );
  XNOR U6508 ( .A(n6704), .B(n6705), .Z(n6701) );
  AND U6509 ( .A(n705), .B(n6700), .Z(n6705) );
  XNOR U6510 ( .A(n6704), .B(n6698), .Z(n6700) );
  XOR U6511 ( .A(n6706), .B(n6707), .Z(n6698) );
  AND U6512 ( .A(n720), .B(n6708), .Z(n6707) );
  XNOR U6513 ( .A(n6709), .B(n6710), .Z(n6704) );
  AND U6514 ( .A(n712), .B(n6711), .Z(n6710) );
  XOR U6515 ( .A(p_input[1915]), .B(n6709), .Z(n6711) );
  XNOR U6516 ( .A(n6712), .B(n6713), .Z(n6709) );
  AND U6517 ( .A(n716), .B(n6708), .Z(n6713) );
  XNOR U6518 ( .A(n6712), .B(n6706), .Z(n6708) );
  XOR U6519 ( .A(n6714), .B(n6715), .Z(n6706) );
  AND U6520 ( .A(n731), .B(n6716), .Z(n6715) );
  XNOR U6521 ( .A(n6717), .B(n6718), .Z(n6712) );
  AND U6522 ( .A(n723), .B(n6719), .Z(n6718) );
  XOR U6523 ( .A(p_input[1947]), .B(n6717), .Z(n6719) );
  XNOR U6524 ( .A(n6720), .B(n6721), .Z(n6717) );
  AND U6525 ( .A(n727), .B(n6716), .Z(n6721) );
  XNOR U6526 ( .A(n6720), .B(n6714), .Z(n6716) );
  XOR U6527 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n6722), .Z(n6714) );
  AND U6528 ( .A(n741), .B(n6723), .Z(n6722) );
  XNOR U6529 ( .A(n6724), .B(n6725), .Z(n6720) );
  AND U6530 ( .A(n734), .B(n6726), .Z(n6725) );
  XOR U6531 ( .A(p_input[1979]), .B(n6724), .Z(n6726) );
  XNOR U6532 ( .A(n6727), .B(n6728), .Z(n6724) );
  AND U6533 ( .A(n738), .B(n6723), .Z(n6728) );
  XOR U6534 ( .A(n6729), .B(n6727), .Z(n6723) );
  IV U6535 ( .A(\knn_comb_/min_val_out[0][27] ), .Z(n6729) );
  IV U6536 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .Z(n6727) );
  XOR U6537 ( .A(n21), .B(n6730), .Z(o[26]) );
  AND U6538 ( .A(n58), .B(n6731), .Z(n21) );
  XOR U6539 ( .A(n22), .B(n6730), .Z(n6731) );
  XOR U6540 ( .A(n6732), .B(n6733), .Z(n6730) );
  AND U6541 ( .A(n70), .B(n6734), .Z(n6733) );
  XOR U6542 ( .A(n6735), .B(n6736), .Z(n22) );
  AND U6543 ( .A(n62), .B(n6737), .Z(n6736) );
  XOR U6544 ( .A(p_input[26]), .B(n6735), .Z(n6737) );
  XNOR U6545 ( .A(n6738), .B(n6739), .Z(n6735) );
  AND U6546 ( .A(n66), .B(n6734), .Z(n6739) );
  XNOR U6547 ( .A(n6738), .B(n6732), .Z(n6734) );
  XOR U6548 ( .A(n6740), .B(n6741), .Z(n6732) );
  AND U6549 ( .A(n82), .B(n6742), .Z(n6741) );
  XNOR U6550 ( .A(n6743), .B(n6744), .Z(n6738) );
  AND U6551 ( .A(n74), .B(n6745), .Z(n6744) );
  XOR U6552 ( .A(p_input[58]), .B(n6743), .Z(n6745) );
  XNOR U6553 ( .A(n6746), .B(n6747), .Z(n6743) );
  AND U6554 ( .A(n78), .B(n6742), .Z(n6747) );
  XNOR U6555 ( .A(n6746), .B(n6740), .Z(n6742) );
  XOR U6556 ( .A(n6748), .B(n6749), .Z(n6740) );
  AND U6557 ( .A(n93), .B(n6750), .Z(n6749) );
  XNOR U6558 ( .A(n6751), .B(n6752), .Z(n6746) );
  AND U6559 ( .A(n85), .B(n6753), .Z(n6752) );
  XOR U6560 ( .A(p_input[90]), .B(n6751), .Z(n6753) );
  XNOR U6561 ( .A(n6754), .B(n6755), .Z(n6751) );
  AND U6562 ( .A(n89), .B(n6750), .Z(n6755) );
  XNOR U6563 ( .A(n6754), .B(n6748), .Z(n6750) );
  XOR U6564 ( .A(n6756), .B(n6757), .Z(n6748) );
  AND U6565 ( .A(n104), .B(n6758), .Z(n6757) );
  XNOR U6566 ( .A(n6759), .B(n6760), .Z(n6754) );
  AND U6567 ( .A(n96), .B(n6761), .Z(n6760) );
  XOR U6568 ( .A(p_input[122]), .B(n6759), .Z(n6761) );
  XNOR U6569 ( .A(n6762), .B(n6763), .Z(n6759) );
  AND U6570 ( .A(n100), .B(n6758), .Z(n6763) );
  XNOR U6571 ( .A(n6762), .B(n6756), .Z(n6758) );
  XOR U6572 ( .A(n6764), .B(n6765), .Z(n6756) );
  AND U6573 ( .A(n115), .B(n6766), .Z(n6765) );
  XNOR U6574 ( .A(n6767), .B(n6768), .Z(n6762) );
  AND U6575 ( .A(n107), .B(n6769), .Z(n6768) );
  XOR U6576 ( .A(p_input[154]), .B(n6767), .Z(n6769) );
  XNOR U6577 ( .A(n6770), .B(n6771), .Z(n6767) );
  AND U6578 ( .A(n111), .B(n6766), .Z(n6771) );
  XNOR U6579 ( .A(n6770), .B(n6764), .Z(n6766) );
  XOR U6580 ( .A(n6772), .B(n6773), .Z(n6764) );
  AND U6581 ( .A(n126), .B(n6774), .Z(n6773) );
  XNOR U6582 ( .A(n6775), .B(n6776), .Z(n6770) );
  AND U6583 ( .A(n118), .B(n6777), .Z(n6776) );
  XOR U6584 ( .A(p_input[186]), .B(n6775), .Z(n6777) );
  XNOR U6585 ( .A(n6778), .B(n6779), .Z(n6775) );
  AND U6586 ( .A(n122), .B(n6774), .Z(n6779) );
  XNOR U6587 ( .A(n6778), .B(n6772), .Z(n6774) );
  XOR U6588 ( .A(n6780), .B(n6781), .Z(n6772) );
  AND U6589 ( .A(n137), .B(n6782), .Z(n6781) );
  XNOR U6590 ( .A(n6783), .B(n6784), .Z(n6778) );
  AND U6591 ( .A(n129), .B(n6785), .Z(n6784) );
  XOR U6592 ( .A(p_input[218]), .B(n6783), .Z(n6785) );
  XNOR U6593 ( .A(n6786), .B(n6787), .Z(n6783) );
  AND U6594 ( .A(n133), .B(n6782), .Z(n6787) );
  XNOR U6595 ( .A(n6786), .B(n6780), .Z(n6782) );
  XOR U6596 ( .A(n6788), .B(n6789), .Z(n6780) );
  AND U6597 ( .A(n148), .B(n6790), .Z(n6789) );
  XNOR U6598 ( .A(n6791), .B(n6792), .Z(n6786) );
  AND U6599 ( .A(n140), .B(n6793), .Z(n6792) );
  XOR U6600 ( .A(p_input[250]), .B(n6791), .Z(n6793) );
  XNOR U6601 ( .A(n6794), .B(n6795), .Z(n6791) );
  AND U6602 ( .A(n144), .B(n6790), .Z(n6795) );
  XNOR U6603 ( .A(n6794), .B(n6788), .Z(n6790) );
  XOR U6604 ( .A(n6796), .B(n6797), .Z(n6788) );
  AND U6605 ( .A(n159), .B(n6798), .Z(n6797) );
  XNOR U6606 ( .A(n6799), .B(n6800), .Z(n6794) );
  AND U6607 ( .A(n151), .B(n6801), .Z(n6800) );
  XOR U6608 ( .A(p_input[282]), .B(n6799), .Z(n6801) );
  XNOR U6609 ( .A(n6802), .B(n6803), .Z(n6799) );
  AND U6610 ( .A(n155), .B(n6798), .Z(n6803) );
  XNOR U6611 ( .A(n6802), .B(n6796), .Z(n6798) );
  XOR U6612 ( .A(n6804), .B(n6805), .Z(n6796) );
  AND U6613 ( .A(n170), .B(n6806), .Z(n6805) );
  XNOR U6614 ( .A(n6807), .B(n6808), .Z(n6802) );
  AND U6615 ( .A(n162), .B(n6809), .Z(n6808) );
  XOR U6616 ( .A(p_input[314]), .B(n6807), .Z(n6809) );
  XNOR U6617 ( .A(n6810), .B(n6811), .Z(n6807) );
  AND U6618 ( .A(n166), .B(n6806), .Z(n6811) );
  XNOR U6619 ( .A(n6810), .B(n6804), .Z(n6806) );
  XOR U6620 ( .A(n6812), .B(n6813), .Z(n6804) );
  AND U6621 ( .A(n181), .B(n6814), .Z(n6813) );
  XNOR U6622 ( .A(n6815), .B(n6816), .Z(n6810) );
  AND U6623 ( .A(n173), .B(n6817), .Z(n6816) );
  XOR U6624 ( .A(p_input[346]), .B(n6815), .Z(n6817) );
  XNOR U6625 ( .A(n6818), .B(n6819), .Z(n6815) );
  AND U6626 ( .A(n177), .B(n6814), .Z(n6819) );
  XNOR U6627 ( .A(n6818), .B(n6812), .Z(n6814) );
  XOR U6628 ( .A(n6820), .B(n6821), .Z(n6812) );
  AND U6629 ( .A(n192), .B(n6822), .Z(n6821) );
  XNOR U6630 ( .A(n6823), .B(n6824), .Z(n6818) );
  AND U6631 ( .A(n184), .B(n6825), .Z(n6824) );
  XOR U6632 ( .A(p_input[378]), .B(n6823), .Z(n6825) );
  XNOR U6633 ( .A(n6826), .B(n6827), .Z(n6823) );
  AND U6634 ( .A(n188), .B(n6822), .Z(n6827) );
  XNOR U6635 ( .A(n6826), .B(n6820), .Z(n6822) );
  XOR U6636 ( .A(n6828), .B(n6829), .Z(n6820) );
  AND U6637 ( .A(n203), .B(n6830), .Z(n6829) );
  XNOR U6638 ( .A(n6831), .B(n6832), .Z(n6826) );
  AND U6639 ( .A(n195), .B(n6833), .Z(n6832) );
  XOR U6640 ( .A(p_input[410]), .B(n6831), .Z(n6833) );
  XNOR U6641 ( .A(n6834), .B(n6835), .Z(n6831) );
  AND U6642 ( .A(n199), .B(n6830), .Z(n6835) );
  XNOR U6643 ( .A(n6834), .B(n6828), .Z(n6830) );
  XOR U6644 ( .A(n6836), .B(n6837), .Z(n6828) );
  AND U6645 ( .A(n214), .B(n6838), .Z(n6837) );
  XNOR U6646 ( .A(n6839), .B(n6840), .Z(n6834) );
  AND U6647 ( .A(n206), .B(n6841), .Z(n6840) );
  XOR U6648 ( .A(p_input[442]), .B(n6839), .Z(n6841) );
  XNOR U6649 ( .A(n6842), .B(n6843), .Z(n6839) );
  AND U6650 ( .A(n210), .B(n6838), .Z(n6843) );
  XNOR U6651 ( .A(n6842), .B(n6836), .Z(n6838) );
  XOR U6652 ( .A(n6844), .B(n6845), .Z(n6836) );
  AND U6653 ( .A(n225), .B(n6846), .Z(n6845) );
  XNOR U6654 ( .A(n6847), .B(n6848), .Z(n6842) );
  AND U6655 ( .A(n217), .B(n6849), .Z(n6848) );
  XOR U6656 ( .A(p_input[474]), .B(n6847), .Z(n6849) );
  XNOR U6657 ( .A(n6850), .B(n6851), .Z(n6847) );
  AND U6658 ( .A(n221), .B(n6846), .Z(n6851) );
  XNOR U6659 ( .A(n6850), .B(n6844), .Z(n6846) );
  XOR U6660 ( .A(n6852), .B(n6853), .Z(n6844) );
  AND U6661 ( .A(n236), .B(n6854), .Z(n6853) );
  XNOR U6662 ( .A(n6855), .B(n6856), .Z(n6850) );
  AND U6663 ( .A(n228), .B(n6857), .Z(n6856) );
  XOR U6664 ( .A(p_input[506]), .B(n6855), .Z(n6857) );
  XNOR U6665 ( .A(n6858), .B(n6859), .Z(n6855) );
  AND U6666 ( .A(n232), .B(n6854), .Z(n6859) );
  XNOR U6667 ( .A(n6858), .B(n6852), .Z(n6854) );
  XOR U6668 ( .A(n6860), .B(n6861), .Z(n6852) );
  AND U6669 ( .A(n247), .B(n6862), .Z(n6861) );
  XNOR U6670 ( .A(n6863), .B(n6864), .Z(n6858) );
  AND U6671 ( .A(n239), .B(n6865), .Z(n6864) );
  XOR U6672 ( .A(p_input[538]), .B(n6863), .Z(n6865) );
  XNOR U6673 ( .A(n6866), .B(n6867), .Z(n6863) );
  AND U6674 ( .A(n243), .B(n6862), .Z(n6867) );
  XNOR U6675 ( .A(n6866), .B(n6860), .Z(n6862) );
  XOR U6676 ( .A(n6868), .B(n6869), .Z(n6860) );
  AND U6677 ( .A(n258), .B(n6870), .Z(n6869) );
  XNOR U6678 ( .A(n6871), .B(n6872), .Z(n6866) );
  AND U6679 ( .A(n250), .B(n6873), .Z(n6872) );
  XOR U6680 ( .A(p_input[570]), .B(n6871), .Z(n6873) );
  XNOR U6681 ( .A(n6874), .B(n6875), .Z(n6871) );
  AND U6682 ( .A(n254), .B(n6870), .Z(n6875) );
  XNOR U6683 ( .A(n6874), .B(n6868), .Z(n6870) );
  XOR U6684 ( .A(n6876), .B(n6877), .Z(n6868) );
  AND U6685 ( .A(n269), .B(n6878), .Z(n6877) );
  XNOR U6686 ( .A(n6879), .B(n6880), .Z(n6874) );
  AND U6687 ( .A(n261), .B(n6881), .Z(n6880) );
  XOR U6688 ( .A(p_input[602]), .B(n6879), .Z(n6881) );
  XNOR U6689 ( .A(n6882), .B(n6883), .Z(n6879) );
  AND U6690 ( .A(n265), .B(n6878), .Z(n6883) );
  XNOR U6691 ( .A(n6882), .B(n6876), .Z(n6878) );
  XOR U6692 ( .A(n6884), .B(n6885), .Z(n6876) );
  AND U6693 ( .A(n280), .B(n6886), .Z(n6885) );
  XNOR U6694 ( .A(n6887), .B(n6888), .Z(n6882) );
  AND U6695 ( .A(n272), .B(n6889), .Z(n6888) );
  XOR U6696 ( .A(p_input[634]), .B(n6887), .Z(n6889) );
  XNOR U6697 ( .A(n6890), .B(n6891), .Z(n6887) );
  AND U6698 ( .A(n276), .B(n6886), .Z(n6891) );
  XNOR U6699 ( .A(n6890), .B(n6884), .Z(n6886) );
  XOR U6700 ( .A(n6892), .B(n6893), .Z(n6884) );
  AND U6701 ( .A(n291), .B(n6894), .Z(n6893) );
  XNOR U6702 ( .A(n6895), .B(n6896), .Z(n6890) );
  AND U6703 ( .A(n283), .B(n6897), .Z(n6896) );
  XOR U6704 ( .A(p_input[666]), .B(n6895), .Z(n6897) );
  XNOR U6705 ( .A(n6898), .B(n6899), .Z(n6895) );
  AND U6706 ( .A(n287), .B(n6894), .Z(n6899) );
  XNOR U6707 ( .A(n6898), .B(n6892), .Z(n6894) );
  XOR U6708 ( .A(n6900), .B(n6901), .Z(n6892) );
  AND U6709 ( .A(n302), .B(n6902), .Z(n6901) );
  XNOR U6710 ( .A(n6903), .B(n6904), .Z(n6898) );
  AND U6711 ( .A(n294), .B(n6905), .Z(n6904) );
  XOR U6712 ( .A(p_input[698]), .B(n6903), .Z(n6905) );
  XNOR U6713 ( .A(n6906), .B(n6907), .Z(n6903) );
  AND U6714 ( .A(n298), .B(n6902), .Z(n6907) );
  XNOR U6715 ( .A(n6906), .B(n6900), .Z(n6902) );
  XOR U6716 ( .A(n6908), .B(n6909), .Z(n6900) );
  AND U6717 ( .A(n313), .B(n6910), .Z(n6909) );
  XNOR U6718 ( .A(n6911), .B(n6912), .Z(n6906) );
  AND U6719 ( .A(n305), .B(n6913), .Z(n6912) );
  XOR U6720 ( .A(p_input[730]), .B(n6911), .Z(n6913) );
  XNOR U6721 ( .A(n6914), .B(n6915), .Z(n6911) );
  AND U6722 ( .A(n309), .B(n6910), .Z(n6915) );
  XNOR U6723 ( .A(n6914), .B(n6908), .Z(n6910) );
  XOR U6724 ( .A(n6916), .B(n6917), .Z(n6908) );
  AND U6725 ( .A(n324), .B(n6918), .Z(n6917) );
  XNOR U6726 ( .A(n6919), .B(n6920), .Z(n6914) );
  AND U6727 ( .A(n316), .B(n6921), .Z(n6920) );
  XOR U6728 ( .A(p_input[762]), .B(n6919), .Z(n6921) );
  XNOR U6729 ( .A(n6922), .B(n6923), .Z(n6919) );
  AND U6730 ( .A(n320), .B(n6918), .Z(n6923) );
  XNOR U6731 ( .A(n6922), .B(n6916), .Z(n6918) );
  XOR U6732 ( .A(n6924), .B(n6925), .Z(n6916) );
  AND U6733 ( .A(n335), .B(n6926), .Z(n6925) );
  XNOR U6734 ( .A(n6927), .B(n6928), .Z(n6922) );
  AND U6735 ( .A(n327), .B(n6929), .Z(n6928) );
  XOR U6736 ( .A(p_input[794]), .B(n6927), .Z(n6929) );
  XNOR U6737 ( .A(n6930), .B(n6931), .Z(n6927) );
  AND U6738 ( .A(n331), .B(n6926), .Z(n6931) );
  XNOR U6739 ( .A(n6930), .B(n6924), .Z(n6926) );
  XOR U6740 ( .A(n6932), .B(n6933), .Z(n6924) );
  AND U6741 ( .A(n346), .B(n6934), .Z(n6933) );
  XNOR U6742 ( .A(n6935), .B(n6936), .Z(n6930) );
  AND U6743 ( .A(n338), .B(n6937), .Z(n6936) );
  XOR U6744 ( .A(p_input[826]), .B(n6935), .Z(n6937) );
  XNOR U6745 ( .A(n6938), .B(n6939), .Z(n6935) );
  AND U6746 ( .A(n342), .B(n6934), .Z(n6939) );
  XNOR U6747 ( .A(n6938), .B(n6932), .Z(n6934) );
  XOR U6748 ( .A(n6940), .B(n6941), .Z(n6932) );
  AND U6749 ( .A(n357), .B(n6942), .Z(n6941) );
  XNOR U6750 ( .A(n6943), .B(n6944), .Z(n6938) );
  AND U6751 ( .A(n349), .B(n6945), .Z(n6944) );
  XOR U6752 ( .A(p_input[858]), .B(n6943), .Z(n6945) );
  XNOR U6753 ( .A(n6946), .B(n6947), .Z(n6943) );
  AND U6754 ( .A(n353), .B(n6942), .Z(n6947) );
  XNOR U6755 ( .A(n6946), .B(n6940), .Z(n6942) );
  XOR U6756 ( .A(n6948), .B(n6949), .Z(n6940) );
  AND U6757 ( .A(n368), .B(n6950), .Z(n6949) );
  XNOR U6758 ( .A(n6951), .B(n6952), .Z(n6946) );
  AND U6759 ( .A(n360), .B(n6953), .Z(n6952) );
  XOR U6760 ( .A(p_input[890]), .B(n6951), .Z(n6953) );
  XNOR U6761 ( .A(n6954), .B(n6955), .Z(n6951) );
  AND U6762 ( .A(n364), .B(n6950), .Z(n6955) );
  XNOR U6763 ( .A(n6954), .B(n6948), .Z(n6950) );
  XOR U6764 ( .A(n6956), .B(n6957), .Z(n6948) );
  AND U6765 ( .A(n379), .B(n6958), .Z(n6957) );
  XNOR U6766 ( .A(n6959), .B(n6960), .Z(n6954) );
  AND U6767 ( .A(n371), .B(n6961), .Z(n6960) );
  XOR U6768 ( .A(p_input[922]), .B(n6959), .Z(n6961) );
  XNOR U6769 ( .A(n6962), .B(n6963), .Z(n6959) );
  AND U6770 ( .A(n375), .B(n6958), .Z(n6963) );
  XNOR U6771 ( .A(n6962), .B(n6956), .Z(n6958) );
  XOR U6772 ( .A(n6964), .B(n6965), .Z(n6956) );
  AND U6773 ( .A(n390), .B(n6966), .Z(n6965) );
  XNOR U6774 ( .A(n6967), .B(n6968), .Z(n6962) );
  AND U6775 ( .A(n382), .B(n6969), .Z(n6968) );
  XOR U6776 ( .A(p_input[954]), .B(n6967), .Z(n6969) );
  XNOR U6777 ( .A(n6970), .B(n6971), .Z(n6967) );
  AND U6778 ( .A(n386), .B(n6966), .Z(n6971) );
  XNOR U6779 ( .A(n6970), .B(n6964), .Z(n6966) );
  XOR U6780 ( .A(n6972), .B(n6973), .Z(n6964) );
  AND U6781 ( .A(n401), .B(n6974), .Z(n6973) );
  XNOR U6782 ( .A(n6975), .B(n6976), .Z(n6970) );
  AND U6783 ( .A(n393), .B(n6977), .Z(n6976) );
  XOR U6784 ( .A(p_input[986]), .B(n6975), .Z(n6977) );
  XNOR U6785 ( .A(n6978), .B(n6979), .Z(n6975) );
  AND U6786 ( .A(n397), .B(n6974), .Z(n6979) );
  XNOR U6787 ( .A(n6978), .B(n6972), .Z(n6974) );
  XOR U6788 ( .A(n6980), .B(n6981), .Z(n6972) );
  AND U6789 ( .A(n412), .B(n6982), .Z(n6981) );
  XNOR U6790 ( .A(n6983), .B(n6984), .Z(n6978) );
  AND U6791 ( .A(n404), .B(n6985), .Z(n6984) );
  XOR U6792 ( .A(p_input[1018]), .B(n6983), .Z(n6985) );
  XNOR U6793 ( .A(n6986), .B(n6987), .Z(n6983) );
  AND U6794 ( .A(n408), .B(n6982), .Z(n6987) );
  XNOR U6795 ( .A(n6986), .B(n6980), .Z(n6982) );
  XOR U6796 ( .A(n6988), .B(n6989), .Z(n6980) );
  AND U6797 ( .A(n423), .B(n6990), .Z(n6989) );
  XNOR U6798 ( .A(n6991), .B(n6992), .Z(n6986) );
  AND U6799 ( .A(n415), .B(n6993), .Z(n6992) );
  XOR U6800 ( .A(p_input[1050]), .B(n6991), .Z(n6993) );
  XNOR U6801 ( .A(n6994), .B(n6995), .Z(n6991) );
  AND U6802 ( .A(n419), .B(n6990), .Z(n6995) );
  XNOR U6803 ( .A(n6994), .B(n6988), .Z(n6990) );
  XOR U6804 ( .A(n6996), .B(n6997), .Z(n6988) );
  AND U6805 ( .A(n434), .B(n6998), .Z(n6997) );
  XNOR U6806 ( .A(n6999), .B(n7000), .Z(n6994) );
  AND U6807 ( .A(n426), .B(n7001), .Z(n7000) );
  XOR U6808 ( .A(p_input[1082]), .B(n6999), .Z(n7001) );
  XNOR U6809 ( .A(n7002), .B(n7003), .Z(n6999) );
  AND U6810 ( .A(n430), .B(n6998), .Z(n7003) );
  XNOR U6811 ( .A(n7002), .B(n6996), .Z(n6998) );
  XOR U6812 ( .A(n7004), .B(n7005), .Z(n6996) );
  AND U6813 ( .A(n445), .B(n7006), .Z(n7005) );
  XNOR U6814 ( .A(n7007), .B(n7008), .Z(n7002) );
  AND U6815 ( .A(n437), .B(n7009), .Z(n7008) );
  XOR U6816 ( .A(p_input[1114]), .B(n7007), .Z(n7009) );
  XNOR U6817 ( .A(n7010), .B(n7011), .Z(n7007) );
  AND U6818 ( .A(n441), .B(n7006), .Z(n7011) );
  XNOR U6819 ( .A(n7010), .B(n7004), .Z(n7006) );
  XOR U6820 ( .A(n7012), .B(n7013), .Z(n7004) );
  AND U6821 ( .A(n456), .B(n7014), .Z(n7013) );
  XNOR U6822 ( .A(n7015), .B(n7016), .Z(n7010) );
  AND U6823 ( .A(n448), .B(n7017), .Z(n7016) );
  XOR U6824 ( .A(p_input[1146]), .B(n7015), .Z(n7017) );
  XNOR U6825 ( .A(n7018), .B(n7019), .Z(n7015) );
  AND U6826 ( .A(n452), .B(n7014), .Z(n7019) );
  XNOR U6827 ( .A(n7018), .B(n7012), .Z(n7014) );
  XOR U6828 ( .A(n7020), .B(n7021), .Z(n7012) );
  AND U6829 ( .A(n467), .B(n7022), .Z(n7021) );
  XNOR U6830 ( .A(n7023), .B(n7024), .Z(n7018) );
  AND U6831 ( .A(n459), .B(n7025), .Z(n7024) );
  XOR U6832 ( .A(p_input[1178]), .B(n7023), .Z(n7025) );
  XNOR U6833 ( .A(n7026), .B(n7027), .Z(n7023) );
  AND U6834 ( .A(n463), .B(n7022), .Z(n7027) );
  XNOR U6835 ( .A(n7026), .B(n7020), .Z(n7022) );
  XOR U6836 ( .A(n7028), .B(n7029), .Z(n7020) );
  AND U6837 ( .A(n478), .B(n7030), .Z(n7029) );
  XNOR U6838 ( .A(n7031), .B(n7032), .Z(n7026) );
  AND U6839 ( .A(n470), .B(n7033), .Z(n7032) );
  XOR U6840 ( .A(p_input[1210]), .B(n7031), .Z(n7033) );
  XNOR U6841 ( .A(n7034), .B(n7035), .Z(n7031) );
  AND U6842 ( .A(n474), .B(n7030), .Z(n7035) );
  XNOR U6843 ( .A(n7034), .B(n7028), .Z(n7030) );
  XOR U6844 ( .A(n7036), .B(n7037), .Z(n7028) );
  AND U6845 ( .A(n489), .B(n7038), .Z(n7037) );
  XNOR U6846 ( .A(n7039), .B(n7040), .Z(n7034) );
  AND U6847 ( .A(n481), .B(n7041), .Z(n7040) );
  XOR U6848 ( .A(p_input[1242]), .B(n7039), .Z(n7041) );
  XNOR U6849 ( .A(n7042), .B(n7043), .Z(n7039) );
  AND U6850 ( .A(n485), .B(n7038), .Z(n7043) );
  XNOR U6851 ( .A(n7042), .B(n7036), .Z(n7038) );
  XOR U6852 ( .A(n7044), .B(n7045), .Z(n7036) );
  AND U6853 ( .A(n500), .B(n7046), .Z(n7045) );
  XNOR U6854 ( .A(n7047), .B(n7048), .Z(n7042) );
  AND U6855 ( .A(n492), .B(n7049), .Z(n7048) );
  XOR U6856 ( .A(p_input[1274]), .B(n7047), .Z(n7049) );
  XNOR U6857 ( .A(n7050), .B(n7051), .Z(n7047) );
  AND U6858 ( .A(n496), .B(n7046), .Z(n7051) );
  XNOR U6859 ( .A(n7050), .B(n7044), .Z(n7046) );
  XOR U6860 ( .A(n7052), .B(n7053), .Z(n7044) );
  AND U6861 ( .A(n511), .B(n7054), .Z(n7053) );
  XNOR U6862 ( .A(n7055), .B(n7056), .Z(n7050) );
  AND U6863 ( .A(n503), .B(n7057), .Z(n7056) );
  XOR U6864 ( .A(p_input[1306]), .B(n7055), .Z(n7057) );
  XNOR U6865 ( .A(n7058), .B(n7059), .Z(n7055) );
  AND U6866 ( .A(n507), .B(n7054), .Z(n7059) );
  XNOR U6867 ( .A(n7058), .B(n7052), .Z(n7054) );
  XOR U6868 ( .A(n7060), .B(n7061), .Z(n7052) );
  AND U6869 ( .A(n522), .B(n7062), .Z(n7061) );
  XNOR U6870 ( .A(n7063), .B(n7064), .Z(n7058) );
  AND U6871 ( .A(n514), .B(n7065), .Z(n7064) );
  XOR U6872 ( .A(p_input[1338]), .B(n7063), .Z(n7065) );
  XNOR U6873 ( .A(n7066), .B(n7067), .Z(n7063) );
  AND U6874 ( .A(n518), .B(n7062), .Z(n7067) );
  XNOR U6875 ( .A(n7066), .B(n7060), .Z(n7062) );
  XOR U6876 ( .A(n7068), .B(n7069), .Z(n7060) );
  AND U6877 ( .A(n533), .B(n7070), .Z(n7069) );
  XNOR U6878 ( .A(n7071), .B(n7072), .Z(n7066) );
  AND U6879 ( .A(n525), .B(n7073), .Z(n7072) );
  XOR U6880 ( .A(p_input[1370]), .B(n7071), .Z(n7073) );
  XNOR U6881 ( .A(n7074), .B(n7075), .Z(n7071) );
  AND U6882 ( .A(n529), .B(n7070), .Z(n7075) );
  XNOR U6883 ( .A(n7074), .B(n7068), .Z(n7070) );
  XOR U6884 ( .A(n7076), .B(n7077), .Z(n7068) );
  AND U6885 ( .A(n544), .B(n7078), .Z(n7077) );
  XNOR U6886 ( .A(n7079), .B(n7080), .Z(n7074) );
  AND U6887 ( .A(n536), .B(n7081), .Z(n7080) );
  XOR U6888 ( .A(p_input[1402]), .B(n7079), .Z(n7081) );
  XNOR U6889 ( .A(n7082), .B(n7083), .Z(n7079) );
  AND U6890 ( .A(n540), .B(n7078), .Z(n7083) );
  XNOR U6891 ( .A(n7082), .B(n7076), .Z(n7078) );
  XOR U6892 ( .A(n7084), .B(n7085), .Z(n7076) );
  AND U6893 ( .A(n555), .B(n7086), .Z(n7085) );
  XNOR U6894 ( .A(n7087), .B(n7088), .Z(n7082) );
  AND U6895 ( .A(n547), .B(n7089), .Z(n7088) );
  XOR U6896 ( .A(p_input[1434]), .B(n7087), .Z(n7089) );
  XNOR U6897 ( .A(n7090), .B(n7091), .Z(n7087) );
  AND U6898 ( .A(n551), .B(n7086), .Z(n7091) );
  XNOR U6899 ( .A(n7090), .B(n7084), .Z(n7086) );
  XOR U6900 ( .A(n7092), .B(n7093), .Z(n7084) );
  AND U6901 ( .A(n566), .B(n7094), .Z(n7093) );
  XNOR U6902 ( .A(n7095), .B(n7096), .Z(n7090) );
  AND U6903 ( .A(n558), .B(n7097), .Z(n7096) );
  XOR U6904 ( .A(p_input[1466]), .B(n7095), .Z(n7097) );
  XNOR U6905 ( .A(n7098), .B(n7099), .Z(n7095) );
  AND U6906 ( .A(n562), .B(n7094), .Z(n7099) );
  XNOR U6907 ( .A(n7098), .B(n7092), .Z(n7094) );
  XOR U6908 ( .A(n7100), .B(n7101), .Z(n7092) );
  AND U6909 ( .A(n577), .B(n7102), .Z(n7101) );
  XNOR U6910 ( .A(n7103), .B(n7104), .Z(n7098) );
  AND U6911 ( .A(n569), .B(n7105), .Z(n7104) );
  XOR U6912 ( .A(p_input[1498]), .B(n7103), .Z(n7105) );
  XNOR U6913 ( .A(n7106), .B(n7107), .Z(n7103) );
  AND U6914 ( .A(n573), .B(n7102), .Z(n7107) );
  XNOR U6915 ( .A(n7106), .B(n7100), .Z(n7102) );
  XOR U6916 ( .A(n7108), .B(n7109), .Z(n7100) );
  AND U6917 ( .A(n588), .B(n7110), .Z(n7109) );
  XNOR U6918 ( .A(n7111), .B(n7112), .Z(n7106) );
  AND U6919 ( .A(n580), .B(n7113), .Z(n7112) );
  XOR U6920 ( .A(p_input[1530]), .B(n7111), .Z(n7113) );
  XNOR U6921 ( .A(n7114), .B(n7115), .Z(n7111) );
  AND U6922 ( .A(n584), .B(n7110), .Z(n7115) );
  XNOR U6923 ( .A(n7114), .B(n7108), .Z(n7110) );
  XOR U6924 ( .A(n7116), .B(n7117), .Z(n7108) );
  AND U6925 ( .A(n599), .B(n7118), .Z(n7117) );
  XNOR U6926 ( .A(n7119), .B(n7120), .Z(n7114) );
  AND U6927 ( .A(n591), .B(n7121), .Z(n7120) );
  XOR U6928 ( .A(p_input[1562]), .B(n7119), .Z(n7121) );
  XNOR U6929 ( .A(n7122), .B(n7123), .Z(n7119) );
  AND U6930 ( .A(n595), .B(n7118), .Z(n7123) );
  XNOR U6931 ( .A(n7122), .B(n7116), .Z(n7118) );
  XOR U6932 ( .A(n7124), .B(n7125), .Z(n7116) );
  AND U6933 ( .A(n610), .B(n7126), .Z(n7125) );
  XNOR U6934 ( .A(n7127), .B(n7128), .Z(n7122) );
  AND U6935 ( .A(n602), .B(n7129), .Z(n7128) );
  XOR U6936 ( .A(p_input[1594]), .B(n7127), .Z(n7129) );
  XNOR U6937 ( .A(n7130), .B(n7131), .Z(n7127) );
  AND U6938 ( .A(n606), .B(n7126), .Z(n7131) );
  XNOR U6939 ( .A(n7130), .B(n7124), .Z(n7126) );
  XOR U6940 ( .A(n7132), .B(n7133), .Z(n7124) );
  AND U6941 ( .A(n621), .B(n7134), .Z(n7133) );
  XNOR U6942 ( .A(n7135), .B(n7136), .Z(n7130) );
  AND U6943 ( .A(n613), .B(n7137), .Z(n7136) );
  XOR U6944 ( .A(p_input[1626]), .B(n7135), .Z(n7137) );
  XNOR U6945 ( .A(n7138), .B(n7139), .Z(n7135) );
  AND U6946 ( .A(n617), .B(n7134), .Z(n7139) );
  XNOR U6947 ( .A(n7138), .B(n7132), .Z(n7134) );
  XOR U6948 ( .A(n7140), .B(n7141), .Z(n7132) );
  AND U6949 ( .A(n632), .B(n7142), .Z(n7141) );
  XNOR U6950 ( .A(n7143), .B(n7144), .Z(n7138) );
  AND U6951 ( .A(n624), .B(n7145), .Z(n7144) );
  XOR U6952 ( .A(p_input[1658]), .B(n7143), .Z(n7145) );
  XNOR U6953 ( .A(n7146), .B(n7147), .Z(n7143) );
  AND U6954 ( .A(n628), .B(n7142), .Z(n7147) );
  XNOR U6955 ( .A(n7146), .B(n7140), .Z(n7142) );
  XOR U6956 ( .A(n7148), .B(n7149), .Z(n7140) );
  AND U6957 ( .A(n643), .B(n7150), .Z(n7149) );
  XNOR U6958 ( .A(n7151), .B(n7152), .Z(n7146) );
  AND U6959 ( .A(n635), .B(n7153), .Z(n7152) );
  XOR U6960 ( .A(p_input[1690]), .B(n7151), .Z(n7153) );
  XNOR U6961 ( .A(n7154), .B(n7155), .Z(n7151) );
  AND U6962 ( .A(n639), .B(n7150), .Z(n7155) );
  XNOR U6963 ( .A(n7154), .B(n7148), .Z(n7150) );
  XOR U6964 ( .A(n7156), .B(n7157), .Z(n7148) );
  AND U6965 ( .A(n654), .B(n7158), .Z(n7157) );
  XNOR U6966 ( .A(n7159), .B(n7160), .Z(n7154) );
  AND U6967 ( .A(n646), .B(n7161), .Z(n7160) );
  XOR U6968 ( .A(p_input[1722]), .B(n7159), .Z(n7161) );
  XNOR U6969 ( .A(n7162), .B(n7163), .Z(n7159) );
  AND U6970 ( .A(n650), .B(n7158), .Z(n7163) );
  XNOR U6971 ( .A(n7162), .B(n7156), .Z(n7158) );
  XOR U6972 ( .A(n7164), .B(n7165), .Z(n7156) );
  AND U6973 ( .A(n665), .B(n7166), .Z(n7165) );
  XNOR U6974 ( .A(n7167), .B(n7168), .Z(n7162) );
  AND U6975 ( .A(n657), .B(n7169), .Z(n7168) );
  XOR U6976 ( .A(p_input[1754]), .B(n7167), .Z(n7169) );
  XNOR U6977 ( .A(n7170), .B(n7171), .Z(n7167) );
  AND U6978 ( .A(n661), .B(n7166), .Z(n7171) );
  XNOR U6979 ( .A(n7170), .B(n7164), .Z(n7166) );
  XOR U6980 ( .A(n7172), .B(n7173), .Z(n7164) );
  AND U6981 ( .A(n676), .B(n7174), .Z(n7173) );
  XNOR U6982 ( .A(n7175), .B(n7176), .Z(n7170) );
  AND U6983 ( .A(n668), .B(n7177), .Z(n7176) );
  XOR U6984 ( .A(p_input[1786]), .B(n7175), .Z(n7177) );
  XNOR U6985 ( .A(n7178), .B(n7179), .Z(n7175) );
  AND U6986 ( .A(n672), .B(n7174), .Z(n7179) );
  XNOR U6987 ( .A(n7178), .B(n7172), .Z(n7174) );
  XOR U6988 ( .A(n7180), .B(n7181), .Z(n7172) );
  AND U6989 ( .A(n687), .B(n7182), .Z(n7181) );
  XNOR U6990 ( .A(n7183), .B(n7184), .Z(n7178) );
  AND U6991 ( .A(n679), .B(n7185), .Z(n7184) );
  XOR U6992 ( .A(p_input[1818]), .B(n7183), .Z(n7185) );
  XNOR U6993 ( .A(n7186), .B(n7187), .Z(n7183) );
  AND U6994 ( .A(n683), .B(n7182), .Z(n7187) );
  XNOR U6995 ( .A(n7186), .B(n7180), .Z(n7182) );
  XOR U6996 ( .A(n7188), .B(n7189), .Z(n7180) );
  AND U6997 ( .A(n698), .B(n7190), .Z(n7189) );
  XNOR U6998 ( .A(n7191), .B(n7192), .Z(n7186) );
  AND U6999 ( .A(n690), .B(n7193), .Z(n7192) );
  XOR U7000 ( .A(p_input[1850]), .B(n7191), .Z(n7193) );
  XNOR U7001 ( .A(n7194), .B(n7195), .Z(n7191) );
  AND U7002 ( .A(n694), .B(n7190), .Z(n7195) );
  XNOR U7003 ( .A(n7194), .B(n7188), .Z(n7190) );
  XOR U7004 ( .A(n7196), .B(n7197), .Z(n7188) );
  AND U7005 ( .A(n709), .B(n7198), .Z(n7197) );
  XNOR U7006 ( .A(n7199), .B(n7200), .Z(n7194) );
  AND U7007 ( .A(n701), .B(n7201), .Z(n7200) );
  XOR U7008 ( .A(p_input[1882]), .B(n7199), .Z(n7201) );
  XNOR U7009 ( .A(n7202), .B(n7203), .Z(n7199) );
  AND U7010 ( .A(n705), .B(n7198), .Z(n7203) );
  XNOR U7011 ( .A(n7202), .B(n7196), .Z(n7198) );
  XOR U7012 ( .A(n7204), .B(n7205), .Z(n7196) );
  AND U7013 ( .A(n720), .B(n7206), .Z(n7205) );
  XNOR U7014 ( .A(n7207), .B(n7208), .Z(n7202) );
  AND U7015 ( .A(n712), .B(n7209), .Z(n7208) );
  XOR U7016 ( .A(p_input[1914]), .B(n7207), .Z(n7209) );
  XNOR U7017 ( .A(n7210), .B(n7211), .Z(n7207) );
  AND U7018 ( .A(n716), .B(n7206), .Z(n7211) );
  XNOR U7019 ( .A(n7210), .B(n7204), .Z(n7206) );
  XOR U7020 ( .A(n7212), .B(n7213), .Z(n7204) );
  AND U7021 ( .A(n731), .B(n7214), .Z(n7213) );
  XNOR U7022 ( .A(n7215), .B(n7216), .Z(n7210) );
  AND U7023 ( .A(n723), .B(n7217), .Z(n7216) );
  XOR U7024 ( .A(p_input[1946]), .B(n7215), .Z(n7217) );
  XNOR U7025 ( .A(n7218), .B(n7219), .Z(n7215) );
  AND U7026 ( .A(n727), .B(n7214), .Z(n7219) );
  XNOR U7027 ( .A(n7218), .B(n7212), .Z(n7214) );
  XOR U7028 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n7220), .Z(n7212) );
  AND U7029 ( .A(n741), .B(n7221), .Z(n7220) );
  XNOR U7030 ( .A(n7222), .B(n7223), .Z(n7218) );
  AND U7031 ( .A(n734), .B(n7224), .Z(n7223) );
  XOR U7032 ( .A(p_input[1978]), .B(n7222), .Z(n7224) );
  XNOR U7033 ( .A(n7225), .B(n7226), .Z(n7222) );
  AND U7034 ( .A(n738), .B(n7221), .Z(n7226) );
  XOR U7035 ( .A(\knn_comb_/min_val_out[0][26] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .Z(n7221) );
  XOR U7036 ( .A(n23), .B(n7227), .Z(o[25]) );
  AND U7037 ( .A(n58), .B(n7228), .Z(n23) );
  XOR U7038 ( .A(n24), .B(n7227), .Z(n7228) );
  XOR U7039 ( .A(n7229), .B(n7230), .Z(n7227) );
  AND U7040 ( .A(n70), .B(n7231), .Z(n7230) );
  XOR U7041 ( .A(n7232), .B(n7233), .Z(n24) );
  AND U7042 ( .A(n62), .B(n7234), .Z(n7233) );
  XOR U7043 ( .A(p_input[25]), .B(n7232), .Z(n7234) );
  XNOR U7044 ( .A(n7235), .B(n7236), .Z(n7232) );
  AND U7045 ( .A(n66), .B(n7231), .Z(n7236) );
  XNOR U7046 ( .A(n7235), .B(n7229), .Z(n7231) );
  XOR U7047 ( .A(n7237), .B(n7238), .Z(n7229) );
  AND U7048 ( .A(n82), .B(n7239), .Z(n7238) );
  XNOR U7049 ( .A(n7240), .B(n7241), .Z(n7235) );
  AND U7050 ( .A(n74), .B(n7242), .Z(n7241) );
  XOR U7051 ( .A(p_input[57]), .B(n7240), .Z(n7242) );
  XNOR U7052 ( .A(n7243), .B(n7244), .Z(n7240) );
  AND U7053 ( .A(n78), .B(n7239), .Z(n7244) );
  XNOR U7054 ( .A(n7243), .B(n7237), .Z(n7239) );
  XOR U7055 ( .A(n7245), .B(n7246), .Z(n7237) );
  AND U7056 ( .A(n93), .B(n7247), .Z(n7246) );
  XNOR U7057 ( .A(n7248), .B(n7249), .Z(n7243) );
  AND U7058 ( .A(n85), .B(n7250), .Z(n7249) );
  XOR U7059 ( .A(p_input[89]), .B(n7248), .Z(n7250) );
  XNOR U7060 ( .A(n7251), .B(n7252), .Z(n7248) );
  AND U7061 ( .A(n89), .B(n7247), .Z(n7252) );
  XNOR U7062 ( .A(n7251), .B(n7245), .Z(n7247) );
  XOR U7063 ( .A(n7253), .B(n7254), .Z(n7245) );
  AND U7064 ( .A(n104), .B(n7255), .Z(n7254) );
  XNOR U7065 ( .A(n7256), .B(n7257), .Z(n7251) );
  AND U7066 ( .A(n96), .B(n7258), .Z(n7257) );
  XOR U7067 ( .A(p_input[121]), .B(n7256), .Z(n7258) );
  XNOR U7068 ( .A(n7259), .B(n7260), .Z(n7256) );
  AND U7069 ( .A(n100), .B(n7255), .Z(n7260) );
  XNOR U7070 ( .A(n7259), .B(n7253), .Z(n7255) );
  XOR U7071 ( .A(n7261), .B(n7262), .Z(n7253) );
  AND U7072 ( .A(n115), .B(n7263), .Z(n7262) );
  XNOR U7073 ( .A(n7264), .B(n7265), .Z(n7259) );
  AND U7074 ( .A(n107), .B(n7266), .Z(n7265) );
  XOR U7075 ( .A(p_input[153]), .B(n7264), .Z(n7266) );
  XNOR U7076 ( .A(n7267), .B(n7268), .Z(n7264) );
  AND U7077 ( .A(n111), .B(n7263), .Z(n7268) );
  XNOR U7078 ( .A(n7267), .B(n7261), .Z(n7263) );
  XOR U7079 ( .A(n7269), .B(n7270), .Z(n7261) );
  AND U7080 ( .A(n126), .B(n7271), .Z(n7270) );
  XNOR U7081 ( .A(n7272), .B(n7273), .Z(n7267) );
  AND U7082 ( .A(n118), .B(n7274), .Z(n7273) );
  XOR U7083 ( .A(p_input[185]), .B(n7272), .Z(n7274) );
  XNOR U7084 ( .A(n7275), .B(n7276), .Z(n7272) );
  AND U7085 ( .A(n122), .B(n7271), .Z(n7276) );
  XNOR U7086 ( .A(n7275), .B(n7269), .Z(n7271) );
  XOR U7087 ( .A(n7277), .B(n7278), .Z(n7269) );
  AND U7088 ( .A(n137), .B(n7279), .Z(n7278) );
  XNOR U7089 ( .A(n7280), .B(n7281), .Z(n7275) );
  AND U7090 ( .A(n129), .B(n7282), .Z(n7281) );
  XOR U7091 ( .A(p_input[217]), .B(n7280), .Z(n7282) );
  XNOR U7092 ( .A(n7283), .B(n7284), .Z(n7280) );
  AND U7093 ( .A(n133), .B(n7279), .Z(n7284) );
  XNOR U7094 ( .A(n7283), .B(n7277), .Z(n7279) );
  XOR U7095 ( .A(n7285), .B(n7286), .Z(n7277) );
  AND U7096 ( .A(n148), .B(n7287), .Z(n7286) );
  XNOR U7097 ( .A(n7288), .B(n7289), .Z(n7283) );
  AND U7098 ( .A(n140), .B(n7290), .Z(n7289) );
  XOR U7099 ( .A(p_input[249]), .B(n7288), .Z(n7290) );
  XNOR U7100 ( .A(n7291), .B(n7292), .Z(n7288) );
  AND U7101 ( .A(n144), .B(n7287), .Z(n7292) );
  XNOR U7102 ( .A(n7291), .B(n7285), .Z(n7287) );
  XOR U7103 ( .A(n7293), .B(n7294), .Z(n7285) );
  AND U7104 ( .A(n159), .B(n7295), .Z(n7294) );
  XNOR U7105 ( .A(n7296), .B(n7297), .Z(n7291) );
  AND U7106 ( .A(n151), .B(n7298), .Z(n7297) );
  XOR U7107 ( .A(p_input[281]), .B(n7296), .Z(n7298) );
  XNOR U7108 ( .A(n7299), .B(n7300), .Z(n7296) );
  AND U7109 ( .A(n155), .B(n7295), .Z(n7300) );
  XNOR U7110 ( .A(n7299), .B(n7293), .Z(n7295) );
  XOR U7111 ( .A(n7301), .B(n7302), .Z(n7293) );
  AND U7112 ( .A(n170), .B(n7303), .Z(n7302) );
  XNOR U7113 ( .A(n7304), .B(n7305), .Z(n7299) );
  AND U7114 ( .A(n162), .B(n7306), .Z(n7305) );
  XOR U7115 ( .A(p_input[313]), .B(n7304), .Z(n7306) );
  XNOR U7116 ( .A(n7307), .B(n7308), .Z(n7304) );
  AND U7117 ( .A(n166), .B(n7303), .Z(n7308) );
  XNOR U7118 ( .A(n7307), .B(n7301), .Z(n7303) );
  XOR U7119 ( .A(n7309), .B(n7310), .Z(n7301) );
  AND U7120 ( .A(n181), .B(n7311), .Z(n7310) );
  XNOR U7121 ( .A(n7312), .B(n7313), .Z(n7307) );
  AND U7122 ( .A(n173), .B(n7314), .Z(n7313) );
  XOR U7123 ( .A(p_input[345]), .B(n7312), .Z(n7314) );
  XNOR U7124 ( .A(n7315), .B(n7316), .Z(n7312) );
  AND U7125 ( .A(n177), .B(n7311), .Z(n7316) );
  XNOR U7126 ( .A(n7315), .B(n7309), .Z(n7311) );
  XOR U7127 ( .A(n7317), .B(n7318), .Z(n7309) );
  AND U7128 ( .A(n192), .B(n7319), .Z(n7318) );
  XNOR U7129 ( .A(n7320), .B(n7321), .Z(n7315) );
  AND U7130 ( .A(n184), .B(n7322), .Z(n7321) );
  XOR U7131 ( .A(p_input[377]), .B(n7320), .Z(n7322) );
  XNOR U7132 ( .A(n7323), .B(n7324), .Z(n7320) );
  AND U7133 ( .A(n188), .B(n7319), .Z(n7324) );
  XNOR U7134 ( .A(n7323), .B(n7317), .Z(n7319) );
  XOR U7135 ( .A(n7325), .B(n7326), .Z(n7317) );
  AND U7136 ( .A(n203), .B(n7327), .Z(n7326) );
  XNOR U7137 ( .A(n7328), .B(n7329), .Z(n7323) );
  AND U7138 ( .A(n195), .B(n7330), .Z(n7329) );
  XOR U7139 ( .A(p_input[409]), .B(n7328), .Z(n7330) );
  XNOR U7140 ( .A(n7331), .B(n7332), .Z(n7328) );
  AND U7141 ( .A(n199), .B(n7327), .Z(n7332) );
  XNOR U7142 ( .A(n7331), .B(n7325), .Z(n7327) );
  XOR U7143 ( .A(n7333), .B(n7334), .Z(n7325) );
  AND U7144 ( .A(n214), .B(n7335), .Z(n7334) );
  XNOR U7145 ( .A(n7336), .B(n7337), .Z(n7331) );
  AND U7146 ( .A(n206), .B(n7338), .Z(n7337) );
  XOR U7147 ( .A(p_input[441]), .B(n7336), .Z(n7338) );
  XNOR U7148 ( .A(n7339), .B(n7340), .Z(n7336) );
  AND U7149 ( .A(n210), .B(n7335), .Z(n7340) );
  XNOR U7150 ( .A(n7339), .B(n7333), .Z(n7335) );
  XOR U7151 ( .A(n7341), .B(n7342), .Z(n7333) );
  AND U7152 ( .A(n225), .B(n7343), .Z(n7342) );
  XNOR U7153 ( .A(n7344), .B(n7345), .Z(n7339) );
  AND U7154 ( .A(n217), .B(n7346), .Z(n7345) );
  XOR U7155 ( .A(p_input[473]), .B(n7344), .Z(n7346) );
  XNOR U7156 ( .A(n7347), .B(n7348), .Z(n7344) );
  AND U7157 ( .A(n221), .B(n7343), .Z(n7348) );
  XNOR U7158 ( .A(n7347), .B(n7341), .Z(n7343) );
  XOR U7159 ( .A(n7349), .B(n7350), .Z(n7341) );
  AND U7160 ( .A(n236), .B(n7351), .Z(n7350) );
  XNOR U7161 ( .A(n7352), .B(n7353), .Z(n7347) );
  AND U7162 ( .A(n228), .B(n7354), .Z(n7353) );
  XOR U7163 ( .A(p_input[505]), .B(n7352), .Z(n7354) );
  XNOR U7164 ( .A(n7355), .B(n7356), .Z(n7352) );
  AND U7165 ( .A(n232), .B(n7351), .Z(n7356) );
  XNOR U7166 ( .A(n7355), .B(n7349), .Z(n7351) );
  XOR U7167 ( .A(n7357), .B(n7358), .Z(n7349) );
  AND U7168 ( .A(n247), .B(n7359), .Z(n7358) );
  XNOR U7169 ( .A(n7360), .B(n7361), .Z(n7355) );
  AND U7170 ( .A(n239), .B(n7362), .Z(n7361) );
  XOR U7171 ( .A(p_input[537]), .B(n7360), .Z(n7362) );
  XNOR U7172 ( .A(n7363), .B(n7364), .Z(n7360) );
  AND U7173 ( .A(n243), .B(n7359), .Z(n7364) );
  XNOR U7174 ( .A(n7363), .B(n7357), .Z(n7359) );
  XOR U7175 ( .A(n7365), .B(n7366), .Z(n7357) );
  AND U7176 ( .A(n258), .B(n7367), .Z(n7366) );
  XNOR U7177 ( .A(n7368), .B(n7369), .Z(n7363) );
  AND U7178 ( .A(n250), .B(n7370), .Z(n7369) );
  XOR U7179 ( .A(p_input[569]), .B(n7368), .Z(n7370) );
  XNOR U7180 ( .A(n7371), .B(n7372), .Z(n7368) );
  AND U7181 ( .A(n254), .B(n7367), .Z(n7372) );
  XNOR U7182 ( .A(n7371), .B(n7365), .Z(n7367) );
  XOR U7183 ( .A(n7373), .B(n7374), .Z(n7365) );
  AND U7184 ( .A(n269), .B(n7375), .Z(n7374) );
  XNOR U7185 ( .A(n7376), .B(n7377), .Z(n7371) );
  AND U7186 ( .A(n261), .B(n7378), .Z(n7377) );
  XOR U7187 ( .A(p_input[601]), .B(n7376), .Z(n7378) );
  XNOR U7188 ( .A(n7379), .B(n7380), .Z(n7376) );
  AND U7189 ( .A(n265), .B(n7375), .Z(n7380) );
  XNOR U7190 ( .A(n7379), .B(n7373), .Z(n7375) );
  XOR U7191 ( .A(n7381), .B(n7382), .Z(n7373) );
  AND U7192 ( .A(n280), .B(n7383), .Z(n7382) );
  XNOR U7193 ( .A(n7384), .B(n7385), .Z(n7379) );
  AND U7194 ( .A(n272), .B(n7386), .Z(n7385) );
  XOR U7195 ( .A(p_input[633]), .B(n7384), .Z(n7386) );
  XNOR U7196 ( .A(n7387), .B(n7388), .Z(n7384) );
  AND U7197 ( .A(n276), .B(n7383), .Z(n7388) );
  XNOR U7198 ( .A(n7387), .B(n7381), .Z(n7383) );
  XOR U7199 ( .A(n7389), .B(n7390), .Z(n7381) );
  AND U7200 ( .A(n291), .B(n7391), .Z(n7390) );
  XNOR U7201 ( .A(n7392), .B(n7393), .Z(n7387) );
  AND U7202 ( .A(n283), .B(n7394), .Z(n7393) );
  XOR U7203 ( .A(p_input[665]), .B(n7392), .Z(n7394) );
  XNOR U7204 ( .A(n7395), .B(n7396), .Z(n7392) );
  AND U7205 ( .A(n287), .B(n7391), .Z(n7396) );
  XNOR U7206 ( .A(n7395), .B(n7389), .Z(n7391) );
  XOR U7207 ( .A(n7397), .B(n7398), .Z(n7389) );
  AND U7208 ( .A(n302), .B(n7399), .Z(n7398) );
  XNOR U7209 ( .A(n7400), .B(n7401), .Z(n7395) );
  AND U7210 ( .A(n294), .B(n7402), .Z(n7401) );
  XOR U7211 ( .A(p_input[697]), .B(n7400), .Z(n7402) );
  XNOR U7212 ( .A(n7403), .B(n7404), .Z(n7400) );
  AND U7213 ( .A(n298), .B(n7399), .Z(n7404) );
  XNOR U7214 ( .A(n7403), .B(n7397), .Z(n7399) );
  XOR U7215 ( .A(n7405), .B(n7406), .Z(n7397) );
  AND U7216 ( .A(n313), .B(n7407), .Z(n7406) );
  XNOR U7217 ( .A(n7408), .B(n7409), .Z(n7403) );
  AND U7218 ( .A(n305), .B(n7410), .Z(n7409) );
  XOR U7219 ( .A(p_input[729]), .B(n7408), .Z(n7410) );
  XNOR U7220 ( .A(n7411), .B(n7412), .Z(n7408) );
  AND U7221 ( .A(n309), .B(n7407), .Z(n7412) );
  XNOR U7222 ( .A(n7411), .B(n7405), .Z(n7407) );
  XOR U7223 ( .A(n7413), .B(n7414), .Z(n7405) );
  AND U7224 ( .A(n324), .B(n7415), .Z(n7414) );
  XNOR U7225 ( .A(n7416), .B(n7417), .Z(n7411) );
  AND U7226 ( .A(n316), .B(n7418), .Z(n7417) );
  XOR U7227 ( .A(p_input[761]), .B(n7416), .Z(n7418) );
  XNOR U7228 ( .A(n7419), .B(n7420), .Z(n7416) );
  AND U7229 ( .A(n320), .B(n7415), .Z(n7420) );
  XNOR U7230 ( .A(n7419), .B(n7413), .Z(n7415) );
  XOR U7231 ( .A(n7421), .B(n7422), .Z(n7413) );
  AND U7232 ( .A(n335), .B(n7423), .Z(n7422) );
  XNOR U7233 ( .A(n7424), .B(n7425), .Z(n7419) );
  AND U7234 ( .A(n327), .B(n7426), .Z(n7425) );
  XOR U7235 ( .A(p_input[793]), .B(n7424), .Z(n7426) );
  XNOR U7236 ( .A(n7427), .B(n7428), .Z(n7424) );
  AND U7237 ( .A(n331), .B(n7423), .Z(n7428) );
  XNOR U7238 ( .A(n7427), .B(n7421), .Z(n7423) );
  XOR U7239 ( .A(n7429), .B(n7430), .Z(n7421) );
  AND U7240 ( .A(n346), .B(n7431), .Z(n7430) );
  XNOR U7241 ( .A(n7432), .B(n7433), .Z(n7427) );
  AND U7242 ( .A(n338), .B(n7434), .Z(n7433) );
  XOR U7243 ( .A(p_input[825]), .B(n7432), .Z(n7434) );
  XNOR U7244 ( .A(n7435), .B(n7436), .Z(n7432) );
  AND U7245 ( .A(n342), .B(n7431), .Z(n7436) );
  XNOR U7246 ( .A(n7435), .B(n7429), .Z(n7431) );
  XOR U7247 ( .A(n7437), .B(n7438), .Z(n7429) );
  AND U7248 ( .A(n357), .B(n7439), .Z(n7438) );
  XNOR U7249 ( .A(n7440), .B(n7441), .Z(n7435) );
  AND U7250 ( .A(n349), .B(n7442), .Z(n7441) );
  XOR U7251 ( .A(p_input[857]), .B(n7440), .Z(n7442) );
  XNOR U7252 ( .A(n7443), .B(n7444), .Z(n7440) );
  AND U7253 ( .A(n353), .B(n7439), .Z(n7444) );
  XNOR U7254 ( .A(n7443), .B(n7437), .Z(n7439) );
  XOR U7255 ( .A(n7445), .B(n7446), .Z(n7437) );
  AND U7256 ( .A(n368), .B(n7447), .Z(n7446) );
  XNOR U7257 ( .A(n7448), .B(n7449), .Z(n7443) );
  AND U7258 ( .A(n360), .B(n7450), .Z(n7449) );
  XOR U7259 ( .A(p_input[889]), .B(n7448), .Z(n7450) );
  XNOR U7260 ( .A(n7451), .B(n7452), .Z(n7448) );
  AND U7261 ( .A(n364), .B(n7447), .Z(n7452) );
  XNOR U7262 ( .A(n7451), .B(n7445), .Z(n7447) );
  XOR U7263 ( .A(n7453), .B(n7454), .Z(n7445) );
  AND U7264 ( .A(n379), .B(n7455), .Z(n7454) );
  XNOR U7265 ( .A(n7456), .B(n7457), .Z(n7451) );
  AND U7266 ( .A(n371), .B(n7458), .Z(n7457) );
  XOR U7267 ( .A(p_input[921]), .B(n7456), .Z(n7458) );
  XNOR U7268 ( .A(n7459), .B(n7460), .Z(n7456) );
  AND U7269 ( .A(n375), .B(n7455), .Z(n7460) );
  XNOR U7270 ( .A(n7459), .B(n7453), .Z(n7455) );
  XOR U7271 ( .A(n7461), .B(n7462), .Z(n7453) );
  AND U7272 ( .A(n390), .B(n7463), .Z(n7462) );
  XNOR U7273 ( .A(n7464), .B(n7465), .Z(n7459) );
  AND U7274 ( .A(n382), .B(n7466), .Z(n7465) );
  XOR U7275 ( .A(p_input[953]), .B(n7464), .Z(n7466) );
  XNOR U7276 ( .A(n7467), .B(n7468), .Z(n7464) );
  AND U7277 ( .A(n386), .B(n7463), .Z(n7468) );
  XNOR U7278 ( .A(n7467), .B(n7461), .Z(n7463) );
  XOR U7279 ( .A(n7469), .B(n7470), .Z(n7461) );
  AND U7280 ( .A(n401), .B(n7471), .Z(n7470) );
  XNOR U7281 ( .A(n7472), .B(n7473), .Z(n7467) );
  AND U7282 ( .A(n393), .B(n7474), .Z(n7473) );
  XOR U7283 ( .A(p_input[985]), .B(n7472), .Z(n7474) );
  XNOR U7284 ( .A(n7475), .B(n7476), .Z(n7472) );
  AND U7285 ( .A(n397), .B(n7471), .Z(n7476) );
  XNOR U7286 ( .A(n7475), .B(n7469), .Z(n7471) );
  XOR U7287 ( .A(n7477), .B(n7478), .Z(n7469) );
  AND U7288 ( .A(n412), .B(n7479), .Z(n7478) );
  XNOR U7289 ( .A(n7480), .B(n7481), .Z(n7475) );
  AND U7290 ( .A(n404), .B(n7482), .Z(n7481) );
  XOR U7291 ( .A(p_input[1017]), .B(n7480), .Z(n7482) );
  XNOR U7292 ( .A(n7483), .B(n7484), .Z(n7480) );
  AND U7293 ( .A(n408), .B(n7479), .Z(n7484) );
  XNOR U7294 ( .A(n7483), .B(n7477), .Z(n7479) );
  XOR U7295 ( .A(n7485), .B(n7486), .Z(n7477) );
  AND U7296 ( .A(n423), .B(n7487), .Z(n7486) );
  XNOR U7297 ( .A(n7488), .B(n7489), .Z(n7483) );
  AND U7298 ( .A(n415), .B(n7490), .Z(n7489) );
  XOR U7299 ( .A(p_input[1049]), .B(n7488), .Z(n7490) );
  XNOR U7300 ( .A(n7491), .B(n7492), .Z(n7488) );
  AND U7301 ( .A(n419), .B(n7487), .Z(n7492) );
  XNOR U7302 ( .A(n7491), .B(n7485), .Z(n7487) );
  XOR U7303 ( .A(n7493), .B(n7494), .Z(n7485) );
  AND U7304 ( .A(n434), .B(n7495), .Z(n7494) );
  XNOR U7305 ( .A(n7496), .B(n7497), .Z(n7491) );
  AND U7306 ( .A(n426), .B(n7498), .Z(n7497) );
  XOR U7307 ( .A(p_input[1081]), .B(n7496), .Z(n7498) );
  XNOR U7308 ( .A(n7499), .B(n7500), .Z(n7496) );
  AND U7309 ( .A(n430), .B(n7495), .Z(n7500) );
  XNOR U7310 ( .A(n7499), .B(n7493), .Z(n7495) );
  XOR U7311 ( .A(n7501), .B(n7502), .Z(n7493) );
  AND U7312 ( .A(n445), .B(n7503), .Z(n7502) );
  XNOR U7313 ( .A(n7504), .B(n7505), .Z(n7499) );
  AND U7314 ( .A(n437), .B(n7506), .Z(n7505) );
  XOR U7315 ( .A(p_input[1113]), .B(n7504), .Z(n7506) );
  XNOR U7316 ( .A(n7507), .B(n7508), .Z(n7504) );
  AND U7317 ( .A(n441), .B(n7503), .Z(n7508) );
  XNOR U7318 ( .A(n7507), .B(n7501), .Z(n7503) );
  XOR U7319 ( .A(n7509), .B(n7510), .Z(n7501) );
  AND U7320 ( .A(n456), .B(n7511), .Z(n7510) );
  XNOR U7321 ( .A(n7512), .B(n7513), .Z(n7507) );
  AND U7322 ( .A(n448), .B(n7514), .Z(n7513) );
  XOR U7323 ( .A(p_input[1145]), .B(n7512), .Z(n7514) );
  XNOR U7324 ( .A(n7515), .B(n7516), .Z(n7512) );
  AND U7325 ( .A(n452), .B(n7511), .Z(n7516) );
  XNOR U7326 ( .A(n7515), .B(n7509), .Z(n7511) );
  XOR U7327 ( .A(n7517), .B(n7518), .Z(n7509) );
  AND U7328 ( .A(n467), .B(n7519), .Z(n7518) );
  XNOR U7329 ( .A(n7520), .B(n7521), .Z(n7515) );
  AND U7330 ( .A(n459), .B(n7522), .Z(n7521) );
  XOR U7331 ( .A(p_input[1177]), .B(n7520), .Z(n7522) );
  XNOR U7332 ( .A(n7523), .B(n7524), .Z(n7520) );
  AND U7333 ( .A(n463), .B(n7519), .Z(n7524) );
  XNOR U7334 ( .A(n7523), .B(n7517), .Z(n7519) );
  XOR U7335 ( .A(n7525), .B(n7526), .Z(n7517) );
  AND U7336 ( .A(n478), .B(n7527), .Z(n7526) );
  XNOR U7337 ( .A(n7528), .B(n7529), .Z(n7523) );
  AND U7338 ( .A(n470), .B(n7530), .Z(n7529) );
  XOR U7339 ( .A(p_input[1209]), .B(n7528), .Z(n7530) );
  XNOR U7340 ( .A(n7531), .B(n7532), .Z(n7528) );
  AND U7341 ( .A(n474), .B(n7527), .Z(n7532) );
  XNOR U7342 ( .A(n7531), .B(n7525), .Z(n7527) );
  XOR U7343 ( .A(n7533), .B(n7534), .Z(n7525) );
  AND U7344 ( .A(n489), .B(n7535), .Z(n7534) );
  XNOR U7345 ( .A(n7536), .B(n7537), .Z(n7531) );
  AND U7346 ( .A(n481), .B(n7538), .Z(n7537) );
  XOR U7347 ( .A(p_input[1241]), .B(n7536), .Z(n7538) );
  XNOR U7348 ( .A(n7539), .B(n7540), .Z(n7536) );
  AND U7349 ( .A(n485), .B(n7535), .Z(n7540) );
  XNOR U7350 ( .A(n7539), .B(n7533), .Z(n7535) );
  XOR U7351 ( .A(n7541), .B(n7542), .Z(n7533) );
  AND U7352 ( .A(n500), .B(n7543), .Z(n7542) );
  XNOR U7353 ( .A(n7544), .B(n7545), .Z(n7539) );
  AND U7354 ( .A(n492), .B(n7546), .Z(n7545) );
  XOR U7355 ( .A(p_input[1273]), .B(n7544), .Z(n7546) );
  XNOR U7356 ( .A(n7547), .B(n7548), .Z(n7544) );
  AND U7357 ( .A(n496), .B(n7543), .Z(n7548) );
  XNOR U7358 ( .A(n7547), .B(n7541), .Z(n7543) );
  XOR U7359 ( .A(n7549), .B(n7550), .Z(n7541) );
  AND U7360 ( .A(n511), .B(n7551), .Z(n7550) );
  XNOR U7361 ( .A(n7552), .B(n7553), .Z(n7547) );
  AND U7362 ( .A(n503), .B(n7554), .Z(n7553) );
  XOR U7363 ( .A(p_input[1305]), .B(n7552), .Z(n7554) );
  XNOR U7364 ( .A(n7555), .B(n7556), .Z(n7552) );
  AND U7365 ( .A(n507), .B(n7551), .Z(n7556) );
  XNOR U7366 ( .A(n7555), .B(n7549), .Z(n7551) );
  XOR U7367 ( .A(n7557), .B(n7558), .Z(n7549) );
  AND U7368 ( .A(n522), .B(n7559), .Z(n7558) );
  XNOR U7369 ( .A(n7560), .B(n7561), .Z(n7555) );
  AND U7370 ( .A(n514), .B(n7562), .Z(n7561) );
  XOR U7371 ( .A(p_input[1337]), .B(n7560), .Z(n7562) );
  XNOR U7372 ( .A(n7563), .B(n7564), .Z(n7560) );
  AND U7373 ( .A(n518), .B(n7559), .Z(n7564) );
  XNOR U7374 ( .A(n7563), .B(n7557), .Z(n7559) );
  XOR U7375 ( .A(n7565), .B(n7566), .Z(n7557) );
  AND U7376 ( .A(n533), .B(n7567), .Z(n7566) );
  XNOR U7377 ( .A(n7568), .B(n7569), .Z(n7563) );
  AND U7378 ( .A(n525), .B(n7570), .Z(n7569) );
  XOR U7379 ( .A(p_input[1369]), .B(n7568), .Z(n7570) );
  XNOR U7380 ( .A(n7571), .B(n7572), .Z(n7568) );
  AND U7381 ( .A(n529), .B(n7567), .Z(n7572) );
  XNOR U7382 ( .A(n7571), .B(n7565), .Z(n7567) );
  XOR U7383 ( .A(n7573), .B(n7574), .Z(n7565) );
  AND U7384 ( .A(n544), .B(n7575), .Z(n7574) );
  XNOR U7385 ( .A(n7576), .B(n7577), .Z(n7571) );
  AND U7386 ( .A(n536), .B(n7578), .Z(n7577) );
  XOR U7387 ( .A(p_input[1401]), .B(n7576), .Z(n7578) );
  XNOR U7388 ( .A(n7579), .B(n7580), .Z(n7576) );
  AND U7389 ( .A(n540), .B(n7575), .Z(n7580) );
  XNOR U7390 ( .A(n7579), .B(n7573), .Z(n7575) );
  XOR U7391 ( .A(n7581), .B(n7582), .Z(n7573) );
  AND U7392 ( .A(n555), .B(n7583), .Z(n7582) );
  XNOR U7393 ( .A(n7584), .B(n7585), .Z(n7579) );
  AND U7394 ( .A(n547), .B(n7586), .Z(n7585) );
  XOR U7395 ( .A(p_input[1433]), .B(n7584), .Z(n7586) );
  XNOR U7396 ( .A(n7587), .B(n7588), .Z(n7584) );
  AND U7397 ( .A(n551), .B(n7583), .Z(n7588) );
  XNOR U7398 ( .A(n7587), .B(n7581), .Z(n7583) );
  XOR U7399 ( .A(n7589), .B(n7590), .Z(n7581) );
  AND U7400 ( .A(n566), .B(n7591), .Z(n7590) );
  XNOR U7401 ( .A(n7592), .B(n7593), .Z(n7587) );
  AND U7402 ( .A(n558), .B(n7594), .Z(n7593) );
  XOR U7403 ( .A(p_input[1465]), .B(n7592), .Z(n7594) );
  XNOR U7404 ( .A(n7595), .B(n7596), .Z(n7592) );
  AND U7405 ( .A(n562), .B(n7591), .Z(n7596) );
  XNOR U7406 ( .A(n7595), .B(n7589), .Z(n7591) );
  XOR U7407 ( .A(n7597), .B(n7598), .Z(n7589) );
  AND U7408 ( .A(n577), .B(n7599), .Z(n7598) );
  XNOR U7409 ( .A(n7600), .B(n7601), .Z(n7595) );
  AND U7410 ( .A(n569), .B(n7602), .Z(n7601) );
  XOR U7411 ( .A(p_input[1497]), .B(n7600), .Z(n7602) );
  XNOR U7412 ( .A(n7603), .B(n7604), .Z(n7600) );
  AND U7413 ( .A(n573), .B(n7599), .Z(n7604) );
  XNOR U7414 ( .A(n7603), .B(n7597), .Z(n7599) );
  XOR U7415 ( .A(n7605), .B(n7606), .Z(n7597) );
  AND U7416 ( .A(n588), .B(n7607), .Z(n7606) );
  XNOR U7417 ( .A(n7608), .B(n7609), .Z(n7603) );
  AND U7418 ( .A(n580), .B(n7610), .Z(n7609) );
  XOR U7419 ( .A(p_input[1529]), .B(n7608), .Z(n7610) );
  XNOR U7420 ( .A(n7611), .B(n7612), .Z(n7608) );
  AND U7421 ( .A(n584), .B(n7607), .Z(n7612) );
  XNOR U7422 ( .A(n7611), .B(n7605), .Z(n7607) );
  XOR U7423 ( .A(n7613), .B(n7614), .Z(n7605) );
  AND U7424 ( .A(n599), .B(n7615), .Z(n7614) );
  XNOR U7425 ( .A(n7616), .B(n7617), .Z(n7611) );
  AND U7426 ( .A(n591), .B(n7618), .Z(n7617) );
  XOR U7427 ( .A(p_input[1561]), .B(n7616), .Z(n7618) );
  XNOR U7428 ( .A(n7619), .B(n7620), .Z(n7616) );
  AND U7429 ( .A(n595), .B(n7615), .Z(n7620) );
  XNOR U7430 ( .A(n7619), .B(n7613), .Z(n7615) );
  XOR U7431 ( .A(n7621), .B(n7622), .Z(n7613) );
  AND U7432 ( .A(n610), .B(n7623), .Z(n7622) );
  XNOR U7433 ( .A(n7624), .B(n7625), .Z(n7619) );
  AND U7434 ( .A(n602), .B(n7626), .Z(n7625) );
  XOR U7435 ( .A(p_input[1593]), .B(n7624), .Z(n7626) );
  XNOR U7436 ( .A(n7627), .B(n7628), .Z(n7624) );
  AND U7437 ( .A(n606), .B(n7623), .Z(n7628) );
  XNOR U7438 ( .A(n7627), .B(n7621), .Z(n7623) );
  XOR U7439 ( .A(n7629), .B(n7630), .Z(n7621) );
  AND U7440 ( .A(n621), .B(n7631), .Z(n7630) );
  XNOR U7441 ( .A(n7632), .B(n7633), .Z(n7627) );
  AND U7442 ( .A(n613), .B(n7634), .Z(n7633) );
  XOR U7443 ( .A(p_input[1625]), .B(n7632), .Z(n7634) );
  XNOR U7444 ( .A(n7635), .B(n7636), .Z(n7632) );
  AND U7445 ( .A(n617), .B(n7631), .Z(n7636) );
  XNOR U7446 ( .A(n7635), .B(n7629), .Z(n7631) );
  XOR U7447 ( .A(n7637), .B(n7638), .Z(n7629) );
  AND U7448 ( .A(n632), .B(n7639), .Z(n7638) );
  XNOR U7449 ( .A(n7640), .B(n7641), .Z(n7635) );
  AND U7450 ( .A(n624), .B(n7642), .Z(n7641) );
  XOR U7451 ( .A(p_input[1657]), .B(n7640), .Z(n7642) );
  XNOR U7452 ( .A(n7643), .B(n7644), .Z(n7640) );
  AND U7453 ( .A(n628), .B(n7639), .Z(n7644) );
  XNOR U7454 ( .A(n7643), .B(n7637), .Z(n7639) );
  XOR U7455 ( .A(n7645), .B(n7646), .Z(n7637) );
  AND U7456 ( .A(n643), .B(n7647), .Z(n7646) );
  XNOR U7457 ( .A(n7648), .B(n7649), .Z(n7643) );
  AND U7458 ( .A(n635), .B(n7650), .Z(n7649) );
  XOR U7459 ( .A(p_input[1689]), .B(n7648), .Z(n7650) );
  XNOR U7460 ( .A(n7651), .B(n7652), .Z(n7648) );
  AND U7461 ( .A(n639), .B(n7647), .Z(n7652) );
  XNOR U7462 ( .A(n7651), .B(n7645), .Z(n7647) );
  XOR U7463 ( .A(n7653), .B(n7654), .Z(n7645) );
  AND U7464 ( .A(n654), .B(n7655), .Z(n7654) );
  XNOR U7465 ( .A(n7656), .B(n7657), .Z(n7651) );
  AND U7466 ( .A(n646), .B(n7658), .Z(n7657) );
  XOR U7467 ( .A(p_input[1721]), .B(n7656), .Z(n7658) );
  XNOR U7468 ( .A(n7659), .B(n7660), .Z(n7656) );
  AND U7469 ( .A(n650), .B(n7655), .Z(n7660) );
  XNOR U7470 ( .A(n7659), .B(n7653), .Z(n7655) );
  XOR U7471 ( .A(n7661), .B(n7662), .Z(n7653) );
  AND U7472 ( .A(n665), .B(n7663), .Z(n7662) );
  XNOR U7473 ( .A(n7664), .B(n7665), .Z(n7659) );
  AND U7474 ( .A(n657), .B(n7666), .Z(n7665) );
  XOR U7475 ( .A(p_input[1753]), .B(n7664), .Z(n7666) );
  XNOR U7476 ( .A(n7667), .B(n7668), .Z(n7664) );
  AND U7477 ( .A(n661), .B(n7663), .Z(n7668) );
  XNOR U7478 ( .A(n7667), .B(n7661), .Z(n7663) );
  XOR U7479 ( .A(n7669), .B(n7670), .Z(n7661) );
  AND U7480 ( .A(n676), .B(n7671), .Z(n7670) );
  XNOR U7481 ( .A(n7672), .B(n7673), .Z(n7667) );
  AND U7482 ( .A(n668), .B(n7674), .Z(n7673) );
  XOR U7483 ( .A(p_input[1785]), .B(n7672), .Z(n7674) );
  XNOR U7484 ( .A(n7675), .B(n7676), .Z(n7672) );
  AND U7485 ( .A(n672), .B(n7671), .Z(n7676) );
  XNOR U7486 ( .A(n7675), .B(n7669), .Z(n7671) );
  XOR U7487 ( .A(n7677), .B(n7678), .Z(n7669) );
  AND U7488 ( .A(n687), .B(n7679), .Z(n7678) );
  XNOR U7489 ( .A(n7680), .B(n7681), .Z(n7675) );
  AND U7490 ( .A(n679), .B(n7682), .Z(n7681) );
  XOR U7491 ( .A(p_input[1817]), .B(n7680), .Z(n7682) );
  XNOR U7492 ( .A(n7683), .B(n7684), .Z(n7680) );
  AND U7493 ( .A(n683), .B(n7679), .Z(n7684) );
  XNOR U7494 ( .A(n7683), .B(n7677), .Z(n7679) );
  XOR U7495 ( .A(n7685), .B(n7686), .Z(n7677) );
  AND U7496 ( .A(n698), .B(n7687), .Z(n7686) );
  XNOR U7497 ( .A(n7688), .B(n7689), .Z(n7683) );
  AND U7498 ( .A(n690), .B(n7690), .Z(n7689) );
  XOR U7499 ( .A(p_input[1849]), .B(n7688), .Z(n7690) );
  XNOR U7500 ( .A(n7691), .B(n7692), .Z(n7688) );
  AND U7501 ( .A(n694), .B(n7687), .Z(n7692) );
  XNOR U7502 ( .A(n7691), .B(n7685), .Z(n7687) );
  XOR U7503 ( .A(n7693), .B(n7694), .Z(n7685) );
  AND U7504 ( .A(n709), .B(n7695), .Z(n7694) );
  XNOR U7505 ( .A(n7696), .B(n7697), .Z(n7691) );
  AND U7506 ( .A(n701), .B(n7698), .Z(n7697) );
  XOR U7507 ( .A(p_input[1881]), .B(n7696), .Z(n7698) );
  XNOR U7508 ( .A(n7699), .B(n7700), .Z(n7696) );
  AND U7509 ( .A(n705), .B(n7695), .Z(n7700) );
  XNOR U7510 ( .A(n7699), .B(n7693), .Z(n7695) );
  XOR U7511 ( .A(n7701), .B(n7702), .Z(n7693) );
  AND U7512 ( .A(n720), .B(n7703), .Z(n7702) );
  XNOR U7513 ( .A(n7704), .B(n7705), .Z(n7699) );
  AND U7514 ( .A(n712), .B(n7706), .Z(n7705) );
  XOR U7515 ( .A(p_input[1913]), .B(n7704), .Z(n7706) );
  XNOR U7516 ( .A(n7707), .B(n7708), .Z(n7704) );
  AND U7517 ( .A(n716), .B(n7703), .Z(n7708) );
  XNOR U7518 ( .A(n7707), .B(n7701), .Z(n7703) );
  XOR U7519 ( .A(n7709), .B(n7710), .Z(n7701) );
  AND U7520 ( .A(n731), .B(n7711), .Z(n7710) );
  XNOR U7521 ( .A(n7712), .B(n7713), .Z(n7707) );
  AND U7522 ( .A(n723), .B(n7714), .Z(n7713) );
  XOR U7523 ( .A(p_input[1945]), .B(n7712), .Z(n7714) );
  XNOR U7524 ( .A(n7715), .B(n7716), .Z(n7712) );
  AND U7525 ( .A(n727), .B(n7711), .Z(n7716) );
  XNOR U7526 ( .A(n7715), .B(n7709), .Z(n7711) );
  XOR U7527 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n7717), .Z(n7709) );
  AND U7528 ( .A(n741), .B(n7718), .Z(n7717) );
  XNOR U7529 ( .A(n7719), .B(n7720), .Z(n7715) );
  AND U7530 ( .A(n734), .B(n7721), .Z(n7720) );
  XOR U7531 ( .A(p_input[1977]), .B(n7719), .Z(n7721) );
  XNOR U7532 ( .A(n7722), .B(n7723), .Z(n7719) );
  AND U7533 ( .A(n738), .B(n7718), .Z(n7723) );
  XOR U7534 ( .A(\knn_comb_/min_val_out[0][25] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .Z(n7718) );
  XOR U7535 ( .A(n25), .B(n7724), .Z(o[24]) );
  AND U7536 ( .A(n58), .B(n7725), .Z(n25) );
  XOR U7537 ( .A(n26), .B(n7724), .Z(n7725) );
  XOR U7538 ( .A(n7726), .B(n7727), .Z(n7724) );
  AND U7539 ( .A(n70), .B(n7728), .Z(n7727) );
  XOR U7540 ( .A(n7729), .B(n7730), .Z(n26) );
  AND U7541 ( .A(n62), .B(n7731), .Z(n7730) );
  XOR U7542 ( .A(p_input[24]), .B(n7729), .Z(n7731) );
  XNOR U7543 ( .A(n7732), .B(n7733), .Z(n7729) );
  AND U7544 ( .A(n66), .B(n7728), .Z(n7733) );
  XNOR U7545 ( .A(n7732), .B(n7726), .Z(n7728) );
  XOR U7546 ( .A(n7734), .B(n7735), .Z(n7726) );
  AND U7547 ( .A(n82), .B(n7736), .Z(n7735) );
  XNOR U7548 ( .A(n7737), .B(n7738), .Z(n7732) );
  AND U7549 ( .A(n74), .B(n7739), .Z(n7738) );
  XOR U7550 ( .A(p_input[56]), .B(n7737), .Z(n7739) );
  XNOR U7551 ( .A(n7740), .B(n7741), .Z(n7737) );
  AND U7552 ( .A(n78), .B(n7736), .Z(n7741) );
  XNOR U7553 ( .A(n7740), .B(n7734), .Z(n7736) );
  XOR U7554 ( .A(n7742), .B(n7743), .Z(n7734) );
  AND U7555 ( .A(n93), .B(n7744), .Z(n7743) );
  XNOR U7556 ( .A(n7745), .B(n7746), .Z(n7740) );
  AND U7557 ( .A(n85), .B(n7747), .Z(n7746) );
  XOR U7558 ( .A(p_input[88]), .B(n7745), .Z(n7747) );
  XNOR U7559 ( .A(n7748), .B(n7749), .Z(n7745) );
  AND U7560 ( .A(n89), .B(n7744), .Z(n7749) );
  XNOR U7561 ( .A(n7748), .B(n7742), .Z(n7744) );
  XOR U7562 ( .A(n7750), .B(n7751), .Z(n7742) );
  AND U7563 ( .A(n104), .B(n7752), .Z(n7751) );
  XNOR U7564 ( .A(n7753), .B(n7754), .Z(n7748) );
  AND U7565 ( .A(n96), .B(n7755), .Z(n7754) );
  XOR U7566 ( .A(p_input[120]), .B(n7753), .Z(n7755) );
  XNOR U7567 ( .A(n7756), .B(n7757), .Z(n7753) );
  AND U7568 ( .A(n100), .B(n7752), .Z(n7757) );
  XNOR U7569 ( .A(n7756), .B(n7750), .Z(n7752) );
  XOR U7570 ( .A(n7758), .B(n7759), .Z(n7750) );
  AND U7571 ( .A(n115), .B(n7760), .Z(n7759) );
  XNOR U7572 ( .A(n7761), .B(n7762), .Z(n7756) );
  AND U7573 ( .A(n107), .B(n7763), .Z(n7762) );
  XOR U7574 ( .A(p_input[152]), .B(n7761), .Z(n7763) );
  XNOR U7575 ( .A(n7764), .B(n7765), .Z(n7761) );
  AND U7576 ( .A(n111), .B(n7760), .Z(n7765) );
  XNOR U7577 ( .A(n7764), .B(n7758), .Z(n7760) );
  XOR U7578 ( .A(n7766), .B(n7767), .Z(n7758) );
  AND U7579 ( .A(n126), .B(n7768), .Z(n7767) );
  XNOR U7580 ( .A(n7769), .B(n7770), .Z(n7764) );
  AND U7581 ( .A(n118), .B(n7771), .Z(n7770) );
  XOR U7582 ( .A(p_input[184]), .B(n7769), .Z(n7771) );
  XNOR U7583 ( .A(n7772), .B(n7773), .Z(n7769) );
  AND U7584 ( .A(n122), .B(n7768), .Z(n7773) );
  XNOR U7585 ( .A(n7772), .B(n7766), .Z(n7768) );
  XOR U7586 ( .A(n7774), .B(n7775), .Z(n7766) );
  AND U7587 ( .A(n137), .B(n7776), .Z(n7775) );
  XNOR U7588 ( .A(n7777), .B(n7778), .Z(n7772) );
  AND U7589 ( .A(n129), .B(n7779), .Z(n7778) );
  XOR U7590 ( .A(p_input[216]), .B(n7777), .Z(n7779) );
  XNOR U7591 ( .A(n7780), .B(n7781), .Z(n7777) );
  AND U7592 ( .A(n133), .B(n7776), .Z(n7781) );
  XNOR U7593 ( .A(n7780), .B(n7774), .Z(n7776) );
  XOR U7594 ( .A(n7782), .B(n7783), .Z(n7774) );
  AND U7595 ( .A(n148), .B(n7784), .Z(n7783) );
  XNOR U7596 ( .A(n7785), .B(n7786), .Z(n7780) );
  AND U7597 ( .A(n140), .B(n7787), .Z(n7786) );
  XOR U7598 ( .A(p_input[248]), .B(n7785), .Z(n7787) );
  XNOR U7599 ( .A(n7788), .B(n7789), .Z(n7785) );
  AND U7600 ( .A(n144), .B(n7784), .Z(n7789) );
  XNOR U7601 ( .A(n7788), .B(n7782), .Z(n7784) );
  XOR U7602 ( .A(n7790), .B(n7791), .Z(n7782) );
  AND U7603 ( .A(n159), .B(n7792), .Z(n7791) );
  XNOR U7604 ( .A(n7793), .B(n7794), .Z(n7788) );
  AND U7605 ( .A(n151), .B(n7795), .Z(n7794) );
  XOR U7606 ( .A(p_input[280]), .B(n7793), .Z(n7795) );
  XNOR U7607 ( .A(n7796), .B(n7797), .Z(n7793) );
  AND U7608 ( .A(n155), .B(n7792), .Z(n7797) );
  XNOR U7609 ( .A(n7796), .B(n7790), .Z(n7792) );
  XOR U7610 ( .A(n7798), .B(n7799), .Z(n7790) );
  AND U7611 ( .A(n170), .B(n7800), .Z(n7799) );
  XNOR U7612 ( .A(n7801), .B(n7802), .Z(n7796) );
  AND U7613 ( .A(n162), .B(n7803), .Z(n7802) );
  XOR U7614 ( .A(p_input[312]), .B(n7801), .Z(n7803) );
  XNOR U7615 ( .A(n7804), .B(n7805), .Z(n7801) );
  AND U7616 ( .A(n166), .B(n7800), .Z(n7805) );
  XNOR U7617 ( .A(n7804), .B(n7798), .Z(n7800) );
  XOR U7618 ( .A(n7806), .B(n7807), .Z(n7798) );
  AND U7619 ( .A(n181), .B(n7808), .Z(n7807) );
  XNOR U7620 ( .A(n7809), .B(n7810), .Z(n7804) );
  AND U7621 ( .A(n173), .B(n7811), .Z(n7810) );
  XOR U7622 ( .A(p_input[344]), .B(n7809), .Z(n7811) );
  XNOR U7623 ( .A(n7812), .B(n7813), .Z(n7809) );
  AND U7624 ( .A(n177), .B(n7808), .Z(n7813) );
  XNOR U7625 ( .A(n7812), .B(n7806), .Z(n7808) );
  XOR U7626 ( .A(n7814), .B(n7815), .Z(n7806) );
  AND U7627 ( .A(n192), .B(n7816), .Z(n7815) );
  XNOR U7628 ( .A(n7817), .B(n7818), .Z(n7812) );
  AND U7629 ( .A(n184), .B(n7819), .Z(n7818) );
  XOR U7630 ( .A(p_input[376]), .B(n7817), .Z(n7819) );
  XNOR U7631 ( .A(n7820), .B(n7821), .Z(n7817) );
  AND U7632 ( .A(n188), .B(n7816), .Z(n7821) );
  XNOR U7633 ( .A(n7820), .B(n7814), .Z(n7816) );
  XOR U7634 ( .A(n7822), .B(n7823), .Z(n7814) );
  AND U7635 ( .A(n203), .B(n7824), .Z(n7823) );
  XNOR U7636 ( .A(n7825), .B(n7826), .Z(n7820) );
  AND U7637 ( .A(n195), .B(n7827), .Z(n7826) );
  XOR U7638 ( .A(p_input[408]), .B(n7825), .Z(n7827) );
  XNOR U7639 ( .A(n7828), .B(n7829), .Z(n7825) );
  AND U7640 ( .A(n199), .B(n7824), .Z(n7829) );
  XNOR U7641 ( .A(n7828), .B(n7822), .Z(n7824) );
  XOR U7642 ( .A(n7830), .B(n7831), .Z(n7822) );
  AND U7643 ( .A(n214), .B(n7832), .Z(n7831) );
  XNOR U7644 ( .A(n7833), .B(n7834), .Z(n7828) );
  AND U7645 ( .A(n206), .B(n7835), .Z(n7834) );
  XOR U7646 ( .A(p_input[440]), .B(n7833), .Z(n7835) );
  XNOR U7647 ( .A(n7836), .B(n7837), .Z(n7833) );
  AND U7648 ( .A(n210), .B(n7832), .Z(n7837) );
  XNOR U7649 ( .A(n7836), .B(n7830), .Z(n7832) );
  XOR U7650 ( .A(n7838), .B(n7839), .Z(n7830) );
  AND U7651 ( .A(n225), .B(n7840), .Z(n7839) );
  XNOR U7652 ( .A(n7841), .B(n7842), .Z(n7836) );
  AND U7653 ( .A(n217), .B(n7843), .Z(n7842) );
  XOR U7654 ( .A(p_input[472]), .B(n7841), .Z(n7843) );
  XNOR U7655 ( .A(n7844), .B(n7845), .Z(n7841) );
  AND U7656 ( .A(n221), .B(n7840), .Z(n7845) );
  XNOR U7657 ( .A(n7844), .B(n7838), .Z(n7840) );
  XOR U7658 ( .A(n7846), .B(n7847), .Z(n7838) );
  AND U7659 ( .A(n236), .B(n7848), .Z(n7847) );
  XNOR U7660 ( .A(n7849), .B(n7850), .Z(n7844) );
  AND U7661 ( .A(n228), .B(n7851), .Z(n7850) );
  XOR U7662 ( .A(p_input[504]), .B(n7849), .Z(n7851) );
  XNOR U7663 ( .A(n7852), .B(n7853), .Z(n7849) );
  AND U7664 ( .A(n232), .B(n7848), .Z(n7853) );
  XNOR U7665 ( .A(n7852), .B(n7846), .Z(n7848) );
  XOR U7666 ( .A(n7854), .B(n7855), .Z(n7846) );
  AND U7667 ( .A(n247), .B(n7856), .Z(n7855) );
  XNOR U7668 ( .A(n7857), .B(n7858), .Z(n7852) );
  AND U7669 ( .A(n239), .B(n7859), .Z(n7858) );
  XOR U7670 ( .A(p_input[536]), .B(n7857), .Z(n7859) );
  XNOR U7671 ( .A(n7860), .B(n7861), .Z(n7857) );
  AND U7672 ( .A(n243), .B(n7856), .Z(n7861) );
  XNOR U7673 ( .A(n7860), .B(n7854), .Z(n7856) );
  XOR U7674 ( .A(n7862), .B(n7863), .Z(n7854) );
  AND U7675 ( .A(n258), .B(n7864), .Z(n7863) );
  XNOR U7676 ( .A(n7865), .B(n7866), .Z(n7860) );
  AND U7677 ( .A(n250), .B(n7867), .Z(n7866) );
  XOR U7678 ( .A(p_input[568]), .B(n7865), .Z(n7867) );
  XNOR U7679 ( .A(n7868), .B(n7869), .Z(n7865) );
  AND U7680 ( .A(n254), .B(n7864), .Z(n7869) );
  XNOR U7681 ( .A(n7868), .B(n7862), .Z(n7864) );
  XOR U7682 ( .A(n7870), .B(n7871), .Z(n7862) );
  AND U7683 ( .A(n269), .B(n7872), .Z(n7871) );
  XNOR U7684 ( .A(n7873), .B(n7874), .Z(n7868) );
  AND U7685 ( .A(n261), .B(n7875), .Z(n7874) );
  XOR U7686 ( .A(p_input[600]), .B(n7873), .Z(n7875) );
  XNOR U7687 ( .A(n7876), .B(n7877), .Z(n7873) );
  AND U7688 ( .A(n265), .B(n7872), .Z(n7877) );
  XNOR U7689 ( .A(n7876), .B(n7870), .Z(n7872) );
  XOR U7690 ( .A(n7878), .B(n7879), .Z(n7870) );
  AND U7691 ( .A(n280), .B(n7880), .Z(n7879) );
  XNOR U7692 ( .A(n7881), .B(n7882), .Z(n7876) );
  AND U7693 ( .A(n272), .B(n7883), .Z(n7882) );
  XOR U7694 ( .A(p_input[632]), .B(n7881), .Z(n7883) );
  XNOR U7695 ( .A(n7884), .B(n7885), .Z(n7881) );
  AND U7696 ( .A(n276), .B(n7880), .Z(n7885) );
  XNOR U7697 ( .A(n7884), .B(n7878), .Z(n7880) );
  XOR U7698 ( .A(n7886), .B(n7887), .Z(n7878) );
  AND U7699 ( .A(n291), .B(n7888), .Z(n7887) );
  XNOR U7700 ( .A(n7889), .B(n7890), .Z(n7884) );
  AND U7701 ( .A(n283), .B(n7891), .Z(n7890) );
  XOR U7702 ( .A(p_input[664]), .B(n7889), .Z(n7891) );
  XNOR U7703 ( .A(n7892), .B(n7893), .Z(n7889) );
  AND U7704 ( .A(n287), .B(n7888), .Z(n7893) );
  XNOR U7705 ( .A(n7892), .B(n7886), .Z(n7888) );
  XOR U7706 ( .A(n7894), .B(n7895), .Z(n7886) );
  AND U7707 ( .A(n302), .B(n7896), .Z(n7895) );
  XNOR U7708 ( .A(n7897), .B(n7898), .Z(n7892) );
  AND U7709 ( .A(n294), .B(n7899), .Z(n7898) );
  XOR U7710 ( .A(p_input[696]), .B(n7897), .Z(n7899) );
  XNOR U7711 ( .A(n7900), .B(n7901), .Z(n7897) );
  AND U7712 ( .A(n298), .B(n7896), .Z(n7901) );
  XNOR U7713 ( .A(n7900), .B(n7894), .Z(n7896) );
  XOR U7714 ( .A(n7902), .B(n7903), .Z(n7894) );
  AND U7715 ( .A(n313), .B(n7904), .Z(n7903) );
  XNOR U7716 ( .A(n7905), .B(n7906), .Z(n7900) );
  AND U7717 ( .A(n305), .B(n7907), .Z(n7906) );
  XOR U7718 ( .A(p_input[728]), .B(n7905), .Z(n7907) );
  XNOR U7719 ( .A(n7908), .B(n7909), .Z(n7905) );
  AND U7720 ( .A(n309), .B(n7904), .Z(n7909) );
  XNOR U7721 ( .A(n7908), .B(n7902), .Z(n7904) );
  XOR U7722 ( .A(n7910), .B(n7911), .Z(n7902) );
  AND U7723 ( .A(n324), .B(n7912), .Z(n7911) );
  XNOR U7724 ( .A(n7913), .B(n7914), .Z(n7908) );
  AND U7725 ( .A(n316), .B(n7915), .Z(n7914) );
  XOR U7726 ( .A(p_input[760]), .B(n7913), .Z(n7915) );
  XNOR U7727 ( .A(n7916), .B(n7917), .Z(n7913) );
  AND U7728 ( .A(n320), .B(n7912), .Z(n7917) );
  XNOR U7729 ( .A(n7916), .B(n7910), .Z(n7912) );
  XOR U7730 ( .A(n7918), .B(n7919), .Z(n7910) );
  AND U7731 ( .A(n335), .B(n7920), .Z(n7919) );
  XNOR U7732 ( .A(n7921), .B(n7922), .Z(n7916) );
  AND U7733 ( .A(n327), .B(n7923), .Z(n7922) );
  XOR U7734 ( .A(p_input[792]), .B(n7921), .Z(n7923) );
  XNOR U7735 ( .A(n7924), .B(n7925), .Z(n7921) );
  AND U7736 ( .A(n331), .B(n7920), .Z(n7925) );
  XNOR U7737 ( .A(n7924), .B(n7918), .Z(n7920) );
  XOR U7738 ( .A(n7926), .B(n7927), .Z(n7918) );
  AND U7739 ( .A(n346), .B(n7928), .Z(n7927) );
  XNOR U7740 ( .A(n7929), .B(n7930), .Z(n7924) );
  AND U7741 ( .A(n338), .B(n7931), .Z(n7930) );
  XOR U7742 ( .A(p_input[824]), .B(n7929), .Z(n7931) );
  XNOR U7743 ( .A(n7932), .B(n7933), .Z(n7929) );
  AND U7744 ( .A(n342), .B(n7928), .Z(n7933) );
  XNOR U7745 ( .A(n7932), .B(n7926), .Z(n7928) );
  XOR U7746 ( .A(n7934), .B(n7935), .Z(n7926) );
  AND U7747 ( .A(n357), .B(n7936), .Z(n7935) );
  XNOR U7748 ( .A(n7937), .B(n7938), .Z(n7932) );
  AND U7749 ( .A(n349), .B(n7939), .Z(n7938) );
  XOR U7750 ( .A(p_input[856]), .B(n7937), .Z(n7939) );
  XNOR U7751 ( .A(n7940), .B(n7941), .Z(n7937) );
  AND U7752 ( .A(n353), .B(n7936), .Z(n7941) );
  XNOR U7753 ( .A(n7940), .B(n7934), .Z(n7936) );
  XOR U7754 ( .A(n7942), .B(n7943), .Z(n7934) );
  AND U7755 ( .A(n368), .B(n7944), .Z(n7943) );
  XNOR U7756 ( .A(n7945), .B(n7946), .Z(n7940) );
  AND U7757 ( .A(n360), .B(n7947), .Z(n7946) );
  XOR U7758 ( .A(p_input[888]), .B(n7945), .Z(n7947) );
  XNOR U7759 ( .A(n7948), .B(n7949), .Z(n7945) );
  AND U7760 ( .A(n364), .B(n7944), .Z(n7949) );
  XNOR U7761 ( .A(n7948), .B(n7942), .Z(n7944) );
  XOR U7762 ( .A(n7950), .B(n7951), .Z(n7942) );
  AND U7763 ( .A(n379), .B(n7952), .Z(n7951) );
  XNOR U7764 ( .A(n7953), .B(n7954), .Z(n7948) );
  AND U7765 ( .A(n371), .B(n7955), .Z(n7954) );
  XOR U7766 ( .A(p_input[920]), .B(n7953), .Z(n7955) );
  XNOR U7767 ( .A(n7956), .B(n7957), .Z(n7953) );
  AND U7768 ( .A(n375), .B(n7952), .Z(n7957) );
  XNOR U7769 ( .A(n7956), .B(n7950), .Z(n7952) );
  XOR U7770 ( .A(n7958), .B(n7959), .Z(n7950) );
  AND U7771 ( .A(n390), .B(n7960), .Z(n7959) );
  XNOR U7772 ( .A(n7961), .B(n7962), .Z(n7956) );
  AND U7773 ( .A(n382), .B(n7963), .Z(n7962) );
  XOR U7774 ( .A(p_input[952]), .B(n7961), .Z(n7963) );
  XNOR U7775 ( .A(n7964), .B(n7965), .Z(n7961) );
  AND U7776 ( .A(n386), .B(n7960), .Z(n7965) );
  XNOR U7777 ( .A(n7964), .B(n7958), .Z(n7960) );
  XOR U7778 ( .A(n7966), .B(n7967), .Z(n7958) );
  AND U7779 ( .A(n401), .B(n7968), .Z(n7967) );
  XNOR U7780 ( .A(n7969), .B(n7970), .Z(n7964) );
  AND U7781 ( .A(n393), .B(n7971), .Z(n7970) );
  XOR U7782 ( .A(p_input[984]), .B(n7969), .Z(n7971) );
  XNOR U7783 ( .A(n7972), .B(n7973), .Z(n7969) );
  AND U7784 ( .A(n397), .B(n7968), .Z(n7973) );
  XNOR U7785 ( .A(n7972), .B(n7966), .Z(n7968) );
  XOR U7786 ( .A(n7974), .B(n7975), .Z(n7966) );
  AND U7787 ( .A(n412), .B(n7976), .Z(n7975) );
  XNOR U7788 ( .A(n7977), .B(n7978), .Z(n7972) );
  AND U7789 ( .A(n404), .B(n7979), .Z(n7978) );
  XOR U7790 ( .A(p_input[1016]), .B(n7977), .Z(n7979) );
  XNOR U7791 ( .A(n7980), .B(n7981), .Z(n7977) );
  AND U7792 ( .A(n408), .B(n7976), .Z(n7981) );
  XNOR U7793 ( .A(n7980), .B(n7974), .Z(n7976) );
  XOR U7794 ( .A(n7982), .B(n7983), .Z(n7974) );
  AND U7795 ( .A(n423), .B(n7984), .Z(n7983) );
  XNOR U7796 ( .A(n7985), .B(n7986), .Z(n7980) );
  AND U7797 ( .A(n415), .B(n7987), .Z(n7986) );
  XOR U7798 ( .A(p_input[1048]), .B(n7985), .Z(n7987) );
  XNOR U7799 ( .A(n7988), .B(n7989), .Z(n7985) );
  AND U7800 ( .A(n419), .B(n7984), .Z(n7989) );
  XNOR U7801 ( .A(n7988), .B(n7982), .Z(n7984) );
  XOR U7802 ( .A(n7990), .B(n7991), .Z(n7982) );
  AND U7803 ( .A(n434), .B(n7992), .Z(n7991) );
  XNOR U7804 ( .A(n7993), .B(n7994), .Z(n7988) );
  AND U7805 ( .A(n426), .B(n7995), .Z(n7994) );
  XOR U7806 ( .A(p_input[1080]), .B(n7993), .Z(n7995) );
  XNOR U7807 ( .A(n7996), .B(n7997), .Z(n7993) );
  AND U7808 ( .A(n430), .B(n7992), .Z(n7997) );
  XNOR U7809 ( .A(n7996), .B(n7990), .Z(n7992) );
  XOR U7810 ( .A(n7998), .B(n7999), .Z(n7990) );
  AND U7811 ( .A(n445), .B(n8000), .Z(n7999) );
  XNOR U7812 ( .A(n8001), .B(n8002), .Z(n7996) );
  AND U7813 ( .A(n437), .B(n8003), .Z(n8002) );
  XOR U7814 ( .A(p_input[1112]), .B(n8001), .Z(n8003) );
  XNOR U7815 ( .A(n8004), .B(n8005), .Z(n8001) );
  AND U7816 ( .A(n441), .B(n8000), .Z(n8005) );
  XNOR U7817 ( .A(n8004), .B(n7998), .Z(n8000) );
  XOR U7818 ( .A(n8006), .B(n8007), .Z(n7998) );
  AND U7819 ( .A(n456), .B(n8008), .Z(n8007) );
  XNOR U7820 ( .A(n8009), .B(n8010), .Z(n8004) );
  AND U7821 ( .A(n448), .B(n8011), .Z(n8010) );
  XOR U7822 ( .A(p_input[1144]), .B(n8009), .Z(n8011) );
  XNOR U7823 ( .A(n8012), .B(n8013), .Z(n8009) );
  AND U7824 ( .A(n452), .B(n8008), .Z(n8013) );
  XNOR U7825 ( .A(n8012), .B(n8006), .Z(n8008) );
  XOR U7826 ( .A(n8014), .B(n8015), .Z(n8006) );
  AND U7827 ( .A(n467), .B(n8016), .Z(n8015) );
  XNOR U7828 ( .A(n8017), .B(n8018), .Z(n8012) );
  AND U7829 ( .A(n459), .B(n8019), .Z(n8018) );
  XOR U7830 ( .A(p_input[1176]), .B(n8017), .Z(n8019) );
  XNOR U7831 ( .A(n8020), .B(n8021), .Z(n8017) );
  AND U7832 ( .A(n463), .B(n8016), .Z(n8021) );
  XNOR U7833 ( .A(n8020), .B(n8014), .Z(n8016) );
  XOR U7834 ( .A(n8022), .B(n8023), .Z(n8014) );
  AND U7835 ( .A(n478), .B(n8024), .Z(n8023) );
  XNOR U7836 ( .A(n8025), .B(n8026), .Z(n8020) );
  AND U7837 ( .A(n470), .B(n8027), .Z(n8026) );
  XOR U7838 ( .A(p_input[1208]), .B(n8025), .Z(n8027) );
  XNOR U7839 ( .A(n8028), .B(n8029), .Z(n8025) );
  AND U7840 ( .A(n474), .B(n8024), .Z(n8029) );
  XNOR U7841 ( .A(n8028), .B(n8022), .Z(n8024) );
  XOR U7842 ( .A(n8030), .B(n8031), .Z(n8022) );
  AND U7843 ( .A(n489), .B(n8032), .Z(n8031) );
  XNOR U7844 ( .A(n8033), .B(n8034), .Z(n8028) );
  AND U7845 ( .A(n481), .B(n8035), .Z(n8034) );
  XOR U7846 ( .A(p_input[1240]), .B(n8033), .Z(n8035) );
  XNOR U7847 ( .A(n8036), .B(n8037), .Z(n8033) );
  AND U7848 ( .A(n485), .B(n8032), .Z(n8037) );
  XNOR U7849 ( .A(n8036), .B(n8030), .Z(n8032) );
  XOR U7850 ( .A(n8038), .B(n8039), .Z(n8030) );
  AND U7851 ( .A(n500), .B(n8040), .Z(n8039) );
  XNOR U7852 ( .A(n8041), .B(n8042), .Z(n8036) );
  AND U7853 ( .A(n492), .B(n8043), .Z(n8042) );
  XOR U7854 ( .A(p_input[1272]), .B(n8041), .Z(n8043) );
  XNOR U7855 ( .A(n8044), .B(n8045), .Z(n8041) );
  AND U7856 ( .A(n496), .B(n8040), .Z(n8045) );
  XNOR U7857 ( .A(n8044), .B(n8038), .Z(n8040) );
  XOR U7858 ( .A(n8046), .B(n8047), .Z(n8038) );
  AND U7859 ( .A(n511), .B(n8048), .Z(n8047) );
  XNOR U7860 ( .A(n8049), .B(n8050), .Z(n8044) );
  AND U7861 ( .A(n503), .B(n8051), .Z(n8050) );
  XOR U7862 ( .A(p_input[1304]), .B(n8049), .Z(n8051) );
  XNOR U7863 ( .A(n8052), .B(n8053), .Z(n8049) );
  AND U7864 ( .A(n507), .B(n8048), .Z(n8053) );
  XNOR U7865 ( .A(n8052), .B(n8046), .Z(n8048) );
  XOR U7866 ( .A(n8054), .B(n8055), .Z(n8046) );
  AND U7867 ( .A(n522), .B(n8056), .Z(n8055) );
  XNOR U7868 ( .A(n8057), .B(n8058), .Z(n8052) );
  AND U7869 ( .A(n514), .B(n8059), .Z(n8058) );
  XOR U7870 ( .A(p_input[1336]), .B(n8057), .Z(n8059) );
  XNOR U7871 ( .A(n8060), .B(n8061), .Z(n8057) );
  AND U7872 ( .A(n518), .B(n8056), .Z(n8061) );
  XNOR U7873 ( .A(n8060), .B(n8054), .Z(n8056) );
  XOR U7874 ( .A(n8062), .B(n8063), .Z(n8054) );
  AND U7875 ( .A(n533), .B(n8064), .Z(n8063) );
  XNOR U7876 ( .A(n8065), .B(n8066), .Z(n8060) );
  AND U7877 ( .A(n525), .B(n8067), .Z(n8066) );
  XOR U7878 ( .A(p_input[1368]), .B(n8065), .Z(n8067) );
  XNOR U7879 ( .A(n8068), .B(n8069), .Z(n8065) );
  AND U7880 ( .A(n529), .B(n8064), .Z(n8069) );
  XNOR U7881 ( .A(n8068), .B(n8062), .Z(n8064) );
  XOR U7882 ( .A(n8070), .B(n8071), .Z(n8062) );
  AND U7883 ( .A(n544), .B(n8072), .Z(n8071) );
  XNOR U7884 ( .A(n8073), .B(n8074), .Z(n8068) );
  AND U7885 ( .A(n536), .B(n8075), .Z(n8074) );
  XOR U7886 ( .A(p_input[1400]), .B(n8073), .Z(n8075) );
  XNOR U7887 ( .A(n8076), .B(n8077), .Z(n8073) );
  AND U7888 ( .A(n540), .B(n8072), .Z(n8077) );
  XNOR U7889 ( .A(n8076), .B(n8070), .Z(n8072) );
  XOR U7890 ( .A(n8078), .B(n8079), .Z(n8070) );
  AND U7891 ( .A(n555), .B(n8080), .Z(n8079) );
  XNOR U7892 ( .A(n8081), .B(n8082), .Z(n8076) );
  AND U7893 ( .A(n547), .B(n8083), .Z(n8082) );
  XOR U7894 ( .A(p_input[1432]), .B(n8081), .Z(n8083) );
  XNOR U7895 ( .A(n8084), .B(n8085), .Z(n8081) );
  AND U7896 ( .A(n551), .B(n8080), .Z(n8085) );
  XNOR U7897 ( .A(n8084), .B(n8078), .Z(n8080) );
  XOR U7898 ( .A(n8086), .B(n8087), .Z(n8078) );
  AND U7899 ( .A(n566), .B(n8088), .Z(n8087) );
  XNOR U7900 ( .A(n8089), .B(n8090), .Z(n8084) );
  AND U7901 ( .A(n558), .B(n8091), .Z(n8090) );
  XOR U7902 ( .A(p_input[1464]), .B(n8089), .Z(n8091) );
  XNOR U7903 ( .A(n8092), .B(n8093), .Z(n8089) );
  AND U7904 ( .A(n562), .B(n8088), .Z(n8093) );
  XNOR U7905 ( .A(n8092), .B(n8086), .Z(n8088) );
  XOR U7906 ( .A(n8094), .B(n8095), .Z(n8086) );
  AND U7907 ( .A(n577), .B(n8096), .Z(n8095) );
  XNOR U7908 ( .A(n8097), .B(n8098), .Z(n8092) );
  AND U7909 ( .A(n569), .B(n8099), .Z(n8098) );
  XOR U7910 ( .A(p_input[1496]), .B(n8097), .Z(n8099) );
  XNOR U7911 ( .A(n8100), .B(n8101), .Z(n8097) );
  AND U7912 ( .A(n573), .B(n8096), .Z(n8101) );
  XNOR U7913 ( .A(n8100), .B(n8094), .Z(n8096) );
  XOR U7914 ( .A(n8102), .B(n8103), .Z(n8094) );
  AND U7915 ( .A(n588), .B(n8104), .Z(n8103) );
  XNOR U7916 ( .A(n8105), .B(n8106), .Z(n8100) );
  AND U7917 ( .A(n580), .B(n8107), .Z(n8106) );
  XOR U7918 ( .A(p_input[1528]), .B(n8105), .Z(n8107) );
  XNOR U7919 ( .A(n8108), .B(n8109), .Z(n8105) );
  AND U7920 ( .A(n584), .B(n8104), .Z(n8109) );
  XNOR U7921 ( .A(n8108), .B(n8102), .Z(n8104) );
  XOR U7922 ( .A(n8110), .B(n8111), .Z(n8102) );
  AND U7923 ( .A(n599), .B(n8112), .Z(n8111) );
  XNOR U7924 ( .A(n8113), .B(n8114), .Z(n8108) );
  AND U7925 ( .A(n591), .B(n8115), .Z(n8114) );
  XOR U7926 ( .A(p_input[1560]), .B(n8113), .Z(n8115) );
  XNOR U7927 ( .A(n8116), .B(n8117), .Z(n8113) );
  AND U7928 ( .A(n595), .B(n8112), .Z(n8117) );
  XNOR U7929 ( .A(n8116), .B(n8110), .Z(n8112) );
  XOR U7930 ( .A(n8118), .B(n8119), .Z(n8110) );
  AND U7931 ( .A(n610), .B(n8120), .Z(n8119) );
  XNOR U7932 ( .A(n8121), .B(n8122), .Z(n8116) );
  AND U7933 ( .A(n602), .B(n8123), .Z(n8122) );
  XOR U7934 ( .A(p_input[1592]), .B(n8121), .Z(n8123) );
  XNOR U7935 ( .A(n8124), .B(n8125), .Z(n8121) );
  AND U7936 ( .A(n606), .B(n8120), .Z(n8125) );
  XNOR U7937 ( .A(n8124), .B(n8118), .Z(n8120) );
  XOR U7938 ( .A(n8126), .B(n8127), .Z(n8118) );
  AND U7939 ( .A(n621), .B(n8128), .Z(n8127) );
  XNOR U7940 ( .A(n8129), .B(n8130), .Z(n8124) );
  AND U7941 ( .A(n613), .B(n8131), .Z(n8130) );
  XOR U7942 ( .A(p_input[1624]), .B(n8129), .Z(n8131) );
  XNOR U7943 ( .A(n8132), .B(n8133), .Z(n8129) );
  AND U7944 ( .A(n617), .B(n8128), .Z(n8133) );
  XNOR U7945 ( .A(n8132), .B(n8126), .Z(n8128) );
  XOR U7946 ( .A(n8134), .B(n8135), .Z(n8126) );
  AND U7947 ( .A(n632), .B(n8136), .Z(n8135) );
  XNOR U7948 ( .A(n8137), .B(n8138), .Z(n8132) );
  AND U7949 ( .A(n624), .B(n8139), .Z(n8138) );
  XOR U7950 ( .A(p_input[1656]), .B(n8137), .Z(n8139) );
  XNOR U7951 ( .A(n8140), .B(n8141), .Z(n8137) );
  AND U7952 ( .A(n628), .B(n8136), .Z(n8141) );
  XNOR U7953 ( .A(n8140), .B(n8134), .Z(n8136) );
  XOR U7954 ( .A(n8142), .B(n8143), .Z(n8134) );
  AND U7955 ( .A(n643), .B(n8144), .Z(n8143) );
  XNOR U7956 ( .A(n8145), .B(n8146), .Z(n8140) );
  AND U7957 ( .A(n635), .B(n8147), .Z(n8146) );
  XOR U7958 ( .A(p_input[1688]), .B(n8145), .Z(n8147) );
  XNOR U7959 ( .A(n8148), .B(n8149), .Z(n8145) );
  AND U7960 ( .A(n639), .B(n8144), .Z(n8149) );
  XNOR U7961 ( .A(n8148), .B(n8142), .Z(n8144) );
  XOR U7962 ( .A(n8150), .B(n8151), .Z(n8142) );
  AND U7963 ( .A(n654), .B(n8152), .Z(n8151) );
  XNOR U7964 ( .A(n8153), .B(n8154), .Z(n8148) );
  AND U7965 ( .A(n646), .B(n8155), .Z(n8154) );
  XOR U7966 ( .A(p_input[1720]), .B(n8153), .Z(n8155) );
  XNOR U7967 ( .A(n8156), .B(n8157), .Z(n8153) );
  AND U7968 ( .A(n650), .B(n8152), .Z(n8157) );
  XNOR U7969 ( .A(n8156), .B(n8150), .Z(n8152) );
  XOR U7970 ( .A(n8158), .B(n8159), .Z(n8150) );
  AND U7971 ( .A(n665), .B(n8160), .Z(n8159) );
  XNOR U7972 ( .A(n8161), .B(n8162), .Z(n8156) );
  AND U7973 ( .A(n657), .B(n8163), .Z(n8162) );
  XOR U7974 ( .A(p_input[1752]), .B(n8161), .Z(n8163) );
  XNOR U7975 ( .A(n8164), .B(n8165), .Z(n8161) );
  AND U7976 ( .A(n661), .B(n8160), .Z(n8165) );
  XNOR U7977 ( .A(n8164), .B(n8158), .Z(n8160) );
  XOR U7978 ( .A(n8166), .B(n8167), .Z(n8158) );
  AND U7979 ( .A(n676), .B(n8168), .Z(n8167) );
  XNOR U7980 ( .A(n8169), .B(n8170), .Z(n8164) );
  AND U7981 ( .A(n668), .B(n8171), .Z(n8170) );
  XOR U7982 ( .A(p_input[1784]), .B(n8169), .Z(n8171) );
  XNOR U7983 ( .A(n8172), .B(n8173), .Z(n8169) );
  AND U7984 ( .A(n672), .B(n8168), .Z(n8173) );
  XNOR U7985 ( .A(n8172), .B(n8166), .Z(n8168) );
  XOR U7986 ( .A(n8174), .B(n8175), .Z(n8166) );
  AND U7987 ( .A(n687), .B(n8176), .Z(n8175) );
  XNOR U7988 ( .A(n8177), .B(n8178), .Z(n8172) );
  AND U7989 ( .A(n679), .B(n8179), .Z(n8178) );
  XOR U7990 ( .A(p_input[1816]), .B(n8177), .Z(n8179) );
  XNOR U7991 ( .A(n8180), .B(n8181), .Z(n8177) );
  AND U7992 ( .A(n683), .B(n8176), .Z(n8181) );
  XNOR U7993 ( .A(n8180), .B(n8174), .Z(n8176) );
  XOR U7994 ( .A(n8182), .B(n8183), .Z(n8174) );
  AND U7995 ( .A(n698), .B(n8184), .Z(n8183) );
  XNOR U7996 ( .A(n8185), .B(n8186), .Z(n8180) );
  AND U7997 ( .A(n690), .B(n8187), .Z(n8186) );
  XOR U7998 ( .A(p_input[1848]), .B(n8185), .Z(n8187) );
  XNOR U7999 ( .A(n8188), .B(n8189), .Z(n8185) );
  AND U8000 ( .A(n694), .B(n8184), .Z(n8189) );
  XNOR U8001 ( .A(n8188), .B(n8182), .Z(n8184) );
  XOR U8002 ( .A(n8190), .B(n8191), .Z(n8182) );
  AND U8003 ( .A(n709), .B(n8192), .Z(n8191) );
  XNOR U8004 ( .A(n8193), .B(n8194), .Z(n8188) );
  AND U8005 ( .A(n701), .B(n8195), .Z(n8194) );
  XOR U8006 ( .A(p_input[1880]), .B(n8193), .Z(n8195) );
  XNOR U8007 ( .A(n8196), .B(n8197), .Z(n8193) );
  AND U8008 ( .A(n705), .B(n8192), .Z(n8197) );
  XNOR U8009 ( .A(n8196), .B(n8190), .Z(n8192) );
  XOR U8010 ( .A(n8198), .B(n8199), .Z(n8190) );
  AND U8011 ( .A(n720), .B(n8200), .Z(n8199) );
  XNOR U8012 ( .A(n8201), .B(n8202), .Z(n8196) );
  AND U8013 ( .A(n712), .B(n8203), .Z(n8202) );
  XOR U8014 ( .A(p_input[1912]), .B(n8201), .Z(n8203) );
  XNOR U8015 ( .A(n8204), .B(n8205), .Z(n8201) );
  AND U8016 ( .A(n716), .B(n8200), .Z(n8205) );
  XNOR U8017 ( .A(n8204), .B(n8198), .Z(n8200) );
  XOR U8018 ( .A(n8206), .B(n8207), .Z(n8198) );
  AND U8019 ( .A(n731), .B(n8208), .Z(n8207) );
  XNOR U8020 ( .A(n8209), .B(n8210), .Z(n8204) );
  AND U8021 ( .A(n723), .B(n8211), .Z(n8210) );
  XOR U8022 ( .A(p_input[1944]), .B(n8209), .Z(n8211) );
  XNOR U8023 ( .A(n8212), .B(n8213), .Z(n8209) );
  AND U8024 ( .A(n727), .B(n8208), .Z(n8213) );
  XNOR U8025 ( .A(n8212), .B(n8206), .Z(n8208) );
  XOR U8026 ( .A(\knn_comb_/min_val_out[0][24] ), .B(n8214), .Z(n8206) );
  AND U8027 ( .A(n741), .B(n8215), .Z(n8214) );
  XNOR U8028 ( .A(n8216), .B(n8217), .Z(n8212) );
  AND U8029 ( .A(n734), .B(n8218), .Z(n8217) );
  XOR U8030 ( .A(p_input[1976]), .B(n8216), .Z(n8218) );
  XNOR U8031 ( .A(n8219), .B(n8220), .Z(n8216) );
  AND U8032 ( .A(n738), .B(n8215), .Z(n8220) );
  XOR U8033 ( .A(\knn_comb_/min_val_out[0][24] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .Z(n8215) );
  XOR U8034 ( .A(n27), .B(n8221), .Z(o[23]) );
  AND U8035 ( .A(n58), .B(n8222), .Z(n27) );
  XOR U8036 ( .A(n28), .B(n8221), .Z(n8222) );
  XOR U8037 ( .A(n8223), .B(n8224), .Z(n8221) );
  AND U8038 ( .A(n70), .B(n8225), .Z(n8224) );
  XOR U8039 ( .A(n8226), .B(n8227), .Z(n28) );
  AND U8040 ( .A(n62), .B(n8228), .Z(n8227) );
  XOR U8041 ( .A(p_input[23]), .B(n8226), .Z(n8228) );
  XNOR U8042 ( .A(n8229), .B(n8230), .Z(n8226) );
  AND U8043 ( .A(n66), .B(n8225), .Z(n8230) );
  XNOR U8044 ( .A(n8229), .B(n8223), .Z(n8225) );
  XOR U8045 ( .A(n8231), .B(n8232), .Z(n8223) );
  AND U8046 ( .A(n82), .B(n8233), .Z(n8232) );
  XNOR U8047 ( .A(n8234), .B(n8235), .Z(n8229) );
  AND U8048 ( .A(n74), .B(n8236), .Z(n8235) );
  XOR U8049 ( .A(p_input[55]), .B(n8234), .Z(n8236) );
  XNOR U8050 ( .A(n8237), .B(n8238), .Z(n8234) );
  AND U8051 ( .A(n78), .B(n8233), .Z(n8238) );
  XNOR U8052 ( .A(n8237), .B(n8231), .Z(n8233) );
  XOR U8053 ( .A(n8239), .B(n8240), .Z(n8231) );
  AND U8054 ( .A(n93), .B(n8241), .Z(n8240) );
  XNOR U8055 ( .A(n8242), .B(n8243), .Z(n8237) );
  AND U8056 ( .A(n85), .B(n8244), .Z(n8243) );
  XOR U8057 ( .A(p_input[87]), .B(n8242), .Z(n8244) );
  XNOR U8058 ( .A(n8245), .B(n8246), .Z(n8242) );
  AND U8059 ( .A(n89), .B(n8241), .Z(n8246) );
  XNOR U8060 ( .A(n8245), .B(n8239), .Z(n8241) );
  XOR U8061 ( .A(n8247), .B(n8248), .Z(n8239) );
  AND U8062 ( .A(n104), .B(n8249), .Z(n8248) );
  XNOR U8063 ( .A(n8250), .B(n8251), .Z(n8245) );
  AND U8064 ( .A(n96), .B(n8252), .Z(n8251) );
  XOR U8065 ( .A(p_input[119]), .B(n8250), .Z(n8252) );
  XNOR U8066 ( .A(n8253), .B(n8254), .Z(n8250) );
  AND U8067 ( .A(n100), .B(n8249), .Z(n8254) );
  XNOR U8068 ( .A(n8253), .B(n8247), .Z(n8249) );
  XOR U8069 ( .A(n8255), .B(n8256), .Z(n8247) );
  AND U8070 ( .A(n115), .B(n8257), .Z(n8256) );
  XNOR U8071 ( .A(n8258), .B(n8259), .Z(n8253) );
  AND U8072 ( .A(n107), .B(n8260), .Z(n8259) );
  XOR U8073 ( .A(p_input[151]), .B(n8258), .Z(n8260) );
  XNOR U8074 ( .A(n8261), .B(n8262), .Z(n8258) );
  AND U8075 ( .A(n111), .B(n8257), .Z(n8262) );
  XNOR U8076 ( .A(n8261), .B(n8255), .Z(n8257) );
  XOR U8077 ( .A(n8263), .B(n8264), .Z(n8255) );
  AND U8078 ( .A(n126), .B(n8265), .Z(n8264) );
  XNOR U8079 ( .A(n8266), .B(n8267), .Z(n8261) );
  AND U8080 ( .A(n118), .B(n8268), .Z(n8267) );
  XOR U8081 ( .A(p_input[183]), .B(n8266), .Z(n8268) );
  XNOR U8082 ( .A(n8269), .B(n8270), .Z(n8266) );
  AND U8083 ( .A(n122), .B(n8265), .Z(n8270) );
  XNOR U8084 ( .A(n8269), .B(n8263), .Z(n8265) );
  XOR U8085 ( .A(n8271), .B(n8272), .Z(n8263) );
  AND U8086 ( .A(n137), .B(n8273), .Z(n8272) );
  XNOR U8087 ( .A(n8274), .B(n8275), .Z(n8269) );
  AND U8088 ( .A(n129), .B(n8276), .Z(n8275) );
  XOR U8089 ( .A(p_input[215]), .B(n8274), .Z(n8276) );
  XNOR U8090 ( .A(n8277), .B(n8278), .Z(n8274) );
  AND U8091 ( .A(n133), .B(n8273), .Z(n8278) );
  XNOR U8092 ( .A(n8277), .B(n8271), .Z(n8273) );
  XOR U8093 ( .A(n8279), .B(n8280), .Z(n8271) );
  AND U8094 ( .A(n148), .B(n8281), .Z(n8280) );
  XNOR U8095 ( .A(n8282), .B(n8283), .Z(n8277) );
  AND U8096 ( .A(n140), .B(n8284), .Z(n8283) );
  XOR U8097 ( .A(p_input[247]), .B(n8282), .Z(n8284) );
  XNOR U8098 ( .A(n8285), .B(n8286), .Z(n8282) );
  AND U8099 ( .A(n144), .B(n8281), .Z(n8286) );
  XNOR U8100 ( .A(n8285), .B(n8279), .Z(n8281) );
  XOR U8101 ( .A(n8287), .B(n8288), .Z(n8279) );
  AND U8102 ( .A(n159), .B(n8289), .Z(n8288) );
  XNOR U8103 ( .A(n8290), .B(n8291), .Z(n8285) );
  AND U8104 ( .A(n151), .B(n8292), .Z(n8291) );
  XOR U8105 ( .A(p_input[279]), .B(n8290), .Z(n8292) );
  XNOR U8106 ( .A(n8293), .B(n8294), .Z(n8290) );
  AND U8107 ( .A(n155), .B(n8289), .Z(n8294) );
  XNOR U8108 ( .A(n8293), .B(n8287), .Z(n8289) );
  XOR U8109 ( .A(n8295), .B(n8296), .Z(n8287) );
  AND U8110 ( .A(n170), .B(n8297), .Z(n8296) );
  XNOR U8111 ( .A(n8298), .B(n8299), .Z(n8293) );
  AND U8112 ( .A(n162), .B(n8300), .Z(n8299) );
  XOR U8113 ( .A(p_input[311]), .B(n8298), .Z(n8300) );
  XNOR U8114 ( .A(n8301), .B(n8302), .Z(n8298) );
  AND U8115 ( .A(n166), .B(n8297), .Z(n8302) );
  XNOR U8116 ( .A(n8301), .B(n8295), .Z(n8297) );
  XOR U8117 ( .A(n8303), .B(n8304), .Z(n8295) );
  AND U8118 ( .A(n181), .B(n8305), .Z(n8304) );
  XNOR U8119 ( .A(n8306), .B(n8307), .Z(n8301) );
  AND U8120 ( .A(n173), .B(n8308), .Z(n8307) );
  XOR U8121 ( .A(p_input[343]), .B(n8306), .Z(n8308) );
  XNOR U8122 ( .A(n8309), .B(n8310), .Z(n8306) );
  AND U8123 ( .A(n177), .B(n8305), .Z(n8310) );
  XNOR U8124 ( .A(n8309), .B(n8303), .Z(n8305) );
  XOR U8125 ( .A(n8311), .B(n8312), .Z(n8303) );
  AND U8126 ( .A(n192), .B(n8313), .Z(n8312) );
  XNOR U8127 ( .A(n8314), .B(n8315), .Z(n8309) );
  AND U8128 ( .A(n184), .B(n8316), .Z(n8315) );
  XOR U8129 ( .A(p_input[375]), .B(n8314), .Z(n8316) );
  XNOR U8130 ( .A(n8317), .B(n8318), .Z(n8314) );
  AND U8131 ( .A(n188), .B(n8313), .Z(n8318) );
  XNOR U8132 ( .A(n8317), .B(n8311), .Z(n8313) );
  XOR U8133 ( .A(n8319), .B(n8320), .Z(n8311) );
  AND U8134 ( .A(n203), .B(n8321), .Z(n8320) );
  XNOR U8135 ( .A(n8322), .B(n8323), .Z(n8317) );
  AND U8136 ( .A(n195), .B(n8324), .Z(n8323) );
  XOR U8137 ( .A(p_input[407]), .B(n8322), .Z(n8324) );
  XNOR U8138 ( .A(n8325), .B(n8326), .Z(n8322) );
  AND U8139 ( .A(n199), .B(n8321), .Z(n8326) );
  XNOR U8140 ( .A(n8325), .B(n8319), .Z(n8321) );
  XOR U8141 ( .A(n8327), .B(n8328), .Z(n8319) );
  AND U8142 ( .A(n214), .B(n8329), .Z(n8328) );
  XNOR U8143 ( .A(n8330), .B(n8331), .Z(n8325) );
  AND U8144 ( .A(n206), .B(n8332), .Z(n8331) );
  XOR U8145 ( .A(p_input[439]), .B(n8330), .Z(n8332) );
  XNOR U8146 ( .A(n8333), .B(n8334), .Z(n8330) );
  AND U8147 ( .A(n210), .B(n8329), .Z(n8334) );
  XNOR U8148 ( .A(n8333), .B(n8327), .Z(n8329) );
  XOR U8149 ( .A(n8335), .B(n8336), .Z(n8327) );
  AND U8150 ( .A(n225), .B(n8337), .Z(n8336) );
  XNOR U8151 ( .A(n8338), .B(n8339), .Z(n8333) );
  AND U8152 ( .A(n217), .B(n8340), .Z(n8339) );
  XOR U8153 ( .A(p_input[471]), .B(n8338), .Z(n8340) );
  XNOR U8154 ( .A(n8341), .B(n8342), .Z(n8338) );
  AND U8155 ( .A(n221), .B(n8337), .Z(n8342) );
  XNOR U8156 ( .A(n8341), .B(n8335), .Z(n8337) );
  XOR U8157 ( .A(n8343), .B(n8344), .Z(n8335) );
  AND U8158 ( .A(n236), .B(n8345), .Z(n8344) );
  XNOR U8159 ( .A(n8346), .B(n8347), .Z(n8341) );
  AND U8160 ( .A(n228), .B(n8348), .Z(n8347) );
  XOR U8161 ( .A(p_input[503]), .B(n8346), .Z(n8348) );
  XNOR U8162 ( .A(n8349), .B(n8350), .Z(n8346) );
  AND U8163 ( .A(n232), .B(n8345), .Z(n8350) );
  XNOR U8164 ( .A(n8349), .B(n8343), .Z(n8345) );
  XOR U8165 ( .A(n8351), .B(n8352), .Z(n8343) );
  AND U8166 ( .A(n247), .B(n8353), .Z(n8352) );
  XNOR U8167 ( .A(n8354), .B(n8355), .Z(n8349) );
  AND U8168 ( .A(n239), .B(n8356), .Z(n8355) );
  XOR U8169 ( .A(p_input[535]), .B(n8354), .Z(n8356) );
  XNOR U8170 ( .A(n8357), .B(n8358), .Z(n8354) );
  AND U8171 ( .A(n243), .B(n8353), .Z(n8358) );
  XNOR U8172 ( .A(n8357), .B(n8351), .Z(n8353) );
  XOR U8173 ( .A(n8359), .B(n8360), .Z(n8351) );
  AND U8174 ( .A(n258), .B(n8361), .Z(n8360) );
  XNOR U8175 ( .A(n8362), .B(n8363), .Z(n8357) );
  AND U8176 ( .A(n250), .B(n8364), .Z(n8363) );
  XOR U8177 ( .A(p_input[567]), .B(n8362), .Z(n8364) );
  XNOR U8178 ( .A(n8365), .B(n8366), .Z(n8362) );
  AND U8179 ( .A(n254), .B(n8361), .Z(n8366) );
  XNOR U8180 ( .A(n8365), .B(n8359), .Z(n8361) );
  XOR U8181 ( .A(n8367), .B(n8368), .Z(n8359) );
  AND U8182 ( .A(n269), .B(n8369), .Z(n8368) );
  XNOR U8183 ( .A(n8370), .B(n8371), .Z(n8365) );
  AND U8184 ( .A(n261), .B(n8372), .Z(n8371) );
  XOR U8185 ( .A(p_input[599]), .B(n8370), .Z(n8372) );
  XNOR U8186 ( .A(n8373), .B(n8374), .Z(n8370) );
  AND U8187 ( .A(n265), .B(n8369), .Z(n8374) );
  XNOR U8188 ( .A(n8373), .B(n8367), .Z(n8369) );
  XOR U8189 ( .A(n8375), .B(n8376), .Z(n8367) );
  AND U8190 ( .A(n280), .B(n8377), .Z(n8376) );
  XNOR U8191 ( .A(n8378), .B(n8379), .Z(n8373) );
  AND U8192 ( .A(n272), .B(n8380), .Z(n8379) );
  XOR U8193 ( .A(p_input[631]), .B(n8378), .Z(n8380) );
  XNOR U8194 ( .A(n8381), .B(n8382), .Z(n8378) );
  AND U8195 ( .A(n276), .B(n8377), .Z(n8382) );
  XNOR U8196 ( .A(n8381), .B(n8375), .Z(n8377) );
  XOR U8197 ( .A(n8383), .B(n8384), .Z(n8375) );
  AND U8198 ( .A(n291), .B(n8385), .Z(n8384) );
  XNOR U8199 ( .A(n8386), .B(n8387), .Z(n8381) );
  AND U8200 ( .A(n283), .B(n8388), .Z(n8387) );
  XOR U8201 ( .A(p_input[663]), .B(n8386), .Z(n8388) );
  XNOR U8202 ( .A(n8389), .B(n8390), .Z(n8386) );
  AND U8203 ( .A(n287), .B(n8385), .Z(n8390) );
  XNOR U8204 ( .A(n8389), .B(n8383), .Z(n8385) );
  XOR U8205 ( .A(n8391), .B(n8392), .Z(n8383) );
  AND U8206 ( .A(n302), .B(n8393), .Z(n8392) );
  XNOR U8207 ( .A(n8394), .B(n8395), .Z(n8389) );
  AND U8208 ( .A(n294), .B(n8396), .Z(n8395) );
  XOR U8209 ( .A(p_input[695]), .B(n8394), .Z(n8396) );
  XNOR U8210 ( .A(n8397), .B(n8398), .Z(n8394) );
  AND U8211 ( .A(n298), .B(n8393), .Z(n8398) );
  XNOR U8212 ( .A(n8397), .B(n8391), .Z(n8393) );
  XOR U8213 ( .A(n8399), .B(n8400), .Z(n8391) );
  AND U8214 ( .A(n313), .B(n8401), .Z(n8400) );
  XNOR U8215 ( .A(n8402), .B(n8403), .Z(n8397) );
  AND U8216 ( .A(n305), .B(n8404), .Z(n8403) );
  XOR U8217 ( .A(p_input[727]), .B(n8402), .Z(n8404) );
  XNOR U8218 ( .A(n8405), .B(n8406), .Z(n8402) );
  AND U8219 ( .A(n309), .B(n8401), .Z(n8406) );
  XNOR U8220 ( .A(n8405), .B(n8399), .Z(n8401) );
  XOR U8221 ( .A(n8407), .B(n8408), .Z(n8399) );
  AND U8222 ( .A(n324), .B(n8409), .Z(n8408) );
  XNOR U8223 ( .A(n8410), .B(n8411), .Z(n8405) );
  AND U8224 ( .A(n316), .B(n8412), .Z(n8411) );
  XOR U8225 ( .A(p_input[759]), .B(n8410), .Z(n8412) );
  XNOR U8226 ( .A(n8413), .B(n8414), .Z(n8410) );
  AND U8227 ( .A(n320), .B(n8409), .Z(n8414) );
  XNOR U8228 ( .A(n8413), .B(n8407), .Z(n8409) );
  XOR U8229 ( .A(n8415), .B(n8416), .Z(n8407) );
  AND U8230 ( .A(n335), .B(n8417), .Z(n8416) );
  XNOR U8231 ( .A(n8418), .B(n8419), .Z(n8413) );
  AND U8232 ( .A(n327), .B(n8420), .Z(n8419) );
  XOR U8233 ( .A(p_input[791]), .B(n8418), .Z(n8420) );
  XNOR U8234 ( .A(n8421), .B(n8422), .Z(n8418) );
  AND U8235 ( .A(n331), .B(n8417), .Z(n8422) );
  XNOR U8236 ( .A(n8421), .B(n8415), .Z(n8417) );
  XOR U8237 ( .A(n8423), .B(n8424), .Z(n8415) );
  AND U8238 ( .A(n346), .B(n8425), .Z(n8424) );
  XNOR U8239 ( .A(n8426), .B(n8427), .Z(n8421) );
  AND U8240 ( .A(n338), .B(n8428), .Z(n8427) );
  XOR U8241 ( .A(p_input[823]), .B(n8426), .Z(n8428) );
  XNOR U8242 ( .A(n8429), .B(n8430), .Z(n8426) );
  AND U8243 ( .A(n342), .B(n8425), .Z(n8430) );
  XNOR U8244 ( .A(n8429), .B(n8423), .Z(n8425) );
  XOR U8245 ( .A(n8431), .B(n8432), .Z(n8423) );
  AND U8246 ( .A(n357), .B(n8433), .Z(n8432) );
  XNOR U8247 ( .A(n8434), .B(n8435), .Z(n8429) );
  AND U8248 ( .A(n349), .B(n8436), .Z(n8435) );
  XOR U8249 ( .A(p_input[855]), .B(n8434), .Z(n8436) );
  XNOR U8250 ( .A(n8437), .B(n8438), .Z(n8434) );
  AND U8251 ( .A(n353), .B(n8433), .Z(n8438) );
  XNOR U8252 ( .A(n8437), .B(n8431), .Z(n8433) );
  XOR U8253 ( .A(n8439), .B(n8440), .Z(n8431) );
  AND U8254 ( .A(n368), .B(n8441), .Z(n8440) );
  XNOR U8255 ( .A(n8442), .B(n8443), .Z(n8437) );
  AND U8256 ( .A(n360), .B(n8444), .Z(n8443) );
  XOR U8257 ( .A(p_input[887]), .B(n8442), .Z(n8444) );
  XNOR U8258 ( .A(n8445), .B(n8446), .Z(n8442) );
  AND U8259 ( .A(n364), .B(n8441), .Z(n8446) );
  XNOR U8260 ( .A(n8445), .B(n8439), .Z(n8441) );
  XOR U8261 ( .A(n8447), .B(n8448), .Z(n8439) );
  AND U8262 ( .A(n379), .B(n8449), .Z(n8448) );
  XNOR U8263 ( .A(n8450), .B(n8451), .Z(n8445) );
  AND U8264 ( .A(n371), .B(n8452), .Z(n8451) );
  XOR U8265 ( .A(p_input[919]), .B(n8450), .Z(n8452) );
  XNOR U8266 ( .A(n8453), .B(n8454), .Z(n8450) );
  AND U8267 ( .A(n375), .B(n8449), .Z(n8454) );
  XNOR U8268 ( .A(n8453), .B(n8447), .Z(n8449) );
  XOR U8269 ( .A(n8455), .B(n8456), .Z(n8447) );
  AND U8270 ( .A(n390), .B(n8457), .Z(n8456) );
  XNOR U8271 ( .A(n8458), .B(n8459), .Z(n8453) );
  AND U8272 ( .A(n382), .B(n8460), .Z(n8459) );
  XOR U8273 ( .A(p_input[951]), .B(n8458), .Z(n8460) );
  XNOR U8274 ( .A(n8461), .B(n8462), .Z(n8458) );
  AND U8275 ( .A(n386), .B(n8457), .Z(n8462) );
  XNOR U8276 ( .A(n8461), .B(n8455), .Z(n8457) );
  XOR U8277 ( .A(n8463), .B(n8464), .Z(n8455) );
  AND U8278 ( .A(n401), .B(n8465), .Z(n8464) );
  XNOR U8279 ( .A(n8466), .B(n8467), .Z(n8461) );
  AND U8280 ( .A(n393), .B(n8468), .Z(n8467) );
  XOR U8281 ( .A(p_input[983]), .B(n8466), .Z(n8468) );
  XNOR U8282 ( .A(n8469), .B(n8470), .Z(n8466) );
  AND U8283 ( .A(n397), .B(n8465), .Z(n8470) );
  XNOR U8284 ( .A(n8469), .B(n8463), .Z(n8465) );
  XOR U8285 ( .A(n8471), .B(n8472), .Z(n8463) );
  AND U8286 ( .A(n412), .B(n8473), .Z(n8472) );
  XNOR U8287 ( .A(n8474), .B(n8475), .Z(n8469) );
  AND U8288 ( .A(n404), .B(n8476), .Z(n8475) );
  XOR U8289 ( .A(p_input[1015]), .B(n8474), .Z(n8476) );
  XNOR U8290 ( .A(n8477), .B(n8478), .Z(n8474) );
  AND U8291 ( .A(n408), .B(n8473), .Z(n8478) );
  XNOR U8292 ( .A(n8477), .B(n8471), .Z(n8473) );
  XOR U8293 ( .A(n8479), .B(n8480), .Z(n8471) );
  AND U8294 ( .A(n423), .B(n8481), .Z(n8480) );
  XNOR U8295 ( .A(n8482), .B(n8483), .Z(n8477) );
  AND U8296 ( .A(n415), .B(n8484), .Z(n8483) );
  XOR U8297 ( .A(p_input[1047]), .B(n8482), .Z(n8484) );
  XNOR U8298 ( .A(n8485), .B(n8486), .Z(n8482) );
  AND U8299 ( .A(n419), .B(n8481), .Z(n8486) );
  XNOR U8300 ( .A(n8485), .B(n8479), .Z(n8481) );
  XOR U8301 ( .A(n8487), .B(n8488), .Z(n8479) );
  AND U8302 ( .A(n434), .B(n8489), .Z(n8488) );
  XNOR U8303 ( .A(n8490), .B(n8491), .Z(n8485) );
  AND U8304 ( .A(n426), .B(n8492), .Z(n8491) );
  XOR U8305 ( .A(p_input[1079]), .B(n8490), .Z(n8492) );
  XNOR U8306 ( .A(n8493), .B(n8494), .Z(n8490) );
  AND U8307 ( .A(n430), .B(n8489), .Z(n8494) );
  XNOR U8308 ( .A(n8493), .B(n8487), .Z(n8489) );
  XOR U8309 ( .A(n8495), .B(n8496), .Z(n8487) );
  AND U8310 ( .A(n445), .B(n8497), .Z(n8496) );
  XNOR U8311 ( .A(n8498), .B(n8499), .Z(n8493) );
  AND U8312 ( .A(n437), .B(n8500), .Z(n8499) );
  XOR U8313 ( .A(p_input[1111]), .B(n8498), .Z(n8500) );
  XNOR U8314 ( .A(n8501), .B(n8502), .Z(n8498) );
  AND U8315 ( .A(n441), .B(n8497), .Z(n8502) );
  XNOR U8316 ( .A(n8501), .B(n8495), .Z(n8497) );
  XOR U8317 ( .A(n8503), .B(n8504), .Z(n8495) );
  AND U8318 ( .A(n456), .B(n8505), .Z(n8504) );
  XNOR U8319 ( .A(n8506), .B(n8507), .Z(n8501) );
  AND U8320 ( .A(n448), .B(n8508), .Z(n8507) );
  XOR U8321 ( .A(p_input[1143]), .B(n8506), .Z(n8508) );
  XNOR U8322 ( .A(n8509), .B(n8510), .Z(n8506) );
  AND U8323 ( .A(n452), .B(n8505), .Z(n8510) );
  XNOR U8324 ( .A(n8509), .B(n8503), .Z(n8505) );
  XOR U8325 ( .A(n8511), .B(n8512), .Z(n8503) );
  AND U8326 ( .A(n467), .B(n8513), .Z(n8512) );
  XNOR U8327 ( .A(n8514), .B(n8515), .Z(n8509) );
  AND U8328 ( .A(n459), .B(n8516), .Z(n8515) );
  XOR U8329 ( .A(p_input[1175]), .B(n8514), .Z(n8516) );
  XNOR U8330 ( .A(n8517), .B(n8518), .Z(n8514) );
  AND U8331 ( .A(n463), .B(n8513), .Z(n8518) );
  XNOR U8332 ( .A(n8517), .B(n8511), .Z(n8513) );
  XOR U8333 ( .A(n8519), .B(n8520), .Z(n8511) );
  AND U8334 ( .A(n478), .B(n8521), .Z(n8520) );
  XNOR U8335 ( .A(n8522), .B(n8523), .Z(n8517) );
  AND U8336 ( .A(n470), .B(n8524), .Z(n8523) );
  XOR U8337 ( .A(p_input[1207]), .B(n8522), .Z(n8524) );
  XNOR U8338 ( .A(n8525), .B(n8526), .Z(n8522) );
  AND U8339 ( .A(n474), .B(n8521), .Z(n8526) );
  XNOR U8340 ( .A(n8525), .B(n8519), .Z(n8521) );
  XOR U8341 ( .A(n8527), .B(n8528), .Z(n8519) );
  AND U8342 ( .A(n489), .B(n8529), .Z(n8528) );
  XNOR U8343 ( .A(n8530), .B(n8531), .Z(n8525) );
  AND U8344 ( .A(n481), .B(n8532), .Z(n8531) );
  XOR U8345 ( .A(p_input[1239]), .B(n8530), .Z(n8532) );
  XNOR U8346 ( .A(n8533), .B(n8534), .Z(n8530) );
  AND U8347 ( .A(n485), .B(n8529), .Z(n8534) );
  XNOR U8348 ( .A(n8533), .B(n8527), .Z(n8529) );
  XOR U8349 ( .A(n8535), .B(n8536), .Z(n8527) );
  AND U8350 ( .A(n500), .B(n8537), .Z(n8536) );
  XNOR U8351 ( .A(n8538), .B(n8539), .Z(n8533) );
  AND U8352 ( .A(n492), .B(n8540), .Z(n8539) );
  XOR U8353 ( .A(p_input[1271]), .B(n8538), .Z(n8540) );
  XNOR U8354 ( .A(n8541), .B(n8542), .Z(n8538) );
  AND U8355 ( .A(n496), .B(n8537), .Z(n8542) );
  XNOR U8356 ( .A(n8541), .B(n8535), .Z(n8537) );
  XOR U8357 ( .A(n8543), .B(n8544), .Z(n8535) );
  AND U8358 ( .A(n511), .B(n8545), .Z(n8544) );
  XNOR U8359 ( .A(n8546), .B(n8547), .Z(n8541) );
  AND U8360 ( .A(n503), .B(n8548), .Z(n8547) );
  XOR U8361 ( .A(p_input[1303]), .B(n8546), .Z(n8548) );
  XNOR U8362 ( .A(n8549), .B(n8550), .Z(n8546) );
  AND U8363 ( .A(n507), .B(n8545), .Z(n8550) );
  XNOR U8364 ( .A(n8549), .B(n8543), .Z(n8545) );
  XOR U8365 ( .A(n8551), .B(n8552), .Z(n8543) );
  AND U8366 ( .A(n522), .B(n8553), .Z(n8552) );
  XNOR U8367 ( .A(n8554), .B(n8555), .Z(n8549) );
  AND U8368 ( .A(n514), .B(n8556), .Z(n8555) );
  XOR U8369 ( .A(p_input[1335]), .B(n8554), .Z(n8556) );
  XNOR U8370 ( .A(n8557), .B(n8558), .Z(n8554) );
  AND U8371 ( .A(n518), .B(n8553), .Z(n8558) );
  XNOR U8372 ( .A(n8557), .B(n8551), .Z(n8553) );
  XOR U8373 ( .A(n8559), .B(n8560), .Z(n8551) );
  AND U8374 ( .A(n533), .B(n8561), .Z(n8560) );
  XNOR U8375 ( .A(n8562), .B(n8563), .Z(n8557) );
  AND U8376 ( .A(n525), .B(n8564), .Z(n8563) );
  XOR U8377 ( .A(p_input[1367]), .B(n8562), .Z(n8564) );
  XNOR U8378 ( .A(n8565), .B(n8566), .Z(n8562) );
  AND U8379 ( .A(n529), .B(n8561), .Z(n8566) );
  XNOR U8380 ( .A(n8565), .B(n8559), .Z(n8561) );
  XOR U8381 ( .A(n8567), .B(n8568), .Z(n8559) );
  AND U8382 ( .A(n544), .B(n8569), .Z(n8568) );
  XNOR U8383 ( .A(n8570), .B(n8571), .Z(n8565) );
  AND U8384 ( .A(n536), .B(n8572), .Z(n8571) );
  XOR U8385 ( .A(p_input[1399]), .B(n8570), .Z(n8572) );
  XNOR U8386 ( .A(n8573), .B(n8574), .Z(n8570) );
  AND U8387 ( .A(n540), .B(n8569), .Z(n8574) );
  XNOR U8388 ( .A(n8573), .B(n8567), .Z(n8569) );
  XOR U8389 ( .A(n8575), .B(n8576), .Z(n8567) );
  AND U8390 ( .A(n555), .B(n8577), .Z(n8576) );
  XNOR U8391 ( .A(n8578), .B(n8579), .Z(n8573) );
  AND U8392 ( .A(n547), .B(n8580), .Z(n8579) );
  XOR U8393 ( .A(p_input[1431]), .B(n8578), .Z(n8580) );
  XNOR U8394 ( .A(n8581), .B(n8582), .Z(n8578) );
  AND U8395 ( .A(n551), .B(n8577), .Z(n8582) );
  XNOR U8396 ( .A(n8581), .B(n8575), .Z(n8577) );
  XOR U8397 ( .A(n8583), .B(n8584), .Z(n8575) );
  AND U8398 ( .A(n566), .B(n8585), .Z(n8584) );
  XNOR U8399 ( .A(n8586), .B(n8587), .Z(n8581) );
  AND U8400 ( .A(n558), .B(n8588), .Z(n8587) );
  XOR U8401 ( .A(p_input[1463]), .B(n8586), .Z(n8588) );
  XNOR U8402 ( .A(n8589), .B(n8590), .Z(n8586) );
  AND U8403 ( .A(n562), .B(n8585), .Z(n8590) );
  XNOR U8404 ( .A(n8589), .B(n8583), .Z(n8585) );
  XOR U8405 ( .A(n8591), .B(n8592), .Z(n8583) );
  AND U8406 ( .A(n577), .B(n8593), .Z(n8592) );
  XNOR U8407 ( .A(n8594), .B(n8595), .Z(n8589) );
  AND U8408 ( .A(n569), .B(n8596), .Z(n8595) );
  XOR U8409 ( .A(p_input[1495]), .B(n8594), .Z(n8596) );
  XNOR U8410 ( .A(n8597), .B(n8598), .Z(n8594) );
  AND U8411 ( .A(n573), .B(n8593), .Z(n8598) );
  XNOR U8412 ( .A(n8597), .B(n8591), .Z(n8593) );
  XOR U8413 ( .A(n8599), .B(n8600), .Z(n8591) );
  AND U8414 ( .A(n588), .B(n8601), .Z(n8600) );
  XNOR U8415 ( .A(n8602), .B(n8603), .Z(n8597) );
  AND U8416 ( .A(n580), .B(n8604), .Z(n8603) );
  XOR U8417 ( .A(p_input[1527]), .B(n8602), .Z(n8604) );
  XNOR U8418 ( .A(n8605), .B(n8606), .Z(n8602) );
  AND U8419 ( .A(n584), .B(n8601), .Z(n8606) );
  XNOR U8420 ( .A(n8605), .B(n8599), .Z(n8601) );
  XOR U8421 ( .A(n8607), .B(n8608), .Z(n8599) );
  AND U8422 ( .A(n599), .B(n8609), .Z(n8608) );
  XNOR U8423 ( .A(n8610), .B(n8611), .Z(n8605) );
  AND U8424 ( .A(n591), .B(n8612), .Z(n8611) );
  XOR U8425 ( .A(p_input[1559]), .B(n8610), .Z(n8612) );
  XNOR U8426 ( .A(n8613), .B(n8614), .Z(n8610) );
  AND U8427 ( .A(n595), .B(n8609), .Z(n8614) );
  XNOR U8428 ( .A(n8613), .B(n8607), .Z(n8609) );
  XOR U8429 ( .A(n8615), .B(n8616), .Z(n8607) );
  AND U8430 ( .A(n610), .B(n8617), .Z(n8616) );
  XNOR U8431 ( .A(n8618), .B(n8619), .Z(n8613) );
  AND U8432 ( .A(n602), .B(n8620), .Z(n8619) );
  XOR U8433 ( .A(p_input[1591]), .B(n8618), .Z(n8620) );
  XNOR U8434 ( .A(n8621), .B(n8622), .Z(n8618) );
  AND U8435 ( .A(n606), .B(n8617), .Z(n8622) );
  XNOR U8436 ( .A(n8621), .B(n8615), .Z(n8617) );
  XOR U8437 ( .A(n8623), .B(n8624), .Z(n8615) );
  AND U8438 ( .A(n621), .B(n8625), .Z(n8624) );
  XNOR U8439 ( .A(n8626), .B(n8627), .Z(n8621) );
  AND U8440 ( .A(n613), .B(n8628), .Z(n8627) );
  XOR U8441 ( .A(p_input[1623]), .B(n8626), .Z(n8628) );
  XNOR U8442 ( .A(n8629), .B(n8630), .Z(n8626) );
  AND U8443 ( .A(n617), .B(n8625), .Z(n8630) );
  XNOR U8444 ( .A(n8629), .B(n8623), .Z(n8625) );
  XOR U8445 ( .A(n8631), .B(n8632), .Z(n8623) );
  AND U8446 ( .A(n632), .B(n8633), .Z(n8632) );
  XNOR U8447 ( .A(n8634), .B(n8635), .Z(n8629) );
  AND U8448 ( .A(n624), .B(n8636), .Z(n8635) );
  XOR U8449 ( .A(p_input[1655]), .B(n8634), .Z(n8636) );
  XNOR U8450 ( .A(n8637), .B(n8638), .Z(n8634) );
  AND U8451 ( .A(n628), .B(n8633), .Z(n8638) );
  XNOR U8452 ( .A(n8637), .B(n8631), .Z(n8633) );
  XOR U8453 ( .A(n8639), .B(n8640), .Z(n8631) );
  AND U8454 ( .A(n643), .B(n8641), .Z(n8640) );
  XNOR U8455 ( .A(n8642), .B(n8643), .Z(n8637) );
  AND U8456 ( .A(n635), .B(n8644), .Z(n8643) );
  XOR U8457 ( .A(p_input[1687]), .B(n8642), .Z(n8644) );
  XNOR U8458 ( .A(n8645), .B(n8646), .Z(n8642) );
  AND U8459 ( .A(n639), .B(n8641), .Z(n8646) );
  XNOR U8460 ( .A(n8645), .B(n8639), .Z(n8641) );
  XOR U8461 ( .A(n8647), .B(n8648), .Z(n8639) );
  AND U8462 ( .A(n654), .B(n8649), .Z(n8648) );
  XNOR U8463 ( .A(n8650), .B(n8651), .Z(n8645) );
  AND U8464 ( .A(n646), .B(n8652), .Z(n8651) );
  XOR U8465 ( .A(p_input[1719]), .B(n8650), .Z(n8652) );
  XNOR U8466 ( .A(n8653), .B(n8654), .Z(n8650) );
  AND U8467 ( .A(n650), .B(n8649), .Z(n8654) );
  XNOR U8468 ( .A(n8653), .B(n8647), .Z(n8649) );
  XOR U8469 ( .A(n8655), .B(n8656), .Z(n8647) );
  AND U8470 ( .A(n665), .B(n8657), .Z(n8656) );
  XNOR U8471 ( .A(n8658), .B(n8659), .Z(n8653) );
  AND U8472 ( .A(n657), .B(n8660), .Z(n8659) );
  XOR U8473 ( .A(p_input[1751]), .B(n8658), .Z(n8660) );
  XNOR U8474 ( .A(n8661), .B(n8662), .Z(n8658) );
  AND U8475 ( .A(n661), .B(n8657), .Z(n8662) );
  XNOR U8476 ( .A(n8661), .B(n8655), .Z(n8657) );
  XOR U8477 ( .A(n8663), .B(n8664), .Z(n8655) );
  AND U8478 ( .A(n676), .B(n8665), .Z(n8664) );
  XNOR U8479 ( .A(n8666), .B(n8667), .Z(n8661) );
  AND U8480 ( .A(n668), .B(n8668), .Z(n8667) );
  XOR U8481 ( .A(p_input[1783]), .B(n8666), .Z(n8668) );
  XNOR U8482 ( .A(n8669), .B(n8670), .Z(n8666) );
  AND U8483 ( .A(n672), .B(n8665), .Z(n8670) );
  XNOR U8484 ( .A(n8669), .B(n8663), .Z(n8665) );
  XOR U8485 ( .A(n8671), .B(n8672), .Z(n8663) );
  AND U8486 ( .A(n687), .B(n8673), .Z(n8672) );
  XNOR U8487 ( .A(n8674), .B(n8675), .Z(n8669) );
  AND U8488 ( .A(n679), .B(n8676), .Z(n8675) );
  XOR U8489 ( .A(p_input[1815]), .B(n8674), .Z(n8676) );
  XNOR U8490 ( .A(n8677), .B(n8678), .Z(n8674) );
  AND U8491 ( .A(n683), .B(n8673), .Z(n8678) );
  XNOR U8492 ( .A(n8677), .B(n8671), .Z(n8673) );
  XOR U8493 ( .A(n8679), .B(n8680), .Z(n8671) );
  AND U8494 ( .A(n698), .B(n8681), .Z(n8680) );
  XNOR U8495 ( .A(n8682), .B(n8683), .Z(n8677) );
  AND U8496 ( .A(n690), .B(n8684), .Z(n8683) );
  XOR U8497 ( .A(p_input[1847]), .B(n8682), .Z(n8684) );
  XNOR U8498 ( .A(n8685), .B(n8686), .Z(n8682) );
  AND U8499 ( .A(n694), .B(n8681), .Z(n8686) );
  XNOR U8500 ( .A(n8685), .B(n8679), .Z(n8681) );
  XOR U8501 ( .A(n8687), .B(n8688), .Z(n8679) );
  AND U8502 ( .A(n709), .B(n8689), .Z(n8688) );
  XNOR U8503 ( .A(n8690), .B(n8691), .Z(n8685) );
  AND U8504 ( .A(n701), .B(n8692), .Z(n8691) );
  XOR U8505 ( .A(p_input[1879]), .B(n8690), .Z(n8692) );
  XNOR U8506 ( .A(n8693), .B(n8694), .Z(n8690) );
  AND U8507 ( .A(n705), .B(n8689), .Z(n8694) );
  XNOR U8508 ( .A(n8693), .B(n8687), .Z(n8689) );
  XOR U8509 ( .A(n8695), .B(n8696), .Z(n8687) );
  AND U8510 ( .A(n720), .B(n8697), .Z(n8696) );
  XNOR U8511 ( .A(n8698), .B(n8699), .Z(n8693) );
  AND U8512 ( .A(n712), .B(n8700), .Z(n8699) );
  XOR U8513 ( .A(p_input[1911]), .B(n8698), .Z(n8700) );
  XNOR U8514 ( .A(n8701), .B(n8702), .Z(n8698) );
  AND U8515 ( .A(n716), .B(n8697), .Z(n8702) );
  XNOR U8516 ( .A(n8701), .B(n8695), .Z(n8697) );
  XOR U8517 ( .A(n8703), .B(n8704), .Z(n8695) );
  AND U8518 ( .A(n731), .B(n8705), .Z(n8704) );
  XNOR U8519 ( .A(n8706), .B(n8707), .Z(n8701) );
  AND U8520 ( .A(n723), .B(n8708), .Z(n8707) );
  XOR U8521 ( .A(p_input[1943]), .B(n8706), .Z(n8708) );
  XNOR U8522 ( .A(n8709), .B(n8710), .Z(n8706) );
  AND U8523 ( .A(n727), .B(n8705), .Z(n8710) );
  XNOR U8524 ( .A(n8709), .B(n8703), .Z(n8705) );
  XOR U8525 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n8711), .Z(n8703) );
  AND U8526 ( .A(n741), .B(n8712), .Z(n8711) );
  XNOR U8527 ( .A(n8713), .B(n8714), .Z(n8709) );
  AND U8528 ( .A(n734), .B(n8715), .Z(n8714) );
  XOR U8529 ( .A(p_input[1975]), .B(n8713), .Z(n8715) );
  XNOR U8530 ( .A(n8716), .B(n8717), .Z(n8713) );
  AND U8531 ( .A(n738), .B(n8712), .Z(n8717) );
  XOR U8532 ( .A(n8718), .B(n8716), .Z(n8712) );
  IV U8533 ( .A(\knn_comb_/min_val_out[0][23] ), .Z(n8718) );
  IV U8534 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .Z(n8716) );
  XOR U8535 ( .A(n29), .B(n8719), .Z(o[22]) );
  AND U8536 ( .A(n58), .B(n8720), .Z(n29) );
  XOR U8537 ( .A(n30), .B(n8719), .Z(n8720) );
  XOR U8538 ( .A(n8721), .B(n8722), .Z(n8719) );
  AND U8539 ( .A(n70), .B(n8723), .Z(n8722) );
  XOR U8540 ( .A(n8724), .B(n8725), .Z(n30) );
  AND U8541 ( .A(n62), .B(n8726), .Z(n8725) );
  XOR U8542 ( .A(p_input[22]), .B(n8724), .Z(n8726) );
  XNOR U8543 ( .A(n8727), .B(n8728), .Z(n8724) );
  AND U8544 ( .A(n66), .B(n8723), .Z(n8728) );
  XNOR U8545 ( .A(n8727), .B(n8721), .Z(n8723) );
  XOR U8546 ( .A(n8729), .B(n8730), .Z(n8721) );
  AND U8547 ( .A(n82), .B(n8731), .Z(n8730) );
  XNOR U8548 ( .A(n8732), .B(n8733), .Z(n8727) );
  AND U8549 ( .A(n74), .B(n8734), .Z(n8733) );
  XOR U8550 ( .A(p_input[54]), .B(n8732), .Z(n8734) );
  XNOR U8551 ( .A(n8735), .B(n8736), .Z(n8732) );
  AND U8552 ( .A(n78), .B(n8731), .Z(n8736) );
  XNOR U8553 ( .A(n8735), .B(n8729), .Z(n8731) );
  XOR U8554 ( .A(n8737), .B(n8738), .Z(n8729) );
  AND U8555 ( .A(n93), .B(n8739), .Z(n8738) );
  XNOR U8556 ( .A(n8740), .B(n8741), .Z(n8735) );
  AND U8557 ( .A(n85), .B(n8742), .Z(n8741) );
  XOR U8558 ( .A(p_input[86]), .B(n8740), .Z(n8742) );
  XNOR U8559 ( .A(n8743), .B(n8744), .Z(n8740) );
  AND U8560 ( .A(n89), .B(n8739), .Z(n8744) );
  XNOR U8561 ( .A(n8743), .B(n8737), .Z(n8739) );
  XOR U8562 ( .A(n8745), .B(n8746), .Z(n8737) );
  AND U8563 ( .A(n104), .B(n8747), .Z(n8746) );
  XNOR U8564 ( .A(n8748), .B(n8749), .Z(n8743) );
  AND U8565 ( .A(n96), .B(n8750), .Z(n8749) );
  XOR U8566 ( .A(p_input[118]), .B(n8748), .Z(n8750) );
  XNOR U8567 ( .A(n8751), .B(n8752), .Z(n8748) );
  AND U8568 ( .A(n100), .B(n8747), .Z(n8752) );
  XNOR U8569 ( .A(n8751), .B(n8745), .Z(n8747) );
  XOR U8570 ( .A(n8753), .B(n8754), .Z(n8745) );
  AND U8571 ( .A(n115), .B(n8755), .Z(n8754) );
  XNOR U8572 ( .A(n8756), .B(n8757), .Z(n8751) );
  AND U8573 ( .A(n107), .B(n8758), .Z(n8757) );
  XOR U8574 ( .A(p_input[150]), .B(n8756), .Z(n8758) );
  XNOR U8575 ( .A(n8759), .B(n8760), .Z(n8756) );
  AND U8576 ( .A(n111), .B(n8755), .Z(n8760) );
  XNOR U8577 ( .A(n8759), .B(n8753), .Z(n8755) );
  XOR U8578 ( .A(n8761), .B(n8762), .Z(n8753) );
  AND U8579 ( .A(n126), .B(n8763), .Z(n8762) );
  XNOR U8580 ( .A(n8764), .B(n8765), .Z(n8759) );
  AND U8581 ( .A(n118), .B(n8766), .Z(n8765) );
  XOR U8582 ( .A(p_input[182]), .B(n8764), .Z(n8766) );
  XNOR U8583 ( .A(n8767), .B(n8768), .Z(n8764) );
  AND U8584 ( .A(n122), .B(n8763), .Z(n8768) );
  XNOR U8585 ( .A(n8767), .B(n8761), .Z(n8763) );
  XOR U8586 ( .A(n8769), .B(n8770), .Z(n8761) );
  AND U8587 ( .A(n137), .B(n8771), .Z(n8770) );
  XNOR U8588 ( .A(n8772), .B(n8773), .Z(n8767) );
  AND U8589 ( .A(n129), .B(n8774), .Z(n8773) );
  XOR U8590 ( .A(p_input[214]), .B(n8772), .Z(n8774) );
  XNOR U8591 ( .A(n8775), .B(n8776), .Z(n8772) );
  AND U8592 ( .A(n133), .B(n8771), .Z(n8776) );
  XNOR U8593 ( .A(n8775), .B(n8769), .Z(n8771) );
  XOR U8594 ( .A(n8777), .B(n8778), .Z(n8769) );
  AND U8595 ( .A(n148), .B(n8779), .Z(n8778) );
  XNOR U8596 ( .A(n8780), .B(n8781), .Z(n8775) );
  AND U8597 ( .A(n140), .B(n8782), .Z(n8781) );
  XOR U8598 ( .A(p_input[246]), .B(n8780), .Z(n8782) );
  XNOR U8599 ( .A(n8783), .B(n8784), .Z(n8780) );
  AND U8600 ( .A(n144), .B(n8779), .Z(n8784) );
  XNOR U8601 ( .A(n8783), .B(n8777), .Z(n8779) );
  XOR U8602 ( .A(n8785), .B(n8786), .Z(n8777) );
  AND U8603 ( .A(n159), .B(n8787), .Z(n8786) );
  XNOR U8604 ( .A(n8788), .B(n8789), .Z(n8783) );
  AND U8605 ( .A(n151), .B(n8790), .Z(n8789) );
  XOR U8606 ( .A(p_input[278]), .B(n8788), .Z(n8790) );
  XNOR U8607 ( .A(n8791), .B(n8792), .Z(n8788) );
  AND U8608 ( .A(n155), .B(n8787), .Z(n8792) );
  XNOR U8609 ( .A(n8791), .B(n8785), .Z(n8787) );
  XOR U8610 ( .A(n8793), .B(n8794), .Z(n8785) );
  AND U8611 ( .A(n170), .B(n8795), .Z(n8794) );
  XNOR U8612 ( .A(n8796), .B(n8797), .Z(n8791) );
  AND U8613 ( .A(n162), .B(n8798), .Z(n8797) );
  XOR U8614 ( .A(p_input[310]), .B(n8796), .Z(n8798) );
  XNOR U8615 ( .A(n8799), .B(n8800), .Z(n8796) );
  AND U8616 ( .A(n166), .B(n8795), .Z(n8800) );
  XNOR U8617 ( .A(n8799), .B(n8793), .Z(n8795) );
  XOR U8618 ( .A(n8801), .B(n8802), .Z(n8793) );
  AND U8619 ( .A(n181), .B(n8803), .Z(n8802) );
  XNOR U8620 ( .A(n8804), .B(n8805), .Z(n8799) );
  AND U8621 ( .A(n173), .B(n8806), .Z(n8805) );
  XOR U8622 ( .A(p_input[342]), .B(n8804), .Z(n8806) );
  XNOR U8623 ( .A(n8807), .B(n8808), .Z(n8804) );
  AND U8624 ( .A(n177), .B(n8803), .Z(n8808) );
  XNOR U8625 ( .A(n8807), .B(n8801), .Z(n8803) );
  XOR U8626 ( .A(n8809), .B(n8810), .Z(n8801) );
  AND U8627 ( .A(n192), .B(n8811), .Z(n8810) );
  XNOR U8628 ( .A(n8812), .B(n8813), .Z(n8807) );
  AND U8629 ( .A(n184), .B(n8814), .Z(n8813) );
  XOR U8630 ( .A(p_input[374]), .B(n8812), .Z(n8814) );
  XNOR U8631 ( .A(n8815), .B(n8816), .Z(n8812) );
  AND U8632 ( .A(n188), .B(n8811), .Z(n8816) );
  XNOR U8633 ( .A(n8815), .B(n8809), .Z(n8811) );
  XOR U8634 ( .A(n8817), .B(n8818), .Z(n8809) );
  AND U8635 ( .A(n203), .B(n8819), .Z(n8818) );
  XNOR U8636 ( .A(n8820), .B(n8821), .Z(n8815) );
  AND U8637 ( .A(n195), .B(n8822), .Z(n8821) );
  XOR U8638 ( .A(p_input[406]), .B(n8820), .Z(n8822) );
  XNOR U8639 ( .A(n8823), .B(n8824), .Z(n8820) );
  AND U8640 ( .A(n199), .B(n8819), .Z(n8824) );
  XNOR U8641 ( .A(n8823), .B(n8817), .Z(n8819) );
  XOR U8642 ( .A(n8825), .B(n8826), .Z(n8817) );
  AND U8643 ( .A(n214), .B(n8827), .Z(n8826) );
  XNOR U8644 ( .A(n8828), .B(n8829), .Z(n8823) );
  AND U8645 ( .A(n206), .B(n8830), .Z(n8829) );
  XOR U8646 ( .A(p_input[438]), .B(n8828), .Z(n8830) );
  XNOR U8647 ( .A(n8831), .B(n8832), .Z(n8828) );
  AND U8648 ( .A(n210), .B(n8827), .Z(n8832) );
  XNOR U8649 ( .A(n8831), .B(n8825), .Z(n8827) );
  XOR U8650 ( .A(n8833), .B(n8834), .Z(n8825) );
  AND U8651 ( .A(n225), .B(n8835), .Z(n8834) );
  XNOR U8652 ( .A(n8836), .B(n8837), .Z(n8831) );
  AND U8653 ( .A(n217), .B(n8838), .Z(n8837) );
  XOR U8654 ( .A(p_input[470]), .B(n8836), .Z(n8838) );
  XNOR U8655 ( .A(n8839), .B(n8840), .Z(n8836) );
  AND U8656 ( .A(n221), .B(n8835), .Z(n8840) );
  XNOR U8657 ( .A(n8839), .B(n8833), .Z(n8835) );
  XOR U8658 ( .A(n8841), .B(n8842), .Z(n8833) );
  AND U8659 ( .A(n236), .B(n8843), .Z(n8842) );
  XNOR U8660 ( .A(n8844), .B(n8845), .Z(n8839) );
  AND U8661 ( .A(n228), .B(n8846), .Z(n8845) );
  XOR U8662 ( .A(p_input[502]), .B(n8844), .Z(n8846) );
  XNOR U8663 ( .A(n8847), .B(n8848), .Z(n8844) );
  AND U8664 ( .A(n232), .B(n8843), .Z(n8848) );
  XNOR U8665 ( .A(n8847), .B(n8841), .Z(n8843) );
  XOR U8666 ( .A(n8849), .B(n8850), .Z(n8841) );
  AND U8667 ( .A(n247), .B(n8851), .Z(n8850) );
  XNOR U8668 ( .A(n8852), .B(n8853), .Z(n8847) );
  AND U8669 ( .A(n239), .B(n8854), .Z(n8853) );
  XOR U8670 ( .A(p_input[534]), .B(n8852), .Z(n8854) );
  XNOR U8671 ( .A(n8855), .B(n8856), .Z(n8852) );
  AND U8672 ( .A(n243), .B(n8851), .Z(n8856) );
  XNOR U8673 ( .A(n8855), .B(n8849), .Z(n8851) );
  XOR U8674 ( .A(n8857), .B(n8858), .Z(n8849) );
  AND U8675 ( .A(n258), .B(n8859), .Z(n8858) );
  XNOR U8676 ( .A(n8860), .B(n8861), .Z(n8855) );
  AND U8677 ( .A(n250), .B(n8862), .Z(n8861) );
  XOR U8678 ( .A(p_input[566]), .B(n8860), .Z(n8862) );
  XNOR U8679 ( .A(n8863), .B(n8864), .Z(n8860) );
  AND U8680 ( .A(n254), .B(n8859), .Z(n8864) );
  XNOR U8681 ( .A(n8863), .B(n8857), .Z(n8859) );
  XOR U8682 ( .A(n8865), .B(n8866), .Z(n8857) );
  AND U8683 ( .A(n269), .B(n8867), .Z(n8866) );
  XNOR U8684 ( .A(n8868), .B(n8869), .Z(n8863) );
  AND U8685 ( .A(n261), .B(n8870), .Z(n8869) );
  XOR U8686 ( .A(p_input[598]), .B(n8868), .Z(n8870) );
  XNOR U8687 ( .A(n8871), .B(n8872), .Z(n8868) );
  AND U8688 ( .A(n265), .B(n8867), .Z(n8872) );
  XNOR U8689 ( .A(n8871), .B(n8865), .Z(n8867) );
  XOR U8690 ( .A(n8873), .B(n8874), .Z(n8865) );
  AND U8691 ( .A(n280), .B(n8875), .Z(n8874) );
  XNOR U8692 ( .A(n8876), .B(n8877), .Z(n8871) );
  AND U8693 ( .A(n272), .B(n8878), .Z(n8877) );
  XOR U8694 ( .A(p_input[630]), .B(n8876), .Z(n8878) );
  XNOR U8695 ( .A(n8879), .B(n8880), .Z(n8876) );
  AND U8696 ( .A(n276), .B(n8875), .Z(n8880) );
  XNOR U8697 ( .A(n8879), .B(n8873), .Z(n8875) );
  XOR U8698 ( .A(n8881), .B(n8882), .Z(n8873) );
  AND U8699 ( .A(n291), .B(n8883), .Z(n8882) );
  XNOR U8700 ( .A(n8884), .B(n8885), .Z(n8879) );
  AND U8701 ( .A(n283), .B(n8886), .Z(n8885) );
  XOR U8702 ( .A(p_input[662]), .B(n8884), .Z(n8886) );
  XNOR U8703 ( .A(n8887), .B(n8888), .Z(n8884) );
  AND U8704 ( .A(n287), .B(n8883), .Z(n8888) );
  XNOR U8705 ( .A(n8887), .B(n8881), .Z(n8883) );
  XOR U8706 ( .A(n8889), .B(n8890), .Z(n8881) );
  AND U8707 ( .A(n302), .B(n8891), .Z(n8890) );
  XNOR U8708 ( .A(n8892), .B(n8893), .Z(n8887) );
  AND U8709 ( .A(n294), .B(n8894), .Z(n8893) );
  XOR U8710 ( .A(p_input[694]), .B(n8892), .Z(n8894) );
  XNOR U8711 ( .A(n8895), .B(n8896), .Z(n8892) );
  AND U8712 ( .A(n298), .B(n8891), .Z(n8896) );
  XNOR U8713 ( .A(n8895), .B(n8889), .Z(n8891) );
  XOR U8714 ( .A(n8897), .B(n8898), .Z(n8889) );
  AND U8715 ( .A(n313), .B(n8899), .Z(n8898) );
  XNOR U8716 ( .A(n8900), .B(n8901), .Z(n8895) );
  AND U8717 ( .A(n305), .B(n8902), .Z(n8901) );
  XOR U8718 ( .A(p_input[726]), .B(n8900), .Z(n8902) );
  XNOR U8719 ( .A(n8903), .B(n8904), .Z(n8900) );
  AND U8720 ( .A(n309), .B(n8899), .Z(n8904) );
  XNOR U8721 ( .A(n8903), .B(n8897), .Z(n8899) );
  XOR U8722 ( .A(n8905), .B(n8906), .Z(n8897) );
  AND U8723 ( .A(n324), .B(n8907), .Z(n8906) );
  XNOR U8724 ( .A(n8908), .B(n8909), .Z(n8903) );
  AND U8725 ( .A(n316), .B(n8910), .Z(n8909) );
  XOR U8726 ( .A(p_input[758]), .B(n8908), .Z(n8910) );
  XNOR U8727 ( .A(n8911), .B(n8912), .Z(n8908) );
  AND U8728 ( .A(n320), .B(n8907), .Z(n8912) );
  XNOR U8729 ( .A(n8911), .B(n8905), .Z(n8907) );
  XOR U8730 ( .A(n8913), .B(n8914), .Z(n8905) );
  AND U8731 ( .A(n335), .B(n8915), .Z(n8914) );
  XNOR U8732 ( .A(n8916), .B(n8917), .Z(n8911) );
  AND U8733 ( .A(n327), .B(n8918), .Z(n8917) );
  XOR U8734 ( .A(p_input[790]), .B(n8916), .Z(n8918) );
  XNOR U8735 ( .A(n8919), .B(n8920), .Z(n8916) );
  AND U8736 ( .A(n331), .B(n8915), .Z(n8920) );
  XNOR U8737 ( .A(n8919), .B(n8913), .Z(n8915) );
  XOR U8738 ( .A(n8921), .B(n8922), .Z(n8913) );
  AND U8739 ( .A(n346), .B(n8923), .Z(n8922) );
  XNOR U8740 ( .A(n8924), .B(n8925), .Z(n8919) );
  AND U8741 ( .A(n338), .B(n8926), .Z(n8925) );
  XOR U8742 ( .A(p_input[822]), .B(n8924), .Z(n8926) );
  XNOR U8743 ( .A(n8927), .B(n8928), .Z(n8924) );
  AND U8744 ( .A(n342), .B(n8923), .Z(n8928) );
  XNOR U8745 ( .A(n8927), .B(n8921), .Z(n8923) );
  XOR U8746 ( .A(n8929), .B(n8930), .Z(n8921) );
  AND U8747 ( .A(n357), .B(n8931), .Z(n8930) );
  XNOR U8748 ( .A(n8932), .B(n8933), .Z(n8927) );
  AND U8749 ( .A(n349), .B(n8934), .Z(n8933) );
  XOR U8750 ( .A(p_input[854]), .B(n8932), .Z(n8934) );
  XNOR U8751 ( .A(n8935), .B(n8936), .Z(n8932) );
  AND U8752 ( .A(n353), .B(n8931), .Z(n8936) );
  XNOR U8753 ( .A(n8935), .B(n8929), .Z(n8931) );
  XOR U8754 ( .A(n8937), .B(n8938), .Z(n8929) );
  AND U8755 ( .A(n368), .B(n8939), .Z(n8938) );
  XNOR U8756 ( .A(n8940), .B(n8941), .Z(n8935) );
  AND U8757 ( .A(n360), .B(n8942), .Z(n8941) );
  XOR U8758 ( .A(p_input[886]), .B(n8940), .Z(n8942) );
  XNOR U8759 ( .A(n8943), .B(n8944), .Z(n8940) );
  AND U8760 ( .A(n364), .B(n8939), .Z(n8944) );
  XNOR U8761 ( .A(n8943), .B(n8937), .Z(n8939) );
  XOR U8762 ( .A(n8945), .B(n8946), .Z(n8937) );
  AND U8763 ( .A(n379), .B(n8947), .Z(n8946) );
  XNOR U8764 ( .A(n8948), .B(n8949), .Z(n8943) );
  AND U8765 ( .A(n371), .B(n8950), .Z(n8949) );
  XOR U8766 ( .A(p_input[918]), .B(n8948), .Z(n8950) );
  XNOR U8767 ( .A(n8951), .B(n8952), .Z(n8948) );
  AND U8768 ( .A(n375), .B(n8947), .Z(n8952) );
  XNOR U8769 ( .A(n8951), .B(n8945), .Z(n8947) );
  XOR U8770 ( .A(n8953), .B(n8954), .Z(n8945) );
  AND U8771 ( .A(n390), .B(n8955), .Z(n8954) );
  XNOR U8772 ( .A(n8956), .B(n8957), .Z(n8951) );
  AND U8773 ( .A(n382), .B(n8958), .Z(n8957) );
  XOR U8774 ( .A(p_input[950]), .B(n8956), .Z(n8958) );
  XNOR U8775 ( .A(n8959), .B(n8960), .Z(n8956) );
  AND U8776 ( .A(n386), .B(n8955), .Z(n8960) );
  XNOR U8777 ( .A(n8959), .B(n8953), .Z(n8955) );
  XOR U8778 ( .A(n8961), .B(n8962), .Z(n8953) );
  AND U8779 ( .A(n401), .B(n8963), .Z(n8962) );
  XNOR U8780 ( .A(n8964), .B(n8965), .Z(n8959) );
  AND U8781 ( .A(n393), .B(n8966), .Z(n8965) );
  XOR U8782 ( .A(p_input[982]), .B(n8964), .Z(n8966) );
  XNOR U8783 ( .A(n8967), .B(n8968), .Z(n8964) );
  AND U8784 ( .A(n397), .B(n8963), .Z(n8968) );
  XNOR U8785 ( .A(n8967), .B(n8961), .Z(n8963) );
  XOR U8786 ( .A(n8969), .B(n8970), .Z(n8961) );
  AND U8787 ( .A(n412), .B(n8971), .Z(n8970) );
  XNOR U8788 ( .A(n8972), .B(n8973), .Z(n8967) );
  AND U8789 ( .A(n404), .B(n8974), .Z(n8973) );
  XOR U8790 ( .A(p_input[1014]), .B(n8972), .Z(n8974) );
  XNOR U8791 ( .A(n8975), .B(n8976), .Z(n8972) );
  AND U8792 ( .A(n408), .B(n8971), .Z(n8976) );
  XNOR U8793 ( .A(n8975), .B(n8969), .Z(n8971) );
  XOR U8794 ( .A(n8977), .B(n8978), .Z(n8969) );
  AND U8795 ( .A(n423), .B(n8979), .Z(n8978) );
  XNOR U8796 ( .A(n8980), .B(n8981), .Z(n8975) );
  AND U8797 ( .A(n415), .B(n8982), .Z(n8981) );
  XOR U8798 ( .A(p_input[1046]), .B(n8980), .Z(n8982) );
  XNOR U8799 ( .A(n8983), .B(n8984), .Z(n8980) );
  AND U8800 ( .A(n419), .B(n8979), .Z(n8984) );
  XNOR U8801 ( .A(n8983), .B(n8977), .Z(n8979) );
  XOR U8802 ( .A(n8985), .B(n8986), .Z(n8977) );
  AND U8803 ( .A(n434), .B(n8987), .Z(n8986) );
  XNOR U8804 ( .A(n8988), .B(n8989), .Z(n8983) );
  AND U8805 ( .A(n426), .B(n8990), .Z(n8989) );
  XOR U8806 ( .A(p_input[1078]), .B(n8988), .Z(n8990) );
  XNOR U8807 ( .A(n8991), .B(n8992), .Z(n8988) );
  AND U8808 ( .A(n430), .B(n8987), .Z(n8992) );
  XNOR U8809 ( .A(n8991), .B(n8985), .Z(n8987) );
  XOR U8810 ( .A(n8993), .B(n8994), .Z(n8985) );
  AND U8811 ( .A(n445), .B(n8995), .Z(n8994) );
  XNOR U8812 ( .A(n8996), .B(n8997), .Z(n8991) );
  AND U8813 ( .A(n437), .B(n8998), .Z(n8997) );
  XOR U8814 ( .A(p_input[1110]), .B(n8996), .Z(n8998) );
  XNOR U8815 ( .A(n8999), .B(n9000), .Z(n8996) );
  AND U8816 ( .A(n441), .B(n8995), .Z(n9000) );
  XNOR U8817 ( .A(n8999), .B(n8993), .Z(n8995) );
  XOR U8818 ( .A(n9001), .B(n9002), .Z(n8993) );
  AND U8819 ( .A(n456), .B(n9003), .Z(n9002) );
  XNOR U8820 ( .A(n9004), .B(n9005), .Z(n8999) );
  AND U8821 ( .A(n448), .B(n9006), .Z(n9005) );
  XOR U8822 ( .A(p_input[1142]), .B(n9004), .Z(n9006) );
  XNOR U8823 ( .A(n9007), .B(n9008), .Z(n9004) );
  AND U8824 ( .A(n452), .B(n9003), .Z(n9008) );
  XNOR U8825 ( .A(n9007), .B(n9001), .Z(n9003) );
  XOR U8826 ( .A(n9009), .B(n9010), .Z(n9001) );
  AND U8827 ( .A(n467), .B(n9011), .Z(n9010) );
  XNOR U8828 ( .A(n9012), .B(n9013), .Z(n9007) );
  AND U8829 ( .A(n459), .B(n9014), .Z(n9013) );
  XOR U8830 ( .A(p_input[1174]), .B(n9012), .Z(n9014) );
  XNOR U8831 ( .A(n9015), .B(n9016), .Z(n9012) );
  AND U8832 ( .A(n463), .B(n9011), .Z(n9016) );
  XNOR U8833 ( .A(n9015), .B(n9009), .Z(n9011) );
  XOR U8834 ( .A(n9017), .B(n9018), .Z(n9009) );
  AND U8835 ( .A(n478), .B(n9019), .Z(n9018) );
  XNOR U8836 ( .A(n9020), .B(n9021), .Z(n9015) );
  AND U8837 ( .A(n470), .B(n9022), .Z(n9021) );
  XOR U8838 ( .A(p_input[1206]), .B(n9020), .Z(n9022) );
  XNOR U8839 ( .A(n9023), .B(n9024), .Z(n9020) );
  AND U8840 ( .A(n474), .B(n9019), .Z(n9024) );
  XNOR U8841 ( .A(n9023), .B(n9017), .Z(n9019) );
  XOR U8842 ( .A(n9025), .B(n9026), .Z(n9017) );
  AND U8843 ( .A(n489), .B(n9027), .Z(n9026) );
  XNOR U8844 ( .A(n9028), .B(n9029), .Z(n9023) );
  AND U8845 ( .A(n481), .B(n9030), .Z(n9029) );
  XOR U8846 ( .A(p_input[1238]), .B(n9028), .Z(n9030) );
  XNOR U8847 ( .A(n9031), .B(n9032), .Z(n9028) );
  AND U8848 ( .A(n485), .B(n9027), .Z(n9032) );
  XNOR U8849 ( .A(n9031), .B(n9025), .Z(n9027) );
  XOR U8850 ( .A(n9033), .B(n9034), .Z(n9025) );
  AND U8851 ( .A(n500), .B(n9035), .Z(n9034) );
  XNOR U8852 ( .A(n9036), .B(n9037), .Z(n9031) );
  AND U8853 ( .A(n492), .B(n9038), .Z(n9037) );
  XOR U8854 ( .A(p_input[1270]), .B(n9036), .Z(n9038) );
  XNOR U8855 ( .A(n9039), .B(n9040), .Z(n9036) );
  AND U8856 ( .A(n496), .B(n9035), .Z(n9040) );
  XNOR U8857 ( .A(n9039), .B(n9033), .Z(n9035) );
  XOR U8858 ( .A(n9041), .B(n9042), .Z(n9033) );
  AND U8859 ( .A(n511), .B(n9043), .Z(n9042) );
  XNOR U8860 ( .A(n9044), .B(n9045), .Z(n9039) );
  AND U8861 ( .A(n503), .B(n9046), .Z(n9045) );
  XOR U8862 ( .A(p_input[1302]), .B(n9044), .Z(n9046) );
  XNOR U8863 ( .A(n9047), .B(n9048), .Z(n9044) );
  AND U8864 ( .A(n507), .B(n9043), .Z(n9048) );
  XNOR U8865 ( .A(n9047), .B(n9041), .Z(n9043) );
  XOR U8866 ( .A(n9049), .B(n9050), .Z(n9041) );
  AND U8867 ( .A(n522), .B(n9051), .Z(n9050) );
  XNOR U8868 ( .A(n9052), .B(n9053), .Z(n9047) );
  AND U8869 ( .A(n514), .B(n9054), .Z(n9053) );
  XOR U8870 ( .A(p_input[1334]), .B(n9052), .Z(n9054) );
  XNOR U8871 ( .A(n9055), .B(n9056), .Z(n9052) );
  AND U8872 ( .A(n518), .B(n9051), .Z(n9056) );
  XNOR U8873 ( .A(n9055), .B(n9049), .Z(n9051) );
  XOR U8874 ( .A(n9057), .B(n9058), .Z(n9049) );
  AND U8875 ( .A(n533), .B(n9059), .Z(n9058) );
  XNOR U8876 ( .A(n9060), .B(n9061), .Z(n9055) );
  AND U8877 ( .A(n525), .B(n9062), .Z(n9061) );
  XOR U8878 ( .A(p_input[1366]), .B(n9060), .Z(n9062) );
  XNOR U8879 ( .A(n9063), .B(n9064), .Z(n9060) );
  AND U8880 ( .A(n529), .B(n9059), .Z(n9064) );
  XNOR U8881 ( .A(n9063), .B(n9057), .Z(n9059) );
  XOR U8882 ( .A(n9065), .B(n9066), .Z(n9057) );
  AND U8883 ( .A(n544), .B(n9067), .Z(n9066) );
  XNOR U8884 ( .A(n9068), .B(n9069), .Z(n9063) );
  AND U8885 ( .A(n536), .B(n9070), .Z(n9069) );
  XOR U8886 ( .A(p_input[1398]), .B(n9068), .Z(n9070) );
  XNOR U8887 ( .A(n9071), .B(n9072), .Z(n9068) );
  AND U8888 ( .A(n540), .B(n9067), .Z(n9072) );
  XNOR U8889 ( .A(n9071), .B(n9065), .Z(n9067) );
  XOR U8890 ( .A(n9073), .B(n9074), .Z(n9065) );
  AND U8891 ( .A(n555), .B(n9075), .Z(n9074) );
  XNOR U8892 ( .A(n9076), .B(n9077), .Z(n9071) );
  AND U8893 ( .A(n547), .B(n9078), .Z(n9077) );
  XOR U8894 ( .A(p_input[1430]), .B(n9076), .Z(n9078) );
  XNOR U8895 ( .A(n9079), .B(n9080), .Z(n9076) );
  AND U8896 ( .A(n551), .B(n9075), .Z(n9080) );
  XNOR U8897 ( .A(n9079), .B(n9073), .Z(n9075) );
  XOR U8898 ( .A(n9081), .B(n9082), .Z(n9073) );
  AND U8899 ( .A(n566), .B(n9083), .Z(n9082) );
  XNOR U8900 ( .A(n9084), .B(n9085), .Z(n9079) );
  AND U8901 ( .A(n558), .B(n9086), .Z(n9085) );
  XOR U8902 ( .A(p_input[1462]), .B(n9084), .Z(n9086) );
  XNOR U8903 ( .A(n9087), .B(n9088), .Z(n9084) );
  AND U8904 ( .A(n562), .B(n9083), .Z(n9088) );
  XNOR U8905 ( .A(n9087), .B(n9081), .Z(n9083) );
  XOR U8906 ( .A(n9089), .B(n9090), .Z(n9081) );
  AND U8907 ( .A(n577), .B(n9091), .Z(n9090) );
  XNOR U8908 ( .A(n9092), .B(n9093), .Z(n9087) );
  AND U8909 ( .A(n569), .B(n9094), .Z(n9093) );
  XOR U8910 ( .A(p_input[1494]), .B(n9092), .Z(n9094) );
  XNOR U8911 ( .A(n9095), .B(n9096), .Z(n9092) );
  AND U8912 ( .A(n573), .B(n9091), .Z(n9096) );
  XNOR U8913 ( .A(n9095), .B(n9089), .Z(n9091) );
  XOR U8914 ( .A(n9097), .B(n9098), .Z(n9089) );
  AND U8915 ( .A(n588), .B(n9099), .Z(n9098) );
  XNOR U8916 ( .A(n9100), .B(n9101), .Z(n9095) );
  AND U8917 ( .A(n580), .B(n9102), .Z(n9101) );
  XOR U8918 ( .A(p_input[1526]), .B(n9100), .Z(n9102) );
  XNOR U8919 ( .A(n9103), .B(n9104), .Z(n9100) );
  AND U8920 ( .A(n584), .B(n9099), .Z(n9104) );
  XNOR U8921 ( .A(n9103), .B(n9097), .Z(n9099) );
  XOR U8922 ( .A(n9105), .B(n9106), .Z(n9097) );
  AND U8923 ( .A(n599), .B(n9107), .Z(n9106) );
  XNOR U8924 ( .A(n9108), .B(n9109), .Z(n9103) );
  AND U8925 ( .A(n591), .B(n9110), .Z(n9109) );
  XOR U8926 ( .A(p_input[1558]), .B(n9108), .Z(n9110) );
  XNOR U8927 ( .A(n9111), .B(n9112), .Z(n9108) );
  AND U8928 ( .A(n595), .B(n9107), .Z(n9112) );
  XNOR U8929 ( .A(n9111), .B(n9105), .Z(n9107) );
  XOR U8930 ( .A(n9113), .B(n9114), .Z(n9105) );
  AND U8931 ( .A(n610), .B(n9115), .Z(n9114) );
  XNOR U8932 ( .A(n9116), .B(n9117), .Z(n9111) );
  AND U8933 ( .A(n602), .B(n9118), .Z(n9117) );
  XOR U8934 ( .A(p_input[1590]), .B(n9116), .Z(n9118) );
  XNOR U8935 ( .A(n9119), .B(n9120), .Z(n9116) );
  AND U8936 ( .A(n606), .B(n9115), .Z(n9120) );
  XNOR U8937 ( .A(n9119), .B(n9113), .Z(n9115) );
  XOR U8938 ( .A(n9121), .B(n9122), .Z(n9113) );
  AND U8939 ( .A(n621), .B(n9123), .Z(n9122) );
  XNOR U8940 ( .A(n9124), .B(n9125), .Z(n9119) );
  AND U8941 ( .A(n613), .B(n9126), .Z(n9125) );
  XOR U8942 ( .A(p_input[1622]), .B(n9124), .Z(n9126) );
  XNOR U8943 ( .A(n9127), .B(n9128), .Z(n9124) );
  AND U8944 ( .A(n617), .B(n9123), .Z(n9128) );
  XNOR U8945 ( .A(n9127), .B(n9121), .Z(n9123) );
  XOR U8946 ( .A(n9129), .B(n9130), .Z(n9121) );
  AND U8947 ( .A(n632), .B(n9131), .Z(n9130) );
  XNOR U8948 ( .A(n9132), .B(n9133), .Z(n9127) );
  AND U8949 ( .A(n624), .B(n9134), .Z(n9133) );
  XOR U8950 ( .A(p_input[1654]), .B(n9132), .Z(n9134) );
  XNOR U8951 ( .A(n9135), .B(n9136), .Z(n9132) );
  AND U8952 ( .A(n628), .B(n9131), .Z(n9136) );
  XNOR U8953 ( .A(n9135), .B(n9129), .Z(n9131) );
  XOR U8954 ( .A(n9137), .B(n9138), .Z(n9129) );
  AND U8955 ( .A(n643), .B(n9139), .Z(n9138) );
  XNOR U8956 ( .A(n9140), .B(n9141), .Z(n9135) );
  AND U8957 ( .A(n635), .B(n9142), .Z(n9141) );
  XOR U8958 ( .A(p_input[1686]), .B(n9140), .Z(n9142) );
  XNOR U8959 ( .A(n9143), .B(n9144), .Z(n9140) );
  AND U8960 ( .A(n639), .B(n9139), .Z(n9144) );
  XNOR U8961 ( .A(n9143), .B(n9137), .Z(n9139) );
  XOR U8962 ( .A(n9145), .B(n9146), .Z(n9137) );
  AND U8963 ( .A(n654), .B(n9147), .Z(n9146) );
  XNOR U8964 ( .A(n9148), .B(n9149), .Z(n9143) );
  AND U8965 ( .A(n646), .B(n9150), .Z(n9149) );
  XOR U8966 ( .A(p_input[1718]), .B(n9148), .Z(n9150) );
  XNOR U8967 ( .A(n9151), .B(n9152), .Z(n9148) );
  AND U8968 ( .A(n650), .B(n9147), .Z(n9152) );
  XNOR U8969 ( .A(n9151), .B(n9145), .Z(n9147) );
  XOR U8970 ( .A(n9153), .B(n9154), .Z(n9145) );
  AND U8971 ( .A(n665), .B(n9155), .Z(n9154) );
  XNOR U8972 ( .A(n9156), .B(n9157), .Z(n9151) );
  AND U8973 ( .A(n657), .B(n9158), .Z(n9157) );
  XOR U8974 ( .A(p_input[1750]), .B(n9156), .Z(n9158) );
  XNOR U8975 ( .A(n9159), .B(n9160), .Z(n9156) );
  AND U8976 ( .A(n661), .B(n9155), .Z(n9160) );
  XNOR U8977 ( .A(n9159), .B(n9153), .Z(n9155) );
  XOR U8978 ( .A(n9161), .B(n9162), .Z(n9153) );
  AND U8979 ( .A(n676), .B(n9163), .Z(n9162) );
  XNOR U8980 ( .A(n9164), .B(n9165), .Z(n9159) );
  AND U8981 ( .A(n668), .B(n9166), .Z(n9165) );
  XOR U8982 ( .A(p_input[1782]), .B(n9164), .Z(n9166) );
  XNOR U8983 ( .A(n9167), .B(n9168), .Z(n9164) );
  AND U8984 ( .A(n672), .B(n9163), .Z(n9168) );
  XNOR U8985 ( .A(n9167), .B(n9161), .Z(n9163) );
  XOR U8986 ( .A(n9169), .B(n9170), .Z(n9161) );
  AND U8987 ( .A(n687), .B(n9171), .Z(n9170) );
  XNOR U8988 ( .A(n9172), .B(n9173), .Z(n9167) );
  AND U8989 ( .A(n679), .B(n9174), .Z(n9173) );
  XOR U8990 ( .A(p_input[1814]), .B(n9172), .Z(n9174) );
  XNOR U8991 ( .A(n9175), .B(n9176), .Z(n9172) );
  AND U8992 ( .A(n683), .B(n9171), .Z(n9176) );
  XNOR U8993 ( .A(n9175), .B(n9169), .Z(n9171) );
  XOR U8994 ( .A(n9177), .B(n9178), .Z(n9169) );
  AND U8995 ( .A(n698), .B(n9179), .Z(n9178) );
  XNOR U8996 ( .A(n9180), .B(n9181), .Z(n9175) );
  AND U8997 ( .A(n690), .B(n9182), .Z(n9181) );
  XOR U8998 ( .A(p_input[1846]), .B(n9180), .Z(n9182) );
  XNOR U8999 ( .A(n9183), .B(n9184), .Z(n9180) );
  AND U9000 ( .A(n694), .B(n9179), .Z(n9184) );
  XNOR U9001 ( .A(n9183), .B(n9177), .Z(n9179) );
  XOR U9002 ( .A(n9185), .B(n9186), .Z(n9177) );
  AND U9003 ( .A(n709), .B(n9187), .Z(n9186) );
  XNOR U9004 ( .A(n9188), .B(n9189), .Z(n9183) );
  AND U9005 ( .A(n701), .B(n9190), .Z(n9189) );
  XOR U9006 ( .A(p_input[1878]), .B(n9188), .Z(n9190) );
  XNOR U9007 ( .A(n9191), .B(n9192), .Z(n9188) );
  AND U9008 ( .A(n705), .B(n9187), .Z(n9192) );
  XNOR U9009 ( .A(n9191), .B(n9185), .Z(n9187) );
  XOR U9010 ( .A(n9193), .B(n9194), .Z(n9185) );
  AND U9011 ( .A(n720), .B(n9195), .Z(n9194) );
  XNOR U9012 ( .A(n9196), .B(n9197), .Z(n9191) );
  AND U9013 ( .A(n712), .B(n9198), .Z(n9197) );
  XOR U9014 ( .A(p_input[1910]), .B(n9196), .Z(n9198) );
  XNOR U9015 ( .A(n9199), .B(n9200), .Z(n9196) );
  AND U9016 ( .A(n716), .B(n9195), .Z(n9200) );
  XNOR U9017 ( .A(n9199), .B(n9193), .Z(n9195) );
  XOR U9018 ( .A(n9201), .B(n9202), .Z(n9193) );
  AND U9019 ( .A(n731), .B(n9203), .Z(n9202) );
  XNOR U9020 ( .A(n9204), .B(n9205), .Z(n9199) );
  AND U9021 ( .A(n723), .B(n9206), .Z(n9205) );
  XOR U9022 ( .A(p_input[1942]), .B(n9204), .Z(n9206) );
  XNOR U9023 ( .A(n9207), .B(n9208), .Z(n9204) );
  AND U9024 ( .A(n727), .B(n9203), .Z(n9208) );
  XNOR U9025 ( .A(n9207), .B(n9201), .Z(n9203) );
  XOR U9026 ( .A(\knn_comb_/min_val_out[0][22] ), .B(n9209), .Z(n9201) );
  AND U9027 ( .A(n741), .B(n9210), .Z(n9209) );
  XNOR U9028 ( .A(n9211), .B(n9212), .Z(n9207) );
  AND U9029 ( .A(n734), .B(n9213), .Z(n9212) );
  XOR U9030 ( .A(p_input[1974]), .B(n9211), .Z(n9213) );
  XNOR U9031 ( .A(n9214), .B(n9215), .Z(n9211) );
  AND U9032 ( .A(n738), .B(n9210), .Z(n9215) );
  XOR U9033 ( .A(\knn_comb_/min_val_out[0][22] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .Z(n9210) );
  XOR U9034 ( .A(n31), .B(n9216), .Z(o[21]) );
  AND U9035 ( .A(n58), .B(n9217), .Z(n31) );
  XOR U9036 ( .A(n32), .B(n9216), .Z(n9217) );
  XOR U9037 ( .A(n9218), .B(n9219), .Z(n9216) );
  AND U9038 ( .A(n70), .B(n9220), .Z(n9219) );
  XOR U9039 ( .A(n9221), .B(n9222), .Z(n32) );
  AND U9040 ( .A(n62), .B(n9223), .Z(n9222) );
  XOR U9041 ( .A(p_input[21]), .B(n9221), .Z(n9223) );
  XNOR U9042 ( .A(n9224), .B(n9225), .Z(n9221) );
  AND U9043 ( .A(n66), .B(n9220), .Z(n9225) );
  XNOR U9044 ( .A(n9224), .B(n9218), .Z(n9220) );
  XOR U9045 ( .A(n9226), .B(n9227), .Z(n9218) );
  AND U9046 ( .A(n82), .B(n9228), .Z(n9227) );
  XNOR U9047 ( .A(n9229), .B(n9230), .Z(n9224) );
  AND U9048 ( .A(n74), .B(n9231), .Z(n9230) );
  XOR U9049 ( .A(p_input[53]), .B(n9229), .Z(n9231) );
  XNOR U9050 ( .A(n9232), .B(n9233), .Z(n9229) );
  AND U9051 ( .A(n78), .B(n9228), .Z(n9233) );
  XNOR U9052 ( .A(n9232), .B(n9226), .Z(n9228) );
  XOR U9053 ( .A(n9234), .B(n9235), .Z(n9226) );
  AND U9054 ( .A(n93), .B(n9236), .Z(n9235) );
  XNOR U9055 ( .A(n9237), .B(n9238), .Z(n9232) );
  AND U9056 ( .A(n85), .B(n9239), .Z(n9238) );
  XOR U9057 ( .A(p_input[85]), .B(n9237), .Z(n9239) );
  XNOR U9058 ( .A(n9240), .B(n9241), .Z(n9237) );
  AND U9059 ( .A(n89), .B(n9236), .Z(n9241) );
  XNOR U9060 ( .A(n9240), .B(n9234), .Z(n9236) );
  XOR U9061 ( .A(n9242), .B(n9243), .Z(n9234) );
  AND U9062 ( .A(n104), .B(n9244), .Z(n9243) );
  XNOR U9063 ( .A(n9245), .B(n9246), .Z(n9240) );
  AND U9064 ( .A(n96), .B(n9247), .Z(n9246) );
  XOR U9065 ( .A(p_input[117]), .B(n9245), .Z(n9247) );
  XNOR U9066 ( .A(n9248), .B(n9249), .Z(n9245) );
  AND U9067 ( .A(n100), .B(n9244), .Z(n9249) );
  XNOR U9068 ( .A(n9248), .B(n9242), .Z(n9244) );
  XOR U9069 ( .A(n9250), .B(n9251), .Z(n9242) );
  AND U9070 ( .A(n115), .B(n9252), .Z(n9251) );
  XNOR U9071 ( .A(n9253), .B(n9254), .Z(n9248) );
  AND U9072 ( .A(n107), .B(n9255), .Z(n9254) );
  XOR U9073 ( .A(p_input[149]), .B(n9253), .Z(n9255) );
  XNOR U9074 ( .A(n9256), .B(n9257), .Z(n9253) );
  AND U9075 ( .A(n111), .B(n9252), .Z(n9257) );
  XNOR U9076 ( .A(n9256), .B(n9250), .Z(n9252) );
  XOR U9077 ( .A(n9258), .B(n9259), .Z(n9250) );
  AND U9078 ( .A(n126), .B(n9260), .Z(n9259) );
  XNOR U9079 ( .A(n9261), .B(n9262), .Z(n9256) );
  AND U9080 ( .A(n118), .B(n9263), .Z(n9262) );
  XOR U9081 ( .A(p_input[181]), .B(n9261), .Z(n9263) );
  XNOR U9082 ( .A(n9264), .B(n9265), .Z(n9261) );
  AND U9083 ( .A(n122), .B(n9260), .Z(n9265) );
  XNOR U9084 ( .A(n9264), .B(n9258), .Z(n9260) );
  XOR U9085 ( .A(n9266), .B(n9267), .Z(n9258) );
  AND U9086 ( .A(n137), .B(n9268), .Z(n9267) );
  XNOR U9087 ( .A(n9269), .B(n9270), .Z(n9264) );
  AND U9088 ( .A(n129), .B(n9271), .Z(n9270) );
  XOR U9089 ( .A(p_input[213]), .B(n9269), .Z(n9271) );
  XNOR U9090 ( .A(n9272), .B(n9273), .Z(n9269) );
  AND U9091 ( .A(n133), .B(n9268), .Z(n9273) );
  XNOR U9092 ( .A(n9272), .B(n9266), .Z(n9268) );
  XOR U9093 ( .A(n9274), .B(n9275), .Z(n9266) );
  AND U9094 ( .A(n148), .B(n9276), .Z(n9275) );
  XNOR U9095 ( .A(n9277), .B(n9278), .Z(n9272) );
  AND U9096 ( .A(n140), .B(n9279), .Z(n9278) );
  XOR U9097 ( .A(p_input[245]), .B(n9277), .Z(n9279) );
  XNOR U9098 ( .A(n9280), .B(n9281), .Z(n9277) );
  AND U9099 ( .A(n144), .B(n9276), .Z(n9281) );
  XNOR U9100 ( .A(n9280), .B(n9274), .Z(n9276) );
  XOR U9101 ( .A(n9282), .B(n9283), .Z(n9274) );
  AND U9102 ( .A(n159), .B(n9284), .Z(n9283) );
  XNOR U9103 ( .A(n9285), .B(n9286), .Z(n9280) );
  AND U9104 ( .A(n151), .B(n9287), .Z(n9286) );
  XOR U9105 ( .A(p_input[277]), .B(n9285), .Z(n9287) );
  XNOR U9106 ( .A(n9288), .B(n9289), .Z(n9285) );
  AND U9107 ( .A(n155), .B(n9284), .Z(n9289) );
  XNOR U9108 ( .A(n9288), .B(n9282), .Z(n9284) );
  XOR U9109 ( .A(n9290), .B(n9291), .Z(n9282) );
  AND U9110 ( .A(n170), .B(n9292), .Z(n9291) );
  XNOR U9111 ( .A(n9293), .B(n9294), .Z(n9288) );
  AND U9112 ( .A(n162), .B(n9295), .Z(n9294) );
  XOR U9113 ( .A(p_input[309]), .B(n9293), .Z(n9295) );
  XNOR U9114 ( .A(n9296), .B(n9297), .Z(n9293) );
  AND U9115 ( .A(n166), .B(n9292), .Z(n9297) );
  XNOR U9116 ( .A(n9296), .B(n9290), .Z(n9292) );
  XOR U9117 ( .A(n9298), .B(n9299), .Z(n9290) );
  AND U9118 ( .A(n181), .B(n9300), .Z(n9299) );
  XNOR U9119 ( .A(n9301), .B(n9302), .Z(n9296) );
  AND U9120 ( .A(n173), .B(n9303), .Z(n9302) );
  XOR U9121 ( .A(p_input[341]), .B(n9301), .Z(n9303) );
  XNOR U9122 ( .A(n9304), .B(n9305), .Z(n9301) );
  AND U9123 ( .A(n177), .B(n9300), .Z(n9305) );
  XNOR U9124 ( .A(n9304), .B(n9298), .Z(n9300) );
  XOR U9125 ( .A(n9306), .B(n9307), .Z(n9298) );
  AND U9126 ( .A(n192), .B(n9308), .Z(n9307) );
  XNOR U9127 ( .A(n9309), .B(n9310), .Z(n9304) );
  AND U9128 ( .A(n184), .B(n9311), .Z(n9310) );
  XOR U9129 ( .A(p_input[373]), .B(n9309), .Z(n9311) );
  XNOR U9130 ( .A(n9312), .B(n9313), .Z(n9309) );
  AND U9131 ( .A(n188), .B(n9308), .Z(n9313) );
  XNOR U9132 ( .A(n9312), .B(n9306), .Z(n9308) );
  XOR U9133 ( .A(n9314), .B(n9315), .Z(n9306) );
  AND U9134 ( .A(n203), .B(n9316), .Z(n9315) );
  XNOR U9135 ( .A(n9317), .B(n9318), .Z(n9312) );
  AND U9136 ( .A(n195), .B(n9319), .Z(n9318) );
  XOR U9137 ( .A(p_input[405]), .B(n9317), .Z(n9319) );
  XNOR U9138 ( .A(n9320), .B(n9321), .Z(n9317) );
  AND U9139 ( .A(n199), .B(n9316), .Z(n9321) );
  XNOR U9140 ( .A(n9320), .B(n9314), .Z(n9316) );
  XOR U9141 ( .A(n9322), .B(n9323), .Z(n9314) );
  AND U9142 ( .A(n214), .B(n9324), .Z(n9323) );
  XNOR U9143 ( .A(n9325), .B(n9326), .Z(n9320) );
  AND U9144 ( .A(n206), .B(n9327), .Z(n9326) );
  XOR U9145 ( .A(p_input[437]), .B(n9325), .Z(n9327) );
  XNOR U9146 ( .A(n9328), .B(n9329), .Z(n9325) );
  AND U9147 ( .A(n210), .B(n9324), .Z(n9329) );
  XNOR U9148 ( .A(n9328), .B(n9322), .Z(n9324) );
  XOR U9149 ( .A(n9330), .B(n9331), .Z(n9322) );
  AND U9150 ( .A(n225), .B(n9332), .Z(n9331) );
  XNOR U9151 ( .A(n9333), .B(n9334), .Z(n9328) );
  AND U9152 ( .A(n217), .B(n9335), .Z(n9334) );
  XOR U9153 ( .A(p_input[469]), .B(n9333), .Z(n9335) );
  XNOR U9154 ( .A(n9336), .B(n9337), .Z(n9333) );
  AND U9155 ( .A(n221), .B(n9332), .Z(n9337) );
  XNOR U9156 ( .A(n9336), .B(n9330), .Z(n9332) );
  XOR U9157 ( .A(n9338), .B(n9339), .Z(n9330) );
  AND U9158 ( .A(n236), .B(n9340), .Z(n9339) );
  XNOR U9159 ( .A(n9341), .B(n9342), .Z(n9336) );
  AND U9160 ( .A(n228), .B(n9343), .Z(n9342) );
  XOR U9161 ( .A(p_input[501]), .B(n9341), .Z(n9343) );
  XNOR U9162 ( .A(n9344), .B(n9345), .Z(n9341) );
  AND U9163 ( .A(n232), .B(n9340), .Z(n9345) );
  XNOR U9164 ( .A(n9344), .B(n9338), .Z(n9340) );
  XOR U9165 ( .A(n9346), .B(n9347), .Z(n9338) );
  AND U9166 ( .A(n247), .B(n9348), .Z(n9347) );
  XNOR U9167 ( .A(n9349), .B(n9350), .Z(n9344) );
  AND U9168 ( .A(n239), .B(n9351), .Z(n9350) );
  XOR U9169 ( .A(p_input[533]), .B(n9349), .Z(n9351) );
  XNOR U9170 ( .A(n9352), .B(n9353), .Z(n9349) );
  AND U9171 ( .A(n243), .B(n9348), .Z(n9353) );
  XNOR U9172 ( .A(n9352), .B(n9346), .Z(n9348) );
  XOR U9173 ( .A(n9354), .B(n9355), .Z(n9346) );
  AND U9174 ( .A(n258), .B(n9356), .Z(n9355) );
  XNOR U9175 ( .A(n9357), .B(n9358), .Z(n9352) );
  AND U9176 ( .A(n250), .B(n9359), .Z(n9358) );
  XOR U9177 ( .A(p_input[565]), .B(n9357), .Z(n9359) );
  XNOR U9178 ( .A(n9360), .B(n9361), .Z(n9357) );
  AND U9179 ( .A(n254), .B(n9356), .Z(n9361) );
  XNOR U9180 ( .A(n9360), .B(n9354), .Z(n9356) );
  XOR U9181 ( .A(n9362), .B(n9363), .Z(n9354) );
  AND U9182 ( .A(n269), .B(n9364), .Z(n9363) );
  XNOR U9183 ( .A(n9365), .B(n9366), .Z(n9360) );
  AND U9184 ( .A(n261), .B(n9367), .Z(n9366) );
  XOR U9185 ( .A(p_input[597]), .B(n9365), .Z(n9367) );
  XNOR U9186 ( .A(n9368), .B(n9369), .Z(n9365) );
  AND U9187 ( .A(n265), .B(n9364), .Z(n9369) );
  XNOR U9188 ( .A(n9368), .B(n9362), .Z(n9364) );
  XOR U9189 ( .A(n9370), .B(n9371), .Z(n9362) );
  AND U9190 ( .A(n280), .B(n9372), .Z(n9371) );
  XNOR U9191 ( .A(n9373), .B(n9374), .Z(n9368) );
  AND U9192 ( .A(n272), .B(n9375), .Z(n9374) );
  XOR U9193 ( .A(p_input[629]), .B(n9373), .Z(n9375) );
  XNOR U9194 ( .A(n9376), .B(n9377), .Z(n9373) );
  AND U9195 ( .A(n276), .B(n9372), .Z(n9377) );
  XNOR U9196 ( .A(n9376), .B(n9370), .Z(n9372) );
  XOR U9197 ( .A(n9378), .B(n9379), .Z(n9370) );
  AND U9198 ( .A(n291), .B(n9380), .Z(n9379) );
  XNOR U9199 ( .A(n9381), .B(n9382), .Z(n9376) );
  AND U9200 ( .A(n283), .B(n9383), .Z(n9382) );
  XOR U9201 ( .A(p_input[661]), .B(n9381), .Z(n9383) );
  XNOR U9202 ( .A(n9384), .B(n9385), .Z(n9381) );
  AND U9203 ( .A(n287), .B(n9380), .Z(n9385) );
  XNOR U9204 ( .A(n9384), .B(n9378), .Z(n9380) );
  XOR U9205 ( .A(n9386), .B(n9387), .Z(n9378) );
  AND U9206 ( .A(n302), .B(n9388), .Z(n9387) );
  XNOR U9207 ( .A(n9389), .B(n9390), .Z(n9384) );
  AND U9208 ( .A(n294), .B(n9391), .Z(n9390) );
  XOR U9209 ( .A(p_input[693]), .B(n9389), .Z(n9391) );
  XNOR U9210 ( .A(n9392), .B(n9393), .Z(n9389) );
  AND U9211 ( .A(n298), .B(n9388), .Z(n9393) );
  XNOR U9212 ( .A(n9392), .B(n9386), .Z(n9388) );
  XOR U9213 ( .A(n9394), .B(n9395), .Z(n9386) );
  AND U9214 ( .A(n313), .B(n9396), .Z(n9395) );
  XNOR U9215 ( .A(n9397), .B(n9398), .Z(n9392) );
  AND U9216 ( .A(n305), .B(n9399), .Z(n9398) );
  XOR U9217 ( .A(p_input[725]), .B(n9397), .Z(n9399) );
  XNOR U9218 ( .A(n9400), .B(n9401), .Z(n9397) );
  AND U9219 ( .A(n309), .B(n9396), .Z(n9401) );
  XNOR U9220 ( .A(n9400), .B(n9394), .Z(n9396) );
  XOR U9221 ( .A(n9402), .B(n9403), .Z(n9394) );
  AND U9222 ( .A(n324), .B(n9404), .Z(n9403) );
  XNOR U9223 ( .A(n9405), .B(n9406), .Z(n9400) );
  AND U9224 ( .A(n316), .B(n9407), .Z(n9406) );
  XOR U9225 ( .A(p_input[757]), .B(n9405), .Z(n9407) );
  XNOR U9226 ( .A(n9408), .B(n9409), .Z(n9405) );
  AND U9227 ( .A(n320), .B(n9404), .Z(n9409) );
  XNOR U9228 ( .A(n9408), .B(n9402), .Z(n9404) );
  XOR U9229 ( .A(n9410), .B(n9411), .Z(n9402) );
  AND U9230 ( .A(n335), .B(n9412), .Z(n9411) );
  XNOR U9231 ( .A(n9413), .B(n9414), .Z(n9408) );
  AND U9232 ( .A(n327), .B(n9415), .Z(n9414) );
  XOR U9233 ( .A(p_input[789]), .B(n9413), .Z(n9415) );
  XNOR U9234 ( .A(n9416), .B(n9417), .Z(n9413) );
  AND U9235 ( .A(n331), .B(n9412), .Z(n9417) );
  XNOR U9236 ( .A(n9416), .B(n9410), .Z(n9412) );
  XOR U9237 ( .A(n9418), .B(n9419), .Z(n9410) );
  AND U9238 ( .A(n346), .B(n9420), .Z(n9419) );
  XNOR U9239 ( .A(n9421), .B(n9422), .Z(n9416) );
  AND U9240 ( .A(n338), .B(n9423), .Z(n9422) );
  XOR U9241 ( .A(p_input[821]), .B(n9421), .Z(n9423) );
  XNOR U9242 ( .A(n9424), .B(n9425), .Z(n9421) );
  AND U9243 ( .A(n342), .B(n9420), .Z(n9425) );
  XNOR U9244 ( .A(n9424), .B(n9418), .Z(n9420) );
  XOR U9245 ( .A(n9426), .B(n9427), .Z(n9418) );
  AND U9246 ( .A(n357), .B(n9428), .Z(n9427) );
  XNOR U9247 ( .A(n9429), .B(n9430), .Z(n9424) );
  AND U9248 ( .A(n349), .B(n9431), .Z(n9430) );
  XOR U9249 ( .A(p_input[853]), .B(n9429), .Z(n9431) );
  XNOR U9250 ( .A(n9432), .B(n9433), .Z(n9429) );
  AND U9251 ( .A(n353), .B(n9428), .Z(n9433) );
  XNOR U9252 ( .A(n9432), .B(n9426), .Z(n9428) );
  XOR U9253 ( .A(n9434), .B(n9435), .Z(n9426) );
  AND U9254 ( .A(n368), .B(n9436), .Z(n9435) );
  XNOR U9255 ( .A(n9437), .B(n9438), .Z(n9432) );
  AND U9256 ( .A(n360), .B(n9439), .Z(n9438) );
  XOR U9257 ( .A(p_input[885]), .B(n9437), .Z(n9439) );
  XNOR U9258 ( .A(n9440), .B(n9441), .Z(n9437) );
  AND U9259 ( .A(n364), .B(n9436), .Z(n9441) );
  XNOR U9260 ( .A(n9440), .B(n9434), .Z(n9436) );
  XOR U9261 ( .A(n9442), .B(n9443), .Z(n9434) );
  AND U9262 ( .A(n379), .B(n9444), .Z(n9443) );
  XNOR U9263 ( .A(n9445), .B(n9446), .Z(n9440) );
  AND U9264 ( .A(n371), .B(n9447), .Z(n9446) );
  XOR U9265 ( .A(p_input[917]), .B(n9445), .Z(n9447) );
  XNOR U9266 ( .A(n9448), .B(n9449), .Z(n9445) );
  AND U9267 ( .A(n375), .B(n9444), .Z(n9449) );
  XNOR U9268 ( .A(n9448), .B(n9442), .Z(n9444) );
  XOR U9269 ( .A(n9450), .B(n9451), .Z(n9442) );
  AND U9270 ( .A(n390), .B(n9452), .Z(n9451) );
  XNOR U9271 ( .A(n9453), .B(n9454), .Z(n9448) );
  AND U9272 ( .A(n382), .B(n9455), .Z(n9454) );
  XOR U9273 ( .A(p_input[949]), .B(n9453), .Z(n9455) );
  XNOR U9274 ( .A(n9456), .B(n9457), .Z(n9453) );
  AND U9275 ( .A(n386), .B(n9452), .Z(n9457) );
  XNOR U9276 ( .A(n9456), .B(n9450), .Z(n9452) );
  XOR U9277 ( .A(n9458), .B(n9459), .Z(n9450) );
  AND U9278 ( .A(n401), .B(n9460), .Z(n9459) );
  XNOR U9279 ( .A(n9461), .B(n9462), .Z(n9456) );
  AND U9280 ( .A(n393), .B(n9463), .Z(n9462) );
  XOR U9281 ( .A(p_input[981]), .B(n9461), .Z(n9463) );
  XNOR U9282 ( .A(n9464), .B(n9465), .Z(n9461) );
  AND U9283 ( .A(n397), .B(n9460), .Z(n9465) );
  XNOR U9284 ( .A(n9464), .B(n9458), .Z(n9460) );
  XOR U9285 ( .A(n9466), .B(n9467), .Z(n9458) );
  AND U9286 ( .A(n412), .B(n9468), .Z(n9467) );
  XNOR U9287 ( .A(n9469), .B(n9470), .Z(n9464) );
  AND U9288 ( .A(n404), .B(n9471), .Z(n9470) );
  XOR U9289 ( .A(p_input[1013]), .B(n9469), .Z(n9471) );
  XNOR U9290 ( .A(n9472), .B(n9473), .Z(n9469) );
  AND U9291 ( .A(n408), .B(n9468), .Z(n9473) );
  XNOR U9292 ( .A(n9472), .B(n9466), .Z(n9468) );
  XOR U9293 ( .A(n9474), .B(n9475), .Z(n9466) );
  AND U9294 ( .A(n423), .B(n9476), .Z(n9475) );
  XNOR U9295 ( .A(n9477), .B(n9478), .Z(n9472) );
  AND U9296 ( .A(n415), .B(n9479), .Z(n9478) );
  XOR U9297 ( .A(p_input[1045]), .B(n9477), .Z(n9479) );
  XNOR U9298 ( .A(n9480), .B(n9481), .Z(n9477) );
  AND U9299 ( .A(n419), .B(n9476), .Z(n9481) );
  XNOR U9300 ( .A(n9480), .B(n9474), .Z(n9476) );
  XOR U9301 ( .A(n9482), .B(n9483), .Z(n9474) );
  AND U9302 ( .A(n434), .B(n9484), .Z(n9483) );
  XNOR U9303 ( .A(n9485), .B(n9486), .Z(n9480) );
  AND U9304 ( .A(n426), .B(n9487), .Z(n9486) );
  XOR U9305 ( .A(p_input[1077]), .B(n9485), .Z(n9487) );
  XNOR U9306 ( .A(n9488), .B(n9489), .Z(n9485) );
  AND U9307 ( .A(n430), .B(n9484), .Z(n9489) );
  XNOR U9308 ( .A(n9488), .B(n9482), .Z(n9484) );
  XOR U9309 ( .A(n9490), .B(n9491), .Z(n9482) );
  AND U9310 ( .A(n445), .B(n9492), .Z(n9491) );
  XNOR U9311 ( .A(n9493), .B(n9494), .Z(n9488) );
  AND U9312 ( .A(n437), .B(n9495), .Z(n9494) );
  XOR U9313 ( .A(p_input[1109]), .B(n9493), .Z(n9495) );
  XNOR U9314 ( .A(n9496), .B(n9497), .Z(n9493) );
  AND U9315 ( .A(n441), .B(n9492), .Z(n9497) );
  XNOR U9316 ( .A(n9496), .B(n9490), .Z(n9492) );
  XOR U9317 ( .A(n9498), .B(n9499), .Z(n9490) );
  AND U9318 ( .A(n456), .B(n9500), .Z(n9499) );
  XNOR U9319 ( .A(n9501), .B(n9502), .Z(n9496) );
  AND U9320 ( .A(n448), .B(n9503), .Z(n9502) );
  XOR U9321 ( .A(p_input[1141]), .B(n9501), .Z(n9503) );
  XNOR U9322 ( .A(n9504), .B(n9505), .Z(n9501) );
  AND U9323 ( .A(n452), .B(n9500), .Z(n9505) );
  XNOR U9324 ( .A(n9504), .B(n9498), .Z(n9500) );
  XOR U9325 ( .A(n9506), .B(n9507), .Z(n9498) );
  AND U9326 ( .A(n467), .B(n9508), .Z(n9507) );
  XNOR U9327 ( .A(n9509), .B(n9510), .Z(n9504) );
  AND U9328 ( .A(n459), .B(n9511), .Z(n9510) );
  XOR U9329 ( .A(p_input[1173]), .B(n9509), .Z(n9511) );
  XNOR U9330 ( .A(n9512), .B(n9513), .Z(n9509) );
  AND U9331 ( .A(n463), .B(n9508), .Z(n9513) );
  XNOR U9332 ( .A(n9512), .B(n9506), .Z(n9508) );
  XOR U9333 ( .A(n9514), .B(n9515), .Z(n9506) );
  AND U9334 ( .A(n478), .B(n9516), .Z(n9515) );
  XNOR U9335 ( .A(n9517), .B(n9518), .Z(n9512) );
  AND U9336 ( .A(n470), .B(n9519), .Z(n9518) );
  XOR U9337 ( .A(p_input[1205]), .B(n9517), .Z(n9519) );
  XNOR U9338 ( .A(n9520), .B(n9521), .Z(n9517) );
  AND U9339 ( .A(n474), .B(n9516), .Z(n9521) );
  XNOR U9340 ( .A(n9520), .B(n9514), .Z(n9516) );
  XOR U9341 ( .A(n9522), .B(n9523), .Z(n9514) );
  AND U9342 ( .A(n489), .B(n9524), .Z(n9523) );
  XNOR U9343 ( .A(n9525), .B(n9526), .Z(n9520) );
  AND U9344 ( .A(n481), .B(n9527), .Z(n9526) );
  XOR U9345 ( .A(p_input[1237]), .B(n9525), .Z(n9527) );
  XNOR U9346 ( .A(n9528), .B(n9529), .Z(n9525) );
  AND U9347 ( .A(n485), .B(n9524), .Z(n9529) );
  XNOR U9348 ( .A(n9528), .B(n9522), .Z(n9524) );
  XOR U9349 ( .A(n9530), .B(n9531), .Z(n9522) );
  AND U9350 ( .A(n500), .B(n9532), .Z(n9531) );
  XNOR U9351 ( .A(n9533), .B(n9534), .Z(n9528) );
  AND U9352 ( .A(n492), .B(n9535), .Z(n9534) );
  XOR U9353 ( .A(p_input[1269]), .B(n9533), .Z(n9535) );
  XNOR U9354 ( .A(n9536), .B(n9537), .Z(n9533) );
  AND U9355 ( .A(n496), .B(n9532), .Z(n9537) );
  XNOR U9356 ( .A(n9536), .B(n9530), .Z(n9532) );
  XOR U9357 ( .A(n9538), .B(n9539), .Z(n9530) );
  AND U9358 ( .A(n511), .B(n9540), .Z(n9539) );
  XNOR U9359 ( .A(n9541), .B(n9542), .Z(n9536) );
  AND U9360 ( .A(n503), .B(n9543), .Z(n9542) );
  XOR U9361 ( .A(p_input[1301]), .B(n9541), .Z(n9543) );
  XNOR U9362 ( .A(n9544), .B(n9545), .Z(n9541) );
  AND U9363 ( .A(n507), .B(n9540), .Z(n9545) );
  XNOR U9364 ( .A(n9544), .B(n9538), .Z(n9540) );
  XOR U9365 ( .A(n9546), .B(n9547), .Z(n9538) );
  AND U9366 ( .A(n522), .B(n9548), .Z(n9547) );
  XNOR U9367 ( .A(n9549), .B(n9550), .Z(n9544) );
  AND U9368 ( .A(n514), .B(n9551), .Z(n9550) );
  XOR U9369 ( .A(p_input[1333]), .B(n9549), .Z(n9551) );
  XNOR U9370 ( .A(n9552), .B(n9553), .Z(n9549) );
  AND U9371 ( .A(n518), .B(n9548), .Z(n9553) );
  XNOR U9372 ( .A(n9552), .B(n9546), .Z(n9548) );
  XOR U9373 ( .A(n9554), .B(n9555), .Z(n9546) );
  AND U9374 ( .A(n533), .B(n9556), .Z(n9555) );
  XNOR U9375 ( .A(n9557), .B(n9558), .Z(n9552) );
  AND U9376 ( .A(n525), .B(n9559), .Z(n9558) );
  XOR U9377 ( .A(p_input[1365]), .B(n9557), .Z(n9559) );
  XNOR U9378 ( .A(n9560), .B(n9561), .Z(n9557) );
  AND U9379 ( .A(n529), .B(n9556), .Z(n9561) );
  XNOR U9380 ( .A(n9560), .B(n9554), .Z(n9556) );
  XOR U9381 ( .A(n9562), .B(n9563), .Z(n9554) );
  AND U9382 ( .A(n544), .B(n9564), .Z(n9563) );
  XNOR U9383 ( .A(n9565), .B(n9566), .Z(n9560) );
  AND U9384 ( .A(n536), .B(n9567), .Z(n9566) );
  XOR U9385 ( .A(p_input[1397]), .B(n9565), .Z(n9567) );
  XNOR U9386 ( .A(n9568), .B(n9569), .Z(n9565) );
  AND U9387 ( .A(n540), .B(n9564), .Z(n9569) );
  XNOR U9388 ( .A(n9568), .B(n9562), .Z(n9564) );
  XOR U9389 ( .A(n9570), .B(n9571), .Z(n9562) );
  AND U9390 ( .A(n555), .B(n9572), .Z(n9571) );
  XNOR U9391 ( .A(n9573), .B(n9574), .Z(n9568) );
  AND U9392 ( .A(n547), .B(n9575), .Z(n9574) );
  XOR U9393 ( .A(p_input[1429]), .B(n9573), .Z(n9575) );
  XNOR U9394 ( .A(n9576), .B(n9577), .Z(n9573) );
  AND U9395 ( .A(n551), .B(n9572), .Z(n9577) );
  XNOR U9396 ( .A(n9576), .B(n9570), .Z(n9572) );
  XOR U9397 ( .A(n9578), .B(n9579), .Z(n9570) );
  AND U9398 ( .A(n566), .B(n9580), .Z(n9579) );
  XNOR U9399 ( .A(n9581), .B(n9582), .Z(n9576) );
  AND U9400 ( .A(n558), .B(n9583), .Z(n9582) );
  XOR U9401 ( .A(p_input[1461]), .B(n9581), .Z(n9583) );
  XNOR U9402 ( .A(n9584), .B(n9585), .Z(n9581) );
  AND U9403 ( .A(n562), .B(n9580), .Z(n9585) );
  XNOR U9404 ( .A(n9584), .B(n9578), .Z(n9580) );
  XOR U9405 ( .A(n9586), .B(n9587), .Z(n9578) );
  AND U9406 ( .A(n577), .B(n9588), .Z(n9587) );
  XNOR U9407 ( .A(n9589), .B(n9590), .Z(n9584) );
  AND U9408 ( .A(n569), .B(n9591), .Z(n9590) );
  XOR U9409 ( .A(p_input[1493]), .B(n9589), .Z(n9591) );
  XNOR U9410 ( .A(n9592), .B(n9593), .Z(n9589) );
  AND U9411 ( .A(n573), .B(n9588), .Z(n9593) );
  XNOR U9412 ( .A(n9592), .B(n9586), .Z(n9588) );
  XOR U9413 ( .A(n9594), .B(n9595), .Z(n9586) );
  AND U9414 ( .A(n588), .B(n9596), .Z(n9595) );
  XNOR U9415 ( .A(n9597), .B(n9598), .Z(n9592) );
  AND U9416 ( .A(n580), .B(n9599), .Z(n9598) );
  XOR U9417 ( .A(p_input[1525]), .B(n9597), .Z(n9599) );
  XNOR U9418 ( .A(n9600), .B(n9601), .Z(n9597) );
  AND U9419 ( .A(n584), .B(n9596), .Z(n9601) );
  XNOR U9420 ( .A(n9600), .B(n9594), .Z(n9596) );
  XOR U9421 ( .A(n9602), .B(n9603), .Z(n9594) );
  AND U9422 ( .A(n599), .B(n9604), .Z(n9603) );
  XNOR U9423 ( .A(n9605), .B(n9606), .Z(n9600) );
  AND U9424 ( .A(n591), .B(n9607), .Z(n9606) );
  XOR U9425 ( .A(p_input[1557]), .B(n9605), .Z(n9607) );
  XNOR U9426 ( .A(n9608), .B(n9609), .Z(n9605) );
  AND U9427 ( .A(n595), .B(n9604), .Z(n9609) );
  XNOR U9428 ( .A(n9608), .B(n9602), .Z(n9604) );
  XOR U9429 ( .A(n9610), .B(n9611), .Z(n9602) );
  AND U9430 ( .A(n610), .B(n9612), .Z(n9611) );
  XNOR U9431 ( .A(n9613), .B(n9614), .Z(n9608) );
  AND U9432 ( .A(n602), .B(n9615), .Z(n9614) );
  XOR U9433 ( .A(p_input[1589]), .B(n9613), .Z(n9615) );
  XNOR U9434 ( .A(n9616), .B(n9617), .Z(n9613) );
  AND U9435 ( .A(n606), .B(n9612), .Z(n9617) );
  XNOR U9436 ( .A(n9616), .B(n9610), .Z(n9612) );
  XOR U9437 ( .A(n9618), .B(n9619), .Z(n9610) );
  AND U9438 ( .A(n621), .B(n9620), .Z(n9619) );
  XNOR U9439 ( .A(n9621), .B(n9622), .Z(n9616) );
  AND U9440 ( .A(n613), .B(n9623), .Z(n9622) );
  XOR U9441 ( .A(p_input[1621]), .B(n9621), .Z(n9623) );
  XNOR U9442 ( .A(n9624), .B(n9625), .Z(n9621) );
  AND U9443 ( .A(n617), .B(n9620), .Z(n9625) );
  XNOR U9444 ( .A(n9624), .B(n9618), .Z(n9620) );
  XOR U9445 ( .A(n9626), .B(n9627), .Z(n9618) );
  AND U9446 ( .A(n632), .B(n9628), .Z(n9627) );
  XNOR U9447 ( .A(n9629), .B(n9630), .Z(n9624) );
  AND U9448 ( .A(n624), .B(n9631), .Z(n9630) );
  XOR U9449 ( .A(p_input[1653]), .B(n9629), .Z(n9631) );
  XNOR U9450 ( .A(n9632), .B(n9633), .Z(n9629) );
  AND U9451 ( .A(n628), .B(n9628), .Z(n9633) );
  XNOR U9452 ( .A(n9632), .B(n9626), .Z(n9628) );
  XOR U9453 ( .A(n9634), .B(n9635), .Z(n9626) );
  AND U9454 ( .A(n643), .B(n9636), .Z(n9635) );
  XNOR U9455 ( .A(n9637), .B(n9638), .Z(n9632) );
  AND U9456 ( .A(n635), .B(n9639), .Z(n9638) );
  XOR U9457 ( .A(p_input[1685]), .B(n9637), .Z(n9639) );
  XNOR U9458 ( .A(n9640), .B(n9641), .Z(n9637) );
  AND U9459 ( .A(n639), .B(n9636), .Z(n9641) );
  XNOR U9460 ( .A(n9640), .B(n9634), .Z(n9636) );
  XOR U9461 ( .A(n9642), .B(n9643), .Z(n9634) );
  AND U9462 ( .A(n654), .B(n9644), .Z(n9643) );
  XNOR U9463 ( .A(n9645), .B(n9646), .Z(n9640) );
  AND U9464 ( .A(n646), .B(n9647), .Z(n9646) );
  XOR U9465 ( .A(p_input[1717]), .B(n9645), .Z(n9647) );
  XNOR U9466 ( .A(n9648), .B(n9649), .Z(n9645) );
  AND U9467 ( .A(n650), .B(n9644), .Z(n9649) );
  XNOR U9468 ( .A(n9648), .B(n9642), .Z(n9644) );
  XOR U9469 ( .A(n9650), .B(n9651), .Z(n9642) );
  AND U9470 ( .A(n665), .B(n9652), .Z(n9651) );
  XNOR U9471 ( .A(n9653), .B(n9654), .Z(n9648) );
  AND U9472 ( .A(n657), .B(n9655), .Z(n9654) );
  XOR U9473 ( .A(p_input[1749]), .B(n9653), .Z(n9655) );
  XNOR U9474 ( .A(n9656), .B(n9657), .Z(n9653) );
  AND U9475 ( .A(n661), .B(n9652), .Z(n9657) );
  XNOR U9476 ( .A(n9656), .B(n9650), .Z(n9652) );
  XOR U9477 ( .A(n9658), .B(n9659), .Z(n9650) );
  AND U9478 ( .A(n676), .B(n9660), .Z(n9659) );
  XNOR U9479 ( .A(n9661), .B(n9662), .Z(n9656) );
  AND U9480 ( .A(n668), .B(n9663), .Z(n9662) );
  XOR U9481 ( .A(p_input[1781]), .B(n9661), .Z(n9663) );
  XNOR U9482 ( .A(n9664), .B(n9665), .Z(n9661) );
  AND U9483 ( .A(n672), .B(n9660), .Z(n9665) );
  XNOR U9484 ( .A(n9664), .B(n9658), .Z(n9660) );
  XOR U9485 ( .A(n9666), .B(n9667), .Z(n9658) );
  AND U9486 ( .A(n687), .B(n9668), .Z(n9667) );
  XNOR U9487 ( .A(n9669), .B(n9670), .Z(n9664) );
  AND U9488 ( .A(n679), .B(n9671), .Z(n9670) );
  XOR U9489 ( .A(p_input[1813]), .B(n9669), .Z(n9671) );
  XNOR U9490 ( .A(n9672), .B(n9673), .Z(n9669) );
  AND U9491 ( .A(n683), .B(n9668), .Z(n9673) );
  XNOR U9492 ( .A(n9672), .B(n9666), .Z(n9668) );
  XOR U9493 ( .A(n9674), .B(n9675), .Z(n9666) );
  AND U9494 ( .A(n698), .B(n9676), .Z(n9675) );
  XNOR U9495 ( .A(n9677), .B(n9678), .Z(n9672) );
  AND U9496 ( .A(n690), .B(n9679), .Z(n9678) );
  XOR U9497 ( .A(p_input[1845]), .B(n9677), .Z(n9679) );
  XNOR U9498 ( .A(n9680), .B(n9681), .Z(n9677) );
  AND U9499 ( .A(n694), .B(n9676), .Z(n9681) );
  XNOR U9500 ( .A(n9680), .B(n9674), .Z(n9676) );
  XOR U9501 ( .A(n9682), .B(n9683), .Z(n9674) );
  AND U9502 ( .A(n709), .B(n9684), .Z(n9683) );
  XNOR U9503 ( .A(n9685), .B(n9686), .Z(n9680) );
  AND U9504 ( .A(n701), .B(n9687), .Z(n9686) );
  XOR U9505 ( .A(p_input[1877]), .B(n9685), .Z(n9687) );
  XNOR U9506 ( .A(n9688), .B(n9689), .Z(n9685) );
  AND U9507 ( .A(n705), .B(n9684), .Z(n9689) );
  XNOR U9508 ( .A(n9688), .B(n9682), .Z(n9684) );
  XOR U9509 ( .A(n9690), .B(n9691), .Z(n9682) );
  AND U9510 ( .A(n720), .B(n9692), .Z(n9691) );
  XNOR U9511 ( .A(n9693), .B(n9694), .Z(n9688) );
  AND U9512 ( .A(n712), .B(n9695), .Z(n9694) );
  XOR U9513 ( .A(p_input[1909]), .B(n9693), .Z(n9695) );
  XNOR U9514 ( .A(n9696), .B(n9697), .Z(n9693) );
  AND U9515 ( .A(n716), .B(n9692), .Z(n9697) );
  XNOR U9516 ( .A(n9696), .B(n9690), .Z(n9692) );
  XOR U9517 ( .A(n9698), .B(n9699), .Z(n9690) );
  AND U9518 ( .A(n731), .B(n9700), .Z(n9699) );
  XNOR U9519 ( .A(n9701), .B(n9702), .Z(n9696) );
  AND U9520 ( .A(n723), .B(n9703), .Z(n9702) );
  XOR U9521 ( .A(p_input[1941]), .B(n9701), .Z(n9703) );
  XNOR U9522 ( .A(n9704), .B(n9705), .Z(n9701) );
  AND U9523 ( .A(n727), .B(n9700), .Z(n9705) );
  XNOR U9524 ( .A(n9704), .B(n9698), .Z(n9700) );
  XOR U9525 ( .A(\knn_comb_/min_val_out[0][21] ), .B(n9706), .Z(n9698) );
  AND U9526 ( .A(n741), .B(n9707), .Z(n9706) );
  XNOR U9527 ( .A(n9708), .B(n9709), .Z(n9704) );
  AND U9528 ( .A(n734), .B(n9710), .Z(n9709) );
  XOR U9529 ( .A(p_input[1973]), .B(n9708), .Z(n9710) );
  XNOR U9530 ( .A(n9711), .B(n9712), .Z(n9708) );
  AND U9531 ( .A(n738), .B(n9707), .Z(n9712) );
  XOR U9532 ( .A(\knn_comb_/min_val_out[0][21] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .Z(n9707) );
  XOR U9533 ( .A(n33), .B(n9713), .Z(o[20]) );
  AND U9534 ( .A(n58), .B(n9714), .Z(n33) );
  XOR U9535 ( .A(n34), .B(n9713), .Z(n9714) );
  XOR U9536 ( .A(n9715), .B(n9716), .Z(n9713) );
  AND U9537 ( .A(n70), .B(n9717), .Z(n9716) );
  XOR U9538 ( .A(n9718), .B(n9719), .Z(n34) );
  AND U9539 ( .A(n62), .B(n9720), .Z(n9719) );
  XOR U9540 ( .A(p_input[20]), .B(n9718), .Z(n9720) );
  XNOR U9541 ( .A(n9721), .B(n9722), .Z(n9718) );
  AND U9542 ( .A(n66), .B(n9717), .Z(n9722) );
  XNOR U9543 ( .A(n9721), .B(n9715), .Z(n9717) );
  XOR U9544 ( .A(n9723), .B(n9724), .Z(n9715) );
  AND U9545 ( .A(n82), .B(n9725), .Z(n9724) );
  XNOR U9546 ( .A(n9726), .B(n9727), .Z(n9721) );
  AND U9547 ( .A(n74), .B(n9728), .Z(n9727) );
  XOR U9548 ( .A(p_input[52]), .B(n9726), .Z(n9728) );
  XNOR U9549 ( .A(n9729), .B(n9730), .Z(n9726) );
  AND U9550 ( .A(n78), .B(n9725), .Z(n9730) );
  XNOR U9551 ( .A(n9729), .B(n9723), .Z(n9725) );
  XOR U9552 ( .A(n9731), .B(n9732), .Z(n9723) );
  AND U9553 ( .A(n93), .B(n9733), .Z(n9732) );
  XNOR U9554 ( .A(n9734), .B(n9735), .Z(n9729) );
  AND U9555 ( .A(n85), .B(n9736), .Z(n9735) );
  XOR U9556 ( .A(p_input[84]), .B(n9734), .Z(n9736) );
  XNOR U9557 ( .A(n9737), .B(n9738), .Z(n9734) );
  AND U9558 ( .A(n89), .B(n9733), .Z(n9738) );
  XNOR U9559 ( .A(n9737), .B(n9731), .Z(n9733) );
  XOR U9560 ( .A(n9739), .B(n9740), .Z(n9731) );
  AND U9561 ( .A(n104), .B(n9741), .Z(n9740) );
  XNOR U9562 ( .A(n9742), .B(n9743), .Z(n9737) );
  AND U9563 ( .A(n96), .B(n9744), .Z(n9743) );
  XOR U9564 ( .A(p_input[116]), .B(n9742), .Z(n9744) );
  XNOR U9565 ( .A(n9745), .B(n9746), .Z(n9742) );
  AND U9566 ( .A(n100), .B(n9741), .Z(n9746) );
  XNOR U9567 ( .A(n9745), .B(n9739), .Z(n9741) );
  XOR U9568 ( .A(n9747), .B(n9748), .Z(n9739) );
  AND U9569 ( .A(n115), .B(n9749), .Z(n9748) );
  XNOR U9570 ( .A(n9750), .B(n9751), .Z(n9745) );
  AND U9571 ( .A(n107), .B(n9752), .Z(n9751) );
  XOR U9572 ( .A(p_input[148]), .B(n9750), .Z(n9752) );
  XNOR U9573 ( .A(n9753), .B(n9754), .Z(n9750) );
  AND U9574 ( .A(n111), .B(n9749), .Z(n9754) );
  XNOR U9575 ( .A(n9753), .B(n9747), .Z(n9749) );
  XOR U9576 ( .A(n9755), .B(n9756), .Z(n9747) );
  AND U9577 ( .A(n126), .B(n9757), .Z(n9756) );
  XNOR U9578 ( .A(n9758), .B(n9759), .Z(n9753) );
  AND U9579 ( .A(n118), .B(n9760), .Z(n9759) );
  XOR U9580 ( .A(p_input[180]), .B(n9758), .Z(n9760) );
  XNOR U9581 ( .A(n9761), .B(n9762), .Z(n9758) );
  AND U9582 ( .A(n122), .B(n9757), .Z(n9762) );
  XNOR U9583 ( .A(n9761), .B(n9755), .Z(n9757) );
  XOR U9584 ( .A(n9763), .B(n9764), .Z(n9755) );
  AND U9585 ( .A(n137), .B(n9765), .Z(n9764) );
  XNOR U9586 ( .A(n9766), .B(n9767), .Z(n9761) );
  AND U9587 ( .A(n129), .B(n9768), .Z(n9767) );
  XOR U9588 ( .A(p_input[212]), .B(n9766), .Z(n9768) );
  XNOR U9589 ( .A(n9769), .B(n9770), .Z(n9766) );
  AND U9590 ( .A(n133), .B(n9765), .Z(n9770) );
  XNOR U9591 ( .A(n9769), .B(n9763), .Z(n9765) );
  XOR U9592 ( .A(n9771), .B(n9772), .Z(n9763) );
  AND U9593 ( .A(n148), .B(n9773), .Z(n9772) );
  XNOR U9594 ( .A(n9774), .B(n9775), .Z(n9769) );
  AND U9595 ( .A(n140), .B(n9776), .Z(n9775) );
  XOR U9596 ( .A(p_input[244]), .B(n9774), .Z(n9776) );
  XNOR U9597 ( .A(n9777), .B(n9778), .Z(n9774) );
  AND U9598 ( .A(n144), .B(n9773), .Z(n9778) );
  XNOR U9599 ( .A(n9777), .B(n9771), .Z(n9773) );
  XOR U9600 ( .A(n9779), .B(n9780), .Z(n9771) );
  AND U9601 ( .A(n159), .B(n9781), .Z(n9780) );
  XNOR U9602 ( .A(n9782), .B(n9783), .Z(n9777) );
  AND U9603 ( .A(n151), .B(n9784), .Z(n9783) );
  XOR U9604 ( .A(p_input[276]), .B(n9782), .Z(n9784) );
  XNOR U9605 ( .A(n9785), .B(n9786), .Z(n9782) );
  AND U9606 ( .A(n155), .B(n9781), .Z(n9786) );
  XNOR U9607 ( .A(n9785), .B(n9779), .Z(n9781) );
  XOR U9608 ( .A(n9787), .B(n9788), .Z(n9779) );
  AND U9609 ( .A(n170), .B(n9789), .Z(n9788) );
  XNOR U9610 ( .A(n9790), .B(n9791), .Z(n9785) );
  AND U9611 ( .A(n162), .B(n9792), .Z(n9791) );
  XOR U9612 ( .A(p_input[308]), .B(n9790), .Z(n9792) );
  XNOR U9613 ( .A(n9793), .B(n9794), .Z(n9790) );
  AND U9614 ( .A(n166), .B(n9789), .Z(n9794) );
  XNOR U9615 ( .A(n9793), .B(n9787), .Z(n9789) );
  XOR U9616 ( .A(n9795), .B(n9796), .Z(n9787) );
  AND U9617 ( .A(n181), .B(n9797), .Z(n9796) );
  XNOR U9618 ( .A(n9798), .B(n9799), .Z(n9793) );
  AND U9619 ( .A(n173), .B(n9800), .Z(n9799) );
  XOR U9620 ( .A(p_input[340]), .B(n9798), .Z(n9800) );
  XNOR U9621 ( .A(n9801), .B(n9802), .Z(n9798) );
  AND U9622 ( .A(n177), .B(n9797), .Z(n9802) );
  XNOR U9623 ( .A(n9801), .B(n9795), .Z(n9797) );
  XOR U9624 ( .A(n9803), .B(n9804), .Z(n9795) );
  AND U9625 ( .A(n192), .B(n9805), .Z(n9804) );
  XNOR U9626 ( .A(n9806), .B(n9807), .Z(n9801) );
  AND U9627 ( .A(n184), .B(n9808), .Z(n9807) );
  XOR U9628 ( .A(p_input[372]), .B(n9806), .Z(n9808) );
  XNOR U9629 ( .A(n9809), .B(n9810), .Z(n9806) );
  AND U9630 ( .A(n188), .B(n9805), .Z(n9810) );
  XNOR U9631 ( .A(n9809), .B(n9803), .Z(n9805) );
  XOR U9632 ( .A(n9811), .B(n9812), .Z(n9803) );
  AND U9633 ( .A(n203), .B(n9813), .Z(n9812) );
  XNOR U9634 ( .A(n9814), .B(n9815), .Z(n9809) );
  AND U9635 ( .A(n195), .B(n9816), .Z(n9815) );
  XOR U9636 ( .A(p_input[404]), .B(n9814), .Z(n9816) );
  XNOR U9637 ( .A(n9817), .B(n9818), .Z(n9814) );
  AND U9638 ( .A(n199), .B(n9813), .Z(n9818) );
  XNOR U9639 ( .A(n9817), .B(n9811), .Z(n9813) );
  XOR U9640 ( .A(n9819), .B(n9820), .Z(n9811) );
  AND U9641 ( .A(n214), .B(n9821), .Z(n9820) );
  XNOR U9642 ( .A(n9822), .B(n9823), .Z(n9817) );
  AND U9643 ( .A(n206), .B(n9824), .Z(n9823) );
  XOR U9644 ( .A(p_input[436]), .B(n9822), .Z(n9824) );
  XNOR U9645 ( .A(n9825), .B(n9826), .Z(n9822) );
  AND U9646 ( .A(n210), .B(n9821), .Z(n9826) );
  XNOR U9647 ( .A(n9825), .B(n9819), .Z(n9821) );
  XOR U9648 ( .A(n9827), .B(n9828), .Z(n9819) );
  AND U9649 ( .A(n225), .B(n9829), .Z(n9828) );
  XNOR U9650 ( .A(n9830), .B(n9831), .Z(n9825) );
  AND U9651 ( .A(n217), .B(n9832), .Z(n9831) );
  XOR U9652 ( .A(p_input[468]), .B(n9830), .Z(n9832) );
  XNOR U9653 ( .A(n9833), .B(n9834), .Z(n9830) );
  AND U9654 ( .A(n221), .B(n9829), .Z(n9834) );
  XNOR U9655 ( .A(n9833), .B(n9827), .Z(n9829) );
  XOR U9656 ( .A(n9835), .B(n9836), .Z(n9827) );
  AND U9657 ( .A(n236), .B(n9837), .Z(n9836) );
  XNOR U9658 ( .A(n9838), .B(n9839), .Z(n9833) );
  AND U9659 ( .A(n228), .B(n9840), .Z(n9839) );
  XOR U9660 ( .A(p_input[500]), .B(n9838), .Z(n9840) );
  XNOR U9661 ( .A(n9841), .B(n9842), .Z(n9838) );
  AND U9662 ( .A(n232), .B(n9837), .Z(n9842) );
  XNOR U9663 ( .A(n9841), .B(n9835), .Z(n9837) );
  XOR U9664 ( .A(n9843), .B(n9844), .Z(n9835) );
  AND U9665 ( .A(n247), .B(n9845), .Z(n9844) );
  XNOR U9666 ( .A(n9846), .B(n9847), .Z(n9841) );
  AND U9667 ( .A(n239), .B(n9848), .Z(n9847) );
  XOR U9668 ( .A(p_input[532]), .B(n9846), .Z(n9848) );
  XNOR U9669 ( .A(n9849), .B(n9850), .Z(n9846) );
  AND U9670 ( .A(n243), .B(n9845), .Z(n9850) );
  XNOR U9671 ( .A(n9849), .B(n9843), .Z(n9845) );
  XOR U9672 ( .A(n9851), .B(n9852), .Z(n9843) );
  AND U9673 ( .A(n258), .B(n9853), .Z(n9852) );
  XNOR U9674 ( .A(n9854), .B(n9855), .Z(n9849) );
  AND U9675 ( .A(n250), .B(n9856), .Z(n9855) );
  XOR U9676 ( .A(p_input[564]), .B(n9854), .Z(n9856) );
  XNOR U9677 ( .A(n9857), .B(n9858), .Z(n9854) );
  AND U9678 ( .A(n254), .B(n9853), .Z(n9858) );
  XNOR U9679 ( .A(n9857), .B(n9851), .Z(n9853) );
  XOR U9680 ( .A(n9859), .B(n9860), .Z(n9851) );
  AND U9681 ( .A(n269), .B(n9861), .Z(n9860) );
  XNOR U9682 ( .A(n9862), .B(n9863), .Z(n9857) );
  AND U9683 ( .A(n261), .B(n9864), .Z(n9863) );
  XOR U9684 ( .A(p_input[596]), .B(n9862), .Z(n9864) );
  XNOR U9685 ( .A(n9865), .B(n9866), .Z(n9862) );
  AND U9686 ( .A(n265), .B(n9861), .Z(n9866) );
  XNOR U9687 ( .A(n9865), .B(n9859), .Z(n9861) );
  XOR U9688 ( .A(n9867), .B(n9868), .Z(n9859) );
  AND U9689 ( .A(n280), .B(n9869), .Z(n9868) );
  XNOR U9690 ( .A(n9870), .B(n9871), .Z(n9865) );
  AND U9691 ( .A(n272), .B(n9872), .Z(n9871) );
  XOR U9692 ( .A(p_input[628]), .B(n9870), .Z(n9872) );
  XNOR U9693 ( .A(n9873), .B(n9874), .Z(n9870) );
  AND U9694 ( .A(n276), .B(n9869), .Z(n9874) );
  XNOR U9695 ( .A(n9873), .B(n9867), .Z(n9869) );
  XOR U9696 ( .A(n9875), .B(n9876), .Z(n9867) );
  AND U9697 ( .A(n291), .B(n9877), .Z(n9876) );
  XNOR U9698 ( .A(n9878), .B(n9879), .Z(n9873) );
  AND U9699 ( .A(n283), .B(n9880), .Z(n9879) );
  XOR U9700 ( .A(p_input[660]), .B(n9878), .Z(n9880) );
  XNOR U9701 ( .A(n9881), .B(n9882), .Z(n9878) );
  AND U9702 ( .A(n287), .B(n9877), .Z(n9882) );
  XNOR U9703 ( .A(n9881), .B(n9875), .Z(n9877) );
  XOR U9704 ( .A(n9883), .B(n9884), .Z(n9875) );
  AND U9705 ( .A(n302), .B(n9885), .Z(n9884) );
  XNOR U9706 ( .A(n9886), .B(n9887), .Z(n9881) );
  AND U9707 ( .A(n294), .B(n9888), .Z(n9887) );
  XOR U9708 ( .A(p_input[692]), .B(n9886), .Z(n9888) );
  XNOR U9709 ( .A(n9889), .B(n9890), .Z(n9886) );
  AND U9710 ( .A(n298), .B(n9885), .Z(n9890) );
  XNOR U9711 ( .A(n9889), .B(n9883), .Z(n9885) );
  XOR U9712 ( .A(n9891), .B(n9892), .Z(n9883) );
  AND U9713 ( .A(n313), .B(n9893), .Z(n9892) );
  XNOR U9714 ( .A(n9894), .B(n9895), .Z(n9889) );
  AND U9715 ( .A(n305), .B(n9896), .Z(n9895) );
  XOR U9716 ( .A(p_input[724]), .B(n9894), .Z(n9896) );
  XNOR U9717 ( .A(n9897), .B(n9898), .Z(n9894) );
  AND U9718 ( .A(n309), .B(n9893), .Z(n9898) );
  XNOR U9719 ( .A(n9897), .B(n9891), .Z(n9893) );
  XOR U9720 ( .A(n9899), .B(n9900), .Z(n9891) );
  AND U9721 ( .A(n324), .B(n9901), .Z(n9900) );
  XNOR U9722 ( .A(n9902), .B(n9903), .Z(n9897) );
  AND U9723 ( .A(n316), .B(n9904), .Z(n9903) );
  XOR U9724 ( .A(p_input[756]), .B(n9902), .Z(n9904) );
  XNOR U9725 ( .A(n9905), .B(n9906), .Z(n9902) );
  AND U9726 ( .A(n320), .B(n9901), .Z(n9906) );
  XNOR U9727 ( .A(n9905), .B(n9899), .Z(n9901) );
  XOR U9728 ( .A(n9907), .B(n9908), .Z(n9899) );
  AND U9729 ( .A(n335), .B(n9909), .Z(n9908) );
  XNOR U9730 ( .A(n9910), .B(n9911), .Z(n9905) );
  AND U9731 ( .A(n327), .B(n9912), .Z(n9911) );
  XOR U9732 ( .A(p_input[788]), .B(n9910), .Z(n9912) );
  XNOR U9733 ( .A(n9913), .B(n9914), .Z(n9910) );
  AND U9734 ( .A(n331), .B(n9909), .Z(n9914) );
  XNOR U9735 ( .A(n9913), .B(n9907), .Z(n9909) );
  XOR U9736 ( .A(n9915), .B(n9916), .Z(n9907) );
  AND U9737 ( .A(n346), .B(n9917), .Z(n9916) );
  XNOR U9738 ( .A(n9918), .B(n9919), .Z(n9913) );
  AND U9739 ( .A(n338), .B(n9920), .Z(n9919) );
  XOR U9740 ( .A(p_input[820]), .B(n9918), .Z(n9920) );
  XNOR U9741 ( .A(n9921), .B(n9922), .Z(n9918) );
  AND U9742 ( .A(n342), .B(n9917), .Z(n9922) );
  XNOR U9743 ( .A(n9921), .B(n9915), .Z(n9917) );
  XOR U9744 ( .A(n9923), .B(n9924), .Z(n9915) );
  AND U9745 ( .A(n357), .B(n9925), .Z(n9924) );
  XNOR U9746 ( .A(n9926), .B(n9927), .Z(n9921) );
  AND U9747 ( .A(n349), .B(n9928), .Z(n9927) );
  XOR U9748 ( .A(p_input[852]), .B(n9926), .Z(n9928) );
  XNOR U9749 ( .A(n9929), .B(n9930), .Z(n9926) );
  AND U9750 ( .A(n353), .B(n9925), .Z(n9930) );
  XNOR U9751 ( .A(n9929), .B(n9923), .Z(n9925) );
  XOR U9752 ( .A(n9931), .B(n9932), .Z(n9923) );
  AND U9753 ( .A(n368), .B(n9933), .Z(n9932) );
  XNOR U9754 ( .A(n9934), .B(n9935), .Z(n9929) );
  AND U9755 ( .A(n360), .B(n9936), .Z(n9935) );
  XOR U9756 ( .A(p_input[884]), .B(n9934), .Z(n9936) );
  XNOR U9757 ( .A(n9937), .B(n9938), .Z(n9934) );
  AND U9758 ( .A(n364), .B(n9933), .Z(n9938) );
  XNOR U9759 ( .A(n9937), .B(n9931), .Z(n9933) );
  XOR U9760 ( .A(n9939), .B(n9940), .Z(n9931) );
  AND U9761 ( .A(n379), .B(n9941), .Z(n9940) );
  XNOR U9762 ( .A(n9942), .B(n9943), .Z(n9937) );
  AND U9763 ( .A(n371), .B(n9944), .Z(n9943) );
  XOR U9764 ( .A(p_input[916]), .B(n9942), .Z(n9944) );
  XNOR U9765 ( .A(n9945), .B(n9946), .Z(n9942) );
  AND U9766 ( .A(n375), .B(n9941), .Z(n9946) );
  XNOR U9767 ( .A(n9945), .B(n9939), .Z(n9941) );
  XOR U9768 ( .A(n9947), .B(n9948), .Z(n9939) );
  AND U9769 ( .A(n390), .B(n9949), .Z(n9948) );
  XNOR U9770 ( .A(n9950), .B(n9951), .Z(n9945) );
  AND U9771 ( .A(n382), .B(n9952), .Z(n9951) );
  XOR U9772 ( .A(p_input[948]), .B(n9950), .Z(n9952) );
  XNOR U9773 ( .A(n9953), .B(n9954), .Z(n9950) );
  AND U9774 ( .A(n386), .B(n9949), .Z(n9954) );
  XNOR U9775 ( .A(n9953), .B(n9947), .Z(n9949) );
  XOR U9776 ( .A(n9955), .B(n9956), .Z(n9947) );
  AND U9777 ( .A(n401), .B(n9957), .Z(n9956) );
  XNOR U9778 ( .A(n9958), .B(n9959), .Z(n9953) );
  AND U9779 ( .A(n393), .B(n9960), .Z(n9959) );
  XOR U9780 ( .A(p_input[980]), .B(n9958), .Z(n9960) );
  XNOR U9781 ( .A(n9961), .B(n9962), .Z(n9958) );
  AND U9782 ( .A(n397), .B(n9957), .Z(n9962) );
  XNOR U9783 ( .A(n9961), .B(n9955), .Z(n9957) );
  XOR U9784 ( .A(n9963), .B(n9964), .Z(n9955) );
  AND U9785 ( .A(n412), .B(n9965), .Z(n9964) );
  XNOR U9786 ( .A(n9966), .B(n9967), .Z(n9961) );
  AND U9787 ( .A(n404), .B(n9968), .Z(n9967) );
  XOR U9788 ( .A(p_input[1012]), .B(n9966), .Z(n9968) );
  XNOR U9789 ( .A(n9969), .B(n9970), .Z(n9966) );
  AND U9790 ( .A(n408), .B(n9965), .Z(n9970) );
  XNOR U9791 ( .A(n9969), .B(n9963), .Z(n9965) );
  XOR U9792 ( .A(n9971), .B(n9972), .Z(n9963) );
  AND U9793 ( .A(n423), .B(n9973), .Z(n9972) );
  XNOR U9794 ( .A(n9974), .B(n9975), .Z(n9969) );
  AND U9795 ( .A(n415), .B(n9976), .Z(n9975) );
  XOR U9796 ( .A(p_input[1044]), .B(n9974), .Z(n9976) );
  XNOR U9797 ( .A(n9977), .B(n9978), .Z(n9974) );
  AND U9798 ( .A(n419), .B(n9973), .Z(n9978) );
  XNOR U9799 ( .A(n9977), .B(n9971), .Z(n9973) );
  XOR U9800 ( .A(n9979), .B(n9980), .Z(n9971) );
  AND U9801 ( .A(n434), .B(n9981), .Z(n9980) );
  XNOR U9802 ( .A(n9982), .B(n9983), .Z(n9977) );
  AND U9803 ( .A(n426), .B(n9984), .Z(n9983) );
  XOR U9804 ( .A(p_input[1076]), .B(n9982), .Z(n9984) );
  XNOR U9805 ( .A(n9985), .B(n9986), .Z(n9982) );
  AND U9806 ( .A(n430), .B(n9981), .Z(n9986) );
  XNOR U9807 ( .A(n9985), .B(n9979), .Z(n9981) );
  XOR U9808 ( .A(n9987), .B(n9988), .Z(n9979) );
  AND U9809 ( .A(n445), .B(n9989), .Z(n9988) );
  XNOR U9810 ( .A(n9990), .B(n9991), .Z(n9985) );
  AND U9811 ( .A(n437), .B(n9992), .Z(n9991) );
  XOR U9812 ( .A(p_input[1108]), .B(n9990), .Z(n9992) );
  XNOR U9813 ( .A(n9993), .B(n9994), .Z(n9990) );
  AND U9814 ( .A(n441), .B(n9989), .Z(n9994) );
  XNOR U9815 ( .A(n9993), .B(n9987), .Z(n9989) );
  XOR U9816 ( .A(n9995), .B(n9996), .Z(n9987) );
  AND U9817 ( .A(n456), .B(n9997), .Z(n9996) );
  XNOR U9818 ( .A(n9998), .B(n9999), .Z(n9993) );
  AND U9819 ( .A(n448), .B(n10000), .Z(n9999) );
  XOR U9820 ( .A(p_input[1140]), .B(n9998), .Z(n10000) );
  XNOR U9821 ( .A(n10001), .B(n10002), .Z(n9998) );
  AND U9822 ( .A(n452), .B(n9997), .Z(n10002) );
  XNOR U9823 ( .A(n10001), .B(n9995), .Z(n9997) );
  XOR U9824 ( .A(n10003), .B(n10004), .Z(n9995) );
  AND U9825 ( .A(n467), .B(n10005), .Z(n10004) );
  XNOR U9826 ( .A(n10006), .B(n10007), .Z(n10001) );
  AND U9827 ( .A(n459), .B(n10008), .Z(n10007) );
  XOR U9828 ( .A(p_input[1172]), .B(n10006), .Z(n10008) );
  XNOR U9829 ( .A(n10009), .B(n10010), .Z(n10006) );
  AND U9830 ( .A(n463), .B(n10005), .Z(n10010) );
  XNOR U9831 ( .A(n10009), .B(n10003), .Z(n10005) );
  XOR U9832 ( .A(n10011), .B(n10012), .Z(n10003) );
  AND U9833 ( .A(n478), .B(n10013), .Z(n10012) );
  XNOR U9834 ( .A(n10014), .B(n10015), .Z(n10009) );
  AND U9835 ( .A(n470), .B(n10016), .Z(n10015) );
  XOR U9836 ( .A(p_input[1204]), .B(n10014), .Z(n10016) );
  XNOR U9837 ( .A(n10017), .B(n10018), .Z(n10014) );
  AND U9838 ( .A(n474), .B(n10013), .Z(n10018) );
  XNOR U9839 ( .A(n10017), .B(n10011), .Z(n10013) );
  XOR U9840 ( .A(n10019), .B(n10020), .Z(n10011) );
  AND U9841 ( .A(n489), .B(n10021), .Z(n10020) );
  XNOR U9842 ( .A(n10022), .B(n10023), .Z(n10017) );
  AND U9843 ( .A(n481), .B(n10024), .Z(n10023) );
  XOR U9844 ( .A(p_input[1236]), .B(n10022), .Z(n10024) );
  XNOR U9845 ( .A(n10025), .B(n10026), .Z(n10022) );
  AND U9846 ( .A(n485), .B(n10021), .Z(n10026) );
  XNOR U9847 ( .A(n10025), .B(n10019), .Z(n10021) );
  XOR U9848 ( .A(n10027), .B(n10028), .Z(n10019) );
  AND U9849 ( .A(n500), .B(n10029), .Z(n10028) );
  XNOR U9850 ( .A(n10030), .B(n10031), .Z(n10025) );
  AND U9851 ( .A(n492), .B(n10032), .Z(n10031) );
  XOR U9852 ( .A(p_input[1268]), .B(n10030), .Z(n10032) );
  XNOR U9853 ( .A(n10033), .B(n10034), .Z(n10030) );
  AND U9854 ( .A(n496), .B(n10029), .Z(n10034) );
  XNOR U9855 ( .A(n10033), .B(n10027), .Z(n10029) );
  XOR U9856 ( .A(n10035), .B(n10036), .Z(n10027) );
  AND U9857 ( .A(n511), .B(n10037), .Z(n10036) );
  XNOR U9858 ( .A(n10038), .B(n10039), .Z(n10033) );
  AND U9859 ( .A(n503), .B(n10040), .Z(n10039) );
  XOR U9860 ( .A(p_input[1300]), .B(n10038), .Z(n10040) );
  XNOR U9861 ( .A(n10041), .B(n10042), .Z(n10038) );
  AND U9862 ( .A(n507), .B(n10037), .Z(n10042) );
  XNOR U9863 ( .A(n10041), .B(n10035), .Z(n10037) );
  XOR U9864 ( .A(n10043), .B(n10044), .Z(n10035) );
  AND U9865 ( .A(n522), .B(n10045), .Z(n10044) );
  XNOR U9866 ( .A(n10046), .B(n10047), .Z(n10041) );
  AND U9867 ( .A(n514), .B(n10048), .Z(n10047) );
  XOR U9868 ( .A(p_input[1332]), .B(n10046), .Z(n10048) );
  XNOR U9869 ( .A(n10049), .B(n10050), .Z(n10046) );
  AND U9870 ( .A(n518), .B(n10045), .Z(n10050) );
  XNOR U9871 ( .A(n10049), .B(n10043), .Z(n10045) );
  XOR U9872 ( .A(n10051), .B(n10052), .Z(n10043) );
  AND U9873 ( .A(n533), .B(n10053), .Z(n10052) );
  XNOR U9874 ( .A(n10054), .B(n10055), .Z(n10049) );
  AND U9875 ( .A(n525), .B(n10056), .Z(n10055) );
  XOR U9876 ( .A(p_input[1364]), .B(n10054), .Z(n10056) );
  XNOR U9877 ( .A(n10057), .B(n10058), .Z(n10054) );
  AND U9878 ( .A(n529), .B(n10053), .Z(n10058) );
  XNOR U9879 ( .A(n10057), .B(n10051), .Z(n10053) );
  XOR U9880 ( .A(n10059), .B(n10060), .Z(n10051) );
  AND U9881 ( .A(n544), .B(n10061), .Z(n10060) );
  XNOR U9882 ( .A(n10062), .B(n10063), .Z(n10057) );
  AND U9883 ( .A(n536), .B(n10064), .Z(n10063) );
  XOR U9884 ( .A(p_input[1396]), .B(n10062), .Z(n10064) );
  XNOR U9885 ( .A(n10065), .B(n10066), .Z(n10062) );
  AND U9886 ( .A(n540), .B(n10061), .Z(n10066) );
  XNOR U9887 ( .A(n10065), .B(n10059), .Z(n10061) );
  XOR U9888 ( .A(n10067), .B(n10068), .Z(n10059) );
  AND U9889 ( .A(n555), .B(n10069), .Z(n10068) );
  XNOR U9890 ( .A(n10070), .B(n10071), .Z(n10065) );
  AND U9891 ( .A(n547), .B(n10072), .Z(n10071) );
  XOR U9892 ( .A(p_input[1428]), .B(n10070), .Z(n10072) );
  XNOR U9893 ( .A(n10073), .B(n10074), .Z(n10070) );
  AND U9894 ( .A(n551), .B(n10069), .Z(n10074) );
  XNOR U9895 ( .A(n10073), .B(n10067), .Z(n10069) );
  XOR U9896 ( .A(n10075), .B(n10076), .Z(n10067) );
  AND U9897 ( .A(n566), .B(n10077), .Z(n10076) );
  XNOR U9898 ( .A(n10078), .B(n10079), .Z(n10073) );
  AND U9899 ( .A(n558), .B(n10080), .Z(n10079) );
  XOR U9900 ( .A(p_input[1460]), .B(n10078), .Z(n10080) );
  XNOR U9901 ( .A(n10081), .B(n10082), .Z(n10078) );
  AND U9902 ( .A(n562), .B(n10077), .Z(n10082) );
  XNOR U9903 ( .A(n10081), .B(n10075), .Z(n10077) );
  XOR U9904 ( .A(n10083), .B(n10084), .Z(n10075) );
  AND U9905 ( .A(n577), .B(n10085), .Z(n10084) );
  XNOR U9906 ( .A(n10086), .B(n10087), .Z(n10081) );
  AND U9907 ( .A(n569), .B(n10088), .Z(n10087) );
  XOR U9908 ( .A(p_input[1492]), .B(n10086), .Z(n10088) );
  XNOR U9909 ( .A(n10089), .B(n10090), .Z(n10086) );
  AND U9910 ( .A(n573), .B(n10085), .Z(n10090) );
  XNOR U9911 ( .A(n10089), .B(n10083), .Z(n10085) );
  XOR U9912 ( .A(n10091), .B(n10092), .Z(n10083) );
  AND U9913 ( .A(n588), .B(n10093), .Z(n10092) );
  XNOR U9914 ( .A(n10094), .B(n10095), .Z(n10089) );
  AND U9915 ( .A(n580), .B(n10096), .Z(n10095) );
  XOR U9916 ( .A(p_input[1524]), .B(n10094), .Z(n10096) );
  XNOR U9917 ( .A(n10097), .B(n10098), .Z(n10094) );
  AND U9918 ( .A(n584), .B(n10093), .Z(n10098) );
  XNOR U9919 ( .A(n10097), .B(n10091), .Z(n10093) );
  XOR U9920 ( .A(n10099), .B(n10100), .Z(n10091) );
  AND U9921 ( .A(n599), .B(n10101), .Z(n10100) );
  XNOR U9922 ( .A(n10102), .B(n10103), .Z(n10097) );
  AND U9923 ( .A(n591), .B(n10104), .Z(n10103) );
  XOR U9924 ( .A(p_input[1556]), .B(n10102), .Z(n10104) );
  XNOR U9925 ( .A(n10105), .B(n10106), .Z(n10102) );
  AND U9926 ( .A(n595), .B(n10101), .Z(n10106) );
  XNOR U9927 ( .A(n10105), .B(n10099), .Z(n10101) );
  XOR U9928 ( .A(n10107), .B(n10108), .Z(n10099) );
  AND U9929 ( .A(n610), .B(n10109), .Z(n10108) );
  XNOR U9930 ( .A(n10110), .B(n10111), .Z(n10105) );
  AND U9931 ( .A(n602), .B(n10112), .Z(n10111) );
  XOR U9932 ( .A(p_input[1588]), .B(n10110), .Z(n10112) );
  XNOR U9933 ( .A(n10113), .B(n10114), .Z(n10110) );
  AND U9934 ( .A(n606), .B(n10109), .Z(n10114) );
  XNOR U9935 ( .A(n10113), .B(n10107), .Z(n10109) );
  XOR U9936 ( .A(n10115), .B(n10116), .Z(n10107) );
  AND U9937 ( .A(n621), .B(n10117), .Z(n10116) );
  XNOR U9938 ( .A(n10118), .B(n10119), .Z(n10113) );
  AND U9939 ( .A(n613), .B(n10120), .Z(n10119) );
  XOR U9940 ( .A(p_input[1620]), .B(n10118), .Z(n10120) );
  XNOR U9941 ( .A(n10121), .B(n10122), .Z(n10118) );
  AND U9942 ( .A(n617), .B(n10117), .Z(n10122) );
  XNOR U9943 ( .A(n10121), .B(n10115), .Z(n10117) );
  XOR U9944 ( .A(n10123), .B(n10124), .Z(n10115) );
  AND U9945 ( .A(n632), .B(n10125), .Z(n10124) );
  XNOR U9946 ( .A(n10126), .B(n10127), .Z(n10121) );
  AND U9947 ( .A(n624), .B(n10128), .Z(n10127) );
  XOR U9948 ( .A(p_input[1652]), .B(n10126), .Z(n10128) );
  XNOR U9949 ( .A(n10129), .B(n10130), .Z(n10126) );
  AND U9950 ( .A(n628), .B(n10125), .Z(n10130) );
  XNOR U9951 ( .A(n10129), .B(n10123), .Z(n10125) );
  XOR U9952 ( .A(n10131), .B(n10132), .Z(n10123) );
  AND U9953 ( .A(n643), .B(n10133), .Z(n10132) );
  XNOR U9954 ( .A(n10134), .B(n10135), .Z(n10129) );
  AND U9955 ( .A(n635), .B(n10136), .Z(n10135) );
  XOR U9956 ( .A(p_input[1684]), .B(n10134), .Z(n10136) );
  XNOR U9957 ( .A(n10137), .B(n10138), .Z(n10134) );
  AND U9958 ( .A(n639), .B(n10133), .Z(n10138) );
  XNOR U9959 ( .A(n10137), .B(n10131), .Z(n10133) );
  XOR U9960 ( .A(n10139), .B(n10140), .Z(n10131) );
  AND U9961 ( .A(n654), .B(n10141), .Z(n10140) );
  XNOR U9962 ( .A(n10142), .B(n10143), .Z(n10137) );
  AND U9963 ( .A(n646), .B(n10144), .Z(n10143) );
  XOR U9964 ( .A(p_input[1716]), .B(n10142), .Z(n10144) );
  XNOR U9965 ( .A(n10145), .B(n10146), .Z(n10142) );
  AND U9966 ( .A(n650), .B(n10141), .Z(n10146) );
  XNOR U9967 ( .A(n10145), .B(n10139), .Z(n10141) );
  XOR U9968 ( .A(n10147), .B(n10148), .Z(n10139) );
  AND U9969 ( .A(n665), .B(n10149), .Z(n10148) );
  XNOR U9970 ( .A(n10150), .B(n10151), .Z(n10145) );
  AND U9971 ( .A(n657), .B(n10152), .Z(n10151) );
  XOR U9972 ( .A(p_input[1748]), .B(n10150), .Z(n10152) );
  XNOR U9973 ( .A(n10153), .B(n10154), .Z(n10150) );
  AND U9974 ( .A(n661), .B(n10149), .Z(n10154) );
  XNOR U9975 ( .A(n10153), .B(n10147), .Z(n10149) );
  XOR U9976 ( .A(n10155), .B(n10156), .Z(n10147) );
  AND U9977 ( .A(n676), .B(n10157), .Z(n10156) );
  XNOR U9978 ( .A(n10158), .B(n10159), .Z(n10153) );
  AND U9979 ( .A(n668), .B(n10160), .Z(n10159) );
  XOR U9980 ( .A(p_input[1780]), .B(n10158), .Z(n10160) );
  XNOR U9981 ( .A(n10161), .B(n10162), .Z(n10158) );
  AND U9982 ( .A(n672), .B(n10157), .Z(n10162) );
  XNOR U9983 ( .A(n10161), .B(n10155), .Z(n10157) );
  XOR U9984 ( .A(n10163), .B(n10164), .Z(n10155) );
  AND U9985 ( .A(n687), .B(n10165), .Z(n10164) );
  XNOR U9986 ( .A(n10166), .B(n10167), .Z(n10161) );
  AND U9987 ( .A(n679), .B(n10168), .Z(n10167) );
  XOR U9988 ( .A(p_input[1812]), .B(n10166), .Z(n10168) );
  XNOR U9989 ( .A(n10169), .B(n10170), .Z(n10166) );
  AND U9990 ( .A(n683), .B(n10165), .Z(n10170) );
  XNOR U9991 ( .A(n10169), .B(n10163), .Z(n10165) );
  XOR U9992 ( .A(n10171), .B(n10172), .Z(n10163) );
  AND U9993 ( .A(n698), .B(n10173), .Z(n10172) );
  XNOR U9994 ( .A(n10174), .B(n10175), .Z(n10169) );
  AND U9995 ( .A(n690), .B(n10176), .Z(n10175) );
  XOR U9996 ( .A(p_input[1844]), .B(n10174), .Z(n10176) );
  XNOR U9997 ( .A(n10177), .B(n10178), .Z(n10174) );
  AND U9998 ( .A(n694), .B(n10173), .Z(n10178) );
  XNOR U9999 ( .A(n10177), .B(n10171), .Z(n10173) );
  XOR U10000 ( .A(n10179), .B(n10180), .Z(n10171) );
  AND U10001 ( .A(n709), .B(n10181), .Z(n10180) );
  XNOR U10002 ( .A(n10182), .B(n10183), .Z(n10177) );
  AND U10003 ( .A(n701), .B(n10184), .Z(n10183) );
  XOR U10004 ( .A(p_input[1876]), .B(n10182), .Z(n10184) );
  XNOR U10005 ( .A(n10185), .B(n10186), .Z(n10182) );
  AND U10006 ( .A(n705), .B(n10181), .Z(n10186) );
  XNOR U10007 ( .A(n10185), .B(n10179), .Z(n10181) );
  XOR U10008 ( .A(n10187), .B(n10188), .Z(n10179) );
  AND U10009 ( .A(n720), .B(n10189), .Z(n10188) );
  XNOR U10010 ( .A(n10190), .B(n10191), .Z(n10185) );
  AND U10011 ( .A(n712), .B(n10192), .Z(n10191) );
  XOR U10012 ( .A(p_input[1908]), .B(n10190), .Z(n10192) );
  XNOR U10013 ( .A(n10193), .B(n10194), .Z(n10190) );
  AND U10014 ( .A(n716), .B(n10189), .Z(n10194) );
  XNOR U10015 ( .A(n10193), .B(n10187), .Z(n10189) );
  XOR U10016 ( .A(n10195), .B(n10196), .Z(n10187) );
  AND U10017 ( .A(n731), .B(n10197), .Z(n10196) );
  XNOR U10018 ( .A(n10198), .B(n10199), .Z(n10193) );
  AND U10019 ( .A(n723), .B(n10200), .Z(n10199) );
  XOR U10020 ( .A(p_input[1940]), .B(n10198), .Z(n10200) );
  XNOR U10021 ( .A(n10201), .B(n10202), .Z(n10198) );
  AND U10022 ( .A(n727), .B(n10197), .Z(n10202) );
  XNOR U10023 ( .A(n10201), .B(n10195), .Z(n10197) );
  XOR U10024 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n10203), .Z(n10195) );
  AND U10025 ( .A(n741), .B(n10204), .Z(n10203) );
  XNOR U10026 ( .A(n10205), .B(n10206), .Z(n10201) );
  AND U10027 ( .A(n734), .B(n10207), .Z(n10206) );
  XOR U10028 ( .A(p_input[1972]), .B(n10205), .Z(n10207) );
  XNOR U10029 ( .A(n10208), .B(n10209), .Z(n10205) );
  AND U10030 ( .A(n738), .B(n10204), .Z(n10209) );
  XOR U10031 ( .A(n10210), .B(n10208), .Z(n10204) );
  IV U10032 ( .A(\knn_comb_/min_val_out[0][20] ), .Z(n10210) );
  IV U10033 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .Z(n10208)
         );
  XOR U10034 ( .A(n3741), .B(n10211), .Z(o[1]) );
  AND U10035 ( .A(n58), .B(n10212), .Z(n3741) );
  XOR U10036 ( .A(n3742), .B(n10211), .Z(n10212) );
  XOR U10037 ( .A(n10213), .B(n10214), .Z(n10211) );
  AND U10038 ( .A(n70), .B(n10215), .Z(n10214) );
  XOR U10039 ( .A(n10216), .B(n10217), .Z(n3742) );
  AND U10040 ( .A(n62), .B(n10218), .Z(n10217) );
  XOR U10041 ( .A(p_input[1]), .B(n10216), .Z(n10218) );
  XNOR U10042 ( .A(n10219), .B(n10220), .Z(n10216) );
  AND U10043 ( .A(n66), .B(n10215), .Z(n10220) );
  XNOR U10044 ( .A(n10219), .B(n10213), .Z(n10215) );
  XOR U10045 ( .A(n10221), .B(n10222), .Z(n10213) );
  AND U10046 ( .A(n82), .B(n10223), .Z(n10222) );
  XNOR U10047 ( .A(n10224), .B(n10225), .Z(n10219) );
  AND U10048 ( .A(n74), .B(n10226), .Z(n10225) );
  XOR U10049 ( .A(p_input[33]), .B(n10224), .Z(n10226) );
  XNOR U10050 ( .A(n10227), .B(n10228), .Z(n10224) );
  AND U10051 ( .A(n78), .B(n10223), .Z(n10228) );
  XNOR U10052 ( .A(n10227), .B(n10221), .Z(n10223) );
  XOR U10053 ( .A(n10229), .B(n10230), .Z(n10221) );
  AND U10054 ( .A(n93), .B(n10231), .Z(n10230) );
  XNOR U10055 ( .A(n10232), .B(n10233), .Z(n10227) );
  AND U10056 ( .A(n85), .B(n10234), .Z(n10233) );
  XOR U10057 ( .A(p_input[65]), .B(n10232), .Z(n10234) );
  XNOR U10058 ( .A(n10235), .B(n10236), .Z(n10232) );
  AND U10059 ( .A(n89), .B(n10231), .Z(n10236) );
  XNOR U10060 ( .A(n10235), .B(n10229), .Z(n10231) );
  XOR U10061 ( .A(n10237), .B(n10238), .Z(n10229) );
  AND U10062 ( .A(n104), .B(n10239), .Z(n10238) );
  XNOR U10063 ( .A(n10240), .B(n10241), .Z(n10235) );
  AND U10064 ( .A(n96), .B(n10242), .Z(n10241) );
  XOR U10065 ( .A(p_input[97]), .B(n10240), .Z(n10242) );
  XNOR U10066 ( .A(n10243), .B(n10244), .Z(n10240) );
  AND U10067 ( .A(n100), .B(n10239), .Z(n10244) );
  XNOR U10068 ( .A(n10243), .B(n10237), .Z(n10239) );
  XOR U10069 ( .A(n10245), .B(n10246), .Z(n10237) );
  AND U10070 ( .A(n115), .B(n10247), .Z(n10246) );
  XNOR U10071 ( .A(n10248), .B(n10249), .Z(n10243) );
  AND U10072 ( .A(n107), .B(n10250), .Z(n10249) );
  XOR U10073 ( .A(p_input[129]), .B(n10248), .Z(n10250) );
  XNOR U10074 ( .A(n10251), .B(n10252), .Z(n10248) );
  AND U10075 ( .A(n111), .B(n10247), .Z(n10252) );
  XNOR U10076 ( .A(n10251), .B(n10245), .Z(n10247) );
  XOR U10077 ( .A(n10253), .B(n10254), .Z(n10245) );
  AND U10078 ( .A(n126), .B(n10255), .Z(n10254) );
  XNOR U10079 ( .A(n10256), .B(n10257), .Z(n10251) );
  AND U10080 ( .A(n118), .B(n10258), .Z(n10257) );
  XOR U10081 ( .A(p_input[161]), .B(n10256), .Z(n10258) );
  XNOR U10082 ( .A(n10259), .B(n10260), .Z(n10256) );
  AND U10083 ( .A(n122), .B(n10255), .Z(n10260) );
  XNOR U10084 ( .A(n10259), .B(n10253), .Z(n10255) );
  XOR U10085 ( .A(n10261), .B(n10262), .Z(n10253) );
  AND U10086 ( .A(n137), .B(n10263), .Z(n10262) );
  XNOR U10087 ( .A(n10264), .B(n10265), .Z(n10259) );
  AND U10088 ( .A(n129), .B(n10266), .Z(n10265) );
  XOR U10089 ( .A(p_input[193]), .B(n10264), .Z(n10266) );
  XNOR U10090 ( .A(n10267), .B(n10268), .Z(n10264) );
  AND U10091 ( .A(n133), .B(n10263), .Z(n10268) );
  XNOR U10092 ( .A(n10267), .B(n10261), .Z(n10263) );
  XOR U10093 ( .A(n10269), .B(n10270), .Z(n10261) );
  AND U10094 ( .A(n148), .B(n10271), .Z(n10270) );
  XNOR U10095 ( .A(n10272), .B(n10273), .Z(n10267) );
  AND U10096 ( .A(n140), .B(n10274), .Z(n10273) );
  XOR U10097 ( .A(p_input[225]), .B(n10272), .Z(n10274) );
  XNOR U10098 ( .A(n10275), .B(n10276), .Z(n10272) );
  AND U10099 ( .A(n144), .B(n10271), .Z(n10276) );
  XNOR U10100 ( .A(n10275), .B(n10269), .Z(n10271) );
  XOR U10101 ( .A(n10277), .B(n10278), .Z(n10269) );
  AND U10102 ( .A(n159), .B(n10279), .Z(n10278) );
  XNOR U10103 ( .A(n10280), .B(n10281), .Z(n10275) );
  AND U10104 ( .A(n151), .B(n10282), .Z(n10281) );
  XOR U10105 ( .A(p_input[257]), .B(n10280), .Z(n10282) );
  XNOR U10106 ( .A(n10283), .B(n10284), .Z(n10280) );
  AND U10107 ( .A(n155), .B(n10279), .Z(n10284) );
  XNOR U10108 ( .A(n10283), .B(n10277), .Z(n10279) );
  XOR U10109 ( .A(n10285), .B(n10286), .Z(n10277) );
  AND U10110 ( .A(n170), .B(n10287), .Z(n10286) );
  XNOR U10111 ( .A(n10288), .B(n10289), .Z(n10283) );
  AND U10112 ( .A(n162), .B(n10290), .Z(n10289) );
  XOR U10113 ( .A(p_input[289]), .B(n10288), .Z(n10290) );
  XNOR U10114 ( .A(n10291), .B(n10292), .Z(n10288) );
  AND U10115 ( .A(n166), .B(n10287), .Z(n10292) );
  XNOR U10116 ( .A(n10291), .B(n10285), .Z(n10287) );
  XOR U10117 ( .A(n10293), .B(n10294), .Z(n10285) );
  AND U10118 ( .A(n181), .B(n10295), .Z(n10294) );
  XNOR U10119 ( .A(n10296), .B(n10297), .Z(n10291) );
  AND U10120 ( .A(n173), .B(n10298), .Z(n10297) );
  XOR U10121 ( .A(p_input[321]), .B(n10296), .Z(n10298) );
  XNOR U10122 ( .A(n10299), .B(n10300), .Z(n10296) );
  AND U10123 ( .A(n177), .B(n10295), .Z(n10300) );
  XNOR U10124 ( .A(n10299), .B(n10293), .Z(n10295) );
  XOR U10125 ( .A(n10301), .B(n10302), .Z(n10293) );
  AND U10126 ( .A(n192), .B(n10303), .Z(n10302) );
  XNOR U10127 ( .A(n10304), .B(n10305), .Z(n10299) );
  AND U10128 ( .A(n184), .B(n10306), .Z(n10305) );
  XOR U10129 ( .A(p_input[353]), .B(n10304), .Z(n10306) );
  XNOR U10130 ( .A(n10307), .B(n10308), .Z(n10304) );
  AND U10131 ( .A(n188), .B(n10303), .Z(n10308) );
  XNOR U10132 ( .A(n10307), .B(n10301), .Z(n10303) );
  XOR U10133 ( .A(n10309), .B(n10310), .Z(n10301) );
  AND U10134 ( .A(n203), .B(n10311), .Z(n10310) );
  XNOR U10135 ( .A(n10312), .B(n10313), .Z(n10307) );
  AND U10136 ( .A(n195), .B(n10314), .Z(n10313) );
  XOR U10137 ( .A(p_input[385]), .B(n10312), .Z(n10314) );
  XNOR U10138 ( .A(n10315), .B(n10316), .Z(n10312) );
  AND U10139 ( .A(n199), .B(n10311), .Z(n10316) );
  XNOR U10140 ( .A(n10315), .B(n10309), .Z(n10311) );
  XOR U10141 ( .A(n10317), .B(n10318), .Z(n10309) );
  AND U10142 ( .A(n214), .B(n10319), .Z(n10318) );
  XNOR U10143 ( .A(n10320), .B(n10321), .Z(n10315) );
  AND U10144 ( .A(n206), .B(n10322), .Z(n10321) );
  XOR U10145 ( .A(p_input[417]), .B(n10320), .Z(n10322) );
  XNOR U10146 ( .A(n10323), .B(n10324), .Z(n10320) );
  AND U10147 ( .A(n210), .B(n10319), .Z(n10324) );
  XNOR U10148 ( .A(n10323), .B(n10317), .Z(n10319) );
  XOR U10149 ( .A(n10325), .B(n10326), .Z(n10317) );
  AND U10150 ( .A(n225), .B(n10327), .Z(n10326) );
  XNOR U10151 ( .A(n10328), .B(n10329), .Z(n10323) );
  AND U10152 ( .A(n217), .B(n10330), .Z(n10329) );
  XOR U10153 ( .A(p_input[449]), .B(n10328), .Z(n10330) );
  XNOR U10154 ( .A(n10331), .B(n10332), .Z(n10328) );
  AND U10155 ( .A(n221), .B(n10327), .Z(n10332) );
  XNOR U10156 ( .A(n10331), .B(n10325), .Z(n10327) );
  XOR U10157 ( .A(n10333), .B(n10334), .Z(n10325) );
  AND U10158 ( .A(n236), .B(n10335), .Z(n10334) );
  XNOR U10159 ( .A(n10336), .B(n10337), .Z(n10331) );
  AND U10160 ( .A(n228), .B(n10338), .Z(n10337) );
  XOR U10161 ( .A(p_input[481]), .B(n10336), .Z(n10338) );
  XNOR U10162 ( .A(n10339), .B(n10340), .Z(n10336) );
  AND U10163 ( .A(n232), .B(n10335), .Z(n10340) );
  XNOR U10164 ( .A(n10339), .B(n10333), .Z(n10335) );
  XOR U10165 ( .A(n10341), .B(n10342), .Z(n10333) );
  AND U10166 ( .A(n247), .B(n10343), .Z(n10342) );
  XNOR U10167 ( .A(n10344), .B(n10345), .Z(n10339) );
  AND U10168 ( .A(n239), .B(n10346), .Z(n10345) );
  XOR U10169 ( .A(p_input[513]), .B(n10344), .Z(n10346) );
  XNOR U10170 ( .A(n10347), .B(n10348), .Z(n10344) );
  AND U10171 ( .A(n243), .B(n10343), .Z(n10348) );
  XNOR U10172 ( .A(n10347), .B(n10341), .Z(n10343) );
  XOR U10173 ( .A(n10349), .B(n10350), .Z(n10341) );
  AND U10174 ( .A(n258), .B(n10351), .Z(n10350) );
  XNOR U10175 ( .A(n10352), .B(n10353), .Z(n10347) );
  AND U10176 ( .A(n250), .B(n10354), .Z(n10353) );
  XOR U10177 ( .A(p_input[545]), .B(n10352), .Z(n10354) );
  XNOR U10178 ( .A(n10355), .B(n10356), .Z(n10352) );
  AND U10179 ( .A(n254), .B(n10351), .Z(n10356) );
  XNOR U10180 ( .A(n10355), .B(n10349), .Z(n10351) );
  XOR U10181 ( .A(n10357), .B(n10358), .Z(n10349) );
  AND U10182 ( .A(n269), .B(n10359), .Z(n10358) );
  XNOR U10183 ( .A(n10360), .B(n10361), .Z(n10355) );
  AND U10184 ( .A(n261), .B(n10362), .Z(n10361) );
  XOR U10185 ( .A(p_input[577]), .B(n10360), .Z(n10362) );
  XNOR U10186 ( .A(n10363), .B(n10364), .Z(n10360) );
  AND U10187 ( .A(n265), .B(n10359), .Z(n10364) );
  XNOR U10188 ( .A(n10363), .B(n10357), .Z(n10359) );
  XOR U10189 ( .A(n10365), .B(n10366), .Z(n10357) );
  AND U10190 ( .A(n280), .B(n10367), .Z(n10366) );
  XNOR U10191 ( .A(n10368), .B(n10369), .Z(n10363) );
  AND U10192 ( .A(n272), .B(n10370), .Z(n10369) );
  XOR U10193 ( .A(p_input[609]), .B(n10368), .Z(n10370) );
  XNOR U10194 ( .A(n10371), .B(n10372), .Z(n10368) );
  AND U10195 ( .A(n276), .B(n10367), .Z(n10372) );
  XNOR U10196 ( .A(n10371), .B(n10365), .Z(n10367) );
  XOR U10197 ( .A(n10373), .B(n10374), .Z(n10365) );
  AND U10198 ( .A(n291), .B(n10375), .Z(n10374) );
  XNOR U10199 ( .A(n10376), .B(n10377), .Z(n10371) );
  AND U10200 ( .A(n283), .B(n10378), .Z(n10377) );
  XOR U10201 ( .A(p_input[641]), .B(n10376), .Z(n10378) );
  XNOR U10202 ( .A(n10379), .B(n10380), .Z(n10376) );
  AND U10203 ( .A(n287), .B(n10375), .Z(n10380) );
  XNOR U10204 ( .A(n10379), .B(n10373), .Z(n10375) );
  XOR U10205 ( .A(n10381), .B(n10382), .Z(n10373) );
  AND U10206 ( .A(n302), .B(n10383), .Z(n10382) );
  XNOR U10207 ( .A(n10384), .B(n10385), .Z(n10379) );
  AND U10208 ( .A(n294), .B(n10386), .Z(n10385) );
  XOR U10209 ( .A(p_input[673]), .B(n10384), .Z(n10386) );
  XNOR U10210 ( .A(n10387), .B(n10388), .Z(n10384) );
  AND U10211 ( .A(n298), .B(n10383), .Z(n10388) );
  XNOR U10212 ( .A(n10387), .B(n10381), .Z(n10383) );
  XOR U10213 ( .A(n10389), .B(n10390), .Z(n10381) );
  AND U10214 ( .A(n313), .B(n10391), .Z(n10390) );
  XNOR U10215 ( .A(n10392), .B(n10393), .Z(n10387) );
  AND U10216 ( .A(n305), .B(n10394), .Z(n10393) );
  XOR U10217 ( .A(p_input[705]), .B(n10392), .Z(n10394) );
  XNOR U10218 ( .A(n10395), .B(n10396), .Z(n10392) );
  AND U10219 ( .A(n309), .B(n10391), .Z(n10396) );
  XNOR U10220 ( .A(n10395), .B(n10389), .Z(n10391) );
  XOR U10221 ( .A(n10397), .B(n10398), .Z(n10389) );
  AND U10222 ( .A(n324), .B(n10399), .Z(n10398) );
  XNOR U10223 ( .A(n10400), .B(n10401), .Z(n10395) );
  AND U10224 ( .A(n316), .B(n10402), .Z(n10401) );
  XOR U10225 ( .A(p_input[737]), .B(n10400), .Z(n10402) );
  XNOR U10226 ( .A(n10403), .B(n10404), .Z(n10400) );
  AND U10227 ( .A(n320), .B(n10399), .Z(n10404) );
  XNOR U10228 ( .A(n10403), .B(n10397), .Z(n10399) );
  XOR U10229 ( .A(n10405), .B(n10406), .Z(n10397) );
  AND U10230 ( .A(n335), .B(n10407), .Z(n10406) );
  XNOR U10231 ( .A(n10408), .B(n10409), .Z(n10403) );
  AND U10232 ( .A(n327), .B(n10410), .Z(n10409) );
  XOR U10233 ( .A(p_input[769]), .B(n10408), .Z(n10410) );
  XNOR U10234 ( .A(n10411), .B(n10412), .Z(n10408) );
  AND U10235 ( .A(n331), .B(n10407), .Z(n10412) );
  XNOR U10236 ( .A(n10411), .B(n10405), .Z(n10407) );
  XOR U10237 ( .A(n10413), .B(n10414), .Z(n10405) );
  AND U10238 ( .A(n346), .B(n10415), .Z(n10414) );
  XNOR U10239 ( .A(n10416), .B(n10417), .Z(n10411) );
  AND U10240 ( .A(n338), .B(n10418), .Z(n10417) );
  XOR U10241 ( .A(p_input[801]), .B(n10416), .Z(n10418) );
  XNOR U10242 ( .A(n10419), .B(n10420), .Z(n10416) );
  AND U10243 ( .A(n342), .B(n10415), .Z(n10420) );
  XNOR U10244 ( .A(n10419), .B(n10413), .Z(n10415) );
  XOR U10245 ( .A(n10421), .B(n10422), .Z(n10413) );
  AND U10246 ( .A(n357), .B(n10423), .Z(n10422) );
  XNOR U10247 ( .A(n10424), .B(n10425), .Z(n10419) );
  AND U10248 ( .A(n349), .B(n10426), .Z(n10425) );
  XOR U10249 ( .A(p_input[833]), .B(n10424), .Z(n10426) );
  XNOR U10250 ( .A(n10427), .B(n10428), .Z(n10424) );
  AND U10251 ( .A(n353), .B(n10423), .Z(n10428) );
  XNOR U10252 ( .A(n10427), .B(n10421), .Z(n10423) );
  XOR U10253 ( .A(n10429), .B(n10430), .Z(n10421) );
  AND U10254 ( .A(n368), .B(n10431), .Z(n10430) );
  XNOR U10255 ( .A(n10432), .B(n10433), .Z(n10427) );
  AND U10256 ( .A(n360), .B(n10434), .Z(n10433) );
  XOR U10257 ( .A(p_input[865]), .B(n10432), .Z(n10434) );
  XNOR U10258 ( .A(n10435), .B(n10436), .Z(n10432) );
  AND U10259 ( .A(n364), .B(n10431), .Z(n10436) );
  XNOR U10260 ( .A(n10435), .B(n10429), .Z(n10431) );
  XOR U10261 ( .A(n10437), .B(n10438), .Z(n10429) );
  AND U10262 ( .A(n379), .B(n10439), .Z(n10438) );
  XNOR U10263 ( .A(n10440), .B(n10441), .Z(n10435) );
  AND U10264 ( .A(n371), .B(n10442), .Z(n10441) );
  XOR U10265 ( .A(p_input[897]), .B(n10440), .Z(n10442) );
  XNOR U10266 ( .A(n10443), .B(n10444), .Z(n10440) );
  AND U10267 ( .A(n375), .B(n10439), .Z(n10444) );
  XNOR U10268 ( .A(n10443), .B(n10437), .Z(n10439) );
  XOR U10269 ( .A(n10445), .B(n10446), .Z(n10437) );
  AND U10270 ( .A(n390), .B(n10447), .Z(n10446) );
  XNOR U10271 ( .A(n10448), .B(n10449), .Z(n10443) );
  AND U10272 ( .A(n382), .B(n10450), .Z(n10449) );
  XOR U10273 ( .A(p_input[929]), .B(n10448), .Z(n10450) );
  XNOR U10274 ( .A(n10451), .B(n10452), .Z(n10448) );
  AND U10275 ( .A(n386), .B(n10447), .Z(n10452) );
  XNOR U10276 ( .A(n10451), .B(n10445), .Z(n10447) );
  XOR U10277 ( .A(n10453), .B(n10454), .Z(n10445) );
  AND U10278 ( .A(n401), .B(n10455), .Z(n10454) );
  XNOR U10279 ( .A(n10456), .B(n10457), .Z(n10451) );
  AND U10280 ( .A(n393), .B(n10458), .Z(n10457) );
  XOR U10281 ( .A(p_input[961]), .B(n10456), .Z(n10458) );
  XNOR U10282 ( .A(n10459), .B(n10460), .Z(n10456) );
  AND U10283 ( .A(n397), .B(n10455), .Z(n10460) );
  XNOR U10284 ( .A(n10459), .B(n10453), .Z(n10455) );
  XOR U10285 ( .A(n10461), .B(n10462), .Z(n10453) );
  AND U10286 ( .A(n412), .B(n10463), .Z(n10462) );
  XNOR U10287 ( .A(n10464), .B(n10465), .Z(n10459) );
  AND U10288 ( .A(n404), .B(n10466), .Z(n10465) );
  XOR U10289 ( .A(p_input[993]), .B(n10464), .Z(n10466) );
  XNOR U10290 ( .A(n10467), .B(n10468), .Z(n10464) );
  AND U10291 ( .A(n408), .B(n10463), .Z(n10468) );
  XNOR U10292 ( .A(n10467), .B(n10461), .Z(n10463) );
  XOR U10293 ( .A(n10469), .B(n10470), .Z(n10461) );
  AND U10294 ( .A(n423), .B(n10471), .Z(n10470) );
  XNOR U10295 ( .A(n10472), .B(n10473), .Z(n10467) );
  AND U10296 ( .A(n415), .B(n10474), .Z(n10473) );
  XOR U10297 ( .A(p_input[1025]), .B(n10472), .Z(n10474) );
  XNOR U10298 ( .A(n10475), .B(n10476), .Z(n10472) );
  AND U10299 ( .A(n419), .B(n10471), .Z(n10476) );
  XNOR U10300 ( .A(n10475), .B(n10469), .Z(n10471) );
  XOR U10301 ( .A(n10477), .B(n10478), .Z(n10469) );
  AND U10302 ( .A(n434), .B(n10479), .Z(n10478) );
  XNOR U10303 ( .A(n10480), .B(n10481), .Z(n10475) );
  AND U10304 ( .A(n426), .B(n10482), .Z(n10481) );
  XOR U10305 ( .A(p_input[1057]), .B(n10480), .Z(n10482) );
  XNOR U10306 ( .A(n10483), .B(n10484), .Z(n10480) );
  AND U10307 ( .A(n430), .B(n10479), .Z(n10484) );
  XNOR U10308 ( .A(n10483), .B(n10477), .Z(n10479) );
  XOR U10309 ( .A(n10485), .B(n10486), .Z(n10477) );
  AND U10310 ( .A(n445), .B(n10487), .Z(n10486) );
  XNOR U10311 ( .A(n10488), .B(n10489), .Z(n10483) );
  AND U10312 ( .A(n437), .B(n10490), .Z(n10489) );
  XOR U10313 ( .A(p_input[1089]), .B(n10488), .Z(n10490) );
  XNOR U10314 ( .A(n10491), .B(n10492), .Z(n10488) );
  AND U10315 ( .A(n441), .B(n10487), .Z(n10492) );
  XNOR U10316 ( .A(n10491), .B(n10485), .Z(n10487) );
  XOR U10317 ( .A(n10493), .B(n10494), .Z(n10485) );
  AND U10318 ( .A(n456), .B(n10495), .Z(n10494) );
  XNOR U10319 ( .A(n10496), .B(n10497), .Z(n10491) );
  AND U10320 ( .A(n448), .B(n10498), .Z(n10497) );
  XOR U10321 ( .A(p_input[1121]), .B(n10496), .Z(n10498) );
  XNOR U10322 ( .A(n10499), .B(n10500), .Z(n10496) );
  AND U10323 ( .A(n452), .B(n10495), .Z(n10500) );
  XNOR U10324 ( .A(n10499), .B(n10493), .Z(n10495) );
  XOR U10325 ( .A(n10501), .B(n10502), .Z(n10493) );
  AND U10326 ( .A(n467), .B(n10503), .Z(n10502) );
  XNOR U10327 ( .A(n10504), .B(n10505), .Z(n10499) );
  AND U10328 ( .A(n459), .B(n10506), .Z(n10505) );
  XOR U10329 ( .A(p_input[1153]), .B(n10504), .Z(n10506) );
  XNOR U10330 ( .A(n10507), .B(n10508), .Z(n10504) );
  AND U10331 ( .A(n463), .B(n10503), .Z(n10508) );
  XNOR U10332 ( .A(n10507), .B(n10501), .Z(n10503) );
  XOR U10333 ( .A(n10509), .B(n10510), .Z(n10501) );
  AND U10334 ( .A(n478), .B(n10511), .Z(n10510) );
  XNOR U10335 ( .A(n10512), .B(n10513), .Z(n10507) );
  AND U10336 ( .A(n470), .B(n10514), .Z(n10513) );
  XOR U10337 ( .A(p_input[1185]), .B(n10512), .Z(n10514) );
  XNOR U10338 ( .A(n10515), .B(n10516), .Z(n10512) );
  AND U10339 ( .A(n474), .B(n10511), .Z(n10516) );
  XNOR U10340 ( .A(n10515), .B(n10509), .Z(n10511) );
  XOR U10341 ( .A(n10517), .B(n10518), .Z(n10509) );
  AND U10342 ( .A(n489), .B(n10519), .Z(n10518) );
  XNOR U10343 ( .A(n10520), .B(n10521), .Z(n10515) );
  AND U10344 ( .A(n481), .B(n10522), .Z(n10521) );
  XOR U10345 ( .A(p_input[1217]), .B(n10520), .Z(n10522) );
  XNOR U10346 ( .A(n10523), .B(n10524), .Z(n10520) );
  AND U10347 ( .A(n485), .B(n10519), .Z(n10524) );
  XNOR U10348 ( .A(n10523), .B(n10517), .Z(n10519) );
  XOR U10349 ( .A(n10525), .B(n10526), .Z(n10517) );
  AND U10350 ( .A(n500), .B(n10527), .Z(n10526) );
  XNOR U10351 ( .A(n10528), .B(n10529), .Z(n10523) );
  AND U10352 ( .A(n492), .B(n10530), .Z(n10529) );
  XOR U10353 ( .A(p_input[1249]), .B(n10528), .Z(n10530) );
  XNOR U10354 ( .A(n10531), .B(n10532), .Z(n10528) );
  AND U10355 ( .A(n496), .B(n10527), .Z(n10532) );
  XNOR U10356 ( .A(n10531), .B(n10525), .Z(n10527) );
  XOR U10357 ( .A(n10533), .B(n10534), .Z(n10525) );
  AND U10358 ( .A(n511), .B(n10535), .Z(n10534) );
  XNOR U10359 ( .A(n10536), .B(n10537), .Z(n10531) );
  AND U10360 ( .A(n503), .B(n10538), .Z(n10537) );
  XOR U10361 ( .A(p_input[1281]), .B(n10536), .Z(n10538) );
  XNOR U10362 ( .A(n10539), .B(n10540), .Z(n10536) );
  AND U10363 ( .A(n507), .B(n10535), .Z(n10540) );
  XNOR U10364 ( .A(n10539), .B(n10533), .Z(n10535) );
  XOR U10365 ( .A(n10541), .B(n10542), .Z(n10533) );
  AND U10366 ( .A(n522), .B(n10543), .Z(n10542) );
  XNOR U10367 ( .A(n10544), .B(n10545), .Z(n10539) );
  AND U10368 ( .A(n514), .B(n10546), .Z(n10545) );
  XOR U10369 ( .A(p_input[1313]), .B(n10544), .Z(n10546) );
  XNOR U10370 ( .A(n10547), .B(n10548), .Z(n10544) );
  AND U10371 ( .A(n518), .B(n10543), .Z(n10548) );
  XNOR U10372 ( .A(n10547), .B(n10541), .Z(n10543) );
  XOR U10373 ( .A(n10549), .B(n10550), .Z(n10541) );
  AND U10374 ( .A(n533), .B(n10551), .Z(n10550) );
  XNOR U10375 ( .A(n10552), .B(n10553), .Z(n10547) );
  AND U10376 ( .A(n525), .B(n10554), .Z(n10553) );
  XOR U10377 ( .A(p_input[1345]), .B(n10552), .Z(n10554) );
  XNOR U10378 ( .A(n10555), .B(n10556), .Z(n10552) );
  AND U10379 ( .A(n529), .B(n10551), .Z(n10556) );
  XNOR U10380 ( .A(n10555), .B(n10549), .Z(n10551) );
  XOR U10381 ( .A(n10557), .B(n10558), .Z(n10549) );
  AND U10382 ( .A(n544), .B(n10559), .Z(n10558) );
  XNOR U10383 ( .A(n10560), .B(n10561), .Z(n10555) );
  AND U10384 ( .A(n536), .B(n10562), .Z(n10561) );
  XOR U10385 ( .A(p_input[1377]), .B(n10560), .Z(n10562) );
  XNOR U10386 ( .A(n10563), .B(n10564), .Z(n10560) );
  AND U10387 ( .A(n540), .B(n10559), .Z(n10564) );
  XNOR U10388 ( .A(n10563), .B(n10557), .Z(n10559) );
  XOR U10389 ( .A(n10565), .B(n10566), .Z(n10557) );
  AND U10390 ( .A(n555), .B(n10567), .Z(n10566) );
  XNOR U10391 ( .A(n10568), .B(n10569), .Z(n10563) );
  AND U10392 ( .A(n547), .B(n10570), .Z(n10569) );
  XOR U10393 ( .A(p_input[1409]), .B(n10568), .Z(n10570) );
  XNOR U10394 ( .A(n10571), .B(n10572), .Z(n10568) );
  AND U10395 ( .A(n551), .B(n10567), .Z(n10572) );
  XNOR U10396 ( .A(n10571), .B(n10565), .Z(n10567) );
  XOR U10397 ( .A(n10573), .B(n10574), .Z(n10565) );
  AND U10398 ( .A(n566), .B(n10575), .Z(n10574) );
  XNOR U10399 ( .A(n10576), .B(n10577), .Z(n10571) );
  AND U10400 ( .A(n558), .B(n10578), .Z(n10577) );
  XOR U10401 ( .A(p_input[1441]), .B(n10576), .Z(n10578) );
  XNOR U10402 ( .A(n10579), .B(n10580), .Z(n10576) );
  AND U10403 ( .A(n562), .B(n10575), .Z(n10580) );
  XNOR U10404 ( .A(n10579), .B(n10573), .Z(n10575) );
  XOR U10405 ( .A(n10581), .B(n10582), .Z(n10573) );
  AND U10406 ( .A(n577), .B(n10583), .Z(n10582) );
  XNOR U10407 ( .A(n10584), .B(n10585), .Z(n10579) );
  AND U10408 ( .A(n569), .B(n10586), .Z(n10585) );
  XOR U10409 ( .A(p_input[1473]), .B(n10584), .Z(n10586) );
  XNOR U10410 ( .A(n10587), .B(n10588), .Z(n10584) );
  AND U10411 ( .A(n573), .B(n10583), .Z(n10588) );
  XNOR U10412 ( .A(n10587), .B(n10581), .Z(n10583) );
  XOR U10413 ( .A(n10589), .B(n10590), .Z(n10581) );
  AND U10414 ( .A(n588), .B(n10591), .Z(n10590) );
  XNOR U10415 ( .A(n10592), .B(n10593), .Z(n10587) );
  AND U10416 ( .A(n580), .B(n10594), .Z(n10593) );
  XOR U10417 ( .A(p_input[1505]), .B(n10592), .Z(n10594) );
  XNOR U10418 ( .A(n10595), .B(n10596), .Z(n10592) );
  AND U10419 ( .A(n584), .B(n10591), .Z(n10596) );
  XNOR U10420 ( .A(n10595), .B(n10589), .Z(n10591) );
  XOR U10421 ( .A(n10597), .B(n10598), .Z(n10589) );
  AND U10422 ( .A(n599), .B(n10599), .Z(n10598) );
  XNOR U10423 ( .A(n10600), .B(n10601), .Z(n10595) );
  AND U10424 ( .A(n591), .B(n10602), .Z(n10601) );
  XOR U10425 ( .A(p_input[1537]), .B(n10600), .Z(n10602) );
  XNOR U10426 ( .A(n10603), .B(n10604), .Z(n10600) );
  AND U10427 ( .A(n595), .B(n10599), .Z(n10604) );
  XNOR U10428 ( .A(n10603), .B(n10597), .Z(n10599) );
  XOR U10429 ( .A(n10605), .B(n10606), .Z(n10597) );
  AND U10430 ( .A(n610), .B(n10607), .Z(n10606) );
  XNOR U10431 ( .A(n10608), .B(n10609), .Z(n10603) );
  AND U10432 ( .A(n602), .B(n10610), .Z(n10609) );
  XOR U10433 ( .A(p_input[1569]), .B(n10608), .Z(n10610) );
  XNOR U10434 ( .A(n10611), .B(n10612), .Z(n10608) );
  AND U10435 ( .A(n606), .B(n10607), .Z(n10612) );
  XNOR U10436 ( .A(n10611), .B(n10605), .Z(n10607) );
  XOR U10437 ( .A(n10613), .B(n10614), .Z(n10605) );
  AND U10438 ( .A(n621), .B(n10615), .Z(n10614) );
  XNOR U10439 ( .A(n10616), .B(n10617), .Z(n10611) );
  AND U10440 ( .A(n613), .B(n10618), .Z(n10617) );
  XOR U10441 ( .A(p_input[1601]), .B(n10616), .Z(n10618) );
  XNOR U10442 ( .A(n10619), .B(n10620), .Z(n10616) );
  AND U10443 ( .A(n617), .B(n10615), .Z(n10620) );
  XNOR U10444 ( .A(n10619), .B(n10613), .Z(n10615) );
  XOR U10445 ( .A(n10621), .B(n10622), .Z(n10613) );
  AND U10446 ( .A(n632), .B(n10623), .Z(n10622) );
  XNOR U10447 ( .A(n10624), .B(n10625), .Z(n10619) );
  AND U10448 ( .A(n624), .B(n10626), .Z(n10625) );
  XOR U10449 ( .A(p_input[1633]), .B(n10624), .Z(n10626) );
  XNOR U10450 ( .A(n10627), .B(n10628), .Z(n10624) );
  AND U10451 ( .A(n628), .B(n10623), .Z(n10628) );
  XNOR U10452 ( .A(n10627), .B(n10621), .Z(n10623) );
  XOR U10453 ( .A(n10629), .B(n10630), .Z(n10621) );
  AND U10454 ( .A(n643), .B(n10631), .Z(n10630) );
  XNOR U10455 ( .A(n10632), .B(n10633), .Z(n10627) );
  AND U10456 ( .A(n635), .B(n10634), .Z(n10633) );
  XOR U10457 ( .A(p_input[1665]), .B(n10632), .Z(n10634) );
  XNOR U10458 ( .A(n10635), .B(n10636), .Z(n10632) );
  AND U10459 ( .A(n639), .B(n10631), .Z(n10636) );
  XNOR U10460 ( .A(n10635), .B(n10629), .Z(n10631) );
  XOR U10461 ( .A(n10637), .B(n10638), .Z(n10629) );
  AND U10462 ( .A(n654), .B(n10639), .Z(n10638) );
  XNOR U10463 ( .A(n10640), .B(n10641), .Z(n10635) );
  AND U10464 ( .A(n646), .B(n10642), .Z(n10641) );
  XOR U10465 ( .A(p_input[1697]), .B(n10640), .Z(n10642) );
  XNOR U10466 ( .A(n10643), .B(n10644), .Z(n10640) );
  AND U10467 ( .A(n650), .B(n10639), .Z(n10644) );
  XNOR U10468 ( .A(n10643), .B(n10637), .Z(n10639) );
  XOR U10469 ( .A(n10645), .B(n10646), .Z(n10637) );
  AND U10470 ( .A(n665), .B(n10647), .Z(n10646) );
  XNOR U10471 ( .A(n10648), .B(n10649), .Z(n10643) );
  AND U10472 ( .A(n657), .B(n10650), .Z(n10649) );
  XOR U10473 ( .A(p_input[1729]), .B(n10648), .Z(n10650) );
  XNOR U10474 ( .A(n10651), .B(n10652), .Z(n10648) );
  AND U10475 ( .A(n661), .B(n10647), .Z(n10652) );
  XNOR U10476 ( .A(n10651), .B(n10645), .Z(n10647) );
  XOR U10477 ( .A(n10653), .B(n10654), .Z(n10645) );
  AND U10478 ( .A(n676), .B(n10655), .Z(n10654) );
  XNOR U10479 ( .A(n10656), .B(n10657), .Z(n10651) );
  AND U10480 ( .A(n668), .B(n10658), .Z(n10657) );
  XOR U10481 ( .A(p_input[1761]), .B(n10656), .Z(n10658) );
  XNOR U10482 ( .A(n10659), .B(n10660), .Z(n10656) );
  AND U10483 ( .A(n672), .B(n10655), .Z(n10660) );
  XNOR U10484 ( .A(n10659), .B(n10653), .Z(n10655) );
  XOR U10485 ( .A(n10661), .B(n10662), .Z(n10653) );
  AND U10486 ( .A(n687), .B(n10663), .Z(n10662) );
  XNOR U10487 ( .A(n10664), .B(n10665), .Z(n10659) );
  AND U10488 ( .A(n679), .B(n10666), .Z(n10665) );
  XOR U10489 ( .A(p_input[1793]), .B(n10664), .Z(n10666) );
  XNOR U10490 ( .A(n10667), .B(n10668), .Z(n10664) );
  AND U10491 ( .A(n683), .B(n10663), .Z(n10668) );
  XNOR U10492 ( .A(n10667), .B(n10661), .Z(n10663) );
  XOR U10493 ( .A(n10669), .B(n10670), .Z(n10661) );
  AND U10494 ( .A(n698), .B(n10671), .Z(n10670) );
  XNOR U10495 ( .A(n10672), .B(n10673), .Z(n10667) );
  AND U10496 ( .A(n690), .B(n10674), .Z(n10673) );
  XOR U10497 ( .A(p_input[1825]), .B(n10672), .Z(n10674) );
  XNOR U10498 ( .A(n10675), .B(n10676), .Z(n10672) );
  AND U10499 ( .A(n694), .B(n10671), .Z(n10676) );
  XNOR U10500 ( .A(n10675), .B(n10669), .Z(n10671) );
  XOR U10501 ( .A(n10677), .B(n10678), .Z(n10669) );
  AND U10502 ( .A(n709), .B(n10679), .Z(n10678) );
  XNOR U10503 ( .A(n10680), .B(n10681), .Z(n10675) );
  AND U10504 ( .A(n701), .B(n10682), .Z(n10681) );
  XOR U10505 ( .A(p_input[1857]), .B(n10680), .Z(n10682) );
  XNOR U10506 ( .A(n10683), .B(n10684), .Z(n10680) );
  AND U10507 ( .A(n705), .B(n10679), .Z(n10684) );
  XNOR U10508 ( .A(n10683), .B(n10677), .Z(n10679) );
  XOR U10509 ( .A(n10685), .B(n10686), .Z(n10677) );
  AND U10510 ( .A(n720), .B(n10687), .Z(n10686) );
  XNOR U10511 ( .A(n10688), .B(n10689), .Z(n10683) );
  AND U10512 ( .A(n712), .B(n10690), .Z(n10689) );
  XOR U10513 ( .A(p_input[1889]), .B(n10688), .Z(n10690) );
  XNOR U10514 ( .A(n10691), .B(n10692), .Z(n10688) );
  AND U10515 ( .A(n716), .B(n10687), .Z(n10692) );
  XNOR U10516 ( .A(n10691), .B(n10685), .Z(n10687) );
  XOR U10517 ( .A(n10693), .B(n10694), .Z(n10685) );
  AND U10518 ( .A(n731), .B(n10695), .Z(n10694) );
  XNOR U10519 ( .A(n10696), .B(n10697), .Z(n10691) );
  AND U10520 ( .A(n723), .B(n10698), .Z(n10697) );
  XOR U10521 ( .A(p_input[1921]), .B(n10696), .Z(n10698) );
  XNOR U10522 ( .A(n10699), .B(n10700), .Z(n10696) );
  AND U10523 ( .A(n727), .B(n10695), .Z(n10700) );
  XNOR U10524 ( .A(n10699), .B(n10693), .Z(n10695) );
  XOR U10525 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n10701), .Z(n10693) );
  AND U10526 ( .A(n741), .B(n10702), .Z(n10701) );
  XNOR U10527 ( .A(n10703), .B(n10704), .Z(n10699) );
  AND U10528 ( .A(n734), .B(n10705), .Z(n10704) );
  XOR U10529 ( .A(p_input[1953]), .B(n10703), .Z(n10705) );
  XNOR U10530 ( .A(n10706), .B(n10707), .Z(n10703) );
  AND U10531 ( .A(n738), .B(n10702), .Z(n10707) );
  XOR U10532 ( .A(\knn_comb_/min_val_out[0][1] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n10702) );
  XOR U10533 ( .A(n35), .B(n10708), .Z(o[19]) );
  AND U10534 ( .A(n58), .B(n10709), .Z(n35) );
  XOR U10535 ( .A(n36), .B(n10708), .Z(n10709) );
  XOR U10536 ( .A(n10710), .B(n10711), .Z(n10708) );
  AND U10537 ( .A(n70), .B(n10712), .Z(n10711) );
  XOR U10538 ( .A(n10713), .B(n10714), .Z(n36) );
  AND U10539 ( .A(n62), .B(n10715), .Z(n10714) );
  XOR U10540 ( .A(p_input[19]), .B(n10713), .Z(n10715) );
  XNOR U10541 ( .A(n10716), .B(n10717), .Z(n10713) );
  AND U10542 ( .A(n66), .B(n10712), .Z(n10717) );
  XNOR U10543 ( .A(n10716), .B(n10710), .Z(n10712) );
  XOR U10544 ( .A(n10718), .B(n10719), .Z(n10710) );
  AND U10545 ( .A(n82), .B(n10720), .Z(n10719) );
  XNOR U10546 ( .A(n10721), .B(n10722), .Z(n10716) );
  AND U10547 ( .A(n74), .B(n10723), .Z(n10722) );
  XOR U10548 ( .A(p_input[51]), .B(n10721), .Z(n10723) );
  XNOR U10549 ( .A(n10724), .B(n10725), .Z(n10721) );
  AND U10550 ( .A(n78), .B(n10720), .Z(n10725) );
  XNOR U10551 ( .A(n10724), .B(n10718), .Z(n10720) );
  XOR U10552 ( .A(n10726), .B(n10727), .Z(n10718) );
  AND U10553 ( .A(n93), .B(n10728), .Z(n10727) );
  XNOR U10554 ( .A(n10729), .B(n10730), .Z(n10724) );
  AND U10555 ( .A(n85), .B(n10731), .Z(n10730) );
  XOR U10556 ( .A(p_input[83]), .B(n10729), .Z(n10731) );
  XNOR U10557 ( .A(n10732), .B(n10733), .Z(n10729) );
  AND U10558 ( .A(n89), .B(n10728), .Z(n10733) );
  XNOR U10559 ( .A(n10732), .B(n10726), .Z(n10728) );
  XOR U10560 ( .A(n10734), .B(n10735), .Z(n10726) );
  AND U10561 ( .A(n104), .B(n10736), .Z(n10735) );
  XNOR U10562 ( .A(n10737), .B(n10738), .Z(n10732) );
  AND U10563 ( .A(n96), .B(n10739), .Z(n10738) );
  XOR U10564 ( .A(p_input[115]), .B(n10737), .Z(n10739) );
  XNOR U10565 ( .A(n10740), .B(n10741), .Z(n10737) );
  AND U10566 ( .A(n100), .B(n10736), .Z(n10741) );
  XNOR U10567 ( .A(n10740), .B(n10734), .Z(n10736) );
  XOR U10568 ( .A(n10742), .B(n10743), .Z(n10734) );
  AND U10569 ( .A(n115), .B(n10744), .Z(n10743) );
  XNOR U10570 ( .A(n10745), .B(n10746), .Z(n10740) );
  AND U10571 ( .A(n107), .B(n10747), .Z(n10746) );
  XOR U10572 ( .A(p_input[147]), .B(n10745), .Z(n10747) );
  XNOR U10573 ( .A(n10748), .B(n10749), .Z(n10745) );
  AND U10574 ( .A(n111), .B(n10744), .Z(n10749) );
  XNOR U10575 ( .A(n10748), .B(n10742), .Z(n10744) );
  XOR U10576 ( .A(n10750), .B(n10751), .Z(n10742) );
  AND U10577 ( .A(n126), .B(n10752), .Z(n10751) );
  XNOR U10578 ( .A(n10753), .B(n10754), .Z(n10748) );
  AND U10579 ( .A(n118), .B(n10755), .Z(n10754) );
  XOR U10580 ( .A(p_input[179]), .B(n10753), .Z(n10755) );
  XNOR U10581 ( .A(n10756), .B(n10757), .Z(n10753) );
  AND U10582 ( .A(n122), .B(n10752), .Z(n10757) );
  XNOR U10583 ( .A(n10756), .B(n10750), .Z(n10752) );
  XOR U10584 ( .A(n10758), .B(n10759), .Z(n10750) );
  AND U10585 ( .A(n137), .B(n10760), .Z(n10759) );
  XNOR U10586 ( .A(n10761), .B(n10762), .Z(n10756) );
  AND U10587 ( .A(n129), .B(n10763), .Z(n10762) );
  XOR U10588 ( .A(p_input[211]), .B(n10761), .Z(n10763) );
  XNOR U10589 ( .A(n10764), .B(n10765), .Z(n10761) );
  AND U10590 ( .A(n133), .B(n10760), .Z(n10765) );
  XNOR U10591 ( .A(n10764), .B(n10758), .Z(n10760) );
  XOR U10592 ( .A(n10766), .B(n10767), .Z(n10758) );
  AND U10593 ( .A(n148), .B(n10768), .Z(n10767) );
  XNOR U10594 ( .A(n10769), .B(n10770), .Z(n10764) );
  AND U10595 ( .A(n140), .B(n10771), .Z(n10770) );
  XOR U10596 ( .A(p_input[243]), .B(n10769), .Z(n10771) );
  XNOR U10597 ( .A(n10772), .B(n10773), .Z(n10769) );
  AND U10598 ( .A(n144), .B(n10768), .Z(n10773) );
  XNOR U10599 ( .A(n10772), .B(n10766), .Z(n10768) );
  XOR U10600 ( .A(n10774), .B(n10775), .Z(n10766) );
  AND U10601 ( .A(n159), .B(n10776), .Z(n10775) );
  XNOR U10602 ( .A(n10777), .B(n10778), .Z(n10772) );
  AND U10603 ( .A(n151), .B(n10779), .Z(n10778) );
  XOR U10604 ( .A(p_input[275]), .B(n10777), .Z(n10779) );
  XNOR U10605 ( .A(n10780), .B(n10781), .Z(n10777) );
  AND U10606 ( .A(n155), .B(n10776), .Z(n10781) );
  XNOR U10607 ( .A(n10780), .B(n10774), .Z(n10776) );
  XOR U10608 ( .A(n10782), .B(n10783), .Z(n10774) );
  AND U10609 ( .A(n170), .B(n10784), .Z(n10783) );
  XNOR U10610 ( .A(n10785), .B(n10786), .Z(n10780) );
  AND U10611 ( .A(n162), .B(n10787), .Z(n10786) );
  XOR U10612 ( .A(p_input[307]), .B(n10785), .Z(n10787) );
  XNOR U10613 ( .A(n10788), .B(n10789), .Z(n10785) );
  AND U10614 ( .A(n166), .B(n10784), .Z(n10789) );
  XNOR U10615 ( .A(n10788), .B(n10782), .Z(n10784) );
  XOR U10616 ( .A(n10790), .B(n10791), .Z(n10782) );
  AND U10617 ( .A(n181), .B(n10792), .Z(n10791) );
  XNOR U10618 ( .A(n10793), .B(n10794), .Z(n10788) );
  AND U10619 ( .A(n173), .B(n10795), .Z(n10794) );
  XOR U10620 ( .A(p_input[339]), .B(n10793), .Z(n10795) );
  XNOR U10621 ( .A(n10796), .B(n10797), .Z(n10793) );
  AND U10622 ( .A(n177), .B(n10792), .Z(n10797) );
  XNOR U10623 ( .A(n10796), .B(n10790), .Z(n10792) );
  XOR U10624 ( .A(n10798), .B(n10799), .Z(n10790) );
  AND U10625 ( .A(n192), .B(n10800), .Z(n10799) );
  XNOR U10626 ( .A(n10801), .B(n10802), .Z(n10796) );
  AND U10627 ( .A(n184), .B(n10803), .Z(n10802) );
  XOR U10628 ( .A(p_input[371]), .B(n10801), .Z(n10803) );
  XNOR U10629 ( .A(n10804), .B(n10805), .Z(n10801) );
  AND U10630 ( .A(n188), .B(n10800), .Z(n10805) );
  XNOR U10631 ( .A(n10804), .B(n10798), .Z(n10800) );
  XOR U10632 ( .A(n10806), .B(n10807), .Z(n10798) );
  AND U10633 ( .A(n203), .B(n10808), .Z(n10807) );
  XNOR U10634 ( .A(n10809), .B(n10810), .Z(n10804) );
  AND U10635 ( .A(n195), .B(n10811), .Z(n10810) );
  XOR U10636 ( .A(p_input[403]), .B(n10809), .Z(n10811) );
  XNOR U10637 ( .A(n10812), .B(n10813), .Z(n10809) );
  AND U10638 ( .A(n199), .B(n10808), .Z(n10813) );
  XNOR U10639 ( .A(n10812), .B(n10806), .Z(n10808) );
  XOR U10640 ( .A(n10814), .B(n10815), .Z(n10806) );
  AND U10641 ( .A(n214), .B(n10816), .Z(n10815) );
  XNOR U10642 ( .A(n10817), .B(n10818), .Z(n10812) );
  AND U10643 ( .A(n206), .B(n10819), .Z(n10818) );
  XOR U10644 ( .A(p_input[435]), .B(n10817), .Z(n10819) );
  XNOR U10645 ( .A(n10820), .B(n10821), .Z(n10817) );
  AND U10646 ( .A(n210), .B(n10816), .Z(n10821) );
  XNOR U10647 ( .A(n10820), .B(n10814), .Z(n10816) );
  XOR U10648 ( .A(n10822), .B(n10823), .Z(n10814) );
  AND U10649 ( .A(n225), .B(n10824), .Z(n10823) );
  XNOR U10650 ( .A(n10825), .B(n10826), .Z(n10820) );
  AND U10651 ( .A(n217), .B(n10827), .Z(n10826) );
  XOR U10652 ( .A(p_input[467]), .B(n10825), .Z(n10827) );
  XNOR U10653 ( .A(n10828), .B(n10829), .Z(n10825) );
  AND U10654 ( .A(n221), .B(n10824), .Z(n10829) );
  XNOR U10655 ( .A(n10828), .B(n10822), .Z(n10824) );
  XOR U10656 ( .A(n10830), .B(n10831), .Z(n10822) );
  AND U10657 ( .A(n236), .B(n10832), .Z(n10831) );
  XNOR U10658 ( .A(n10833), .B(n10834), .Z(n10828) );
  AND U10659 ( .A(n228), .B(n10835), .Z(n10834) );
  XOR U10660 ( .A(p_input[499]), .B(n10833), .Z(n10835) );
  XNOR U10661 ( .A(n10836), .B(n10837), .Z(n10833) );
  AND U10662 ( .A(n232), .B(n10832), .Z(n10837) );
  XNOR U10663 ( .A(n10836), .B(n10830), .Z(n10832) );
  XOR U10664 ( .A(n10838), .B(n10839), .Z(n10830) );
  AND U10665 ( .A(n247), .B(n10840), .Z(n10839) );
  XNOR U10666 ( .A(n10841), .B(n10842), .Z(n10836) );
  AND U10667 ( .A(n239), .B(n10843), .Z(n10842) );
  XOR U10668 ( .A(p_input[531]), .B(n10841), .Z(n10843) );
  XNOR U10669 ( .A(n10844), .B(n10845), .Z(n10841) );
  AND U10670 ( .A(n243), .B(n10840), .Z(n10845) );
  XNOR U10671 ( .A(n10844), .B(n10838), .Z(n10840) );
  XOR U10672 ( .A(n10846), .B(n10847), .Z(n10838) );
  AND U10673 ( .A(n258), .B(n10848), .Z(n10847) );
  XNOR U10674 ( .A(n10849), .B(n10850), .Z(n10844) );
  AND U10675 ( .A(n250), .B(n10851), .Z(n10850) );
  XOR U10676 ( .A(p_input[563]), .B(n10849), .Z(n10851) );
  XNOR U10677 ( .A(n10852), .B(n10853), .Z(n10849) );
  AND U10678 ( .A(n254), .B(n10848), .Z(n10853) );
  XNOR U10679 ( .A(n10852), .B(n10846), .Z(n10848) );
  XOR U10680 ( .A(n10854), .B(n10855), .Z(n10846) );
  AND U10681 ( .A(n269), .B(n10856), .Z(n10855) );
  XNOR U10682 ( .A(n10857), .B(n10858), .Z(n10852) );
  AND U10683 ( .A(n261), .B(n10859), .Z(n10858) );
  XOR U10684 ( .A(p_input[595]), .B(n10857), .Z(n10859) );
  XNOR U10685 ( .A(n10860), .B(n10861), .Z(n10857) );
  AND U10686 ( .A(n265), .B(n10856), .Z(n10861) );
  XNOR U10687 ( .A(n10860), .B(n10854), .Z(n10856) );
  XOR U10688 ( .A(n10862), .B(n10863), .Z(n10854) );
  AND U10689 ( .A(n280), .B(n10864), .Z(n10863) );
  XNOR U10690 ( .A(n10865), .B(n10866), .Z(n10860) );
  AND U10691 ( .A(n272), .B(n10867), .Z(n10866) );
  XOR U10692 ( .A(p_input[627]), .B(n10865), .Z(n10867) );
  XNOR U10693 ( .A(n10868), .B(n10869), .Z(n10865) );
  AND U10694 ( .A(n276), .B(n10864), .Z(n10869) );
  XNOR U10695 ( .A(n10868), .B(n10862), .Z(n10864) );
  XOR U10696 ( .A(n10870), .B(n10871), .Z(n10862) );
  AND U10697 ( .A(n291), .B(n10872), .Z(n10871) );
  XNOR U10698 ( .A(n10873), .B(n10874), .Z(n10868) );
  AND U10699 ( .A(n283), .B(n10875), .Z(n10874) );
  XOR U10700 ( .A(p_input[659]), .B(n10873), .Z(n10875) );
  XNOR U10701 ( .A(n10876), .B(n10877), .Z(n10873) );
  AND U10702 ( .A(n287), .B(n10872), .Z(n10877) );
  XNOR U10703 ( .A(n10876), .B(n10870), .Z(n10872) );
  XOR U10704 ( .A(n10878), .B(n10879), .Z(n10870) );
  AND U10705 ( .A(n302), .B(n10880), .Z(n10879) );
  XNOR U10706 ( .A(n10881), .B(n10882), .Z(n10876) );
  AND U10707 ( .A(n294), .B(n10883), .Z(n10882) );
  XOR U10708 ( .A(p_input[691]), .B(n10881), .Z(n10883) );
  XNOR U10709 ( .A(n10884), .B(n10885), .Z(n10881) );
  AND U10710 ( .A(n298), .B(n10880), .Z(n10885) );
  XNOR U10711 ( .A(n10884), .B(n10878), .Z(n10880) );
  XOR U10712 ( .A(n10886), .B(n10887), .Z(n10878) );
  AND U10713 ( .A(n313), .B(n10888), .Z(n10887) );
  XNOR U10714 ( .A(n10889), .B(n10890), .Z(n10884) );
  AND U10715 ( .A(n305), .B(n10891), .Z(n10890) );
  XOR U10716 ( .A(p_input[723]), .B(n10889), .Z(n10891) );
  XNOR U10717 ( .A(n10892), .B(n10893), .Z(n10889) );
  AND U10718 ( .A(n309), .B(n10888), .Z(n10893) );
  XNOR U10719 ( .A(n10892), .B(n10886), .Z(n10888) );
  XOR U10720 ( .A(n10894), .B(n10895), .Z(n10886) );
  AND U10721 ( .A(n324), .B(n10896), .Z(n10895) );
  XNOR U10722 ( .A(n10897), .B(n10898), .Z(n10892) );
  AND U10723 ( .A(n316), .B(n10899), .Z(n10898) );
  XOR U10724 ( .A(p_input[755]), .B(n10897), .Z(n10899) );
  XNOR U10725 ( .A(n10900), .B(n10901), .Z(n10897) );
  AND U10726 ( .A(n320), .B(n10896), .Z(n10901) );
  XNOR U10727 ( .A(n10900), .B(n10894), .Z(n10896) );
  XOR U10728 ( .A(n10902), .B(n10903), .Z(n10894) );
  AND U10729 ( .A(n335), .B(n10904), .Z(n10903) );
  XNOR U10730 ( .A(n10905), .B(n10906), .Z(n10900) );
  AND U10731 ( .A(n327), .B(n10907), .Z(n10906) );
  XOR U10732 ( .A(p_input[787]), .B(n10905), .Z(n10907) );
  XNOR U10733 ( .A(n10908), .B(n10909), .Z(n10905) );
  AND U10734 ( .A(n331), .B(n10904), .Z(n10909) );
  XNOR U10735 ( .A(n10908), .B(n10902), .Z(n10904) );
  XOR U10736 ( .A(n10910), .B(n10911), .Z(n10902) );
  AND U10737 ( .A(n346), .B(n10912), .Z(n10911) );
  XNOR U10738 ( .A(n10913), .B(n10914), .Z(n10908) );
  AND U10739 ( .A(n338), .B(n10915), .Z(n10914) );
  XOR U10740 ( .A(p_input[819]), .B(n10913), .Z(n10915) );
  XNOR U10741 ( .A(n10916), .B(n10917), .Z(n10913) );
  AND U10742 ( .A(n342), .B(n10912), .Z(n10917) );
  XNOR U10743 ( .A(n10916), .B(n10910), .Z(n10912) );
  XOR U10744 ( .A(n10918), .B(n10919), .Z(n10910) );
  AND U10745 ( .A(n357), .B(n10920), .Z(n10919) );
  XNOR U10746 ( .A(n10921), .B(n10922), .Z(n10916) );
  AND U10747 ( .A(n349), .B(n10923), .Z(n10922) );
  XOR U10748 ( .A(p_input[851]), .B(n10921), .Z(n10923) );
  XNOR U10749 ( .A(n10924), .B(n10925), .Z(n10921) );
  AND U10750 ( .A(n353), .B(n10920), .Z(n10925) );
  XNOR U10751 ( .A(n10924), .B(n10918), .Z(n10920) );
  XOR U10752 ( .A(n10926), .B(n10927), .Z(n10918) );
  AND U10753 ( .A(n368), .B(n10928), .Z(n10927) );
  XNOR U10754 ( .A(n10929), .B(n10930), .Z(n10924) );
  AND U10755 ( .A(n360), .B(n10931), .Z(n10930) );
  XOR U10756 ( .A(p_input[883]), .B(n10929), .Z(n10931) );
  XNOR U10757 ( .A(n10932), .B(n10933), .Z(n10929) );
  AND U10758 ( .A(n364), .B(n10928), .Z(n10933) );
  XNOR U10759 ( .A(n10932), .B(n10926), .Z(n10928) );
  XOR U10760 ( .A(n10934), .B(n10935), .Z(n10926) );
  AND U10761 ( .A(n379), .B(n10936), .Z(n10935) );
  XNOR U10762 ( .A(n10937), .B(n10938), .Z(n10932) );
  AND U10763 ( .A(n371), .B(n10939), .Z(n10938) );
  XOR U10764 ( .A(p_input[915]), .B(n10937), .Z(n10939) );
  XNOR U10765 ( .A(n10940), .B(n10941), .Z(n10937) );
  AND U10766 ( .A(n375), .B(n10936), .Z(n10941) );
  XNOR U10767 ( .A(n10940), .B(n10934), .Z(n10936) );
  XOR U10768 ( .A(n10942), .B(n10943), .Z(n10934) );
  AND U10769 ( .A(n390), .B(n10944), .Z(n10943) );
  XNOR U10770 ( .A(n10945), .B(n10946), .Z(n10940) );
  AND U10771 ( .A(n382), .B(n10947), .Z(n10946) );
  XOR U10772 ( .A(p_input[947]), .B(n10945), .Z(n10947) );
  XNOR U10773 ( .A(n10948), .B(n10949), .Z(n10945) );
  AND U10774 ( .A(n386), .B(n10944), .Z(n10949) );
  XNOR U10775 ( .A(n10948), .B(n10942), .Z(n10944) );
  XOR U10776 ( .A(n10950), .B(n10951), .Z(n10942) );
  AND U10777 ( .A(n401), .B(n10952), .Z(n10951) );
  XNOR U10778 ( .A(n10953), .B(n10954), .Z(n10948) );
  AND U10779 ( .A(n393), .B(n10955), .Z(n10954) );
  XOR U10780 ( .A(p_input[979]), .B(n10953), .Z(n10955) );
  XNOR U10781 ( .A(n10956), .B(n10957), .Z(n10953) );
  AND U10782 ( .A(n397), .B(n10952), .Z(n10957) );
  XNOR U10783 ( .A(n10956), .B(n10950), .Z(n10952) );
  XOR U10784 ( .A(n10958), .B(n10959), .Z(n10950) );
  AND U10785 ( .A(n412), .B(n10960), .Z(n10959) );
  XNOR U10786 ( .A(n10961), .B(n10962), .Z(n10956) );
  AND U10787 ( .A(n404), .B(n10963), .Z(n10962) );
  XOR U10788 ( .A(p_input[1011]), .B(n10961), .Z(n10963) );
  XNOR U10789 ( .A(n10964), .B(n10965), .Z(n10961) );
  AND U10790 ( .A(n408), .B(n10960), .Z(n10965) );
  XNOR U10791 ( .A(n10964), .B(n10958), .Z(n10960) );
  XOR U10792 ( .A(n10966), .B(n10967), .Z(n10958) );
  AND U10793 ( .A(n423), .B(n10968), .Z(n10967) );
  XNOR U10794 ( .A(n10969), .B(n10970), .Z(n10964) );
  AND U10795 ( .A(n415), .B(n10971), .Z(n10970) );
  XOR U10796 ( .A(p_input[1043]), .B(n10969), .Z(n10971) );
  XNOR U10797 ( .A(n10972), .B(n10973), .Z(n10969) );
  AND U10798 ( .A(n419), .B(n10968), .Z(n10973) );
  XNOR U10799 ( .A(n10972), .B(n10966), .Z(n10968) );
  XOR U10800 ( .A(n10974), .B(n10975), .Z(n10966) );
  AND U10801 ( .A(n434), .B(n10976), .Z(n10975) );
  XNOR U10802 ( .A(n10977), .B(n10978), .Z(n10972) );
  AND U10803 ( .A(n426), .B(n10979), .Z(n10978) );
  XOR U10804 ( .A(p_input[1075]), .B(n10977), .Z(n10979) );
  XNOR U10805 ( .A(n10980), .B(n10981), .Z(n10977) );
  AND U10806 ( .A(n430), .B(n10976), .Z(n10981) );
  XNOR U10807 ( .A(n10980), .B(n10974), .Z(n10976) );
  XOR U10808 ( .A(n10982), .B(n10983), .Z(n10974) );
  AND U10809 ( .A(n445), .B(n10984), .Z(n10983) );
  XNOR U10810 ( .A(n10985), .B(n10986), .Z(n10980) );
  AND U10811 ( .A(n437), .B(n10987), .Z(n10986) );
  XOR U10812 ( .A(p_input[1107]), .B(n10985), .Z(n10987) );
  XNOR U10813 ( .A(n10988), .B(n10989), .Z(n10985) );
  AND U10814 ( .A(n441), .B(n10984), .Z(n10989) );
  XNOR U10815 ( .A(n10988), .B(n10982), .Z(n10984) );
  XOR U10816 ( .A(n10990), .B(n10991), .Z(n10982) );
  AND U10817 ( .A(n456), .B(n10992), .Z(n10991) );
  XNOR U10818 ( .A(n10993), .B(n10994), .Z(n10988) );
  AND U10819 ( .A(n448), .B(n10995), .Z(n10994) );
  XOR U10820 ( .A(p_input[1139]), .B(n10993), .Z(n10995) );
  XNOR U10821 ( .A(n10996), .B(n10997), .Z(n10993) );
  AND U10822 ( .A(n452), .B(n10992), .Z(n10997) );
  XNOR U10823 ( .A(n10996), .B(n10990), .Z(n10992) );
  XOR U10824 ( .A(n10998), .B(n10999), .Z(n10990) );
  AND U10825 ( .A(n467), .B(n11000), .Z(n10999) );
  XNOR U10826 ( .A(n11001), .B(n11002), .Z(n10996) );
  AND U10827 ( .A(n459), .B(n11003), .Z(n11002) );
  XOR U10828 ( .A(p_input[1171]), .B(n11001), .Z(n11003) );
  XNOR U10829 ( .A(n11004), .B(n11005), .Z(n11001) );
  AND U10830 ( .A(n463), .B(n11000), .Z(n11005) );
  XNOR U10831 ( .A(n11004), .B(n10998), .Z(n11000) );
  XOR U10832 ( .A(n11006), .B(n11007), .Z(n10998) );
  AND U10833 ( .A(n478), .B(n11008), .Z(n11007) );
  XNOR U10834 ( .A(n11009), .B(n11010), .Z(n11004) );
  AND U10835 ( .A(n470), .B(n11011), .Z(n11010) );
  XOR U10836 ( .A(p_input[1203]), .B(n11009), .Z(n11011) );
  XNOR U10837 ( .A(n11012), .B(n11013), .Z(n11009) );
  AND U10838 ( .A(n474), .B(n11008), .Z(n11013) );
  XNOR U10839 ( .A(n11012), .B(n11006), .Z(n11008) );
  XOR U10840 ( .A(n11014), .B(n11015), .Z(n11006) );
  AND U10841 ( .A(n489), .B(n11016), .Z(n11015) );
  XNOR U10842 ( .A(n11017), .B(n11018), .Z(n11012) );
  AND U10843 ( .A(n481), .B(n11019), .Z(n11018) );
  XOR U10844 ( .A(p_input[1235]), .B(n11017), .Z(n11019) );
  XNOR U10845 ( .A(n11020), .B(n11021), .Z(n11017) );
  AND U10846 ( .A(n485), .B(n11016), .Z(n11021) );
  XNOR U10847 ( .A(n11020), .B(n11014), .Z(n11016) );
  XOR U10848 ( .A(n11022), .B(n11023), .Z(n11014) );
  AND U10849 ( .A(n500), .B(n11024), .Z(n11023) );
  XNOR U10850 ( .A(n11025), .B(n11026), .Z(n11020) );
  AND U10851 ( .A(n492), .B(n11027), .Z(n11026) );
  XOR U10852 ( .A(p_input[1267]), .B(n11025), .Z(n11027) );
  XNOR U10853 ( .A(n11028), .B(n11029), .Z(n11025) );
  AND U10854 ( .A(n496), .B(n11024), .Z(n11029) );
  XNOR U10855 ( .A(n11028), .B(n11022), .Z(n11024) );
  XOR U10856 ( .A(n11030), .B(n11031), .Z(n11022) );
  AND U10857 ( .A(n511), .B(n11032), .Z(n11031) );
  XNOR U10858 ( .A(n11033), .B(n11034), .Z(n11028) );
  AND U10859 ( .A(n503), .B(n11035), .Z(n11034) );
  XOR U10860 ( .A(p_input[1299]), .B(n11033), .Z(n11035) );
  XNOR U10861 ( .A(n11036), .B(n11037), .Z(n11033) );
  AND U10862 ( .A(n507), .B(n11032), .Z(n11037) );
  XNOR U10863 ( .A(n11036), .B(n11030), .Z(n11032) );
  XOR U10864 ( .A(n11038), .B(n11039), .Z(n11030) );
  AND U10865 ( .A(n522), .B(n11040), .Z(n11039) );
  XNOR U10866 ( .A(n11041), .B(n11042), .Z(n11036) );
  AND U10867 ( .A(n514), .B(n11043), .Z(n11042) );
  XOR U10868 ( .A(p_input[1331]), .B(n11041), .Z(n11043) );
  XNOR U10869 ( .A(n11044), .B(n11045), .Z(n11041) );
  AND U10870 ( .A(n518), .B(n11040), .Z(n11045) );
  XNOR U10871 ( .A(n11044), .B(n11038), .Z(n11040) );
  XOR U10872 ( .A(n11046), .B(n11047), .Z(n11038) );
  AND U10873 ( .A(n533), .B(n11048), .Z(n11047) );
  XNOR U10874 ( .A(n11049), .B(n11050), .Z(n11044) );
  AND U10875 ( .A(n525), .B(n11051), .Z(n11050) );
  XOR U10876 ( .A(p_input[1363]), .B(n11049), .Z(n11051) );
  XNOR U10877 ( .A(n11052), .B(n11053), .Z(n11049) );
  AND U10878 ( .A(n529), .B(n11048), .Z(n11053) );
  XNOR U10879 ( .A(n11052), .B(n11046), .Z(n11048) );
  XOR U10880 ( .A(n11054), .B(n11055), .Z(n11046) );
  AND U10881 ( .A(n544), .B(n11056), .Z(n11055) );
  XNOR U10882 ( .A(n11057), .B(n11058), .Z(n11052) );
  AND U10883 ( .A(n536), .B(n11059), .Z(n11058) );
  XOR U10884 ( .A(p_input[1395]), .B(n11057), .Z(n11059) );
  XNOR U10885 ( .A(n11060), .B(n11061), .Z(n11057) );
  AND U10886 ( .A(n540), .B(n11056), .Z(n11061) );
  XNOR U10887 ( .A(n11060), .B(n11054), .Z(n11056) );
  XOR U10888 ( .A(n11062), .B(n11063), .Z(n11054) );
  AND U10889 ( .A(n555), .B(n11064), .Z(n11063) );
  XNOR U10890 ( .A(n11065), .B(n11066), .Z(n11060) );
  AND U10891 ( .A(n547), .B(n11067), .Z(n11066) );
  XOR U10892 ( .A(p_input[1427]), .B(n11065), .Z(n11067) );
  XNOR U10893 ( .A(n11068), .B(n11069), .Z(n11065) );
  AND U10894 ( .A(n551), .B(n11064), .Z(n11069) );
  XNOR U10895 ( .A(n11068), .B(n11062), .Z(n11064) );
  XOR U10896 ( .A(n11070), .B(n11071), .Z(n11062) );
  AND U10897 ( .A(n566), .B(n11072), .Z(n11071) );
  XNOR U10898 ( .A(n11073), .B(n11074), .Z(n11068) );
  AND U10899 ( .A(n558), .B(n11075), .Z(n11074) );
  XOR U10900 ( .A(p_input[1459]), .B(n11073), .Z(n11075) );
  XNOR U10901 ( .A(n11076), .B(n11077), .Z(n11073) );
  AND U10902 ( .A(n562), .B(n11072), .Z(n11077) );
  XNOR U10903 ( .A(n11076), .B(n11070), .Z(n11072) );
  XOR U10904 ( .A(n11078), .B(n11079), .Z(n11070) );
  AND U10905 ( .A(n577), .B(n11080), .Z(n11079) );
  XNOR U10906 ( .A(n11081), .B(n11082), .Z(n11076) );
  AND U10907 ( .A(n569), .B(n11083), .Z(n11082) );
  XOR U10908 ( .A(p_input[1491]), .B(n11081), .Z(n11083) );
  XNOR U10909 ( .A(n11084), .B(n11085), .Z(n11081) );
  AND U10910 ( .A(n573), .B(n11080), .Z(n11085) );
  XNOR U10911 ( .A(n11084), .B(n11078), .Z(n11080) );
  XOR U10912 ( .A(n11086), .B(n11087), .Z(n11078) );
  AND U10913 ( .A(n588), .B(n11088), .Z(n11087) );
  XNOR U10914 ( .A(n11089), .B(n11090), .Z(n11084) );
  AND U10915 ( .A(n580), .B(n11091), .Z(n11090) );
  XOR U10916 ( .A(p_input[1523]), .B(n11089), .Z(n11091) );
  XNOR U10917 ( .A(n11092), .B(n11093), .Z(n11089) );
  AND U10918 ( .A(n584), .B(n11088), .Z(n11093) );
  XNOR U10919 ( .A(n11092), .B(n11086), .Z(n11088) );
  XOR U10920 ( .A(n11094), .B(n11095), .Z(n11086) );
  AND U10921 ( .A(n599), .B(n11096), .Z(n11095) );
  XNOR U10922 ( .A(n11097), .B(n11098), .Z(n11092) );
  AND U10923 ( .A(n591), .B(n11099), .Z(n11098) );
  XOR U10924 ( .A(p_input[1555]), .B(n11097), .Z(n11099) );
  XNOR U10925 ( .A(n11100), .B(n11101), .Z(n11097) );
  AND U10926 ( .A(n595), .B(n11096), .Z(n11101) );
  XNOR U10927 ( .A(n11100), .B(n11094), .Z(n11096) );
  XOR U10928 ( .A(n11102), .B(n11103), .Z(n11094) );
  AND U10929 ( .A(n610), .B(n11104), .Z(n11103) );
  XNOR U10930 ( .A(n11105), .B(n11106), .Z(n11100) );
  AND U10931 ( .A(n602), .B(n11107), .Z(n11106) );
  XOR U10932 ( .A(p_input[1587]), .B(n11105), .Z(n11107) );
  XNOR U10933 ( .A(n11108), .B(n11109), .Z(n11105) );
  AND U10934 ( .A(n606), .B(n11104), .Z(n11109) );
  XNOR U10935 ( .A(n11108), .B(n11102), .Z(n11104) );
  XOR U10936 ( .A(n11110), .B(n11111), .Z(n11102) );
  AND U10937 ( .A(n621), .B(n11112), .Z(n11111) );
  XNOR U10938 ( .A(n11113), .B(n11114), .Z(n11108) );
  AND U10939 ( .A(n613), .B(n11115), .Z(n11114) );
  XOR U10940 ( .A(p_input[1619]), .B(n11113), .Z(n11115) );
  XNOR U10941 ( .A(n11116), .B(n11117), .Z(n11113) );
  AND U10942 ( .A(n617), .B(n11112), .Z(n11117) );
  XNOR U10943 ( .A(n11116), .B(n11110), .Z(n11112) );
  XOR U10944 ( .A(n11118), .B(n11119), .Z(n11110) );
  AND U10945 ( .A(n632), .B(n11120), .Z(n11119) );
  XNOR U10946 ( .A(n11121), .B(n11122), .Z(n11116) );
  AND U10947 ( .A(n624), .B(n11123), .Z(n11122) );
  XOR U10948 ( .A(p_input[1651]), .B(n11121), .Z(n11123) );
  XNOR U10949 ( .A(n11124), .B(n11125), .Z(n11121) );
  AND U10950 ( .A(n628), .B(n11120), .Z(n11125) );
  XNOR U10951 ( .A(n11124), .B(n11118), .Z(n11120) );
  XOR U10952 ( .A(n11126), .B(n11127), .Z(n11118) );
  AND U10953 ( .A(n643), .B(n11128), .Z(n11127) );
  XNOR U10954 ( .A(n11129), .B(n11130), .Z(n11124) );
  AND U10955 ( .A(n635), .B(n11131), .Z(n11130) );
  XOR U10956 ( .A(p_input[1683]), .B(n11129), .Z(n11131) );
  XNOR U10957 ( .A(n11132), .B(n11133), .Z(n11129) );
  AND U10958 ( .A(n639), .B(n11128), .Z(n11133) );
  XNOR U10959 ( .A(n11132), .B(n11126), .Z(n11128) );
  XOR U10960 ( .A(n11134), .B(n11135), .Z(n11126) );
  AND U10961 ( .A(n654), .B(n11136), .Z(n11135) );
  XNOR U10962 ( .A(n11137), .B(n11138), .Z(n11132) );
  AND U10963 ( .A(n646), .B(n11139), .Z(n11138) );
  XOR U10964 ( .A(p_input[1715]), .B(n11137), .Z(n11139) );
  XNOR U10965 ( .A(n11140), .B(n11141), .Z(n11137) );
  AND U10966 ( .A(n650), .B(n11136), .Z(n11141) );
  XNOR U10967 ( .A(n11140), .B(n11134), .Z(n11136) );
  XOR U10968 ( .A(n11142), .B(n11143), .Z(n11134) );
  AND U10969 ( .A(n665), .B(n11144), .Z(n11143) );
  XNOR U10970 ( .A(n11145), .B(n11146), .Z(n11140) );
  AND U10971 ( .A(n657), .B(n11147), .Z(n11146) );
  XOR U10972 ( .A(p_input[1747]), .B(n11145), .Z(n11147) );
  XNOR U10973 ( .A(n11148), .B(n11149), .Z(n11145) );
  AND U10974 ( .A(n661), .B(n11144), .Z(n11149) );
  XNOR U10975 ( .A(n11148), .B(n11142), .Z(n11144) );
  XOR U10976 ( .A(n11150), .B(n11151), .Z(n11142) );
  AND U10977 ( .A(n676), .B(n11152), .Z(n11151) );
  XNOR U10978 ( .A(n11153), .B(n11154), .Z(n11148) );
  AND U10979 ( .A(n668), .B(n11155), .Z(n11154) );
  XOR U10980 ( .A(p_input[1779]), .B(n11153), .Z(n11155) );
  XNOR U10981 ( .A(n11156), .B(n11157), .Z(n11153) );
  AND U10982 ( .A(n672), .B(n11152), .Z(n11157) );
  XNOR U10983 ( .A(n11156), .B(n11150), .Z(n11152) );
  XOR U10984 ( .A(n11158), .B(n11159), .Z(n11150) );
  AND U10985 ( .A(n687), .B(n11160), .Z(n11159) );
  XNOR U10986 ( .A(n11161), .B(n11162), .Z(n11156) );
  AND U10987 ( .A(n679), .B(n11163), .Z(n11162) );
  XOR U10988 ( .A(p_input[1811]), .B(n11161), .Z(n11163) );
  XNOR U10989 ( .A(n11164), .B(n11165), .Z(n11161) );
  AND U10990 ( .A(n683), .B(n11160), .Z(n11165) );
  XNOR U10991 ( .A(n11164), .B(n11158), .Z(n11160) );
  XOR U10992 ( .A(n11166), .B(n11167), .Z(n11158) );
  AND U10993 ( .A(n698), .B(n11168), .Z(n11167) );
  XNOR U10994 ( .A(n11169), .B(n11170), .Z(n11164) );
  AND U10995 ( .A(n690), .B(n11171), .Z(n11170) );
  XOR U10996 ( .A(p_input[1843]), .B(n11169), .Z(n11171) );
  XNOR U10997 ( .A(n11172), .B(n11173), .Z(n11169) );
  AND U10998 ( .A(n694), .B(n11168), .Z(n11173) );
  XNOR U10999 ( .A(n11172), .B(n11166), .Z(n11168) );
  XOR U11000 ( .A(n11174), .B(n11175), .Z(n11166) );
  AND U11001 ( .A(n709), .B(n11176), .Z(n11175) );
  XNOR U11002 ( .A(n11177), .B(n11178), .Z(n11172) );
  AND U11003 ( .A(n701), .B(n11179), .Z(n11178) );
  XOR U11004 ( .A(p_input[1875]), .B(n11177), .Z(n11179) );
  XNOR U11005 ( .A(n11180), .B(n11181), .Z(n11177) );
  AND U11006 ( .A(n705), .B(n11176), .Z(n11181) );
  XNOR U11007 ( .A(n11180), .B(n11174), .Z(n11176) );
  XOR U11008 ( .A(n11182), .B(n11183), .Z(n11174) );
  AND U11009 ( .A(n720), .B(n11184), .Z(n11183) );
  XNOR U11010 ( .A(n11185), .B(n11186), .Z(n11180) );
  AND U11011 ( .A(n712), .B(n11187), .Z(n11186) );
  XOR U11012 ( .A(p_input[1907]), .B(n11185), .Z(n11187) );
  XNOR U11013 ( .A(n11188), .B(n11189), .Z(n11185) );
  AND U11014 ( .A(n716), .B(n11184), .Z(n11189) );
  XNOR U11015 ( .A(n11188), .B(n11182), .Z(n11184) );
  XOR U11016 ( .A(n11190), .B(n11191), .Z(n11182) );
  AND U11017 ( .A(n731), .B(n11192), .Z(n11191) );
  XNOR U11018 ( .A(n11193), .B(n11194), .Z(n11188) );
  AND U11019 ( .A(n723), .B(n11195), .Z(n11194) );
  XOR U11020 ( .A(p_input[1939]), .B(n11193), .Z(n11195) );
  XNOR U11021 ( .A(n11196), .B(n11197), .Z(n11193) );
  AND U11022 ( .A(n727), .B(n11192), .Z(n11197) );
  XNOR U11023 ( .A(n11196), .B(n11190), .Z(n11192) );
  XOR U11024 ( .A(\knn_comb_/min_val_out[0][19] ), .B(n11198), .Z(n11190) );
  AND U11025 ( .A(n741), .B(n11199), .Z(n11198) );
  XNOR U11026 ( .A(n11200), .B(n11201), .Z(n11196) );
  AND U11027 ( .A(n734), .B(n11202), .Z(n11201) );
  XOR U11028 ( .A(p_input[1971]), .B(n11200), .Z(n11202) );
  XNOR U11029 ( .A(n11203), .B(n11204), .Z(n11200) );
  AND U11030 ( .A(n738), .B(n11199), .Z(n11204) );
  XOR U11031 ( .A(\knn_comb_/min_val_out[0][19] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .Z(n11199) );
  XOR U11032 ( .A(n37), .B(n11205), .Z(o[18]) );
  AND U11033 ( .A(n58), .B(n11206), .Z(n37) );
  XOR U11034 ( .A(n38), .B(n11205), .Z(n11206) );
  XOR U11035 ( .A(n11207), .B(n11208), .Z(n11205) );
  AND U11036 ( .A(n70), .B(n11209), .Z(n11208) );
  XOR U11037 ( .A(n11210), .B(n11211), .Z(n38) );
  AND U11038 ( .A(n62), .B(n11212), .Z(n11211) );
  XOR U11039 ( .A(p_input[18]), .B(n11210), .Z(n11212) );
  XNOR U11040 ( .A(n11213), .B(n11214), .Z(n11210) );
  AND U11041 ( .A(n66), .B(n11209), .Z(n11214) );
  XNOR U11042 ( .A(n11213), .B(n11207), .Z(n11209) );
  XOR U11043 ( .A(n11215), .B(n11216), .Z(n11207) );
  AND U11044 ( .A(n82), .B(n11217), .Z(n11216) );
  XNOR U11045 ( .A(n11218), .B(n11219), .Z(n11213) );
  AND U11046 ( .A(n74), .B(n11220), .Z(n11219) );
  XOR U11047 ( .A(p_input[50]), .B(n11218), .Z(n11220) );
  XNOR U11048 ( .A(n11221), .B(n11222), .Z(n11218) );
  AND U11049 ( .A(n78), .B(n11217), .Z(n11222) );
  XNOR U11050 ( .A(n11221), .B(n11215), .Z(n11217) );
  XOR U11051 ( .A(n11223), .B(n11224), .Z(n11215) );
  AND U11052 ( .A(n93), .B(n11225), .Z(n11224) );
  XNOR U11053 ( .A(n11226), .B(n11227), .Z(n11221) );
  AND U11054 ( .A(n85), .B(n11228), .Z(n11227) );
  XOR U11055 ( .A(p_input[82]), .B(n11226), .Z(n11228) );
  XNOR U11056 ( .A(n11229), .B(n11230), .Z(n11226) );
  AND U11057 ( .A(n89), .B(n11225), .Z(n11230) );
  XNOR U11058 ( .A(n11229), .B(n11223), .Z(n11225) );
  XOR U11059 ( .A(n11231), .B(n11232), .Z(n11223) );
  AND U11060 ( .A(n104), .B(n11233), .Z(n11232) );
  XNOR U11061 ( .A(n11234), .B(n11235), .Z(n11229) );
  AND U11062 ( .A(n96), .B(n11236), .Z(n11235) );
  XOR U11063 ( .A(p_input[114]), .B(n11234), .Z(n11236) );
  XNOR U11064 ( .A(n11237), .B(n11238), .Z(n11234) );
  AND U11065 ( .A(n100), .B(n11233), .Z(n11238) );
  XNOR U11066 ( .A(n11237), .B(n11231), .Z(n11233) );
  XOR U11067 ( .A(n11239), .B(n11240), .Z(n11231) );
  AND U11068 ( .A(n115), .B(n11241), .Z(n11240) );
  XNOR U11069 ( .A(n11242), .B(n11243), .Z(n11237) );
  AND U11070 ( .A(n107), .B(n11244), .Z(n11243) );
  XOR U11071 ( .A(p_input[146]), .B(n11242), .Z(n11244) );
  XNOR U11072 ( .A(n11245), .B(n11246), .Z(n11242) );
  AND U11073 ( .A(n111), .B(n11241), .Z(n11246) );
  XNOR U11074 ( .A(n11245), .B(n11239), .Z(n11241) );
  XOR U11075 ( .A(n11247), .B(n11248), .Z(n11239) );
  AND U11076 ( .A(n126), .B(n11249), .Z(n11248) );
  XNOR U11077 ( .A(n11250), .B(n11251), .Z(n11245) );
  AND U11078 ( .A(n118), .B(n11252), .Z(n11251) );
  XOR U11079 ( .A(p_input[178]), .B(n11250), .Z(n11252) );
  XNOR U11080 ( .A(n11253), .B(n11254), .Z(n11250) );
  AND U11081 ( .A(n122), .B(n11249), .Z(n11254) );
  XNOR U11082 ( .A(n11253), .B(n11247), .Z(n11249) );
  XOR U11083 ( .A(n11255), .B(n11256), .Z(n11247) );
  AND U11084 ( .A(n137), .B(n11257), .Z(n11256) );
  XNOR U11085 ( .A(n11258), .B(n11259), .Z(n11253) );
  AND U11086 ( .A(n129), .B(n11260), .Z(n11259) );
  XOR U11087 ( .A(p_input[210]), .B(n11258), .Z(n11260) );
  XNOR U11088 ( .A(n11261), .B(n11262), .Z(n11258) );
  AND U11089 ( .A(n133), .B(n11257), .Z(n11262) );
  XNOR U11090 ( .A(n11261), .B(n11255), .Z(n11257) );
  XOR U11091 ( .A(n11263), .B(n11264), .Z(n11255) );
  AND U11092 ( .A(n148), .B(n11265), .Z(n11264) );
  XNOR U11093 ( .A(n11266), .B(n11267), .Z(n11261) );
  AND U11094 ( .A(n140), .B(n11268), .Z(n11267) );
  XOR U11095 ( .A(p_input[242]), .B(n11266), .Z(n11268) );
  XNOR U11096 ( .A(n11269), .B(n11270), .Z(n11266) );
  AND U11097 ( .A(n144), .B(n11265), .Z(n11270) );
  XNOR U11098 ( .A(n11269), .B(n11263), .Z(n11265) );
  XOR U11099 ( .A(n11271), .B(n11272), .Z(n11263) );
  AND U11100 ( .A(n159), .B(n11273), .Z(n11272) );
  XNOR U11101 ( .A(n11274), .B(n11275), .Z(n11269) );
  AND U11102 ( .A(n151), .B(n11276), .Z(n11275) );
  XOR U11103 ( .A(p_input[274]), .B(n11274), .Z(n11276) );
  XNOR U11104 ( .A(n11277), .B(n11278), .Z(n11274) );
  AND U11105 ( .A(n155), .B(n11273), .Z(n11278) );
  XNOR U11106 ( .A(n11277), .B(n11271), .Z(n11273) );
  XOR U11107 ( .A(n11279), .B(n11280), .Z(n11271) );
  AND U11108 ( .A(n170), .B(n11281), .Z(n11280) );
  XNOR U11109 ( .A(n11282), .B(n11283), .Z(n11277) );
  AND U11110 ( .A(n162), .B(n11284), .Z(n11283) );
  XOR U11111 ( .A(p_input[306]), .B(n11282), .Z(n11284) );
  XNOR U11112 ( .A(n11285), .B(n11286), .Z(n11282) );
  AND U11113 ( .A(n166), .B(n11281), .Z(n11286) );
  XNOR U11114 ( .A(n11285), .B(n11279), .Z(n11281) );
  XOR U11115 ( .A(n11287), .B(n11288), .Z(n11279) );
  AND U11116 ( .A(n181), .B(n11289), .Z(n11288) );
  XNOR U11117 ( .A(n11290), .B(n11291), .Z(n11285) );
  AND U11118 ( .A(n173), .B(n11292), .Z(n11291) );
  XOR U11119 ( .A(p_input[338]), .B(n11290), .Z(n11292) );
  XNOR U11120 ( .A(n11293), .B(n11294), .Z(n11290) );
  AND U11121 ( .A(n177), .B(n11289), .Z(n11294) );
  XNOR U11122 ( .A(n11293), .B(n11287), .Z(n11289) );
  XOR U11123 ( .A(n11295), .B(n11296), .Z(n11287) );
  AND U11124 ( .A(n192), .B(n11297), .Z(n11296) );
  XNOR U11125 ( .A(n11298), .B(n11299), .Z(n11293) );
  AND U11126 ( .A(n184), .B(n11300), .Z(n11299) );
  XOR U11127 ( .A(p_input[370]), .B(n11298), .Z(n11300) );
  XNOR U11128 ( .A(n11301), .B(n11302), .Z(n11298) );
  AND U11129 ( .A(n188), .B(n11297), .Z(n11302) );
  XNOR U11130 ( .A(n11301), .B(n11295), .Z(n11297) );
  XOR U11131 ( .A(n11303), .B(n11304), .Z(n11295) );
  AND U11132 ( .A(n203), .B(n11305), .Z(n11304) );
  XNOR U11133 ( .A(n11306), .B(n11307), .Z(n11301) );
  AND U11134 ( .A(n195), .B(n11308), .Z(n11307) );
  XOR U11135 ( .A(p_input[402]), .B(n11306), .Z(n11308) );
  XNOR U11136 ( .A(n11309), .B(n11310), .Z(n11306) );
  AND U11137 ( .A(n199), .B(n11305), .Z(n11310) );
  XNOR U11138 ( .A(n11309), .B(n11303), .Z(n11305) );
  XOR U11139 ( .A(n11311), .B(n11312), .Z(n11303) );
  AND U11140 ( .A(n214), .B(n11313), .Z(n11312) );
  XNOR U11141 ( .A(n11314), .B(n11315), .Z(n11309) );
  AND U11142 ( .A(n206), .B(n11316), .Z(n11315) );
  XOR U11143 ( .A(p_input[434]), .B(n11314), .Z(n11316) );
  XNOR U11144 ( .A(n11317), .B(n11318), .Z(n11314) );
  AND U11145 ( .A(n210), .B(n11313), .Z(n11318) );
  XNOR U11146 ( .A(n11317), .B(n11311), .Z(n11313) );
  XOR U11147 ( .A(n11319), .B(n11320), .Z(n11311) );
  AND U11148 ( .A(n225), .B(n11321), .Z(n11320) );
  XNOR U11149 ( .A(n11322), .B(n11323), .Z(n11317) );
  AND U11150 ( .A(n217), .B(n11324), .Z(n11323) );
  XOR U11151 ( .A(p_input[466]), .B(n11322), .Z(n11324) );
  XNOR U11152 ( .A(n11325), .B(n11326), .Z(n11322) );
  AND U11153 ( .A(n221), .B(n11321), .Z(n11326) );
  XNOR U11154 ( .A(n11325), .B(n11319), .Z(n11321) );
  XOR U11155 ( .A(n11327), .B(n11328), .Z(n11319) );
  AND U11156 ( .A(n236), .B(n11329), .Z(n11328) );
  XNOR U11157 ( .A(n11330), .B(n11331), .Z(n11325) );
  AND U11158 ( .A(n228), .B(n11332), .Z(n11331) );
  XOR U11159 ( .A(p_input[498]), .B(n11330), .Z(n11332) );
  XNOR U11160 ( .A(n11333), .B(n11334), .Z(n11330) );
  AND U11161 ( .A(n232), .B(n11329), .Z(n11334) );
  XNOR U11162 ( .A(n11333), .B(n11327), .Z(n11329) );
  XOR U11163 ( .A(n11335), .B(n11336), .Z(n11327) );
  AND U11164 ( .A(n247), .B(n11337), .Z(n11336) );
  XNOR U11165 ( .A(n11338), .B(n11339), .Z(n11333) );
  AND U11166 ( .A(n239), .B(n11340), .Z(n11339) );
  XOR U11167 ( .A(p_input[530]), .B(n11338), .Z(n11340) );
  XNOR U11168 ( .A(n11341), .B(n11342), .Z(n11338) );
  AND U11169 ( .A(n243), .B(n11337), .Z(n11342) );
  XNOR U11170 ( .A(n11341), .B(n11335), .Z(n11337) );
  XOR U11171 ( .A(n11343), .B(n11344), .Z(n11335) );
  AND U11172 ( .A(n258), .B(n11345), .Z(n11344) );
  XNOR U11173 ( .A(n11346), .B(n11347), .Z(n11341) );
  AND U11174 ( .A(n250), .B(n11348), .Z(n11347) );
  XOR U11175 ( .A(p_input[562]), .B(n11346), .Z(n11348) );
  XNOR U11176 ( .A(n11349), .B(n11350), .Z(n11346) );
  AND U11177 ( .A(n254), .B(n11345), .Z(n11350) );
  XNOR U11178 ( .A(n11349), .B(n11343), .Z(n11345) );
  XOR U11179 ( .A(n11351), .B(n11352), .Z(n11343) );
  AND U11180 ( .A(n269), .B(n11353), .Z(n11352) );
  XNOR U11181 ( .A(n11354), .B(n11355), .Z(n11349) );
  AND U11182 ( .A(n261), .B(n11356), .Z(n11355) );
  XOR U11183 ( .A(p_input[594]), .B(n11354), .Z(n11356) );
  XNOR U11184 ( .A(n11357), .B(n11358), .Z(n11354) );
  AND U11185 ( .A(n265), .B(n11353), .Z(n11358) );
  XNOR U11186 ( .A(n11357), .B(n11351), .Z(n11353) );
  XOR U11187 ( .A(n11359), .B(n11360), .Z(n11351) );
  AND U11188 ( .A(n280), .B(n11361), .Z(n11360) );
  XNOR U11189 ( .A(n11362), .B(n11363), .Z(n11357) );
  AND U11190 ( .A(n272), .B(n11364), .Z(n11363) );
  XOR U11191 ( .A(p_input[626]), .B(n11362), .Z(n11364) );
  XNOR U11192 ( .A(n11365), .B(n11366), .Z(n11362) );
  AND U11193 ( .A(n276), .B(n11361), .Z(n11366) );
  XNOR U11194 ( .A(n11365), .B(n11359), .Z(n11361) );
  XOR U11195 ( .A(n11367), .B(n11368), .Z(n11359) );
  AND U11196 ( .A(n291), .B(n11369), .Z(n11368) );
  XNOR U11197 ( .A(n11370), .B(n11371), .Z(n11365) );
  AND U11198 ( .A(n283), .B(n11372), .Z(n11371) );
  XOR U11199 ( .A(p_input[658]), .B(n11370), .Z(n11372) );
  XNOR U11200 ( .A(n11373), .B(n11374), .Z(n11370) );
  AND U11201 ( .A(n287), .B(n11369), .Z(n11374) );
  XNOR U11202 ( .A(n11373), .B(n11367), .Z(n11369) );
  XOR U11203 ( .A(n11375), .B(n11376), .Z(n11367) );
  AND U11204 ( .A(n302), .B(n11377), .Z(n11376) );
  XNOR U11205 ( .A(n11378), .B(n11379), .Z(n11373) );
  AND U11206 ( .A(n294), .B(n11380), .Z(n11379) );
  XOR U11207 ( .A(p_input[690]), .B(n11378), .Z(n11380) );
  XNOR U11208 ( .A(n11381), .B(n11382), .Z(n11378) );
  AND U11209 ( .A(n298), .B(n11377), .Z(n11382) );
  XNOR U11210 ( .A(n11381), .B(n11375), .Z(n11377) );
  XOR U11211 ( .A(n11383), .B(n11384), .Z(n11375) );
  AND U11212 ( .A(n313), .B(n11385), .Z(n11384) );
  XNOR U11213 ( .A(n11386), .B(n11387), .Z(n11381) );
  AND U11214 ( .A(n305), .B(n11388), .Z(n11387) );
  XOR U11215 ( .A(p_input[722]), .B(n11386), .Z(n11388) );
  XNOR U11216 ( .A(n11389), .B(n11390), .Z(n11386) );
  AND U11217 ( .A(n309), .B(n11385), .Z(n11390) );
  XNOR U11218 ( .A(n11389), .B(n11383), .Z(n11385) );
  XOR U11219 ( .A(n11391), .B(n11392), .Z(n11383) );
  AND U11220 ( .A(n324), .B(n11393), .Z(n11392) );
  XNOR U11221 ( .A(n11394), .B(n11395), .Z(n11389) );
  AND U11222 ( .A(n316), .B(n11396), .Z(n11395) );
  XOR U11223 ( .A(p_input[754]), .B(n11394), .Z(n11396) );
  XNOR U11224 ( .A(n11397), .B(n11398), .Z(n11394) );
  AND U11225 ( .A(n320), .B(n11393), .Z(n11398) );
  XNOR U11226 ( .A(n11397), .B(n11391), .Z(n11393) );
  XOR U11227 ( .A(n11399), .B(n11400), .Z(n11391) );
  AND U11228 ( .A(n335), .B(n11401), .Z(n11400) );
  XNOR U11229 ( .A(n11402), .B(n11403), .Z(n11397) );
  AND U11230 ( .A(n327), .B(n11404), .Z(n11403) );
  XOR U11231 ( .A(p_input[786]), .B(n11402), .Z(n11404) );
  XNOR U11232 ( .A(n11405), .B(n11406), .Z(n11402) );
  AND U11233 ( .A(n331), .B(n11401), .Z(n11406) );
  XNOR U11234 ( .A(n11405), .B(n11399), .Z(n11401) );
  XOR U11235 ( .A(n11407), .B(n11408), .Z(n11399) );
  AND U11236 ( .A(n346), .B(n11409), .Z(n11408) );
  XNOR U11237 ( .A(n11410), .B(n11411), .Z(n11405) );
  AND U11238 ( .A(n338), .B(n11412), .Z(n11411) );
  XOR U11239 ( .A(p_input[818]), .B(n11410), .Z(n11412) );
  XNOR U11240 ( .A(n11413), .B(n11414), .Z(n11410) );
  AND U11241 ( .A(n342), .B(n11409), .Z(n11414) );
  XNOR U11242 ( .A(n11413), .B(n11407), .Z(n11409) );
  XOR U11243 ( .A(n11415), .B(n11416), .Z(n11407) );
  AND U11244 ( .A(n357), .B(n11417), .Z(n11416) );
  XNOR U11245 ( .A(n11418), .B(n11419), .Z(n11413) );
  AND U11246 ( .A(n349), .B(n11420), .Z(n11419) );
  XOR U11247 ( .A(p_input[850]), .B(n11418), .Z(n11420) );
  XNOR U11248 ( .A(n11421), .B(n11422), .Z(n11418) );
  AND U11249 ( .A(n353), .B(n11417), .Z(n11422) );
  XNOR U11250 ( .A(n11421), .B(n11415), .Z(n11417) );
  XOR U11251 ( .A(n11423), .B(n11424), .Z(n11415) );
  AND U11252 ( .A(n368), .B(n11425), .Z(n11424) );
  XNOR U11253 ( .A(n11426), .B(n11427), .Z(n11421) );
  AND U11254 ( .A(n360), .B(n11428), .Z(n11427) );
  XOR U11255 ( .A(p_input[882]), .B(n11426), .Z(n11428) );
  XNOR U11256 ( .A(n11429), .B(n11430), .Z(n11426) );
  AND U11257 ( .A(n364), .B(n11425), .Z(n11430) );
  XNOR U11258 ( .A(n11429), .B(n11423), .Z(n11425) );
  XOR U11259 ( .A(n11431), .B(n11432), .Z(n11423) );
  AND U11260 ( .A(n379), .B(n11433), .Z(n11432) );
  XNOR U11261 ( .A(n11434), .B(n11435), .Z(n11429) );
  AND U11262 ( .A(n371), .B(n11436), .Z(n11435) );
  XOR U11263 ( .A(p_input[914]), .B(n11434), .Z(n11436) );
  XNOR U11264 ( .A(n11437), .B(n11438), .Z(n11434) );
  AND U11265 ( .A(n375), .B(n11433), .Z(n11438) );
  XNOR U11266 ( .A(n11437), .B(n11431), .Z(n11433) );
  XOR U11267 ( .A(n11439), .B(n11440), .Z(n11431) );
  AND U11268 ( .A(n390), .B(n11441), .Z(n11440) );
  XNOR U11269 ( .A(n11442), .B(n11443), .Z(n11437) );
  AND U11270 ( .A(n382), .B(n11444), .Z(n11443) );
  XOR U11271 ( .A(p_input[946]), .B(n11442), .Z(n11444) );
  XNOR U11272 ( .A(n11445), .B(n11446), .Z(n11442) );
  AND U11273 ( .A(n386), .B(n11441), .Z(n11446) );
  XNOR U11274 ( .A(n11445), .B(n11439), .Z(n11441) );
  XOR U11275 ( .A(n11447), .B(n11448), .Z(n11439) );
  AND U11276 ( .A(n401), .B(n11449), .Z(n11448) );
  XNOR U11277 ( .A(n11450), .B(n11451), .Z(n11445) );
  AND U11278 ( .A(n393), .B(n11452), .Z(n11451) );
  XOR U11279 ( .A(p_input[978]), .B(n11450), .Z(n11452) );
  XNOR U11280 ( .A(n11453), .B(n11454), .Z(n11450) );
  AND U11281 ( .A(n397), .B(n11449), .Z(n11454) );
  XNOR U11282 ( .A(n11453), .B(n11447), .Z(n11449) );
  XOR U11283 ( .A(n11455), .B(n11456), .Z(n11447) );
  AND U11284 ( .A(n412), .B(n11457), .Z(n11456) );
  XNOR U11285 ( .A(n11458), .B(n11459), .Z(n11453) );
  AND U11286 ( .A(n404), .B(n11460), .Z(n11459) );
  XOR U11287 ( .A(p_input[1010]), .B(n11458), .Z(n11460) );
  XNOR U11288 ( .A(n11461), .B(n11462), .Z(n11458) );
  AND U11289 ( .A(n408), .B(n11457), .Z(n11462) );
  XNOR U11290 ( .A(n11461), .B(n11455), .Z(n11457) );
  XOR U11291 ( .A(n11463), .B(n11464), .Z(n11455) );
  AND U11292 ( .A(n423), .B(n11465), .Z(n11464) );
  XNOR U11293 ( .A(n11466), .B(n11467), .Z(n11461) );
  AND U11294 ( .A(n415), .B(n11468), .Z(n11467) );
  XOR U11295 ( .A(p_input[1042]), .B(n11466), .Z(n11468) );
  XNOR U11296 ( .A(n11469), .B(n11470), .Z(n11466) );
  AND U11297 ( .A(n419), .B(n11465), .Z(n11470) );
  XNOR U11298 ( .A(n11469), .B(n11463), .Z(n11465) );
  XOR U11299 ( .A(n11471), .B(n11472), .Z(n11463) );
  AND U11300 ( .A(n434), .B(n11473), .Z(n11472) );
  XNOR U11301 ( .A(n11474), .B(n11475), .Z(n11469) );
  AND U11302 ( .A(n426), .B(n11476), .Z(n11475) );
  XOR U11303 ( .A(p_input[1074]), .B(n11474), .Z(n11476) );
  XNOR U11304 ( .A(n11477), .B(n11478), .Z(n11474) );
  AND U11305 ( .A(n430), .B(n11473), .Z(n11478) );
  XNOR U11306 ( .A(n11477), .B(n11471), .Z(n11473) );
  XOR U11307 ( .A(n11479), .B(n11480), .Z(n11471) );
  AND U11308 ( .A(n445), .B(n11481), .Z(n11480) );
  XNOR U11309 ( .A(n11482), .B(n11483), .Z(n11477) );
  AND U11310 ( .A(n437), .B(n11484), .Z(n11483) );
  XOR U11311 ( .A(p_input[1106]), .B(n11482), .Z(n11484) );
  XNOR U11312 ( .A(n11485), .B(n11486), .Z(n11482) );
  AND U11313 ( .A(n441), .B(n11481), .Z(n11486) );
  XNOR U11314 ( .A(n11485), .B(n11479), .Z(n11481) );
  XOR U11315 ( .A(n11487), .B(n11488), .Z(n11479) );
  AND U11316 ( .A(n456), .B(n11489), .Z(n11488) );
  XNOR U11317 ( .A(n11490), .B(n11491), .Z(n11485) );
  AND U11318 ( .A(n448), .B(n11492), .Z(n11491) );
  XOR U11319 ( .A(p_input[1138]), .B(n11490), .Z(n11492) );
  XNOR U11320 ( .A(n11493), .B(n11494), .Z(n11490) );
  AND U11321 ( .A(n452), .B(n11489), .Z(n11494) );
  XNOR U11322 ( .A(n11493), .B(n11487), .Z(n11489) );
  XOR U11323 ( .A(n11495), .B(n11496), .Z(n11487) );
  AND U11324 ( .A(n467), .B(n11497), .Z(n11496) );
  XNOR U11325 ( .A(n11498), .B(n11499), .Z(n11493) );
  AND U11326 ( .A(n459), .B(n11500), .Z(n11499) );
  XOR U11327 ( .A(p_input[1170]), .B(n11498), .Z(n11500) );
  XNOR U11328 ( .A(n11501), .B(n11502), .Z(n11498) );
  AND U11329 ( .A(n463), .B(n11497), .Z(n11502) );
  XNOR U11330 ( .A(n11501), .B(n11495), .Z(n11497) );
  XOR U11331 ( .A(n11503), .B(n11504), .Z(n11495) );
  AND U11332 ( .A(n478), .B(n11505), .Z(n11504) );
  XNOR U11333 ( .A(n11506), .B(n11507), .Z(n11501) );
  AND U11334 ( .A(n470), .B(n11508), .Z(n11507) );
  XOR U11335 ( .A(p_input[1202]), .B(n11506), .Z(n11508) );
  XNOR U11336 ( .A(n11509), .B(n11510), .Z(n11506) );
  AND U11337 ( .A(n474), .B(n11505), .Z(n11510) );
  XNOR U11338 ( .A(n11509), .B(n11503), .Z(n11505) );
  XOR U11339 ( .A(n11511), .B(n11512), .Z(n11503) );
  AND U11340 ( .A(n489), .B(n11513), .Z(n11512) );
  XNOR U11341 ( .A(n11514), .B(n11515), .Z(n11509) );
  AND U11342 ( .A(n481), .B(n11516), .Z(n11515) );
  XOR U11343 ( .A(p_input[1234]), .B(n11514), .Z(n11516) );
  XNOR U11344 ( .A(n11517), .B(n11518), .Z(n11514) );
  AND U11345 ( .A(n485), .B(n11513), .Z(n11518) );
  XNOR U11346 ( .A(n11517), .B(n11511), .Z(n11513) );
  XOR U11347 ( .A(n11519), .B(n11520), .Z(n11511) );
  AND U11348 ( .A(n500), .B(n11521), .Z(n11520) );
  XNOR U11349 ( .A(n11522), .B(n11523), .Z(n11517) );
  AND U11350 ( .A(n492), .B(n11524), .Z(n11523) );
  XOR U11351 ( .A(p_input[1266]), .B(n11522), .Z(n11524) );
  XNOR U11352 ( .A(n11525), .B(n11526), .Z(n11522) );
  AND U11353 ( .A(n496), .B(n11521), .Z(n11526) );
  XNOR U11354 ( .A(n11525), .B(n11519), .Z(n11521) );
  XOR U11355 ( .A(n11527), .B(n11528), .Z(n11519) );
  AND U11356 ( .A(n511), .B(n11529), .Z(n11528) );
  XNOR U11357 ( .A(n11530), .B(n11531), .Z(n11525) );
  AND U11358 ( .A(n503), .B(n11532), .Z(n11531) );
  XOR U11359 ( .A(p_input[1298]), .B(n11530), .Z(n11532) );
  XNOR U11360 ( .A(n11533), .B(n11534), .Z(n11530) );
  AND U11361 ( .A(n507), .B(n11529), .Z(n11534) );
  XNOR U11362 ( .A(n11533), .B(n11527), .Z(n11529) );
  XOR U11363 ( .A(n11535), .B(n11536), .Z(n11527) );
  AND U11364 ( .A(n522), .B(n11537), .Z(n11536) );
  XNOR U11365 ( .A(n11538), .B(n11539), .Z(n11533) );
  AND U11366 ( .A(n514), .B(n11540), .Z(n11539) );
  XOR U11367 ( .A(p_input[1330]), .B(n11538), .Z(n11540) );
  XNOR U11368 ( .A(n11541), .B(n11542), .Z(n11538) );
  AND U11369 ( .A(n518), .B(n11537), .Z(n11542) );
  XNOR U11370 ( .A(n11541), .B(n11535), .Z(n11537) );
  XOR U11371 ( .A(n11543), .B(n11544), .Z(n11535) );
  AND U11372 ( .A(n533), .B(n11545), .Z(n11544) );
  XNOR U11373 ( .A(n11546), .B(n11547), .Z(n11541) );
  AND U11374 ( .A(n525), .B(n11548), .Z(n11547) );
  XOR U11375 ( .A(p_input[1362]), .B(n11546), .Z(n11548) );
  XNOR U11376 ( .A(n11549), .B(n11550), .Z(n11546) );
  AND U11377 ( .A(n529), .B(n11545), .Z(n11550) );
  XNOR U11378 ( .A(n11549), .B(n11543), .Z(n11545) );
  XOR U11379 ( .A(n11551), .B(n11552), .Z(n11543) );
  AND U11380 ( .A(n544), .B(n11553), .Z(n11552) );
  XNOR U11381 ( .A(n11554), .B(n11555), .Z(n11549) );
  AND U11382 ( .A(n536), .B(n11556), .Z(n11555) );
  XOR U11383 ( .A(p_input[1394]), .B(n11554), .Z(n11556) );
  XNOR U11384 ( .A(n11557), .B(n11558), .Z(n11554) );
  AND U11385 ( .A(n540), .B(n11553), .Z(n11558) );
  XNOR U11386 ( .A(n11557), .B(n11551), .Z(n11553) );
  XOR U11387 ( .A(n11559), .B(n11560), .Z(n11551) );
  AND U11388 ( .A(n555), .B(n11561), .Z(n11560) );
  XNOR U11389 ( .A(n11562), .B(n11563), .Z(n11557) );
  AND U11390 ( .A(n547), .B(n11564), .Z(n11563) );
  XOR U11391 ( .A(p_input[1426]), .B(n11562), .Z(n11564) );
  XNOR U11392 ( .A(n11565), .B(n11566), .Z(n11562) );
  AND U11393 ( .A(n551), .B(n11561), .Z(n11566) );
  XNOR U11394 ( .A(n11565), .B(n11559), .Z(n11561) );
  XOR U11395 ( .A(n11567), .B(n11568), .Z(n11559) );
  AND U11396 ( .A(n566), .B(n11569), .Z(n11568) );
  XNOR U11397 ( .A(n11570), .B(n11571), .Z(n11565) );
  AND U11398 ( .A(n558), .B(n11572), .Z(n11571) );
  XOR U11399 ( .A(p_input[1458]), .B(n11570), .Z(n11572) );
  XNOR U11400 ( .A(n11573), .B(n11574), .Z(n11570) );
  AND U11401 ( .A(n562), .B(n11569), .Z(n11574) );
  XNOR U11402 ( .A(n11573), .B(n11567), .Z(n11569) );
  XOR U11403 ( .A(n11575), .B(n11576), .Z(n11567) );
  AND U11404 ( .A(n577), .B(n11577), .Z(n11576) );
  XNOR U11405 ( .A(n11578), .B(n11579), .Z(n11573) );
  AND U11406 ( .A(n569), .B(n11580), .Z(n11579) );
  XOR U11407 ( .A(p_input[1490]), .B(n11578), .Z(n11580) );
  XNOR U11408 ( .A(n11581), .B(n11582), .Z(n11578) );
  AND U11409 ( .A(n573), .B(n11577), .Z(n11582) );
  XNOR U11410 ( .A(n11581), .B(n11575), .Z(n11577) );
  XOR U11411 ( .A(n11583), .B(n11584), .Z(n11575) );
  AND U11412 ( .A(n588), .B(n11585), .Z(n11584) );
  XNOR U11413 ( .A(n11586), .B(n11587), .Z(n11581) );
  AND U11414 ( .A(n580), .B(n11588), .Z(n11587) );
  XOR U11415 ( .A(p_input[1522]), .B(n11586), .Z(n11588) );
  XNOR U11416 ( .A(n11589), .B(n11590), .Z(n11586) );
  AND U11417 ( .A(n584), .B(n11585), .Z(n11590) );
  XNOR U11418 ( .A(n11589), .B(n11583), .Z(n11585) );
  XOR U11419 ( .A(n11591), .B(n11592), .Z(n11583) );
  AND U11420 ( .A(n599), .B(n11593), .Z(n11592) );
  XNOR U11421 ( .A(n11594), .B(n11595), .Z(n11589) );
  AND U11422 ( .A(n591), .B(n11596), .Z(n11595) );
  XOR U11423 ( .A(p_input[1554]), .B(n11594), .Z(n11596) );
  XNOR U11424 ( .A(n11597), .B(n11598), .Z(n11594) );
  AND U11425 ( .A(n595), .B(n11593), .Z(n11598) );
  XNOR U11426 ( .A(n11597), .B(n11591), .Z(n11593) );
  XOR U11427 ( .A(n11599), .B(n11600), .Z(n11591) );
  AND U11428 ( .A(n610), .B(n11601), .Z(n11600) );
  XNOR U11429 ( .A(n11602), .B(n11603), .Z(n11597) );
  AND U11430 ( .A(n602), .B(n11604), .Z(n11603) );
  XOR U11431 ( .A(p_input[1586]), .B(n11602), .Z(n11604) );
  XNOR U11432 ( .A(n11605), .B(n11606), .Z(n11602) );
  AND U11433 ( .A(n606), .B(n11601), .Z(n11606) );
  XNOR U11434 ( .A(n11605), .B(n11599), .Z(n11601) );
  XOR U11435 ( .A(n11607), .B(n11608), .Z(n11599) );
  AND U11436 ( .A(n621), .B(n11609), .Z(n11608) );
  XNOR U11437 ( .A(n11610), .B(n11611), .Z(n11605) );
  AND U11438 ( .A(n613), .B(n11612), .Z(n11611) );
  XOR U11439 ( .A(p_input[1618]), .B(n11610), .Z(n11612) );
  XNOR U11440 ( .A(n11613), .B(n11614), .Z(n11610) );
  AND U11441 ( .A(n617), .B(n11609), .Z(n11614) );
  XNOR U11442 ( .A(n11613), .B(n11607), .Z(n11609) );
  XOR U11443 ( .A(n11615), .B(n11616), .Z(n11607) );
  AND U11444 ( .A(n632), .B(n11617), .Z(n11616) );
  XNOR U11445 ( .A(n11618), .B(n11619), .Z(n11613) );
  AND U11446 ( .A(n624), .B(n11620), .Z(n11619) );
  XOR U11447 ( .A(p_input[1650]), .B(n11618), .Z(n11620) );
  XNOR U11448 ( .A(n11621), .B(n11622), .Z(n11618) );
  AND U11449 ( .A(n628), .B(n11617), .Z(n11622) );
  XNOR U11450 ( .A(n11621), .B(n11615), .Z(n11617) );
  XOR U11451 ( .A(n11623), .B(n11624), .Z(n11615) );
  AND U11452 ( .A(n643), .B(n11625), .Z(n11624) );
  XNOR U11453 ( .A(n11626), .B(n11627), .Z(n11621) );
  AND U11454 ( .A(n635), .B(n11628), .Z(n11627) );
  XOR U11455 ( .A(p_input[1682]), .B(n11626), .Z(n11628) );
  XNOR U11456 ( .A(n11629), .B(n11630), .Z(n11626) );
  AND U11457 ( .A(n639), .B(n11625), .Z(n11630) );
  XNOR U11458 ( .A(n11629), .B(n11623), .Z(n11625) );
  XOR U11459 ( .A(n11631), .B(n11632), .Z(n11623) );
  AND U11460 ( .A(n654), .B(n11633), .Z(n11632) );
  XNOR U11461 ( .A(n11634), .B(n11635), .Z(n11629) );
  AND U11462 ( .A(n646), .B(n11636), .Z(n11635) );
  XOR U11463 ( .A(p_input[1714]), .B(n11634), .Z(n11636) );
  XNOR U11464 ( .A(n11637), .B(n11638), .Z(n11634) );
  AND U11465 ( .A(n650), .B(n11633), .Z(n11638) );
  XNOR U11466 ( .A(n11637), .B(n11631), .Z(n11633) );
  XOR U11467 ( .A(n11639), .B(n11640), .Z(n11631) );
  AND U11468 ( .A(n665), .B(n11641), .Z(n11640) );
  XNOR U11469 ( .A(n11642), .B(n11643), .Z(n11637) );
  AND U11470 ( .A(n657), .B(n11644), .Z(n11643) );
  XOR U11471 ( .A(p_input[1746]), .B(n11642), .Z(n11644) );
  XNOR U11472 ( .A(n11645), .B(n11646), .Z(n11642) );
  AND U11473 ( .A(n661), .B(n11641), .Z(n11646) );
  XNOR U11474 ( .A(n11645), .B(n11639), .Z(n11641) );
  XOR U11475 ( .A(n11647), .B(n11648), .Z(n11639) );
  AND U11476 ( .A(n676), .B(n11649), .Z(n11648) );
  XNOR U11477 ( .A(n11650), .B(n11651), .Z(n11645) );
  AND U11478 ( .A(n668), .B(n11652), .Z(n11651) );
  XOR U11479 ( .A(p_input[1778]), .B(n11650), .Z(n11652) );
  XNOR U11480 ( .A(n11653), .B(n11654), .Z(n11650) );
  AND U11481 ( .A(n672), .B(n11649), .Z(n11654) );
  XNOR U11482 ( .A(n11653), .B(n11647), .Z(n11649) );
  XOR U11483 ( .A(n11655), .B(n11656), .Z(n11647) );
  AND U11484 ( .A(n687), .B(n11657), .Z(n11656) );
  XNOR U11485 ( .A(n11658), .B(n11659), .Z(n11653) );
  AND U11486 ( .A(n679), .B(n11660), .Z(n11659) );
  XOR U11487 ( .A(p_input[1810]), .B(n11658), .Z(n11660) );
  XNOR U11488 ( .A(n11661), .B(n11662), .Z(n11658) );
  AND U11489 ( .A(n683), .B(n11657), .Z(n11662) );
  XNOR U11490 ( .A(n11661), .B(n11655), .Z(n11657) );
  XOR U11491 ( .A(n11663), .B(n11664), .Z(n11655) );
  AND U11492 ( .A(n698), .B(n11665), .Z(n11664) );
  XNOR U11493 ( .A(n11666), .B(n11667), .Z(n11661) );
  AND U11494 ( .A(n690), .B(n11668), .Z(n11667) );
  XOR U11495 ( .A(p_input[1842]), .B(n11666), .Z(n11668) );
  XNOR U11496 ( .A(n11669), .B(n11670), .Z(n11666) );
  AND U11497 ( .A(n694), .B(n11665), .Z(n11670) );
  XNOR U11498 ( .A(n11669), .B(n11663), .Z(n11665) );
  XOR U11499 ( .A(n11671), .B(n11672), .Z(n11663) );
  AND U11500 ( .A(n709), .B(n11673), .Z(n11672) );
  XNOR U11501 ( .A(n11674), .B(n11675), .Z(n11669) );
  AND U11502 ( .A(n701), .B(n11676), .Z(n11675) );
  XOR U11503 ( .A(p_input[1874]), .B(n11674), .Z(n11676) );
  XNOR U11504 ( .A(n11677), .B(n11678), .Z(n11674) );
  AND U11505 ( .A(n705), .B(n11673), .Z(n11678) );
  XNOR U11506 ( .A(n11677), .B(n11671), .Z(n11673) );
  XOR U11507 ( .A(n11679), .B(n11680), .Z(n11671) );
  AND U11508 ( .A(n720), .B(n11681), .Z(n11680) );
  XNOR U11509 ( .A(n11682), .B(n11683), .Z(n11677) );
  AND U11510 ( .A(n712), .B(n11684), .Z(n11683) );
  XOR U11511 ( .A(p_input[1906]), .B(n11682), .Z(n11684) );
  XNOR U11512 ( .A(n11685), .B(n11686), .Z(n11682) );
  AND U11513 ( .A(n716), .B(n11681), .Z(n11686) );
  XNOR U11514 ( .A(n11685), .B(n11679), .Z(n11681) );
  XOR U11515 ( .A(n11687), .B(n11688), .Z(n11679) );
  AND U11516 ( .A(n731), .B(n11689), .Z(n11688) );
  XNOR U11517 ( .A(n11690), .B(n11691), .Z(n11685) );
  AND U11518 ( .A(n723), .B(n11692), .Z(n11691) );
  XOR U11519 ( .A(p_input[1938]), .B(n11690), .Z(n11692) );
  XNOR U11520 ( .A(n11693), .B(n11694), .Z(n11690) );
  AND U11521 ( .A(n727), .B(n11689), .Z(n11694) );
  XNOR U11522 ( .A(n11693), .B(n11687), .Z(n11689) );
  XOR U11523 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n11695), .Z(n11687) );
  AND U11524 ( .A(n741), .B(n11696), .Z(n11695) );
  XNOR U11525 ( .A(n11697), .B(n11698), .Z(n11693) );
  AND U11526 ( .A(n734), .B(n11699), .Z(n11698) );
  XOR U11527 ( .A(p_input[1970]), .B(n11697), .Z(n11699) );
  XNOR U11528 ( .A(n11700), .B(n11701), .Z(n11697) );
  AND U11529 ( .A(n738), .B(n11696), .Z(n11701) );
  XOR U11530 ( .A(\knn_comb_/min_val_out[0][18] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .Z(n11696) );
  XOR U11531 ( .A(n41), .B(n11702), .Z(o[17]) );
  AND U11532 ( .A(n58), .B(n11703), .Z(n41) );
  XOR U11533 ( .A(n42), .B(n11702), .Z(n11703) );
  XOR U11534 ( .A(n11704), .B(n11705), .Z(n11702) );
  AND U11535 ( .A(n70), .B(n11706), .Z(n11705) );
  XOR U11536 ( .A(n11707), .B(n11708), .Z(n42) );
  AND U11537 ( .A(n62), .B(n11709), .Z(n11708) );
  XOR U11538 ( .A(p_input[17]), .B(n11707), .Z(n11709) );
  XNOR U11539 ( .A(n11710), .B(n11711), .Z(n11707) );
  AND U11540 ( .A(n66), .B(n11706), .Z(n11711) );
  XNOR U11541 ( .A(n11710), .B(n11704), .Z(n11706) );
  XOR U11542 ( .A(n11712), .B(n11713), .Z(n11704) );
  AND U11543 ( .A(n82), .B(n11714), .Z(n11713) );
  XNOR U11544 ( .A(n11715), .B(n11716), .Z(n11710) );
  AND U11545 ( .A(n74), .B(n11717), .Z(n11716) );
  XOR U11546 ( .A(p_input[49]), .B(n11715), .Z(n11717) );
  XNOR U11547 ( .A(n11718), .B(n11719), .Z(n11715) );
  AND U11548 ( .A(n78), .B(n11714), .Z(n11719) );
  XNOR U11549 ( .A(n11718), .B(n11712), .Z(n11714) );
  XOR U11550 ( .A(n11720), .B(n11721), .Z(n11712) );
  AND U11551 ( .A(n93), .B(n11722), .Z(n11721) );
  XNOR U11552 ( .A(n11723), .B(n11724), .Z(n11718) );
  AND U11553 ( .A(n85), .B(n11725), .Z(n11724) );
  XOR U11554 ( .A(p_input[81]), .B(n11723), .Z(n11725) );
  XNOR U11555 ( .A(n11726), .B(n11727), .Z(n11723) );
  AND U11556 ( .A(n89), .B(n11722), .Z(n11727) );
  XNOR U11557 ( .A(n11726), .B(n11720), .Z(n11722) );
  XOR U11558 ( .A(n11728), .B(n11729), .Z(n11720) );
  AND U11559 ( .A(n104), .B(n11730), .Z(n11729) );
  XNOR U11560 ( .A(n11731), .B(n11732), .Z(n11726) );
  AND U11561 ( .A(n96), .B(n11733), .Z(n11732) );
  XOR U11562 ( .A(p_input[113]), .B(n11731), .Z(n11733) );
  XNOR U11563 ( .A(n11734), .B(n11735), .Z(n11731) );
  AND U11564 ( .A(n100), .B(n11730), .Z(n11735) );
  XNOR U11565 ( .A(n11734), .B(n11728), .Z(n11730) );
  XOR U11566 ( .A(n11736), .B(n11737), .Z(n11728) );
  AND U11567 ( .A(n115), .B(n11738), .Z(n11737) );
  XNOR U11568 ( .A(n11739), .B(n11740), .Z(n11734) );
  AND U11569 ( .A(n107), .B(n11741), .Z(n11740) );
  XOR U11570 ( .A(p_input[145]), .B(n11739), .Z(n11741) );
  XNOR U11571 ( .A(n11742), .B(n11743), .Z(n11739) );
  AND U11572 ( .A(n111), .B(n11738), .Z(n11743) );
  XNOR U11573 ( .A(n11742), .B(n11736), .Z(n11738) );
  XOR U11574 ( .A(n11744), .B(n11745), .Z(n11736) );
  AND U11575 ( .A(n126), .B(n11746), .Z(n11745) );
  XNOR U11576 ( .A(n11747), .B(n11748), .Z(n11742) );
  AND U11577 ( .A(n118), .B(n11749), .Z(n11748) );
  XOR U11578 ( .A(p_input[177]), .B(n11747), .Z(n11749) );
  XNOR U11579 ( .A(n11750), .B(n11751), .Z(n11747) );
  AND U11580 ( .A(n122), .B(n11746), .Z(n11751) );
  XNOR U11581 ( .A(n11750), .B(n11744), .Z(n11746) );
  XOR U11582 ( .A(n11752), .B(n11753), .Z(n11744) );
  AND U11583 ( .A(n137), .B(n11754), .Z(n11753) );
  XNOR U11584 ( .A(n11755), .B(n11756), .Z(n11750) );
  AND U11585 ( .A(n129), .B(n11757), .Z(n11756) );
  XOR U11586 ( .A(p_input[209]), .B(n11755), .Z(n11757) );
  XNOR U11587 ( .A(n11758), .B(n11759), .Z(n11755) );
  AND U11588 ( .A(n133), .B(n11754), .Z(n11759) );
  XNOR U11589 ( .A(n11758), .B(n11752), .Z(n11754) );
  XOR U11590 ( .A(n11760), .B(n11761), .Z(n11752) );
  AND U11591 ( .A(n148), .B(n11762), .Z(n11761) );
  XNOR U11592 ( .A(n11763), .B(n11764), .Z(n11758) );
  AND U11593 ( .A(n140), .B(n11765), .Z(n11764) );
  XOR U11594 ( .A(p_input[241]), .B(n11763), .Z(n11765) );
  XNOR U11595 ( .A(n11766), .B(n11767), .Z(n11763) );
  AND U11596 ( .A(n144), .B(n11762), .Z(n11767) );
  XNOR U11597 ( .A(n11766), .B(n11760), .Z(n11762) );
  XOR U11598 ( .A(n11768), .B(n11769), .Z(n11760) );
  AND U11599 ( .A(n159), .B(n11770), .Z(n11769) );
  XNOR U11600 ( .A(n11771), .B(n11772), .Z(n11766) );
  AND U11601 ( .A(n151), .B(n11773), .Z(n11772) );
  XOR U11602 ( .A(p_input[273]), .B(n11771), .Z(n11773) );
  XNOR U11603 ( .A(n11774), .B(n11775), .Z(n11771) );
  AND U11604 ( .A(n155), .B(n11770), .Z(n11775) );
  XNOR U11605 ( .A(n11774), .B(n11768), .Z(n11770) );
  XOR U11606 ( .A(n11776), .B(n11777), .Z(n11768) );
  AND U11607 ( .A(n170), .B(n11778), .Z(n11777) );
  XNOR U11608 ( .A(n11779), .B(n11780), .Z(n11774) );
  AND U11609 ( .A(n162), .B(n11781), .Z(n11780) );
  XOR U11610 ( .A(p_input[305]), .B(n11779), .Z(n11781) );
  XNOR U11611 ( .A(n11782), .B(n11783), .Z(n11779) );
  AND U11612 ( .A(n166), .B(n11778), .Z(n11783) );
  XNOR U11613 ( .A(n11782), .B(n11776), .Z(n11778) );
  XOR U11614 ( .A(n11784), .B(n11785), .Z(n11776) );
  AND U11615 ( .A(n181), .B(n11786), .Z(n11785) );
  XNOR U11616 ( .A(n11787), .B(n11788), .Z(n11782) );
  AND U11617 ( .A(n173), .B(n11789), .Z(n11788) );
  XOR U11618 ( .A(p_input[337]), .B(n11787), .Z(n11789) );
  XNOR U11619 ( .A(n11790), .B(n11791), .Z(n11787) );
  AND U11620 ( .A(n177), .B(n11786), .Z(n11791) );
  XNOR U11621 ( .A(n11790), .B(n11784), .Z(n11786) );
  XOR U11622 ( .A(n11792), .B(n11793), .Z(n11784) );
  AND U11623 ( .A(n192), .B(n11794), .Z(n11793) );
  XNOR U11624 ( .A(n11795), .B(n11796), .Z(n11790) );
  AND U11625 ( .A(n184), .B(n11797), .Z(n11796) );
  XOR U11626 ( .A(p_input[369]), .B(n11795), .Z(n11797) );
  XNOR U11627 ( .A(n11798), .B(n11799), .Z(n11795) );
  AND U11628 ( .A(n188), .B(n11794), .Z(n11799) );
  XNOR U11629 ( .A(n11798), .B(n11792), .Z(n11794) );
  XOR U11630 ( .A(n11800), .B(n11801), .Z(n11792) );
  AND U11631 ( .A(n203), .B(n11802), .Z(n11801) );
  XNOR U11632 ( .A(n11803), .B(n11804), .Z(n11798) );
  AND U11633 ( .A(n195), .B(n11805), .Z(n11804) );
  XOR U11634 ( .A(p_input[401]), .B(n11803), .Z(n11805) );
  XNOR U11635 ( .A(n11806), .B(n11807), .Z(n11803) );
  AND U11636 ( .A(n199), .B(n11802), .Z(n11807) );
  XNOR U11637 ( .A(n11806), .B(n11800), .Z(n11802) );
  XOR U11638 ( .A(n11808), .B(n11809), .Z(n11800) );
  AND U11639 ( .A(n214), .B(n11810), .Z(n11809) );
  XNOR U11640 ( .A(n11811), .B(n11812), .Z(n11806) );
  AND U11641 ( .A(n206), .B(n11813), .Z(n11812) );
  XOR U11642 ( .A(p_input[433]), .B(n11811), .Z(n11813) );
  XNOR U11643 ( .A(n11814), .B(n11815), .Z(n11811) );
  AND U11644 ( .A(n210), .B(n11810), .Z(n11815) );
  XNOR U11645 ( .A(n11814), .B(n11808), .Z(n11810) );
  XOR U11646 ( .A(n11816), .B(n11817), .Z(n11808) );
  AND U11647 ( .A(n225), .B(n11818), .Z(n11817) );
  XNOR U11648 ( .A(n11819), .B(n11820), .Z(n11814) );
  AND U11649 ( .A(n217), .B(n11821), .Z(n11820) );
  XOR U11650 ( .A(p_input[465]), .B(n11819), .Z(n11821) );
  XNOR U11651 ( .A(n11822), .B(n11823), .Z(n11819) );
  AND U11652 ( .A(n221), .B(n11818), .Z(n11823) );
  XNOR U11653 ( .A(n11822), .B(n11816), .Z(n11818) );
  XOR U11654 ( .A(n11824), .B(n11825), .Z(n11816) );
  AND U11655 ( .A(n236), .B(n11826), .Z(n11825) );
  XNOR U11656 ( .A(n11827), .B(n11828), .Z(n11822) );
  AND U11657 ( .A(n228), .B(n11829), .Z(n11828) );
  XOR U11658 ( .A(p_input[497]), .B(n11827), .Z(n11829) );
  XNOR U11659 ( .A(n11830), .B(n11831), .Z(n11827) );
  AND U11660 ( .A(n232), .B(n11826), .Z(n11831) );
  XNOR U11661 ( .A(n11830), .B(n11824), .Z(n11826) );
  XOR U11662 ( .A(n11832), .B(n11833), .Z(n11824) );
  AND U11663 ( .A(n247), .B(n11834), .Z(n11833) );
  XNOR U11664 ( .A(n11835), .B(n11836), .Z(n11830) );
  AND U11665 ( .A(n239), .B(n11837), .Z(n11836) );
  XOR U11666 ( .A(p_input[529]), .B(n11835), .Z(n11837) );
  XNOR U11667 ( .A(n11838), .B(n11839), .Z(n11835) );
  AND U11668 ( .A(n243), .B(n11834), .Z(n11839) );
  XNOR U11669 ( .A(n11838), .B(n11832), .Z(n11834) );
  XOR U11670 ( .A(n11840), .B(n11841), .Z(n11832) );
  AND U11671 ( .A(n258), .B(n11842), .Z(n11841) );
  XNOR U11672 ( .A(n11843), .B(n11844), .Z(n11838) );
  AND U11673 ( .A(n250), .B(n11845), .Z(n11844) );
  XOR U11674 ( .A(p_input[561]), .B(n11843), .Z(n11845) );
  XNOR U11675 ( .A(n11846), .B(n11847), .Z(n11843) );
  AND U11676 ( .A(n254), .B(n11842), .Z(n11847) );
  XNOR U11677 ( .A(n11846), .B(n11840), .Z(n11842) );
  XOR U11678 ( .A(n11848), .B(n11849), .Z(n11840) );
  AND U11679 ( .A(n269), .B(n11850), .Z(n11849) );
  XNOR U11680 ( .A(n11851), .B(n11852), .Z(n11846) );
  AND U11681 ( .A(n261), .B(n11853), .Z(n11852) );
  XOR U11682 ( .A(p_input[593]), .B(n11851), .Z(n11853) );
  XNOR U11683 ( .A(n11854), .B(n11855), .Z(n11851) );
  AND U11684 ( .A(n265), .B(n11850), .Z(n11855) );
  XNOR U11685 ( .A(n11854), .B(n11848), .Z(n11850) );
  XOR U11686 ( .A(n11856), .B(n11857), .Z(n11848) );
  AND U11687 ( .A(n280), .B(n11858), .Z(n11857) );
  XNOR U11688 ( .A(n11859), .B(n11860), .Z(n11854) );
  AND U11689 ( .A(n272), .B(n11861), .Z(n11860) );
  XOR U11690 ( .A(p_input[625]), .B(n11859), .Z(n11861) );
  XNOR U11691 ( .A(n11862), .B(n11863), .Z(n11859) );
  AND U11692 ( .A(n276), .B(n11858), .Z(n11863) );
  XNOR U11693 ( .A(n11862), .B(n11856), .Z(n11858) );
  XOR U11694 ( .A(n11864), .B(n11865), .Z(n11856) );
  AND U11695 ( .A(n291), .B(n11866), .Z(n11865) );
  XNOR U11696 ( .A(n11867), .B(n11868), .Z(n11862) );
  AND U11697 ( .A(n283), .B(n11869), .Z(n11868) );
  XOR U11698 ( .A(p_input[657]), .B(n11867), .Z(n11869) );
  XNOR U11699 ( .A(n11870), .B(n11871), .Z(n11867) );
  AND U11700 ( .A(n287), .B(n11866), .Z(n11871) );
  XNOR U11701 ( .A(n11870), .B(n11864), .Z(n11866) );
  XOR U11702 ( .A(n11872), .B(n11873), .Z(n11864) );
  AND U11703 ( .A(n302), .B(n11874), .Z(n11873) );
  XNOR U11704 ( .A(n11875), .B(n11876), .Z(n11870) );
  AND U11705 ( .A(n294), .B(n11877), .Z(n11876) );
  XOR U11706 ( .A(p_input[689]), .B(n11875), .Z(n11877) );
  XNOR U11707 ( .A(n11878), .B(n11879), .Z(n11875) );
  AND U11708 ( .A(n298), .B(n11874), .Z(n11879) );
  XNOR U11709 ( .A(n11878), .B(n11872), .Z(n11874) );
  XOR U11710 ( .A(n11880), .B(n11881), .Z(n11872) );
  AND U11711 ( .A(n313), .B(n11882), .Z(n11881) );
  XNOR U11712 ( .A(n11883), .B(n11884), .Z(n11878) );
  AND U11713 ( .A(n305), .B(n11885), .Z(n11884) );
  XOR U11714 ( .A(p_input[721]), .B(n11883), .Z(n11885) );
  XNOR U11715 ( .A(n11886), .B(n11887), .Z(n11883) );
  AND U11716 ( .A(n309), .B(n11882), .Z(n11887) );
  XNOR U11717 ( .A(n11886), .B(n11880), .Z(n11882) );
  XOR U11718 ( .A(n11888), .B(n11889), .Z(n11880) );
  AND U11719 ( .A(n324), .B(n11890), .Z(n11889) );
  XNOR U11720 ( .A(n11891), .B(n11892), .Z(n11886) );
  AND U11721 ( .A(n316), .B(n11893), .Z(n11892) );
  XOR U11722 ( .A(p_input[753]), .B(n11891), .Z(n11893) );
  XNOR U11723 ( .A(n11894), .B(n11895), .Z(n11891) );
  AND U11724 ( .A(n320), .B(n11890), .Z(n11895) );
  XNOR U11725 ( .A(n11894), .B(n11888), .Z(n11890) );
  XOR U11726 ( .A(n11896), .B(n11897), .Z(n11888) );
  AND U11727 ( .A(n335), .B(n11898), .Z(n11897) );
  XNOR U11728 ( .A(n11899), .B(n11900), .Z(n11894) );
  AND U11729 ( .A(n327), .B(n11901), .Z(n11900) );
  XOR U11730 ( .A(p_input[785]), .B(n11899), .Z(n11901) );
  XNOR U11731 ( .A(n11902), .B(n11903), .Z(n11899) );
  AND U11732 ( .A(n331), .B(n11898), .Z(n11903) );
  XNOR U11733 ( .A(n11902), .B(n11896), .Z(n11898) );
  XOR U11734 ( .A(n11904), .B(n11905), .Z(n11896) );
  AND U11735 ( .A(n346), .B(n11906), .Z(n11905) );
  XNOR U11736 ( .A(n11907), .B(n11908), .Z(n11902) );
  AND U11737 ( .A(n338), .B(n11909), .Z(n11908) );
  XOR U11738 ( .A(p_input[817]), .B(n11907), .Z(n11909) );
  XNOR U11739 ( .A(n11910), .B(n11911), .Z(n11907) );
  AND U11740 ( .A(n342), .B(n11906), .Z(n11911) );
  XNOR U11741 ( .A(n11910), .B(n11904), .Z(n11906) );
  XOR U11742 ( .A(n11912), .B(n11913), .Z(n11904) );
  AND U11743 ( .A(n357), .B(n11914), .Z(n11913) );
  XNOR U11744 ( .A(n11915), .B(n11916), .Z(n11910) );
  AND U11745 ( .A(n349), .B(n11917), .Z(n11916) );
  XOR U11746 ( .A(p_input[849]), .B(n11915), .Z(n11917) );
  XNOR U11747 ( .A(n11918), .B(n11919), .Z(n11915) );
  AND U11748 ( .A(n353), .B(n11914), .Z(n11919) );
  XNOR U11749 ( .A(n11918), .B(n11912), .Z(n11914) );
  XOR U11750 ( .A(n11920), .B(n11921), .Z(n11912) );
  AND U11751 ( .A(n368), .B(n11922), .Z(n11921) );
  XNOR U11752 ( .A(n11923), .B(n11924), .Z(n11918) );
  AND U11753 ( .A(n360), .B(n11925), .Z(n11924) );
  XOR U11754 ( .A(p_input[881]), .B(n11923), .Z(n11925) );
  XNOR U11755 ( .A(n11926), .B(n11927), .Z(n11923) );
  AND U11756 ( .A(n364), .B(n11922), .Z(n11927) );
  XNOR U11757 ( .A(n11926), .B(n11920), .Z(n11922) );
  XOR U11758 ( .A(n11928), .B(n11929), .Z(n11920) );
  AND U11759 ( .A(n379), .B(n11930), .Z(n11929) );
  XNOR U11760 ( .A(n11931), .B(n11932), .Z(n11926) );
  AND U11761 ( .A(n371), .B(n11933), .Z(n11932) );
  XOR U11762 ( .A(p_input[913]), .B(n11931), .Z(n11933) );
  XNOR U11763 ( .A(n11934), .B(n11935), .Z(n11931) );
  AND U11764 ( .A(n375), .B(n11930), .Z(n11935) );
  XNOR U11765 ( .A(n11934), .B(n11928), .Z(n11930) );
  XOR U11766 ( .A(n11936), .B(n11937), .Z(n11928) );
  AND U11767 ( .A(n390), .B(n11938), .Z(n11937) );
  XNOR U11768 ( .A(n11939), .B(n11940), .Z(n11934) );
  AND U11769 ( .A(n382), .B(n11941), .Z(n11940) );
  XOR U11770 ( .A(p_input[945]), .B(n11939), .Z(n11941) );
  XNOR U11771 ( .A(n11942), .B(n11943), .Z(n11939) );
  AND U11772 ( .A(n386), .B(n11938), .Z(n11943) );
  XNOR U11773 ( .A(n11942), .B(n11936), .Z(n11938) );
  XOR U11774 ( .A(n11944), .B(n11945), .Z(n11936) );
  AND U11775 ( .A(n401), .B(n11946), .Z(n11945) );
  XNOR U11776 ( .A(n11947), .B(n11948), .Z(n11942) );
  AND U11777 ( .A(n393), .B(n11949), .Z(n11948) );
  XOR U11778 ( .A(p_input[977]), .B(n11947), .Z(n11949) );
  XNOR U11779 ( .A(n11950), .B(n11951), .Z(n11947) );
  AND U11780 ( .A(n397), .B(n11946), .Z(n11951) );
  XNOR U11781 ( .A(n11950), .B(n11944), .Z(n11946) );
  XOR U11782 ( .A(n11952), .B(n11953), .Z(n11944) );
  AND U11783 ( .A(n412), .B(n11954), .Z(n11953) );
  XNOR U11784 ( .A(n11955), .B(n11956), .Z(n11950) );
  AND U11785 ( .A(n404), .B(n11957), .Z(n11956) );
  XOR U11786 ( .A(p_input[1009]), .B(n11955), .Z(n11957) );
  XNOR U11787 ( .A(n11958), .B(n11959), .Z(n11955) );
  AND U11788 ( .A(n408), .B(n11954), .Z(n11959) );
  XNOR U11789 ( .A(n11958), .B(n11952), .Z(n11954) );
  XOR U11790 ( .A(n11960), .B(n11961), .Z(n11952) );
  AND U11791 ( .A(n423), .B(n11962), .Z(n11961) );
  XNOR U11792 ( .A(n11963), .B(n11964), .Z(n11958) );
  AND U11793 ( .A(n415), .B(n11965), .Z(n11964) );
  XOR U11794 ( .A(p_input[1041]), .B(n11963), .Z(n11965) );
  XNOR U11795 ( .A(n11966), .B(n11967), .Z(n11963) );
  AND U11796 ( .A(n419), .B(n11962), .Z(n11967) );
  XNOR U11797 ( .A(n11966), .B(n11960), .Z(n11962) );
  XOR U11798 ( .A(n11968), .B(n11969), .Z(n11960) );
  AND U11799 ( .A(n434), .B(n11970), .Z(n11969) );
  XNOR U11800 ( .A(n11971), .B(n11972), .Z(n11966) );
  AND U11801 ( .A(n426), .B(n11973), .Z(n11972) );
  XOR U11802 ( .A(p_input[1073]), .B(n11971), .Z(n11973) );
  XNOR U11803 ( .A(n11974), .B(n11975), .Z(n11971) );
  AND U11804 ( .A(n430), .B(n11970), .Z(n11975) );
  XNOR U11805 ( .A(n11974), .B(n11968), .Z(n11970) );
  XOR U11806 ( .A(n11976), .B(n11977), .Z(n11968) );
  AND U11807 ( .A(n445), .B(n11978), .Z(n11977) );
  XNOR U11808 ( .A(n11979), .B(n11980), .Z(n11974) );
  AND U11809 ( .A(n437), .B(n11981), .Z(n11980) );
  XOR U11810 ( .A(p_input[1105]), .B(n11979), .Z(n11981) );
  XNOR U11811 ( .A(n11982), .B(n11983), .Z(n11979) );
  AND U11812 ( .A(n441), .B(n11978), .Z(n11983) );
  XNOR U11813 ( .A(n11982), .B(n11976), .Z(n11978) );
  XOR U11814 ( .A(n11984), .B(n11985), .Z(n11976) );
  AND U11815 ( .A(n456), .B(n11986), .Z(n11985) );
  XNOR U11816 ( .A(n11987), .B(n11988), .Z(n11982) );
  AND U11817 ( .A(n448), .B(n11989), .Z(n11988) );
  XOR U11818 ( .A(p_input[1137]), .B(n11987), .Z(n11989) );
  XNOR U11819 ( .A(n11990), .B(n11991), .Z(n11987) );
  AND U11820 ( .A(n452), .B(n11986), .Z(n11991) );
  XNOR U11821 ( .A(n11990), .B(n11984), .Z(n11986) );
  XOR U11822 ( .A(n11992), .B(n11993), .Z(n11984) );
  AND U11823 ( .A(n467), .B(n11994), .Z(n11993) );
  XNOR U11824 ( .A(n11995), .B(n11996), .Z(n11990) );
  AND U11825 ( .A(n459), .B(n11997), .Z(n11996) );
  XOR U11826 ( .A(p_input[1169]), .B(n11995), .Z(n11997) );
  XNOR U11827 ( .A(n11998), .B(n11999), .Z(n11995) );
  AND U11828 ( .A(n463), .B(n11994), .Z(n11999) );
  XNOR U11829 ( .A(n11998), .B(n11992), .Z(n11994) );
  XOR U11830 ( .A(n12000), .B(n12001), .Z(n11992) );
  AND U11831 ( .A(n478), .B(n12002), .Z(n12001) );
  XNOR U11832 ( .A(n12003), .B(n12004), .Z(n11998) );
  AND U11833 ( .A(n470), .B(n12005), .Z(n12004) );
  XOR U11834 ( .A(p_input[1201]), .B(n12003), .Z(n12005) );
  XNOR U11835 ( .A(n12006), .B(n12007), .Z(n12003) );
  AND U11836 ( .A(n474), .B(n12002), .Z(n12007) );
  XNOR U11837 ( .A(n12006), .B(n12000), .Z(n12002) );
  XOR U11838 ( .A(n12008), .B(n12009), .Z(n12000) );
  AND U11839 ( .A(n489), .B(n12010), .Z(n12009) );
  XNOR U11840 ( .A(n12011), .B(n12012), .Z(n12006) );
  AND U11841 ( .A(n481), .B(n12013), .Z(n12012) );
  XOR U11842 ( .A(p_input[1233]), .B(n12011), .Z(n12013) );
  XNOR U11843 ( .A(n12014), .B(n12015), .Z(n12011) );
  AND U11844 ( .A(n485), .B(n12010), .Z(n12015) );
  XNOR U11845 ( .A(n12014), .B(n12008), .Z(n12010) );
  XOR U11846 ( .A(n12016), .B(n12017), .Z(n12008) );
  AND U11847 ( .A(n500), .B(n12018), .Z(n12017) );
  XNOR U11848 ( .A(n12019), .B(n12020), .Z(n12014) );
  AND U11849 ( .A(n492), .B(n12021), .Z(n12020) );
  XOR U11850 ( .A(p_input[1265]), .B(n12019), .Z(n12021) );
  XNOR U11851 ( .A(n12022), .B(n12023), .Z(n12019) );
  AND U11852 ( .A(n496), .B(n12018), .Z(n12023) );
  XNOR U11853 ( .A(n12022), .B(n12016), .Z(n12018) );
  XOR U11854 ( .A(n12024), .B(n12025), .Z(n12016) );
  AND U11855 ( .A(n511), .B(n12026), .Z(n12025) );
  XNOR U11856 ( .A(n12027), .B(n12028), .Z(n12022) );
  AND U11857 ( .A(n503), .B(n12029), .Z(n12028) );
  XOR U11858 ( .A(p_input[1297]), .B(n12027), .Z(n12029) );
  XNOR U11859 ( .A(n12030), .B(n12031), .Z(n12027) );
  AND U11860 ( .A(n507), .B(n12026), .Z(n12031) );
  XNOR U11861 ( .A(n12030), .B(n12024), .Z(n12026) );
  XOR U11862 ( .A(n12032), .B(n12033), .Z(n12024) );
  AND U11863 ( .A(n522), .B(n12034), .Z(n12033) );
  XNOR U11864 ( .A(n12035), .B(n12036), .Z(n12030) );
  AND U11865 ( .A(n514), .B(n12037), .Z(n12036) );
  XOR U11866 ( .A(p_input[1329]), .B(n12035), .Z(n12037) );
  XNOR U11867 ( .A(n12038), .B(n12039), .Z(n12035) );
  AND U11868 ( .A(n518), .B(n12034), .Z(n12039) );
  XNOR U11869 ( .A(n12038), .B(n12032), .Z(n12034) );
  XOR U11870 ( .A(n12040), .B(n12041), .Z(n12032) );
  AND U11871 ( .A(n533), .B(n12042), .Z(n12041) );
  XNOR U11872 ( .A(n12043), .B(n12044), .Z(n12038) );
  AND U11873 ( .A(n525), .B(n12045), .Z(n12044) );
  XOR U11874 ( .A(p_input[1361]), .B(n12043), .Z(n12045) );
  XNOR U11875 ( .A(n12046), .B(n12047), .Z(n12043) );
  AND U11876 ( .A(n529), .B(n12042), .Z(n12047) );
  XNOR U11877 ( .A(n12046), .B(n12040), .Z(n12042) );
  XOR U11878 ( .A(n12048), .B(n12049), .Z(n12040) );
  AND U11879 ( .A(n544), .B(n12050), .Z(n12049) );
  XNOR U11880 ( .A(n12051), .B(n12052), .Z(n12046) );
  AND U11881 ( .A(n536), .B(n12053), .Z(n12052) );
  XOR U11882 ( .A(p_input[1393]), .B(n12051), .Z(n12053) );
  XNOR U11883 ( .A(n12054), .B(n12055), .Z(n12051) );
  AND U11884 ( .A(n540), .B(n12050), .Z(n12055) );
  XNOR U11885 ( .A(n12054), .B(n12048), .Z(n12050) );
  XOR U11886 ( .A(n12056), .B(n12057), .Z(n12048) );
  AND U11887 ( .A(n555), .B(n12058), .Z(n12057) );
  XNOR U11888 ( .A(n12059), .B(n12060), .Z(n12054) );
  AND U11889 ( .A(n547), .B(n12061), .Z(n12060) );
  XOR U11890 ( .A(p_input[1425]), .B(n12059), .Z(n12061) );
  XNOR U11891 ( .A(n12062), .B(n12063), .Z(n12059) );
  AND U11892 ( .A(n551), .B(n12058), .Z(n12063) );
  XNOR U11893 ( .A(n12062), .B(n12056), .Z(n12058) );
  XOR U11894 ( .A(n12064), .B(n12065), .Z(n12056) );
  AND U11895 ( .A(n566), .B(n12066), .Z(n12065) );
  XNOR U11896 ( .A(n12067), .B(n12068), .Z(n12062) );
  AND U11897 ( .A(n558), .B(n12069), .Z(n12068) );
  XOR U11898 ( .A(p_input[1457]), .B(n12067), .Z(n12069) );
  XNOR U11899 ( .A(n12070), .B(n12071), .Z(n12067) );
  AND U11900 ( .A(n562), .B(n12066), .Z(n12071) );
  XNOR U11901 ( .A(n12070), .B(n12064), .Z(n12066) );
  XOR U11902 ( .A(n12072), .B(n12073), .Z(n12064) );
  AND U11903 ( .A(n577), .B(n12074), .Z(n12073) );
  XNOR U11904 ( .A(n12075), .B(n12076), .Z(n12070) );
  AND U11905 ( .A(n569), .B(n12077), .Z(n12076) );
  XOR U11906 ( .A(p_input[1489]), .B(n12075), .Z(n12077) );
  XNOR U11907 ( .A(n12078), .B(n12079), .Z(n12075) );
  AND U11908 ( .A(n573), .B(n12074), .Z(n12079) );
  XNOR U11909 ( .A(n12078), .B(n12072), .Z(n12074) );
  XOR U11910 ( .A(n12080), .B(n12081), .Z(n12072) );
  AND U11911 ( .A(n588), .B(n12082), .Z(n12081) );
  XNOR U11912 ( .A(n12083), .B(n12084), .Z(n12078) );
  AND U11913 ( .A(n580), .B(n12085), .Z(n12084) );
  XOR U11914 ( .A(p_input[1521]), .B(n12083), .Z(n12085) );
  XNOR U11915 ( .A(n12086), .B(n12087), .Z(n12083) );
  AND U11916 ( .A(n584), .B(n12082), .Z(n12087) );
  XNOR U11917 ( .A(n12086), .B(n12080), .Z(n12082) );
  XOR U11918 ( .A(n12088), .B(n12089), .Z(n12080) );
  AND U11919 ( .A(n599), .B(n12090), .Z(n12089) );
  XNOR U11920 ( .A(n12091), .B(n12092), .Z(n12086) );
  AND U11921 ( .A(n591), .B(n12093), .Z(n12092) );
  XOR U11922 ( .A(p_input[1553]), .B(n12091), .Z(n12093) );
  XNOR U11923 ( .A(n12094), .B(n12095), .Z(n12091) );
  AND U11924 ( .A(n595), .B(n12090), .Z(n12095) );
  XNOR U11925 ( .A(n12094), .B(n12088), .Z(n12090) );
  XOR U11926 ( .A(n12096), .B(n12097), .Z(n12088) );
  AND U11927 ( .A(n610), .B(n12098), .Z(n12097) );
  XNOR U11928 ( .A(n12099), .B(n12100), .Z(n12094) );
  AND U11929 ( .A(n602), .B(n12101), .Z(n12100) );
  XOR U11930 ( .A(p_input[1585]), .B(n12099), .Z(n12101) );
  XNOR U11931 ( .A(n12102), .B(n12103), .Z(n12099) );
  AND U11932 ( .A(n606), .B(n12098), .Z(n12103) );
  XNOR U11933 ( .A(n12102), .B(n12096), .Z(n12098) );
  XOR U11934 ( .A(n12104), .B(n12105), .Z(n12096) );
  AND U11935 ( .A(n621), .B(n12106), .Z(n12105) );
  XNOR U11936 ( .A(n12107), .B(n12108), .Z(n12102) );
  AND U11937 ( .A(n613), .B(n12109), .Z(n12108) );
  XOR U11938 ( .A(p_input[1617]), .B(n12107), .Z(n12109) );
  XNOR U11939 ( .A(n12110), .B(n12111), .Z(n12107) );
  AND U11940 ( .A(n617), .B(n12106), .Z(n12111) );
  XNOR U11941 ( .A(n12110), .B(n12104), .Z(n12106) );
  XOR U11942 ( .A(n12112), .B(n12113), .Z(n12104) );
  AND U11943 ( .A(n632), .B(n12114), .Z(n12113) );
  XNOR U11944 ( .A(n12115), .B(n12116), .Z(n12110) );
  AND U11945 ( .A(n624), .B(n12117), .Z(n12116) );
  XOR U11946 ( .A(p_input[1649]), .B(n12115), .Z(n12117) );
  XNOR U11947 ( .A(n12118), .B(n12119), .Z(n12115) );
  AND U11948 ( .A(n628), .B(n12114), .Z(n12119) );
  XNOR U11949 ( .A(n12118), .B(n12112), .Z(n12114) );
  XOR U11950 ( .A(n12120), .B(n12121), .Z(n12112) );
  AND U11951 ( .A(n643), .B(n12122), .Z(n12121) );
  XNOR U11952 ( .A(n12123), .B(n12124), .Z(n12118) );
  AND U11953 ( .A(n635), .B(n12125), .Z(n12124) );
  XOR U11954 ( .A(p_input[1681]), .B(n12123), .Z(n12125) );
  XNOR U11955 ( .A(n12126), .B(n12127), .Z(n12123) );
  AND U11956 ( .A(n639), .B(n12122), .Z(n12127) );
  XNOR U11957 ( .A(n12126), .B(n12120), .Z(n12122) );
  XOR U11958 ( .A(n12128), .B(n12129), .Z(n12120) );
  AND U11959 ( .A(n654), .B(n12130), .Z(n12129) );
  XNOR U11960 ( .A(n12131), .B(n12132), .Z(n12126) );
  AND U11961 ( .A(n646), .B(n12133), .Z(n12132) );
  XOR U11962 ( .A(p_input[1713]), .B(n12131), .Z(n12133) );
  XNOR U11963 ( .A(n12134), .B(n12135), .Z(n12131) );
  AND U11964 ( .A(n650), .B(n12130), .Z(n12135) );
  XNOR U11965 ( .A(n12134), .B(n12128), .Z(n12130) );
  XOR U11966 ( .A(n12136), .B(n12137), .Z(n12128) );
  AND U11967 ( .A(n665), .B(n12138), .Z(n12137) );
  XNOR U11968 ( .A(n12139), .B(n12140), .Z(n12134) );
  AND U11969 ( .A(n657), .B(n12141), .Z(n12140) );
  XOR U11970 ( .A(p_input[1745]), .B(n12139), .Z(n12141) );
  XNOR U11971 ( .A(n12142), .B(n12143), .Z(n12139) );
  AND U11972 ( .A(n661), .B(n12138), .Z(n12143) );
  XNOR U11973 ( .A(n12142), .B(n12136), .Z(n12138) );
  XOR U11974 ( .A(n12144), .B(n12145), .Z(n12136) );
  AND U11975 ( .A(n676), .B(n12146), .Z(n12145) );
  XNOR U11976 ( .A(n12147), .B(n12148), .Z(n12142) );
  AND U11977 ( .A(n668), .B(n12149), .Z(n12148) );
  XOR U11978 ( .A(p_input[1777]), .B(n12147), .Z(n12149) );
  XNOR U11979 ( .A(n12150), .B(n12151), .Z(n12147) );
  AND U11980 ( .A(n672), .B(n12146), .Z(n12151) );
  XNOR U11981 ( .A(n12150), .B(n12144), .Z(n12146) );
  XOR U11982 ( .A(n12152), .B(n12153), .Z(n12144) );
  AND U11983 ( .A(n687), .B(n12154), .Z(n12153) );
  XNOR U11984 ( .A(n12155), .B(n12156), .Z(n12150) );
  AND U11985 ( .A(n679), .B(n12157), .Z(n12156) );
  XOR U11986 ( .A(p_input[1809]), .B(n12155), .Z(n12157) );
  XNOR U11987 ( .A(n12158), .B(n12159), .Z(n12155) );
  AND U11988 ( .A(n683), .B(n12154), .Z(n12159) );
  XNOR U11989 ( .A(n12158), .B(n12152), .Z(n12154) );
  XOR U11990 ( .A(n12160), .B(n12161), .Z(n12152) );
  AND U11991 ( .A(n698), .B(n12162), .Z(n12161) );
  XNOR U11992 ( .A(n12163), .B(n12164), .Z(n12158) );
  AND U11993 ( .A(n690), .B(n12165), .Z(n12164) );
  XOR U11994 ( .A(p_input[1841]), .B(n12163), .Z(n12165) );
  XNOR U11995 ( .A(n12166), .B(n12167), .Z(n12163) );
  AND U11996 ( .A(n694), .B(n12162), .Z(n12167) );
  XNOR U11997 ( .A(n12166), .B(n12160), .Z(n12162) );
  XOR U11998 ( .A(n12168), .B(n12169), .Z(n12160) );
  AND U11999 ( .A(n709), .B(n12170), .Z(n12169) );
  XNOR U12000 ( .A(n12171), .B(n12172), .Z(n12166) );
  AND U12001 ( .A(n701), .B(n12173), .Z(n12172) );
  XOR U12002 ( .A(p_input[1873]), .B(n12171), .Z(n12173) );
  XNOR U12003 ( .A(n12174), .B(n12175), .Z(n12171) );
  AND U12004 ( .A(n705), .B(n12170), .Z(n12175) );
  XNOR U12005 ( .A(n12174), .B(n12168), .Z(n12170) );
  XOR U12006 ( .A(n12176), .B(n12177), .Z(n12168) );
  AND U12007 ( .A(n720), .B(n12178), .Z(n12177) );
  XNOR U12008 ( .A(n12179), .B(n12180), .Z(n12174) );
  AND U12009 ( .A(n712), .B(n12181), .Z(n12180) );
  XOR U12010 ( .A(p_input[1905]), .B(n12179), .Z(n12181) );
  XNOR U12011 ( .A(n12182), .B(n12183), .Z(n12179) );
  AND U12012 ( .A(n716), .B(n12178), .Z(n12183) );
  XNOR U12013 ( .A(n12182), .B(n12176), .Z(n12178) );
  XOR U12014 ( .A(n12184), .B(n12185), .Z(n12176) );
  AND U12015 ( .A(n731), .B(n12186), .Z(n12185) );
  XNOR U12016 ( .A(n12187), .B(n12188), .Z(n12182) );
  AND U12017 ( .A(n723), .B(n12189), .Z(n12188) );
  XOR U12018 ( .A(p_input[1937]), .B(n12187), .Z(n12189) );
  XNOR U12019 ( .A(n12190), .B(n12191), .Z(n12187) );
  AND U12020 ( .A(n727), .B(n12186), .Z(n12191) );
  XNOR U12021 ( .A(n12190), .B(n12184), .Z(n12186) );
  XOR U12022 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n12192), .Z(n12184) );
  AND U12023 ( .A(n741), .B(n12193), .Z(n12192) );
  XNOR U12024 ( .A(n12194), .B(n12195), .Z(n12190) );
  AND U12025 ( .A(n734), .B(n12196), .Z(n12195) );
  XOR U12026 ( .A(p_input[1969]), .B(n12194), .Z(n12196) );
  XNOR U12027 ( .A(n12197), .B(n12198), .Z(n12194) );
  AND U12028 ( .A(n738), .B(n12193), .Z(n12198) );
  XOR U12029 ( .A(\knn_comb_/min_val_out[0][17] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .Z(n12193) );
  XOR U12030 ( .A(n43), .B(n12199), .Z(o[16]) );
  AND U12031 ( .A(n58), .B(n12200), .Z(n43) );
  XOR U12032 ( .A(n44), .B(n12199), .Z(n12200) );
  XOR U12033 ( .A(n12201), .B(n12202), .Z(n12199) );
  AND U12034 ( .A(n70), .B(n12203), .Z(n12202) );
  XOR U12035 ( .A(n12204), .B(n12205), .Z(n44) );
  AND U12036 ( .A(n62), .B(n12206), .Z(n12205) );
  XOR U12037 ( .A(p_input[16]), .B(n12204), .Z(n12206) );
  XNOR U12038 ( .A(n12207), .B(n12208), .Z(n12204) );
  AND U12039 ( .A(n66), .B(n12203), .Z(n12208) );
  XNOR U12040 ( .A(n12207), .B(n12201), .Z(n12203) );
  XOR U12041 ( .A(n12209), .B(n12210), .Z(n12201) );
  AND U12042 ( .A(n82), .B(n12211), .Z(n12210) );
  XNOR U12043 ( .A(n12212), .B(n12213), .Z(n12207) );
  AND U12044 ( .A(n74), .B(n12214), .Z(n12213) );
  XOR U12045 ( .A(p_input[48]), .B(n12212), .Z(n12214) );
  XNOR U12046 ( .A(n12215), .B(n12216), .Z(n12212) );
  AND U12047 ( .A(n78), .B(n12211), .Z(n12216) );
  XNOR U12048 ( .A(n12215), .B(n12209), .Z(n12211) );
  XOR U12049 ( .A(n12217), .B(n12218), .Z(n12209) );
  AND U12050 ( .A(n93), .B(n12219), .Z(n12218) );
  XNOR U12051 ( .A(n12220), .B(n12221), .Z(n12215) );
  AND U12052 ( .A(n85), .B(n12222), .Z(n12221) );
  XOR U12053 ( .A(p_input[80]), .B(n12220), .Z(n12222) );
  XNOR U12054 ( .A(n12223), .B(n12224), .Z(n12220) );
  AND U12055 ( .A(n89), .B(n12219), .Z(n12224) );
  XNOR U12056 ( .A(n12223), .B(n12217), .Z(n12219) );
  XOR U12057 ( .A(n12225), .B(n12226), .Z(n12217) );
  AND U12058 ( .A(n104), .B(n12227), .Z(n12226) );
  XNOR U12059 ( .A(n12228), .B(n12229), .Z(n12223) );
  AND U12060 ( .A(n96), .B(n12230), .Z(n12229) );
  XOR U12061 ( .A(p_input[112]), .B(n12228), .Z(n12230) );
  XNOR U12062 ( .A(n12231), .B(n12232), .Z(n12228) );
  AND U12063 ( .A(n100), .B(n12227), .Z(n12232) );
  XNOR U12064 ( .A(n12231), .B(n12225), .Z(n12227) );
  XOR U12065 ( .A(n12233), .B(n12234), .Z(n12225) );
  AND U12066 ( .A(n115), .B(n12235), .Z(n12234) );
  XNOR U12067 ( .A(n12236), .B(n12237), .Z(n12231) );
  AND U12068 ( .A(n107), .B(n12238), .Z(n12237) );
  XOR U12069 ( .A(p_input[144]), .B(n12236), .Z(n12238) );
  XNOR U12070 ( .A(n12239), .B(n12240), .Z(n12236) );
  AND U12071 ( .A(n111), .B(n12235), .Z(n12240) );
  XNOR U12072 ( .A(n12239), .B(n12233), .Z(n12235) );
  XOR U12073 ( .A(n12241), .B(n12242), .Z(n12233) );
  AND U12074 ( .A(n126), .B(n12243), .Z(n12242) );
  XNOR U12075 ( .A(n12244), .B(n12245), .Z(n12239) );
  AND U12076 ( .A(n118), .B(n12246), .Z(n12245) );
  XOR U12077 ( .A(p_input[176]), .B(n12244), .Z(n12246) );
  XNOR U12078 ( .A(n12247), .B(n12248), .Z(n12244) );
  AND U12079 ( .A(n122), .B(n12243), .Z(n12248) );
  XNOR U12080 ( .A(n12247), .B(n12241), .Z(n12243) );
  XOR U12081 ( .A(n12249), .B(n12250), .Z(n12241) );
  AND U12082 ( .A(n137), .B(n12251), .Z(n12250) );
  XNOR U12083 ( .A(n12252), .B(n12253), .Z(n12247) );
  AND U12084 ( .A(n129), .B(n12254), .Z(n12253) );
  XOR U12085 ( .A(p_input[208]), .B(n12252), .Z(n12254) );
  XNOR U12086 ( .A(n12255), .B(n12256), .Z(n12252) );
  AND U12087 ( .A(n133), .B(n12251), .Z(n12256) );
  XNOR U12088 ( .A(n12255), .B(n12249), .Z(n12251) );
  XOR U12089 ( .A(n12257), .B(n12258), .Z(n12249) );
  AND U12090 ( .A(n148), .B(n12259), .Z(n12258) );
  XNOR U12091 ( .A(n12260), .B(n12261), .Z(n12255) );
  AND U12092 ( .A(n140), .B(n12262), .Z(n12261) );
  XOR U12093 ( .A(p_input[240]), .B(n12260), .Z(n12262) );
  XNOR U12094 ( .A(n12263), .B(n12264), .Z(n12260) );
  AND U12095 ( .A(n144), .B(n12259), .Z(n12264) );
  XNOR U12096 ( .A(n12263), .B(n12257), .Z(n12259) );
  XOR U12097 ( .A(n12265), .B(n12266), .Z(n12257) );
  AND U12098 ( .A(n159), .B(n12267), .Z(n12266) );
  XNOR U12099 ( .A(n12268), .B(n12269), .Z(n12263) );
  AND U12100 ( .A(n151), .B(n12270), .Z(n12269) );
  XOR U12101 ( .A(p_input[272]), .B(n12268), .Z(n12270) );
  XNOR U12102 ( .A(n12271), .B(n12272), .Z(n12268) );
  AND U12103 ( .A(n155), .B(n12267), .Z(n12272) );
  XNOR U12104 ( .A(n12271), .B(n12265), .Z(n12267) );
  XOR U12105 ( .A(n12273), .B(n12274), .Z(n12265) );
  AND U12106 ( .A(n170), .B(n12275), .Z(n12274) );
  XNOR U12107 ( .A(n12276), .B(n12277), .Z(n12271) );
  AND U12108 ( .A(n162), .B(n12278), .Z(n12277) );
  XOR U12109 ( .A(p_input[304]), .B(n12276), .Z(n12278) );
  XNOR U12110 ( .A(n12279), .B(n12280), .Z(n12276) );
  AND U12111 ( .A(n166), .B(n12275), .Z(n12280) );
  XNOR U12112 ( .A(n12279), .B(n12273), .Z(n12275) );
  XOR U12113 ( .A(n12281), .B(n12282), .Z(n12273) );
  AND U12114 ( .A(n181), .B(n12283), .Z(n12282) );
  XNOR U12115 ( .A(n12284), .B(n12285), .Z(n12279) );
  AND U12116 ( .A(n173), .B(n12286), .Z(n12285) );
  XOR U12117 ( .A(p_input[336]), .B(n12284), .Z(n12286) );
  XNOR U12118 ( .A(n12287), .B(n12288), .Z(n12284) );
  AND U12119 ( .A(n177), .B(n12283), .Z(n12288) );
  XNOR U12120 ( .A(n12287), .B(n12281), .Z(n12283) );
  XOR U12121 ( .A(n12289), .B(n12290), .Z(n12281) );
  AND U12122 ( .A(n192), .B(n12291), .Z(n12290) );
  XNOR U12123 ( .A(n12292), .B(n12293), .Z(n12287) );
  AND U12124 ( .A(n184), .B(n12294), .Z(n12293) );
  XOR U12125 ( .A(p_input[368]), .B(n12292), .Z(n12294) );
  XNOR U12126 ( .A(n12295), .B(n12296), .Z(n12292) );
  AND U12127 ( .A(n188), .B(n12291), .Z(n12296) );
  XNOR U12128 ( .A(n12295), .B(n12289), .Z(n12291) );
  XOR U12129 ( .A(n12297), .B(n12298), .Z(n12289) );
  AND U12130 ( .A(n203), .B(n12299), .Z(n12298) );
  XNOR U12131 ( .A(n12300), .B(n12301), .Z(n12295) );
  AND U12132 ( .A(n195), .B(n12302), .Z(n12301) );
  XOR U12133 ( .A(p_input[400]), .B(n12300), .Z(n12302) );
  XNOR U12134 ( .A(n12303), .B(n12304), .Z(n12300) );
  AND U12135 ( .A(n199), .B(n12299), .Z(n12304) );
  XNOR U12136 ( .A(n12303), .B(n12297), .Z(n12299) );
  XOR U12137 ( .A(n12305), .B(n12306), .Z(n12297) );
  AND U12138 ( .A(n214), .B(n12307), .Z(n12306) );
  XNOR U12139 ( .A(n12308), .B(n12309), .Z(n12303) );
  AND U12140 ( .A(n206), .B(n12310), .Z(n12309) );
  XOR U12141 ( .A(p_input[432]), .B(n12308), .Z(n12310) );
  XNOR U12142 ( .A(n12311), .B(n12312), .Z(n12308) );
  AND U12143 ( .A(n210), .B(n12307), .Z(n12312) );
  XNOR U12144 ( .A(n12311), .B(n12305), .Z(n12307) );
  XOR U12145 ( .A(n12313), .B(n12314), .Z(n12305) );
  AND U12146 ( .A(n225), .B(n12315), .Z(n12314) );
  XNOR U12147 ( .A(n12316), .B(n12317), .Z(n12311) );
  AND U12148 ( .A(n217), .B(n12318), .Z(n12317) );
  XOR U12149 ( .A(p_input[464]), .B(n12316), .Z(n12318) );
  XNOR U12150 ( .A(n12319), .B(n12320), .Z(n12316) );
  AND U12151 ( .A(n221), .B(n12315), .Z(n12320) );
  XNOR U12152 ( .A(n12319), .B(n12313), .Z(n12315) );
  XOR U12153 ( .A(n12321), .B(n12322), .Z(n12313) );
  AND U12154 ( .A(n236), .B(n12323), .Z(n12322) );
  XNOR U12155 ( .A(n12324), .B(n12325), .Z(n12319) );
  AND U12156 ( .A(n228), .B(n12326), .Z(n12325) );
  XOR U12157 ( .A(p_input[496]), .B(n12324), .Z(n12326) );
  XNOR U12158 ( .A(n12327), .B(n12328), .Z(n12324) );
  AND U12159 ( .A(n232), .B(n12323), .Z(n12328) );
  XNOR U12160 ( .A(n12327), .B(n12321), .Z(n12323) );
  XOR U12161 ( .A(n12329), .B(n12330), .Z(n12321) );
  AND U12162 ( .A(n247), .B(n12331), .Z(n12330) );
  XNOR U12163 ( .A(n12332), .B(n12333), .Z(n12327) );
  AND U12164 ( .A(n239), .B(n12334), .Z(n12333) );
  XOR U12165 ( .A(p_input[528]), .B(n12332), .Z(n12334) );
  XNOR U12166 ( .A(n12335), .B(n12336), .Z(n12332) );
  AND U12167 ( .A(n243), .B(n12331), .Z(n12336) );
  XNOR U12168 ( .A(n12335), .B(n12329), .Z(n12331) );
  XOR U12169 ( .A(n12337), .B(n12338), .Z(n12329) );
  AND U12170 ( .A(n258), .B(n12339), .Z(n12338) );
  XNOR U12171 ( .A(n12340), .B(n12341), .Z(n12335) );
  AND U12172 ( .A(n250), .B(n12342), .Z(n12341) );
  XOR U12173 ( .A(p_input[560]), .B(n12340), .Z(n12342) );
  XNOR U12174 ( .A(n12343), .B(n12344), .Z(n12340) );
  AND U12175 ( .A(n254), .B(n12339), .Z(n12344) );
  XNOR U12176 ( .A(n12343), .B(n12337), .Z(n12339) );
  XOR U12177 ( .A(n12345), .B(n12346), .Z(n12337) );
  AND U12178 ( .A(n269), .B(n12347), .Z(n12346) );
  XNOR U12179 ( .A(n12348), .B(n12349), .Z(n12343) );
  AND U12180 ( .A(n261), .B(n12350), .Z(n12349) );
  XOR U12181 ( .A(p_input[592]), .B(n12348), .Z(n12350) );
  XNOR U12182 ( .A(n12351), .B(n12352), .Z(n12348) );
  AND U12183 ( .A(n265), .B(n12347), .Z(n12352) );
  XNOR U12184 ( .A(n12351), .B(n12345), .Z(n12347) );
  XOR U12185 ( .A(n12353), .B(n12354), .Z(n12345) );
  AND U12186 ( .A(n280), .B(n12355), .Z(n12354) );
  XNOR U12187 ( .A(n12356), .B(n12357), .Z(n12351) );
  AND U12188 ( .A(n272), .B(n12358), .Z(n12357) );
  XOR U12189 ( .A(p_input[624]), .B(n12356), .Z(n12358) );
  XNOR U12190 ( .A(n12359), .B(n12360), .Z(n12356) );
  AND U12191 ( .A(n276), .B(n12355), .Z(n12360) );
  XNOR U12192 ( .A(n12359), .B(n12353), .Z(n12355) );
  XOR U12193 ( .A(n12361), .B(n12362), .Z(n12353) );
  AND U12194 ( .A(n291), .B(n12363), .Z(n12362) );
  XNOR U12195 ( .A(n12364), .B(n12365), .Z(n12359) );
  AND U12196 ( .A(n283), .B(n12366), .Z(n12365) );
  XOR U12197 ( .A(p_input[656]), .B(n12364), .Z(n12366) );
  XNOR U12198 ( .A(n12367), .B(n12368), .Z(n12364) );
  AND U12199 ( .A(n287), .B(n12363), .Z(n12368) );
  XNOR U12200 ( .A(n12367), .B(n12361), .Z(n12363) );
  XOR U12201 ( .A(n12369), .B(n12370), .Z(n12361) );
  AND U12202 ( .A(n302), .B(n12371), .Z(n12370) );
  XNOR U12203 ( .A(n12372), .B(n12373), .Z(n12367) );
  AND U12204 ( .A(n294), .B(n12374), .Z(n12373) );
  XOR U12205 ( .A(p_input[688]), .B(n12372), .Z(n12374) );
  XNOR U12206 ( .A(n12375), .B(n12376), .Z(n12372) );
  AND U12207 ( .A(n298), .B(n12371), .Z(n12376) );
  XNOR U12208 ( .A(n12375), .B(n12369), .Z(n12371) );
  XOR U12209 ( .A(n12377), .B(n12378), .Z(n12369) );
  AND U12210 ( .A(n313), .B(n12379), .Z(n12378) );
  XNOR U12211 ( .A(n12380), .B(n12381), .Z(n12375) );
  AND U12212 ( .A(n305), .B(n12382), .Z(n12381) );
  XOR U12213 ( .A(p_input[720]), .B(n12380), .Z(n12382) );
  XNOR U12214 ( .A(n12383), .B(n12384), .Z(n12380) );
  AND U12215 ( .A(n309), .B(n12379), .Z(n12384) );
  XNOR U12216 ( .A(n12383), .B(n12377), .Z(n12379) );
  XOR U12217 ( .A(n12385), .B(n12386), .Z(n12377) );
  AND U12218 ( .A(n324), .B(n12387), .Z(n12386) );
  XNOR U12219 ( .A(n12388), .B(n12389), .Z(n12383) );
  AND U12220 ( .A(n316), .B(n12390), .Z(n12389) );
  XOR U12221 ( .A(p_input[752]), .B(n12388), .Z(n12390) );
  XNOR U12222 ( .A(n12391), .B(n12392), .Z(n12388) );
  AND U12223 ( .A(n320), .B(n12387), .Z(n12392) );
  XNOR U12224 ( .A(n12391), .B(n12385), .Z(n12387) );
  XOR U12225 ( .A(n12393), .B(n12394), .Z(n12385) );
  AND U12226 ( .A(n335), .B(n12395), .Z(n12394) );
  XNOR U12227 ( .A(n12396), .B(n12397), .Z(n12391) );
  AND U12228 ( .A(n327), .B(n12398), .Z(n12397) );
  XOR U12229 ( .A(p_input[784]), .B(n12396), .Z(n12398) );
  XNOR U12230 ( .A(n12399), .B(n12400), .Z(n12396) );
  AND U12231 ( .A(n331), .B(n12395), .Z(n12400) );
  XNOR U12232 ( .A(n12399), .B(n12393), .Z(n12395) );
  XOR U12233 ( .A(n12401), .B(n12402), .Z(n12393) );
  AND U12234 ( .A(n346), .B(n12403), .Z(n12402) );
  XNOR U12235 ( .A(n12404), .B(n12405), .Z(n12399) );
  AND U12236 ( .A(n338), .B(n12406), .Z(n12405) );
  XOR U12237 ( .A(p_input[816]), .B(n12404), .Z(n12406) );
  XNOR U12238 ( .A(n12407), .B(n12408), .Z(n12404) );
  AND U12239 ( .A(n342), .B(n12403), .Z(n12408) );
  XNOR U12240 ( .A(n12407), .B(n12401), .Z(n12403) );
  XOR U12241 ( .A(n12409), .B(n12410), .Z(n12401) );
  AND U12242 ( .A(n357), .B(n12411), .Z(n12410) );
  XNOR U12243 ( .A(n12412), .B(n12413), .Z(n12407) );
  AND U12244 ( .A(n349), .B(n12414), .Z(n12413) );
  XOR U12245 ( .A(p_input[848]), .B(n12412), .Z(n12414) );
  XNOR U12246 ( .A(n12415), .B(n12416), .Z(n12412) );
  AND U12247 ( .A(n353), .B(n12411), .Z(n12416) );
  XNOR U12248 ( .A(n12415), .B(n12409), .Z(n12411) );
  XOR U12249 ( .A(n12417), .B(n12418), .Z(n12409) );
  AND U12250 ( .A(n368), .B(n12419), .Z(n12418) );
  XNOR U12251 ( .A(n12420), .B(n12421), .Z(n12415) );
  AND U12252 ( .A(n360), .B(n12422), .Z(n12421) );
  XOR U12253 ( .A(p_input[880]), .B(n12420), .Z(n12422) );
  XNOR U12254 ( .A(n12423), .B(n12424), .Z(n12420) );
  AND U12255 ( .A(n364), .B(n12419), .Z(n12424) );
  XNOR U12256 ( .A(n12423), .B(n12417), .Z(n12419) );
  XOR U12257 ( .A(n12425), .B(n12426), .Z(n12417) );
  AND U12258 ( .A(n379), .B(n12427), .Z(n12426) );
  XNOR U12259 ( .A(n12428), .B(n12429), .Z(n12423) );
  AND U12260 ( .A(n371), .B(n12430), .Z(n12429) );
  XOR U12261 ( .A(p_input[912]), .B(n12428), .Z(n12430) );
  XNOR U12262 ( .A(n12431), .B(n12432), .Z(n12428) );
  AND U12263 ( .A(n375), .B(n12427), .Z(n12432) );
  XNOR U12264 ( .A(n12431), .B(n12425), .Z(n12427) );
  XOR U12265 ( .A(n12433), .B(n12434), .Z(n12425) );
  AND U12266 ( .A(n390), .B(n12435), .Z(n12434) );
  XNOR U12267 ( .A(n12436), .B(n12437), .Z(n12431) );
  AND U12268 ( .A(n382), .B(n12438), .Z(n12437) );
  XOR U12269 ( .A(p_input[944]), .B(n12436), .Z(n12438) );
  XNOR U12270 ( .A(n12439), .B(n12440), .Z(n12436) );
  AND U12271 ( .A(n386), .B(n12435), .Z(n12440) );
  XNOR U12272 ( .A(n12439), .B(n12433), .Z(n12435) );
  XOR U12273 ( .A(n12441), .B(n12442), .Z(n12433) );
  AND U12274 ( .A(n401), .B(n12443), .Z(n12442) );
  XNOR U12275 ( .A(n12444), .B(n12445), .Z(n12439) );
  AND U12276 ( .A(n393), .B(n12446), .Z(n12445) );
  XOR U12277 ( .A(p_input[976]), .B(n12444), .Z(n12446) );
  XNOR U12278 ( .A(n12447), .B(n12448), .Z(n12444) );
  AND U12279 ( .A(n397), .B(n12443), .Z(n12448) );
  XNOR U12280 ( .A(n12447), .B(n12441), .Z(n12443) );
  XOR U12281 ( .A(n12449), .B(n12450), .Z(n12441) );
  AND U12282 ( .A(n412), .B(n12451), .Z(n12450) );
  XNOR U12283 ( .A(n12452), .B(n12453), .Z(n12447) );
  AND U12284 ( .A(n404), .B(n12454), .Z(n12453) );
  XOR U12285 ( .A(p_input[1008]), .B(n12452), .Z(n12454) );
  XNOR U12286 ( .A(n12455), .B(n12456), .Z(n12452) );
  AND U12287 ( .A(n408), .B(n12451), .Z(n12456) );
  XNOR U12288 ( .A(n12455), .B(n12449), .Z(n12451) );
  XOR U12289 ( .A(n12457), .B(n12458), .Z(n12449) );
  AND U12290 ( .A(n423), .B(n12459), .Z(n12458) );
  XNOR U12291 ( .A(n12460), .B(n12461), .Z(n12455) );
  AND U12292 ( .A(n415), .B(n12462), .Z(n12461) );
  XOR U12293 ( .A(p_input[1040]), .B(n12460), .Z(n12462) );
  XNOR U12294 ( .A(n12463), .B(n12464), .Z(n12460) );
  AND U12295 ( .A(n419), .B(n12459), .Z(n12464) );
  XNOR U12296 ( .A(n12463), .B(n12457), .Z(n12459) );
  XOR U12297 ( .A(n12465), .B(n12466), .Z(n12457) );
  AND U12298 ( .A(n434), .B(n12467), .Z(n12466) );
  XNOR U12299 ( .A(n12468), .B(n12469), .Z(n12463) );
  AND U12300 ( .A(n426), .B(n12470), .Z(n12469) );
  XOR U12301 ( .A(p_input[1072]), .B(n12468), .Z(n12470) );
  XNOR U12302 ( .A(n12471), .B(n12472), .Z(n12468) );
  AND U12303 ( .A(n430), .B(n12467), .Z(n12472) );
  XNOR U12304 ( .A(n12471), .B(n12465), .Z(n12467) );
  XOR U12305 ( .A(n12473), .B(n12474), .Z(n12465) );
  AND U12306 ( .A(n445), .B(n12475), .Z(n12474) );
  XNOR U12307 ( .A(n12476), .B(n12477), .Z(n12471) );
  AND U12308 ( .A(n437), .B(n12478), .Z(n12477) );
  XOR U12309 ( .A(p_input[1104]), .B(n12476), .Z(n12478) );
  XNOR U12310 ( .A(n12479), .B(n12480), .Z(n12476) );
  AND U12311 ( .A(n441), .B(n12475), .Z(n12480) );
  XNOR U12312 ( .A(n12479), .B(n12473), .Z(n12475) );
  XOR U12313 ( .A(n12481), .B(n12482), .Z(n12473) );
  AND U12314 ( .A(n456), .B(n12483), .Z(n12482) );
  XNOR U12315 ( .A(n12484), .B(n12485), .Z(n12479) );
  AND U12316 ( .A(n448), .B(n12486), .Z(n12485) );
  XOR U12317 ( .A(p_input[1136]), .B(n12484), .Z(n12486) );
  XNOR U12318 ( .A(n12487), .B(n12488), .Z(n12484) );
  AND U12319 ( .A(n452), .B(n12483), .Z(n12488) );
  XNOR U12320 ( .A(n12487), .B(n12481), .Z(n12483) );
  XOR U12321 ( .A(n12489), .B(n12490), .Z(n12481) );
  AND U12322 ( .A(n467), .B(n12491), .Z(n12490) );
  XNOR U12323 ( .A(n12492), .B(n12493), .Z(n12487) );
  AND U12324 ( .A(n459), .B(n12494), .Z(n12493) );
  XOR U12325 ( .A(p_input[1168]), .B(n12492), .Z(n12494) );
  XNOR U12326 ( .A(n12495), .B(n12496), .Z(n12492) );
  AND U12327 ( .A(n463), .B(n12491), .Z(n12496) );
  XNOR U12328 ( .A(n12495), .B(n12489), .Z(n12491) );
  XOR U12329 ( .A(n12497), .B(n12498), .Z(n12489) );
  AND U12330 ( .A(n478), .B(n12499), .Z(n12498) );
  XNOR U12331 ( .A(n12500), .B(n12501), .Z(n12495) );
  AND U12332 ( .A(n470), .B(n12502), .Z(n12501) );
  XOR U12333 ( .A(p_input[1200]), .B(n12500), .Z(n12502) );
  XNOR U12334 ( .A(n12503), .B(n12504), .Z(n12500) );
  AND U12335 ( .A(n474), .B(n12499), .Z(n12504) );
  XNOR U12336 ( .A(n12503), .B(n12497), .Z(n12499) );
  XOR U12337 ( .A(n12505), .B(n12506), .Z(n12497) );
  AND U12338 ( .A(n489), .B(n12507), .Z(n12506) );
  XNOR U12339 ( .A(n12508), .B(n12509), .Z(n12503) );
  AND U12340 ( .A(n481), .B(n12510), .Z(n12509) );
  XOR U12341 ( .A(p_input[1232]), .B(n12508), .Z(n12510) );
  XNOR U12342 ( .A(n12511), .B(n12512), .Z(n12508) );
  AND U12343 ( .A(n485), .B(n12507), .Z(n12512) );
  XNOR U12344 ( .A(n12511), .B(n12505), .Z(n12507) );
  XOR U12345 ( .A(n12513), .B(n12514), .Z(n12505) );
  AND U12346 ( .A(n500), .B(n12515), .Z(n12514) );
  XNOR U12347 ( .A(n12516), .B(n12517), .Z(n12511) );
  AND U12348 ( .A(n492), .B(n12518), .Z(n12517) );
  XOR U12349 ( .A(p_input[1264]), .B(n12516), .Z(n12518) );
  XNOR U12350 ( .A(n12519), .B(n12520), .Z(n12516) );
  AND U12351 ( .A(n496), .B(n12515), .Z(n12520) );
  XNOR U12352 ( .A(n12519), .B(n12513), .Z(n12515) );
  XOR U12353 ( .A(n12521), .B(n12522), .Z(n12513) );
  AND U12354 ( .A(n511), .B(n12523), .Z(n12522) );
  XNOR U12355 ( .A(n12524), .B(n12525), .Z(n12519) );
  AND U12356 ( .A(n503), .B(n12526), .Z(n12525) );
  XOR U12357 ( .A(p_input[1296]), .B(n12524), .Z(n12526) );
  XNOR U12358 ( .A(n12527), .B(n12528), .Z(n12524) );
  AND U12359 ( .A(n507), .B(n12523), .Z(n12528) );
  XNOR U12360 ( .A(n12527), .B(n12521), .Z(n12523) );
  XOR U12361 ( .A(n12529), .B(n12530), .Z(n12521) );
  AND U12362 ( .A(n522), .B(n12531), .Z(n12530) );
  XNOR U12363 ( .A(n12532), .B(n12533), .Z(n12527) );
  AND U12364 ( .A(n514), .B(n12534), .Z(n12533) );
  XOR U12365 ( .A(p_input[1328]), .B(n12532), .Z(n12534) );
  XNOR U12366 ( .A(n12535), .B(n12536), .Z(n12532) );
  AND U12367 ( .A(n518), .B(n12531), .Z(n12536) );
  XNOR U12368 ( .A(n12535), .B(n12529), .Z(n12531) );
  XOR U12369 ( .A(n12537), .B(n12538), .Z(n12529) );
  AND U12370 ( .A(n533), .B(n12539), .Z(n12538) );
  XNOR U12371 ( .A(n12540), .B(n12541), .Z(n12535) );
  AND U12372 ( .A(n525), .B(n12542), .Z(n12541) );
  XOR U12373 ( .A(p_input[1360]), .B(n12540), .Z(n12542) );
  XNOR U12374 ( .A(n12543), .B(n12544), .Z(n12540) );
  AND U12375 ( .A(n529), .B(n12539), .Z(n12544) );
  XNOR U12376 ( .A(n12543), .B(n12537), .Z(n12539) );
  XOR U12377 ( .A(n12545), .B(n12546), .Z(n12537) );
  AND U12378 ( .A(n544), .B(n12547), .Z(n12546) );
  XNOR U12379 ( .A(n12548), .B(n12549), .Z(n12543) );
  AND U12380 ( .A(n536), .B(n12550), .Z(n12549) );
  XOR U12381 ( .A(p_input[1392]), .B(n12548), .Z(n12550) );
  XNOR U12382 ( .A(n12551), .B(n12552), .Z(n12548) );
  AND U12383 ( .A(n540), .B(n12547), .Z(n12552) );
  XNOR U12384 ( .A(n12551), .B(n12545), .Z(n12547) );
  XOR U12385 ( .A(n12553), .B(n12554), .Z(n12545) );
  AND U12386 ( .A(n555), .B(n12555), .Z(n12554) );
  XNOR U12387 ( .A(n12556), .B(n12557), .Z(n12551) );
  AND U12388 ( .A(n547), .B(n12558), .Z(n12557) );
  XOR U12389 ( .A(p_input[1424]), .B(n12556), .Z(n12558) );
  XNOR U12390 ( .A(n12559), .B(n12560), .Z(n12556) );
  AND U12391 ( .A(n551), .B(n12555), .Z(n12560) );
  XNOR U12392 ( .A(n12559), .B(n12553), .Z(n12555) );
  XOR U12393 ( .A(n12561), .B(n12562), .Z(n12553) );
  AND U12394 ( .A(n566), .B(n12563), .Z(n12562) );
  XNOR U12395 ( .A(n12564), .B(n12565), .Z(n12559) );
  AND U12396 ( .A(n558), .B(n12566), .Z(n12565) );
  XOR U12397 ( .A(p_input[1456]), .B(n12564), .Z(n12566) );
  XNOR U12398 ( .A(n12567), .B(n12568), .Z(n12564) );
  AND U12399 ( .A(n562), .B(n12563), .Z(n12568) );
  XNOR U12400 ( .A(n12567), .B(n12561), .Z(n12563) );
  XOR U12401 ( .A(n12569), .B(n12570), .Z(n12561) );
  AND U12402 ( .A(n577), .B(n12571), .Z(n12570) );
  XNOR U12403 ( .A(n12572), .B(n12573), .Z(n12567) );
  AND U12404 ( .A(n569), .B(n12574), .Z(n12573) );
  XOR U12405 ( .A(p_input[1488]), .B(n12572), .Z(n12574) );
  XNOR U12406 ( .A(n12575), .B(n12576), .Z(n12572) );
  AND U12407 ( .A(n573), .B(n12571), .Z(n12576) );
  XNOR U12408 ( .A(n12575), .B(n12569), .Z(n12571) );
  XOR U12409 ( .A(n12577), .B(n12578), .Z(n12569) );
  AND U12410 ( .A(n588), .B(n12579), .Z(n12578) );
  XNOR U12411 ( .A(n12580), .B(n12581), .Z(n12575) );
  AND U12412 ( .A(n580), .B(n12582), .Z(n12581) );
  XOR U12413 ( .A(p_input[1520]), .B(n12580), .Z(n12582) );
  XNOR U12414 ( .A(n12583), .B(n12584), .Z(n12580) );
  AND U12415 ( .A(n584), .B(n12579), .Z(n12584) );
  XNOR U12416 ( .A(n12583), .B(n12577), .Z(n12579) );
  XOR U12417 ( .A(n12585), .B(n12586), .Z(n12577) );
  AND U12418 ( .A(n599), .B(n12587), .Z(n12586) );
  XNOR U12419 ( .A(n12588), .B(n12589), .Z(n12583) );
  AND U12420 ( .A(n591), .B(n12590), .Z(n12589) );
  XOR U12421 ( .A(p_input[1552]), .B(n12588), .Z(n12590) );
  XNOR U12422 ( .A(n12591), .B(n12592), .Z(n12588) );
  AND U12423 ( .A(n595), .B(n12587), .Z(n12592) );
  XNOR U12424 ( .A(n12591), .B(n12585), .Z(n12587) );
  XOR U12425 ( .A(n12593), .B(n12594), .Z(n12585) );
  AND U12426 ( .A(n610), .B(n12595), .Z(n12594) );
  XNOR U12427 ( .A(n12596), .B(n12597), .Z(n12591) );
  AND U12428 ( .A(n602), .B(n12598), .Z(n12597) );
  XOR U12429 ( .A(p_input[1584]), .B(n12596), .Z(n12598) );
  XNOR U12430 ( .A(n12599), .B(n12600), .Z(n12596) );
  AND U12431 ( .A(n606), .B(n12595), .Z(n12600) );
  XNOR U12432 ( .A(n12599), .B(n12593), .Z(n12595) );
  XOR U12433 ( .A(n12601), .B(n12602), .Z(n12593) );
  AND U12434 ( .A(n621), .B(n12603), .Z(n12602) );
  XNOR U12435 ( .A(n12604), .B(n12605), .Z(n12599) );
  AND U12436 ( .A(n613), .B(n12606), .Z(n12605) );
  XOR U12437 ( .A(p_input[1616]), .B(n12604), .Z(n12606) );
  XNOR U12438 ( .A(n12607), .B(n12608), .Z(n12604) );
  AND U12439 ( .A(n617), .B(n12603), .Z(n12608) );
  XNOR U12440 ( .A(n12607), .B(n12601), .Z(n12603) );
  XOR U12441 ( .A(n12609), .B(n12610), .Z(n12601) );
  AND U12442 ( .A(n632), .B(n12611), .Z(n12610) );
  XNOR U12443 ( .A(n12612), .B(n12613), .Z(n12607) );
  AND U12444 ( .A(n624), .B(n12614), .Z(n12613) );
  XOR U12445 ( .A(p_input[1648]), .B(n12612), .Z(n12614) );
  XNOR U12446 ( .A(n12615), .B(n12616), .Z(n12612) );
  AND U12447 ( .A(n628), .B(n12611), .Z(n12616) );
  XNOR U12448 ( .A(n12615), .B(n12609), .Z(n12611) );
  XOR U12449 ( .A(n12617), .B(n12618), .Z(n12609) );
  AND U12450 ( .A(n643), .B(n12619), .Z(n12618) );
  XNOR U12451 ( .A(n12620), .B(n12621), .Z(n12615) );
  AND U12452 ( .A(n635), .B(n12622), .Z(n12621) );
  XOR U12453 ( .A(p_input[1680]), .B(n12620), .Z(n12622) );
  XNOR U12454 ( .A(n12623), .B(n12624), .Z(n12620) );
  AND U12455 ( .A(n639), .B(n12619), .Z(n12624) );
  XNOR U12456 ( .A(n12623), .B(n12617), .Z(n12619) );
  XOR U12457 ( .A(n12625), .B(n12626), .Z(n12617) );
  AND U12458 ( .A(n654), .B(n12627), .Z(n12626) );
  XNOR U12459 ( .A(n12628), .B(n12629), .Z(n12623) );
  AND U12460 ( .A(n646), .B(n12630), .Z(n12629) );
  XOR U12461 ( .A(p_input[1712]), .B(n12628), .Z(n12630) );
  XNOR U12462 ( .A(n12631), .B(n12632), .Z(n12628) );
  AND U12463 ( .A(n650), .B(n12627), .Z(n12632) );
  XNOR U12464 ( .A(n12631), .B(n12625), .Z(n12627) );
  XOR U12465 ( .A(n12633), .B(n12634), .Z(n12625) );
  AND U12466 ( .A(n665), .B(n12635), .Z(n12634) );
  XNOR U12467 ( .A(n12636), .B(n12637), .Z(n12631) );
  AND U12468 ( .A(n657), .B(n12638), .Z(n12637) );
  XOR U12469 ( .A(p_input[1744]), .B(n12636), .Z(n12638) );
  XNOR U12470 ( .A(n12639), .B(n12640), .Z(n12636) );
  AND U12471 ( .A(n661), .B(n12635), .Z(n12640) );
  XNOR U12472 ( .A(n12639), .B(n12633), .Z(n12635) );
  XOR U12473 ( .A(n12641), .B(n12642), .Z(n12633) );
  AND U12474 ( .A(n676), .B(n12643), .Z(n12642) );
  XNOR U12475 ( .A(n12644), .B(n12645), .Z(n12639) );
  AND U12476 ( .A(n668), .B(n12646), .Z(n12645) );
  XOR U12477 ( .A(p_input[1776]), .B(n12644), .Z(n12646) );
  XNOR U12478 ( .A(n12647), .B(n12648), .Z(n12644) );
  AND U12479 ( .A(n672), .B(n12643), .Z(n12648) );
  XNOR U12480 ( .A(n12647), .B(n12641), .Z(n12643) );
  XOR U12481 ( .A(n12649), .B(n12650), .Z(n12641) );
  AND U12482 ( .A(n687), .B(n12651), .Z(n12650) );
  XNOR U12483 ( .A(n12652), .B(n12653), .Z(n12647) );
  AND U12484 ( .A(n679), .B(n12654), .Z(n12653) );
  XOR U12485 ( .A(p_input[1808]), .B(n12652), .Z(n12654) );
  XNOR U12486 ( .A(n12655), .B(n12656), .Z(n12652) );
  AND U12487 ( .A(n683), .B(n12651), .Z(n12656) );
  XNOR U12488 ( .A(n12655), .B(n12649), .Z(n12651) );
  XOR U12489 ( .A(n12657), .B(n12658), .Z(n12649) );
  AND U12490 ( .A(n698), .B(n12659), .Z(n12658) );
  XNOR U12491 ( .A(n12660), .B(n12661), .Z(n12655) );
  AND U12492 ( .A(n690), .B(n12662), .Z(n12661) );
  XOR U12493 ( .A(p_input[1840]), .B(n12660), .Z(n12662) );
  XNOR U12494 ( .A(n12663), .B(n12664), .Z(n12660) );
  AND U12495 ( .A(n694), .B(n12659), .Z(n12664) );
  XNOR U12496 ( .A(n12663), .B(n12657), .Z(n12659) );
  XOR U12497 ( .A(n12665), .B(n12666), .Z(n12657) );
  AND U12498 ( .A(n709), .B(n12667), .Z(n12666) );
  XNOR U12499 ( .A(n12668), .B(n12669), .Z(n12663) );
  AND U12500 ( .A(n701), .B(n12670), .Z(n12669) );
  XOR U12501 ( .A(p_input[1872]), .B(n12668), .Z(n12670) );
  XNOR U12502 ( .A(n12671), .B(n12672), .Z(n12668) );
  AND U12503 ( .A(n705), .B(n12667), .Z(n12672) );
  XNOR U12504 ( .A(n12671), .B(n12665), .Z(n12667) );
  XOR U12505 ( .A(n12673), .B(n12674), .Z(n12665) );
  AND U12506 ( .A(n720), .B(n12675), .Z(n12674) );
  XNOR U12507 ( .A(n12676), .B(n12677), .Z(n12671) );
  AND U12508 ( .A(n712), .B(n12678), .Z(n12677) );
  XOR U12509 ( .A(p_input[1904]), .B(n12676), .Z(n12678) );
  XNOR U12510 ( .A(n12679), .B(n12680), .Z(n12676) );
  AND U12511 ( .A(n716), .B(n12675), .Z(n12680) );
  XNOR U12512 ( .A(n12679), .B(n12673), .Z(n12675) );
  XOR U12513 ( .A(n12681), .B(n12682), .Z(n12673) );
  AND U12514 ( .A(n731), .B(n12683), .Z(n12682) );
  XNOR U12515 ( .A(n12684), .B(n12685), .Z(n12679) );
  AND U12516 ( .A(n723), .B(n12686), .Z(n12685) );
  XOR U12517 ( .A(p_input[1936]), .B(n12684), .Z(n12686) );
  XNOR U12518 ( .A(n12687), .B(n12688), .Z(n12684) );
  AND U12519 ( .A(n727), .B(n12683), .Z(n12688) );
  XNOR U12520 ( .A(n12687), .B(n12681), .Z(n12683) );
  XOR U12521 ( .A(\knn_comb_/min_val_out[0][16] ), .B(n12689), .Z(n12681) );
  AND U12522 ( .A(n741), .B(n12690), .Z(n12689) );
  XNOR U12523 ( .A(n12691), .B(n12692), .Z(n12687) );
  AND U12524 ( .A(n734), .B(n12693), .Z(n12692) );
  XOR U12525 ( .A(p_input[1968]), .B(n12691), .Z(n12693) );
  XNOR U12526 ( .A(n12694), .B(n12695), .Z(n12691) );
  AND U12527 ( .A(n738), .B(n12690), .Z(n12695) );
  XOR U12528 ( .A(n12696), .B(n12694), .Z(n12690) );
  IV U12529 ( .A(\knn_comb_/min_val_out[0][16] ), .Z(n12696) );
  IV U12530 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .Z(n12694)
         );
  XOR U12531 ( .A(n45), .B(n12697), .Z(o[15]) );
  AND U12532 ( .A(n58), .B(n12698), .Z(n45) );
  XOR U12533 ( .A(n46), .B(n12697), .Z(n12698) );
  XOR U12534 ( .A(n12699), .B(n12700), .Z(n12697) );
  AND U12535 ( .A(n70), .B(n12701), .Z(n12700) );
  XOR U12536 ( .A(n12702), .B(n12703), .Z(n46) );
  AND U12537 ( .A(n62), .B(n12704), .Z(n12703) );
  XOR U12538 ( .A(p_input[15]), .B(n12702), .Z(n12704) );
  XNOR U12539 ( .A(n12705), .B(n12706), .Z(n12702) );
  AND U12540 ( .A(n66), .B(n12701), .Z(n12706) );
  XNOR U12541 ( .A(n12705), .B(n12699), .Z(n12701) );
  XOR U12542 ( .A(n12707), .B(n12708), .Z(n12699) );
  AND U12543 ( .A(n82), .B(n12709), .Z(n12708) );
  XNOR U12544 ( .A(n12710), .B(n12711), .Z(n12705) );
  AND U12545 ( .A(n74), .B(n12712), .Z(n12711) );
  XOR U12546 ( .A(p_input[47]), .B(n12710), .Z(n12712) );
  XNOR U12547 ( .A(n12713), .B(n12714), .Z(n12710) );
  AND U12548 ( .A(n78), .B(n12709), .Z(n12714) );
  XNOR U12549 ( .A(n12713), .B(n12707), .Z(n12709) );
  XOR U12550 ( .A(n12715), .B(n12716), .Z(n12707) );
  AND U12551 ( .A(n93), .B(n12717), .Z(n12716) );
  XNOR U12552 ( .A(n12718), .B(n12719), .Z(n12713) );
  AND U12553 ( .A(n85), .B(n12720), .Z(n12719) );
  XOR U12554 ( .A(p_input[79]), .B(n12718), .Z(n12720) );
  XNOR U12555 ( .A(n12721), .B(n12722), .Z(n12718) );
  AND U12556 ( .A(n89), .B(n12717), .Z(n12722) );
  XNOR U12557 ( .A(n12721), .B(n12715), .Z(n12717) );
  XOR U12558 ( .A(n12723), .B(n12724), .Z(n12715) );
  AND U12559 ( .A(n104), .B(n12725), .Z(n12724) );
  XNOR U12560 ( .A(n12726), .B(n12727), .Z(n12721) );
  AND U12561 ( .A(n96), .B(n12728), .Z(n12727) );
  XOR U12562 ( .A(p_input[111]), .B(n12726), .Z(n12728) );
  XNOR U12563 ( .A(n12729), .B(n12730), .Z(n12726) );
  AND U12564 ( .A(n100), .B(n12725), .Z(n12730) );
  XNOR U12565 ( .A(n12729), .B(n12723), .Z(n12725) );
  XOR U12566 ( .A(n12731), .B(n12732), .Z(n12723) );
  AND U12567 ( .A(n115), .B(n12733), .Z(n12732) );
  XNOR U12568 ( .A(n12734), .B(n12735), .Z(n12729) );
  AND U12569 ( .A(n107), .B(n12736), .Z(n12735) );
  XOR U12570 ( .A(p_input[143]), .B(n12734), .Z(n12736) );
  XNOR U12571 ( .A(n12737), .B(n12738), .Z(n12734) );
  AND U12572 ( .A(n111), .B(n12733), .Z(n12738) );
  XNOR U12573 ( .A(n12737), .B(n12731), .Z(n12733) );
  XOR U12574 ( .A(n12739), .B(n12740), .Z(n12731) );
  AND U12575 ( .A(n126), .B(n12741), .Z(n12740) );
  XNOR U12576 ( .A(n12742), .B(n12743), .Z(n12737) );
  AND U12577 ( .A(n118), .B(n12744), .Z(n12743) );
  XOR U12578 ( .A(p_input[175]), .B(n12742), .Z(n12744) );
  XNOR U12579 ( .A(n12745), .B(n12746), .Z(n12742) );
  AND U12580 ( .A(n122), .B(n12741), .Z(n12746) );
  XNOR U12581 ( .A(n12745), .B(n12739), .Z(n12741) );
  XOR U12582 ( .A(n12747), .B(n12748), .Z(n12739) );
  AND U12583 ( .A(n137), .B(n12749), .Z(n12748) );
  XNOR U12584 ( .A(n12750), .B(n12751), .Z(n12745) );
  AND U12585 ( .A(n129), .B(n12752), .Z(n12751) );
  XOR U12586 ( .A(p_input[207]), .B(n12750), .Z(n12752) );
  XNOR U12587 ( .A(n12753), .B(n12754), .Z(n12750) );
  AND U12588 ( .A(n133), .B(n12749), .Z(n12754) );
  XNOR U12589 ( .A(n12753), .B(n12747), .Z(n12749) );
  XOR U12590 ( .A(n12755), .B(n12756), .Z(n12747) );
  AND U12591 ( .A(n148), .B(n12757), .Z(n12756) );
  XNOR U12592 ( .A(n12758), .B(n12759), .Z(n12753) );
  AND U12593 ( .A(n140), .B(n12760), .Z(n12759) );
  XOR U12594 ( .A(p_input[239]), .B(n12758), .Z(n12760) );
  XNOR U12595 ( .A(n12761), .B(n12762), .Z(n12758) );
  AND U12596 ( .A(n144), .B(n12757), .Z(n12762) );
  XNOR U12597 ( .A(n12761), .B(n12755), .Z(n12757) );
  XOR U12598 ( .A(n12763), .B(n12764), .Z(n12755) );
  AND U12599 ( .A(n159), .B(n12765), .Z(n12764) );
  XNOR U12600 ( .A(n12766), .B(n12767), .Z(n12761) );
  AND U12601 ( .A(n151), .B(n12768), .Z(n12767) );
  XOR U12602 ( .A(p_input[271]), .B(n12766), .Z(n12768) );
  XNOR U12603 ( .A(n12769), .B(n12770), .Z(n12766) );
  AND U12604 ( .A(n155), .B(n12765), .Z(n12770) );
  XNOR U12605 ( .A(n12769), .B(n12763), .Z(n12765) );
  XOR U12606 ( .A(n12771), .B(n12772), .Z(n12763) );
  AND U12607 ( .A(n170), .B(n12773), .Z(n12772) );
  XNOR U12608 ( .A(n12774), .B(n12775), .Z(n12769) );
  AND U12609 ( .A(n162), .B(n12776), .Z(n12775) );
  XOR U12610 ( .A(p_input[303]), .B(n12774), .Z(n12776) );
  XNOR U12611 ( .A(n12777), .B(n12778), .Z(n12774) );
  AND U12612 ( .A(n166), .B(n12773), .Z(n12778) );
  XNOR U12613 ( .A(n12777), .B(n12771), .Z(n12773) );
  XOR U12614 ( .A(n12779), .B(n12780), .Z(n12771) );
  AND U12615 ( .A(n181), .B(n12781), .Z(n12780) );
  XNOR U12616 ( .A(n12782), .B(n12783), .Z(n12777) );
  AND U12617 ( .A(n173), .B(n12784), .Z(n12783) );
  XOR U12618 ( .A(p_input[335]), .B(n12782), .Z(n12784) );
  XNOR U12619 ( .A(n12785), .B(n12786), .Z(n12782) );
  AND U12620 ( .A(n177), .B(n12781), .Z(n12786) );
  XNOR U12621 ( .A(n12785), .B(n12779), .Z(n12781) );
  XOR U12622 ( .A(n12787), .B(n12788), .Z(n12779) );
  AND U12623 ( .A(n192), .B(n12789), .Z(n12788) );
  XNOR U12624 ( .A(n12790), .B(n12791), .Z(n12785) );
  AND U12625 ( .A(n184), .B(n12792), .Z(n12791) );
  XOR U12626 ( .A(p_input[367]), .B(n12790), .Z(n12792) );
  XNOR U12627 ( .A(n12793), .B(n12794), .Z(n12790) );
  AND U12628 ( .A(n188), .B(n12789), .Z(n12794) );
  XNOR U12629 ( .A(n12793), .B(n12787), .Z(n12789) );
  XOR U12630 ( .A(n12795), .B(n12796), .Z(n12787) );
  AND U12631 ( .A(n203), .B(n12797), .Z(n12796) );
  XNOR U12632 ( .A(n12798), .B(n12799), .Z(n12793) );
  AND U12633 ( .A(n195), .B(n12800), .Z(n12799) );
  XOR U12634 ( .A(p_input[399]), .B(n12798), .Z(n12800) );
  XNOR U12635 ( .A(n12801), .B(n12802), .Z(n12798) );
  AND U12636 ( .A(n199), .B(n12797), .Z(n12802) );
  XNOR U12637 ( .A(n12801), .B(n12795), .Z(n12797) );
  XOR U12638 ( .A(n12803), .B(n12804), .Z(n12795) );
  AND U12639 ( .A(n214), .B(n12805), .Z(n12804) );
  XNOR U12640 ( .A(n12806), .B(n12807), .Z(n12801) );
  AND U12641 ( .A(n206), .B(n12808), .Z(n12807) );
  XOR U12642 ( .A(p_input[431]), .B(n12806), .Z(n12808) );
  XNOR U12643 ( .A(n12809), .B(n12810), .Z(n12806) );
  AND U12644 ( .A(n210), .B(n12805), .Z(n12810) );
  XNOR U12645 ( .A(n12809), .B(n12803), .Z(n12805) );
  XOR U12646 ( .A(n12811), .B(n12812), .Z(n12803) );
  AND U12647 ( .A(n225), .B(n12813), .Z(n12812) );
  XNOR U12648 ( .A(n12814), .B(n12815), .Z(n12809) );
  AND U12649 ( .A(n217), .B(n12816), .Z(n12815) );
  XOR U12650 ( .A(p_input[463]), .B(n12814), .Z(n12816) );
  XNOR U12651 ( .A(n12817), .B(n12818), .Z(n12814) );
  AND U12652 ( .A(n221), .B(n12813), .Z(n12818) );
  XNOR U12653 ( .A(n12817), .B(n12811), .Z(n12813) );
  XOR U12654 ( .A(n12819), .B(n12820), .Z(n12811) );
  AND U12655 ( .A(n236), .B(n12821), .Z(n12820) );
  XNOR U12656 ( .A(n12822), .B(n12823), .Z(n12817) );
  AND U12657 ( .A(n228), .B(n12824), .Z(n12823) );
  XOR U12658 ( .A(p_input[495]), .B(n12822), .Z(n12824) );
  XNOR U12659 ( .A(n12825), .B(n12826), .Z(n12822) );
  AND U12660 ( .A(n232), .B(n12821), .Z(n12826) );
  XNOR U12661 ( .A(n12825), .B(n12819), .Z(n12821) );
  XOR U12662 ( .A(n12827), .B(n12828), .Z(n12819) );
  AND U12663 ( .A(n247), .B(n12829), .Z(n12828) );
  XNOR U12664 ( .A(n12830), .B(n12831), .Z(n12825) );
  AND U12665 ( .A(n239), .B(n12832), .Z(n12831) );
  XOR U12666 ( .A(p_input[527]), .B(n12830), .Z(n12832) );
  XNOR U12667 ( .A(n12833), .B(n12834), .Z(n12830) );
  AND U12668 ( .A(n243), .B(n12829), .Z(n12834) );
  XNOR U12669 ( .A(n12833), .B(n12827), .Z(n12829) );
  XOR U12670 ( .A(n12835), .B(n12836), .Z(n12827) );
  AND U12671 ( .A(n258), .B(n12837), .Z(n12836) );
  XNOR U12672 ( .A(n12838), .B(n12839), .Z(n12833) );
  AND U12673 ( .A(n250), .B(n12840), .Z(n12839) );
  XOR U12674 ( .A(p_input[559]), .B(n12838), .Z(n12840) );
  XNOR U12675 ( .A(n12841), .B(n12842), .Z(n12838) );
  AND U12676 ( .A(n254), .B(n12837), .Z(n12842) );
  XNOR U12677 ( .A(n12841), .B(n12835), .Z(n12837) );
  XOR U12678 ( .A(n12843), .B(n12844), .Z(n12835) );
  AND U12679 ( .A(n269), .B(n12845), .Z(n12844) );
  XNOR U12680 ( .A(n12846), .B(n12847), .Z(n12841) );
  AND U12681 ( .A(n261), .B(n12848), .Z(n12847) );
  XOR U12682 ( .A(p_input[591]), .B(n12846), .Z(n12848) );
  XNOR U12683 ( .A(n12849), .B(n12850), .Z(n12846) );
  AND U12684 ( .A(n265), .B(n12845), .Z(n12850) );
  XNOR U12685 ( .A(n12849), .B(n12843), .Z(n12845) );
  XOR U12686 ( .A(n12851), .B(n12852), .Z(n12843) );
  AND U12687 ( .A(n280), .B(n12853), .Z(n12852) );
  XNOR U12688 ( .A(n12854), .B(n12855), .Z(n12849) );
  AND U12689 ( .A(n272), .B(n12856), .Z(n12855) );
  XOR U12690 ( .A(p_input[623]), .B(n12854), .Z(n12856) );
  XNOR U12691 ( .A(n12857), .B(n12858), .Z(n12854) );
  AND U12692 ( .A(n276), .B(n12853), .Z(n12858) );
  XNOR U12693 ( .A(n12857), .B(n12851), .Z(n12853) );
  XOR U12694 ( .A(n12859), .B(n12860), .Z(n12851) );
  AND U12695 ( .A(n291), .B(n12861), .Z(n12860) );
  XNOR U12696 ( .A(n12862), .B(n12863), .Z(n12857) );
  AND U12697 ( .A(n283), .B(n12864), .Z(n12863) );
  XOR U12698 ( .A(p_input[655]), .B(n12862), .Z(n12864) );
  XNOR U12699 ( .A(n12865), .B(n12866), .Z(n12862) );
  AND U12700 ( .A(n287), .B(n12861), .Z(n12866) );
  XNOR U12701 ( .A(n12865), .B(n12859), .Z(n12861) );
  XOR U12702 ( .A(n12867), .B(n12868), .Z(n12859) );
  AND U12703 ( .A(n302), .B(n12869), .Z(n12868) );
  XNOR U12704 ( .A(n12870), .B(n12871), .Z(n12865) );
  AND U12705 ( .A(n294), .B(n12872), .Z(n12871) );
  XOR U12706 ( .A(p_input[687]), .B(n12870), .Z(n12872) );
  XNOR U12707 ( .A(n12873), .B(n12874), .Z(n12870) );
  AND U12708 ( .A(n298), .B(n12869), .Z(n12874) );
  XNOR U12709 ( .A(n12873), .B(n12867), .Z(n12869) );
  XOR U12710 ( .A(n12875), .B(n12876), .Z(n12867) );
  AND U12711 ( .A(n313), .B(n12877), .Z(n12876) );
  XNOR U12712 ( .A(n12878), .B(n12879), .Z(n12873) );
  AND U12713 ( .A(n305), .B(n12880), .Z(n12879) );
  XOR U12714 ( .A(p_input[719]), .B(n12878), .Z(n12880) );
  XNOR U12715 ( .A(n12881), .B(n12882), .Z(n12878) );
  AND U12716 ( .A(n309), .B(n12877), .Z(n12882) );
  XNOR U12717 ( .A(n12881), .B(n12875), .Z(n12877) );
  XOR U12718 ( .A(n12883), .B(n12884), .Z(n12875) );
  AND U12719 ( .A(n324), .B(n12885), .Z(n12884) );
  XNOR U12720 ( .A(n12886), .B(n12887), .Z(n12881) );
  AND U12721 ( .A(n316), .B(n12888), .Z(n12887) );
  XOR U12722 ( .A(p_input[751]), .B(n12886), .Z(n12888) );
  XNOR U12723 ( .A(n12889), .B(n12890), .Z(n12886) );
  AND U12724 ( .A(n320), .B(n12885), .Z(n12890) );
  XNOR U12725 ( .A(n12889), .B(n12883), .Z(n12885) );
  XOR U12726 ( .A(n12891), .B(n12892), .Z(n12883) );
  AND U12727 ( .A(n335), .B(n12893), .Z(n12892) );
  XNOR U12728 ( .A(n12894), .B(n12895), .Z(n12889) );
  AND U12729 ( .A(n327), .B(n12896), .Z(n12895) );
  XOR U12730 ( .A(p_input[783]), .B(n12894), .Z(n12896) );
  XNOR U12731 ( .A(n12897), .B(n12898), .Z(n12894) );
  AND U12732 ( .A(n331), .B(n12893), .Z(n12898) );
  XNOR U12733 ( .A(n12897), .B(n12891), .Z(n12893) );
  XOR U12734 ( .A(n12899), .B(n12900), .Z(n12891) );
  AND U12735 ( .A(n346), .B(n12901), .Z(n12900) );
  XNOR U12736 ( .A(n12902), .B(n12903), .Z(n12897) );
  AND U12737 ( .A(n338), .B(n12904), .Z(n12903) );
  XOR U12738 ( .A(p_input[815]), .B(n12902), .Z(n12904) );
  XNOR U12739 ( .A(n12905), .B(n12906), .Z(n12902) );
  AND U12740 ( .A(n342), .B(n12901), .Z(n12906) );
  XNOR U12741 ( .A(n12905), .B(n12899), .Z(n12901) );
  XOR U12742 ( .A(n12907), .B(n12908), .Z(n12899) );
  AND U12743 ( .A(n357), .B(n12909), .Z(n12908) );
  XNOR U12744 ( .A(n12910), .B(n12911), .Z(n12905) );
  AND U12745 ( .A(n349), .B(n12912), .Z(n12911) );
  XOR U12746 ( .A(p_input[847]), .B(n12910), .Z(n12912) );
  XNOR U12747 ( .A(n12913), .B(n12914), .Z(n12910) );
  AND U12748 ( .A(n353), .B(n12909), .Z(n12914) );
  XNOR U12749 ( .A(n12913), .B(n12907), .Z(n12909) );
  XOR U12750 ( .A(n12915), .B(n12916), .Z(n12907) );
  AND U12751 ( .A(n368), .B(n12917), .Z(n12916) );
  XNOR U12752 ( .A(n12918), .B(n12919), .Z(n12913) );
  AND U12753 ( .A(n360), .B(n12920), .Z(n12919) );
  XOR U12754 ( .A(p_input[879]), .B(n12918), .Z(n12920) );
  XNOR U12755 ( .A(n12921), .B(n12922), .Z(n12918) );
  AND U12756 ( .A(n364), .B(n12917), .Z(n12922) );
  XNOR U12757 ( .A(n12921), .B(n12915), .Z(n12917) );
  XOR U12758 ( .A(n12923), .B(n12924), .Z(n12915) );
  AND U12759 ( .A(n379), .B(n12925), .Z(n12924) );
  XNOR U12760 ( .A(n12926), .B(n12927), .Z(n12921) );
  AND U12761 ( .A(n371), .B(n12928), .Z(n12927) );
  XOR U12762 ( .A(p_input[911]), .B(n12926), .Z(n12928) );
  XNOR U12763 ( .A(n12929), .B(n12930), .Z(n12926) );
  AND U12764 ( .A(n375), .B(n12925), .Z(n12930) );
  XNOR U12765 ( .A(n12929), .B(n12923), .Z(n12925) );
  XOR U12766 ( .A(n12931), .B(n12932), .Z(n12923) );
  AND U12767 ( .A(n390), .B(n12933), .Z(n12932) );
  XNOR U12768 ( .A(n12934), .B(n12935), .Z(n12929) );
  AND U12769 ( .A(n382), .B(n12936), .Z(n12935) );
  XOR U12770 ( .A(p_input[943]), .B(n12934), .Z(n12936) );
  XNOR U12771 ( .A(n12937), .B(n12938), .Z(n12934) );
  AND U12772 ( .A(n386), .B(n12933), .Z(n12938) );
  XNOR U12773 ( .A(n12937), .B(n12931), .Z(n12933) );
  XOR U12774 ( .A(n12939), .B(n12940), .Z(n12931) );
  AND U12775 ( .A(n401), .B(n12941), .Z(n12940) );
  XNOR U12776 ( .A(n12942), .B(n12943), .Z(n12937) );
  AND U12777 ( .A(n393), .B(n12944), .Z(n12943) );
  XOR U12778 ( .A(p_input[975]), .B(n12942), .Z(n12944) );
  XNOR U12779 ( .A(n12945), .B(n12946), .Z(n12942) );
  AND U12780 ( .A(n397), .B(n12941), .Z(n12946) );
  XNOR U12781 ( .A(n12945), .B(n12939), .Z(n12941) );
  XOR U12782 ( .A(n12947), .B(n12948), .Z(n12939) );
  AND U12783 ( .A(n412), .B(n12949), .Z(n12948) );
  XNOR U12784 ( .A(n12950), .B(n12951), .Z(n12945) );
  AND U12785 ( .A(n404), .B(n12952), .Z(n12951) );
  XOR U12786 ( .A(p_input[1007]), .B(n12950), .Z(n12952) );
  XNOR U12787 ( .A(n12953), .B(n12954), .Z(n12950) );
  AND U12788 ( .A(n408), .B(n12949), .Z(n12954) );
  XNOR U12789 ( .A(n12953), .B(n12947), .Z(n12949) );
  XOR U12790 ( .A(n12955), .B(n12956), .Z(n12947) );
  AND U12791 ( .A(n423), .B(n12957), .Z(n12956) );
  XNOR U12792 ( .A(n12958), .B(n12959), .Z(n12953) );
  AND U12793 ( .A(n415), .B(n12960), .Z(n12959) );
  XOR U12794 ( .A(p_input[1039]), .B(n12958), .Z(n12960) );
  XNOR U12795 ( .A(n12961), .B(n12962), .Z(n12958) );
  AND U12796 ( .A(n419), .B(n12957), .Z(n12962) );
  XNOR U12797 ( .A(n12961), .B(n12955), .Z(n12957) );
  XOR U12798 ( .A(n12963), .B(n12964), .Z(n12955) );
  AND U12799 ( .A(n434), .B(n12965), .Z(n12964) );
  XNOR U12800 ( .A(n12966), .B(n12967), .Z(n12961) );
  AND U12801 ( .A(n426), .B(n12968), .Z(n12967) );
  XOR U12802 ( .A(p_input[1071]), .B(n12966), .Z(n12968) );
  XNOR U12803 ( .A(n12969), .B(n12970), .Z(n12966) );
  AND U12804 ( .A(n430), .B(n12965), .Z(n12970) );
  XNOR U12805 ( .A(n12969), .B(n12963), .Z(n12965) );
  XOR U12806 ( .A(n12971), .B(n12972), .Z(n12963) );
  AND U12807 ( .A(n445), .B(n12973), .Z(n12972) );
  XNOR U12808 ( .A(n12974), .B(n12975), .Z(n12969) );
  AND U12809 ( .A(n437), .B(n12976), .Z(n12975) );
  XOR U12810 ( .A(p_input[1103]), .B(n12974), .Z(n12976) );
  XNOR U12811 ( .A(n12977), .B(n12978), .Z(n12974) );
  AND U12812 ( .A(n441), .B(n12973), .Z(n12978) );
  XNOR U12813 ( .A(n12977), .B(n12971), .Z(n12973) );
  XOR U12814 ( .A(n12979), .B(n12980), .Z(n12971) );
  AND U12815 ( .A(n456), .B(n12981), .Z(n12980) );
  XNOR U12816 ( .A(n12982), .B(n12983), .Z(n12977) );
  AND U12817 ( .A(n448), .B(n12984), .Z(n12983) );
  XOR U12818 ( .A(p_input[1135]), .B(n12982), .Z(n12984) );
  XNOR U12819 ( .A(n12985), .B(n12986), .Z(n12982) );
  AND U12820 ( .A(n452), .B(n12981), .Z(n12986) );
  XNOR U12821 ( .A(n12985), .B(n12979), .Z(n12981) );
  XOR U12822 ( .A(n12987), .B(n12988), .Z(n12979) );
  AND U12823 ( .A(n467), .B(n12989), .Z(n12988) );
  XNOR U12824 ( .A(n12990), .B(n12991), .Z(n12985) );
  AND U12825 ( .A(n459), .B(n12992), .Z(n12991) );
  XOR U12826 ( .A(p_input[1167]), .B(n12990), .Z(n12992) );
  XNOR U12827 ( .A(n12993), .B(n12994), .Z(n12990) );
  AND U12828 ( .A(n463), .B(n12989), .Z(n12994) );
  XNOR U12829 ( .A(n12993), .B(n12987), .Z(n12989) );
  XOR U12830 ( .A(n12995), .B(n12996), .Z(n12987) );
  AND U12831 ( .A(n478), .B(n12997), .Z(n12996) );
  XNOR U12832 ( .A(n12998), .B(n12999), .Z(n12993) );
  AND U12833 ( .A(n470), .B(n13000), .Z(n12999) );
  XOR U12834 ( .A(p_input[1199]), .B(n12998), .Z(n13000) );
  XNOR U12835 ( .A(n13001), .B(n13002), .Z(n12998) );
  AND U12836 ( .A(n474), .B(n12997), .Z(n13002) );
  XNOR U12837 ( .A(n13001), .B(n12995), .Z(n12997) );
  XOR U12838 ( .A(n13003), .B(n13004), .Z(n12995) );
  AND U12839 ( .A(n489), .B(n13005), .Z(n13004) );
  XNOR U12840 ( .A(n13006), .B(n13007), .Z(n13001) );
  AND U12841 ( .A(n481), .B(n13008), .Z(n13007) );
  XOR U12842 ( .A(p_input[1231]), .B(n13006), .Z(n13008) );
  XNOR U12843 ( .A(n13009), .B(n13010), .Z(n13006) );
  AND U12844 ( .A(n485), .B(n13005), .Z(n13010) );
  XNOR U12845 ( .A(n13009), .B(n13003), .Z(n13005) );
  XOR U12846 ( .A(n13011), .B(n13012), .Z(n13003) );
  AND U12847 ( .A(n500), .B(n13013), .Z(n13012) );
  XNOR U12848 ( .A(n13014), .B(n13015), .Z(n13009) );
  AND U12849 ( .A(n492), .B(n13016), .Z(n13015) );
  XOR U12850 ( .A(p_input[1263]), .B(n13014), .Z(n13016) );
  XNOR U12851 ( .A(n13017), .B(n13018), .Z(n13014) );
  AND U12852 ( .A(n496), .B(n13013), .Z(n13018) );
  XNOR U12853 ( .A(n13017), .B(n13011), .Z(n13013) );
  XOR U12854 ( .A(n13019), .B(n13020), .Z(n13011) );
  AND U12855 ( .A(n511), .B(n13021), .Z(n13020) );
  XNOR U12856 ( .A(n13022), .B(n13023), .Z(n13017) );
  AND U12857 ( .A(n503), .B(n13024), .Z(n13023) );
  XOR U12858 ( .A(p_input[1295]), .B(n13022), .Z(n13024) );
  XNOR U12859 ( .A(n13025), .B(n13026), .Z(n13022) );
  AND U12860 ( .A(n507), .B(n13021), .Z(n13026) );
  XNOR U12861 ( .A(n13025), .B(n13019), .Z(n13021) );
  XOR U12862 ( .A(n13027), .B(n13028), .Z(n13019) );
  AND U12863 ( .A(n522), .B(n13029), .Z(n13028) );
  XNOR U12864 ( .A(n13030), .B(n13031), .Z(n13025) );
  AND U12865 ( .A(n514), .B(n13032), .Z(n13031) );
  XOR U12866 ( .A(p_input[1327]), .B(n13030), .Z(n13032) );
  XNOR U12867 ( .A(n13033), .B(n13034), .Z(n13030) );
  AND U12868 ( .A(n518), .B(n13029), .Z(n13034) );
  XNOR U12869 ( .A(n13033), .B(n13027), .Z(n13029) );
  XOR U12870 ( .A(n13035), .B(n13036), .Z(n13027) );
  AND U12871 ( .A(n533), .B(n13037), .Z(n13036) );
  XNOR U12872 ( .A(n13038), .B(n13039), .Z(n13033) );
  AND U12873 ( .A(n525), .B(n13040), .Z(n13039) );
  XOR U12874 ( .A(p_input[1359]), .B(n13038), .Z(n13040) );
  XNOR U12875 ( .A(n13041), .B(n13042), .Z(n13038) );
  AND U12876 ( .A(n529), .B(n13037), .Z(n13042) );
  XNOR U12877 ( .A(n13041), .B(n13035), .Z(n13037) );
  XOR U12878 ( .A(n13043), .B(n13044), .Z(n13035) );
  AND U12879 ( .A(n544), .B(n13045), .Z(n13044) );
  XNOR U12880 ( .A(n13046), .B(n13047), .Z(n13041) );
  AND U12881 ( .A(n536), .B(n13048), .Z(n13047) );
  XOR U12882 ( .A(p_input[1391]), .B(n13046), .Z(n13048) );
  XNOR U12883 ( .A(n13049), .B(n13050), .Z(n13046) );
  AND U12884 ( .A(n540), .B(n13045), .Z(n13050) );
  XNOR U12885 ( .A(n13049), .B(n13043), .Z(n13045) );
  XOR U12886 ( .A(n13051), .B(n13052), .Z(n13043) );
  AND U12887 ( .A(n555), .B(n13053), .Z(n13052) );
  XNOR U12888 ( .A(n13054), .B(n13055), .Z(n13049) );
  AND U12889 ( .A(n547), .B(n13056), .Z(n13055) );
  XOR U12890 ( .A(p_input[1423]), .B(n13054), .Z(n13056) );
  XNOR U12891 ( .A(n13057), .B(n13058), .Z(n13054) );
  AND U12892 ( .A(n551), .B(n13053), .Z(n13058) );
  XNOR U12893 ( .A(n13057), .B(n13051), .Z(n13053) );
  XOR U12894 ( .A(n13059), .B(n13060), .Z(n13051) );
  AND U12895 ( .A(n566), .B(n13061), .Z(n13060) );
  XNOR U12896 ( .A(n13062), .B(n13063), .Z(n13057) );
  AND U12897 ( .A(n558), .B(n13064), .Z(n13063) );
  XOR U12898 ( .A(p_input[1455]), .B(n13062), .Z(n13064) );
  XNOR U12899 ( .A(n13065), .B(n13066), .Z(n13062) );
  AND U12900 ( .A(n562), .B(n13061), .Z(n13066) );
  XNOR U12901 ( .A(n13065), .B(n13059), .Z(n13061) );
  XOR U12902 ( .A(n13067), .B(n13068), .Z(n13059) );
  AND U12903 ( .A(n577), .B(n13069), .Z(n13068) );
  XNOR U12904 ( .A(n13070), .B(n13071), .Z(n13065) );
  AND U12905 ( .A(n569), .B(n13072), .Z(n13071) );
  XOR U12906 ( .A(p_input[1487]), .B(n13070), .Z(n13072) );
  XNOR U12907 ( .A(n13073), .B(n13074), .Z(n13070) );
  AND U12908 ( .A(n573), .B(n13069), .Z(n13074) );
  XNOR U12909 ( .A(n13073), .B(n13067), .Z(n13069) );
  XOR U12910 ( .A(n13075), .B(n13076), .Z(n13067) );
  AND U12911 ( .A(n588), .B(n13077), .Z(n13076) );
  XNOR U12912 ( .A(n13078), .B(n13079), .Z(n13073) );
  AND U12913 ( .A(n580), .B(n13080), .Z(n13079) );
  XOR U12914 ( .A(p_input[1519]), .B(n13078), .Z(n13080) );
  XNOR U12915 ( .A(n13081), .B(n13082), .Z(n13078) );
  AND U12916 ( .A(n584), .B(n13077), .Z(n13082) );
  XNOR U12917 ( .A(n13081), .B(n13075), .Z(n13077) );
  XOR U12918 ( .A(n13083), .B(n13084), .Z(n13075) );
  AND U12919 ( .A(n599), .B(n13085), .Z(n13084) );
  XNOR U12920 ( .A(n13086), .B(n13087), .Z(n13081) );
  AND U12921 ( .A(n591), .B(n13088), .Z(n13087) );
  XOR U12922 ( .A(p_input[1551]), .B(n13086), .Z(n13088) );
  XNOR U12923 ( .A(n13089), .B(n13090), .Z(n13086) );
  AND U12924 ( .A(n595), .B(n13085), .Z(n13090) );
  XNOR U12925 ( .A(n13089), .B(n13083), .Z(n13085) );
  XOR U12926 ( .A(n13091), .B(n13092), .Z(n13083) );
  AND U12927 ( .A(n610), .B(n13093), .Z(n13092) );
  XNOR U12928 ( .A(n13094), .B(n13095), .Z(n13089) );
  AND U12929 ( .A(n602), .B(n13096), .Z(n13095) );
  XOR U12930 ( .A(p_input[1583]), .B(n13094), .Z(n13096) );
  XNOR U12931 ( .A(n13097), .B(n13098), .Z(n13094) );
  AND U12932 ( .A(n606), .B(n13093), .Z(n13098) );
  XNOR U12933 ( .A(n13097), .B(n13091), .Z(n13093) );
  XOR U12934 ( .A(n13099), .B(n13100), .Z(n13091) );
  AND U12935 ( .A(n621), .B(n13101), .Z(n13100) );
  XNOR U12936 ( .A(n13102), .B(n13103), .Z(n13097) );
  AND U12937 ( .A(n613), .B(n13104), .Z(n13103) );
  XOR U12938 ( .A(p_input[1615]), .B(n13102), .Z(n13104) );
  XNOR U12939 ( .A(n13105), .B(n13106), .Z(n13102) );
  AND U12940 ( .A(n617), .B(n13101), .Z(n13106) );
  XNOR U12941 ( .A(n13105), .B(n13099), .Z(n13101) );
  XOR U12942 ( .A(n13107), .B(n13108), .Z(n13099) );
  AND U12943 ( .A(n632), .B(n13109), .Z(n13108) );
  XNOR U12944 ( .A(n13110), .B(n13111), .Z(n13105) );
  AND U12945 ( .A(n624), .B(n13112), .Z(n13111) );
  XOR U12946 ( .A(p_input[1647]), .B(n13110), .Z(n13112) );
  XNOR U12947 ( .A(n13113), .B(n13114), .Z(n13110) );
  AND U12948 ( .A(n628), .B(n13109), .Z(n13114) );
  XNOR U12949 ( .A(n13113), .B(n13107), .Z(n13109) );
  XOR U12950 ( .A(n13115), .B(n13116), .Z(n13107) );
  AND U12951 ( .A(n643), .B(n13117), .Z(n13116) );
  XNOR U12952 ( .A(n13118), .B(n13119), .Z(n13113) );
  AND U12953 ( .A(n635), .B(n13120), .Z(n13119) );
  XOR U12954 ( .A(p_input[1679]), .B(n13118), .Z(n13120) );
  XNOR U12955 ( .A(n13121), .B(n13122), .Z(n13118) );
  AND U12956 ( .A(n639), .B(n13117), .Z(n13122) );
  XNOR U12957 ( .A(n13121), .B(n13115), .Z(n13117) );
  XOR U12958 ( .A(n13123), .B(n13124), .Z(n13115) );
  AND U12959 ( .A(n654), .B(n13125), .Z(n13124) );
  XNOR U12960 ( .A(n13126), .B(n13127), .Z(n13121) );
  AND U12961 ( .A(n646), .B(n13128), .Z(n13127) );
  XOR U12962 ( .A(p_input[1711]), .B(n13126), .Z(n13128) );
  XNOR U12963 ( .A(n13129), .B(n13130), .Z(n13126) );
  AND U12964 ( .A(n650), .B(n13125), .Z(n13130) );
  XNOR U12965 ( .A(n13129), .B(n13123), .Z(n13125) );
  XOR U12966 ( .A(n13131), .B(n13132), .Z(n13123) );
  AND U12967 ( .A(n665), .B(n13133), .Z(n13132) );
  XNOR U12968 ( .A(n13134), .B(n13135), .Z(n13129) );
  AND U12969 ( .A(n657), .B(n13136), .Z(n13135) );
  XOR U12970 ( .A(p_input[1743]), .B(n13134), .Z(n13136) );
  XNOR U12971 ( .A(n13137), .B(n13138), .Z(n13134) );
  AND U12972 ( .A(n661), .B(n13133), .Z(n13138) );
  XNOR U12973 ( .A(n13137), .B(n13131), .Z(n13133) );
  XOR U12974 ( .A(n13139), .B(n13140), .Z(n13131) );
  AND U12975 ( .A(n676), .B(n13141), .Z(n13140) );
  XNOR U12976 ( .A(n13142), .B(n13143), .Z(n13137) );
  AND U12977 ( .A(n668), .B(n13144), .Z(n13143) );
  XOR U12978 ( .A(p_input[1775]), .B(n13142), .Z(n13144) );
  XNOR U12979 ( .A(n13145), .B(n13146), .Z(n13142) );
  AND U12980 ( .A(n672), .B(n13141), .Z(n13146) );
  XNOR U12981 ( .A(n13145), .B(n13139), .Z(n13141) );
  XOR U12982 ( .A(n13147), .B(n13148), .Z(n13139) );
  AND U12983 ( .A(n687), .B(n13149), .Z(n13148) );
  XNOR U12984 ( .A(n13150), .B(n13151), .Z(n13145) );
  AND U12985 ( .A(n679), .B(n13152), .Z(n13151) );
  XOR U12986 ( .A(p_input[1807]), .B(n13150), .Z(n13152) );
  XNOR U12987 ( .A(n13153), .B(n13154), .Z(n13150) );
  AND U12988 ( .A(n683), .B(n13149), .Z(n13154) );
  XNOR U12989 ( .A(n13153), .B(n13147), .Z(n13149) );
  XOR U12990 ( .A(n13155), .B(n13156), .Z(n13147) );
  AND U12991 ( .A(n698), .B(n13157), .Z(n13156) );
  XNOR U12992 ( .A(n13158), .B(n13159), .Z(n13153) );
  AND U12993 ( .A(n690), .B(n13160), .Z(n13159) );
  XOR U12994 ( .A(p_input[1839]), .B(n13158), .Z(n13160) );
  XNOR U12995 ( .A(n13161), .B(n13162), .Z(n13158) );
  AND U12996 ( .A(n694), .B(n13157), .Z(n13162) );
  XNOR U12997 ( .A(n13161), .B(n13155), .Z(n13157) );
  XOR U12998 ( .A(n13163), .B(n13164), .Z(n13155) );
  AND U12999 ( .A(n709), .B(n13165), .Z(n13164) );
  XNOR U13000 ( .A(n13166), .B(n13167), .Z(n13161) );
  AND U13001 ( .A(n701), .B(n13168), .Z(n13167) );
  XOR U13002 ( .A(p_input[1871]), .B(n13166), .Z(n13168) );
  XNOR U13003 ( .A(n13169), .B(n13170), .Z(n13166) );
  AND U13004 ( .A(n705), .B(n13165), .Z(n13170) );
  XNOR U13005 ( .A(n13169), .B(n13163), .Z(n13165) );
  XOR U13006 ( .A(n13171), .B(n13172), .Z(n13163) );
  AND U13007 ( .A(n720), .B(n13173), .Z(n13172) );
  XNOR U13008 ( .A(n13174), .B(n13175), .Z(n13169) );
  AND U13009 ( .A(n712), .B(n13176), .Z(n13175) );
  XOR U13010 ( .A(p_input[1903]), .B(n13174), .Z(n13176) );
  XNOR U13011 ( .A(n13177), .B(n13178), .Z(n13174) );
  AND U13012 ( .A(n716), .B(n13173), .Z(n13178) );
  XNOR U13013 ( .A(n13177), .B(n13171), .Z(n13173) );
  XOR U13014 ( .A(n13179), .B(n13180), .Z(n13171) );
  AND U13015 ( .A(n731), .B(n13181), .Z(n13180) );
  XNOR U13016 ( .A(n13182), .B(n13183), .Z(n13177) );
  AND U13017 ( .A(n723), .B(n13184), .Z(n13183) );
  XOR U13018 ( .A(p_input[1935]), .B(n13182), .Z(n13184) );
  XNOR U13019 ( .A(n13185), .B(n13186), .Z(n13182) );
  AND U13020 ( .A(n727), .B(n13181), .Z(n13186) );
  XNOR U13021 ( .A(n13185), .B(n13179), .Z(n13181) );
  XOR U13022 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n13187), .Z(n13179) );
  AND U13023 ( .A(n741), .B(n13188), .Z(n13187) );
  XNOR U13024 ( .A(n13189), .B(n13190), .Z(n13185) );
  AND U13025 ( .A(n734), .B(n13191), .Z(n13190) );
  XOR U13026 ( .A(p_input[1967]), .B(n13189), .Z(n13191) );
  XNOR U13027 ( .A(n13192), .B(n13193), .Z(n13189) );
  AND U13028 ( .A(n738), .B(n13188), .Z(n13193) );
  XOR U13029 ( .A(n13194), .B(n13192), .Z(n13188) );
  IV U13030 ( .A(\knn_comb_/min_val_out[0][15] ), .Z(n13194) );
  IV U13031 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .Z(n13192)
         );
  XOR U13032 ( .A(n47), .B(n13195), .Z(o[14]) );
  AND U13033 ( .A(n58), .B(n13196), .Z(n47) );
  XOR U13034 ( .A(n48), .B(n13195), .Z(n13196) );
  XOR U13035 ( .A(n13197), .B(n13198), .Z(n13195) );
  AND U13036 ( .A(n70), .B(n13199), .Z(n13198) );
  XOR U13037 ( .A(n13200), .B(n13201), .Z(n48) );
  AND U13038 ( .A(n62), .B(n13202), .Z(n13201) );
  XOR U13039 ( .A(p_input[14]), .B(n13200), .Z(n13202) );
  XNOR U13040 ( .A(n13203), .B(n13204), .Z(n13200) );
  AND U13041 ( .A(n66), .B(n13199), .Z(n13204) );
  XNOR U13042 ( .A(n13203), .B(n13197), .Z(n13199) );
  XOR U13043 ( .A(n13205), .B(n13206), .Z(n13197) );
  AND U13044 ( .A(n82), .B(n13207), .Z(n13206) );
  XNOR U13045 ( .A(n13208), .B(n13209), .Z(n13203) );
  AND U13046 ( .A(n74), .B(n13210), .Z(n13209) );
  XOR U13047 ( .A(p_input[46]), .B(n13208), .Z(n13210) );
  XNOR U13048 ( .A(n13211), .B(n13212), .Z(n13208) );
  AND U13049 ( .A(n78), .B(n13207), .Z(n13212) );
  XNOR U13050 ( .A(n13211), .B(n13205), .Z(n13207) );
  XOR U13051 ( .A(n13213), .B(n13214), .Z(n13205) );
  AND U13052 ( .A(n93), .B(n13215), .Z(n13214) );
  XNOR U13053 ( .A(n13216), .B(n13217), .Z(n13211) );
  AND U13054 ( .A(n85), .B(n13218), .Z(n13217) );
  XOR U13055 ( .A(p_input[78]), .B(n13216), .Z(n13218) );
  XNOR U13056 ( .A(n13219), .B(n13220), .Z(n13216) );
  AND U13057 ( .A(n89), .B(n13215), .Z(n13220) );
  XNOR U13058 ( .A(n13219), .B(n13213), .Z(n13215) );
  XOR U13059 ( .A(n13221), .B(n13222), .Z(n13213) );
  AND U13060 ( .A(n104), .B(n13223), .Z(n13222) );
  XNOR U13061 ( .A(n13224), .B(n13225), .Z(n13219) );
  AND U13062 ( .A(n96), .B(n13226), .Z(n13225) );
  XOR U13063 ( .A(p_input[110]), .B(n13224), .Z(n13226) );
  XNOR U13064 ( .A(n13227), .B(n13228), .Z(n13224) );
  AND U13065 ( .A(n100), .B(n13223), .Z(n13228) );
  XNOR U13066 ( .A(n13227), .B(n13221), .Z(n13223) );
  XOR U13067 ( .A(n13229), .B(n13230), .Z(n13221) );
  AND U13068 ( .A(n115), .B(n13231), .Z(n13230) );
  XNOR U13069 ( .A(n13232), .B(n13233), .Z(n13227) );
  AND U13070 ( .A(n107), .B(n13234), .Z(n13233) );
  XOR U13071 ( .A(p_input[142]), .B(n13232), .Z(n13234) );
  XNOR U13072 ( .A(n13235), .B(n13236), .Z(n13232) );
  AND U13073 ( .A(n111), .B(n13231), .Z(n13236) );
  XNOR U13074 ( .A(n13235), .B(n13229), .Z(n13231) );
  XOR U13075 ( .A(n13237), .B(n13238), .Z(n13229) );
  AND U13076 ( .A(n126), .B(n13239), .Z(n13238) );
  XNOR U13077 ( .A(n13240), .B(n13241), .Z(n13235) );
  AND U13078 ( .A(n118), .B(n13242), .Z(n13241) );
  XOR U13079 ( .A(p_input[174]), .B(n13240), .Z(n13242) );
  XNOR U13080 ( .A(n13243), .B(n13244), .Z(n13240) );
  AND U13081 ( .A(n122), .B(n13239), .Z(n13244) );
  XNOR U13082 ( .A(n13243), .B(n13237), .Z(n13239) );
  XOR U13083 ( .A(n13245), .B(n13246), .Z(n13237) );
  AND U13084 ( .A(n137), .B(n13247), .Z(n13246) );
  XNOR U13085 ( .A(n13248), .B(n13249), .Z(n13243) );
  AND U13086 ( .A(n129), .B(n13250), .Z(n13249) );
  XOR U13087 ( .A(p_input[206]), .B(n13248), .Z(n13250) );
  XNOR U13088 ( .A(n13251), .B(n13252), .Z(n13248) );
  AND U13089 ( .A(n133), .B(n13247), .Z(n13252) );
  XNOR U13090 ( .A(n13251), .B(n13245), .Z(n13247) );
  XOR U13091 ( .A(n13253), .B(n13254), .Z(n13245) );
  AND U13092 ( .A(n148), .B(n13255), .Z(n13254) );
  XNOR U13093 ( .A(n13256), .B(n13257), .Z(n13251) );
  AND U13094 ( .A(n140), .B(n13258), .Z(n13257) );
  XOR U13095 ( .A(p_input[238]), .B(n13256), .Z(n13258) );
  XNOR U13096 ( .A(n13259), .B(n13260), .Z(n13256) );
  AND U13097 ( .A(n144), .B(n13255), .Z(n13260) );
  XNOR U13098 ( .A(n13259), .B(n13253), .Z(n13255) );
  XOR U13099 ( .A(n13261), .B(n13262), .Z(n13253) );
  AND U13100 ( .A(n159), .B(n13263), .Z(n13262) );
  XNOR U13101 ( .A(n13264), .B(n13265), .Z(n13259) );
  AND U13102 ( .A(n151), .B(n13266), .Z(n13265) );
  XOR U13103 ( .A(p_input[270]), .B(n13264), .Z(n13266) );
  XNOR U13104 ( .A(n13267), .B(n13268), .Z(n13264) );
  AND U13105 ( .A(n155), .B(n13263), .Z(n13268) );
  XNOR U13106 ( .A(n13267), .B(n13261), .Z(n13263) );
  XOR U13107 ( .A(n13269), .B(n13270), .Z(n13261) );
  AND U13108 ( .A(n170), .B(n13271), .Z(n13270) );
  XNOR U13109 ( .A(n13272), .B(n13273), .Z(n13267) );
  AND U13110 ( .A(n162), .B(n13274), .Z(n13273) );
  XOR U13111 ( .A(p_input[302]), .B(n13272), .Z(n13274) );
  XNOR U13112 ( .A(n13275), .B(n13276), .Z(n13272) );
  AND U13113 ( .A(n166), .B(n13271), .Z(n13276) );
  XNOR U13114 ( .A(n13275), .B(n13269), .Z(n13271) );
  XOR U13115 ( .A(n13277), .B(n13278), .Z(n13269) );
  AND U13116 ( .A(n181), .B(n13279), .Z(n13278) );
  XNOR U13117 ( .A(n13280), .B(n13281), .Z(n13275) );
  AND U13118 ( .A(n173), .B(n13282), .Z(n13281) );
  XOR U13119 ( .A(p_input[334]), .B(n13280), .Z(n13282) );
  XNOR U13120 ( .A(n13283), .B(n13284), .Z(n13280) );
  AND U13121 ( .A(n177), .B(n13279), .Z(n13284) );
  XNOR U13122 ( .A(n13283), .B(n13277), .Z(n13279) );
  XOR U13123 ( .A(n13285), .B(n13286), .Z(n13277) );
  AND U13124 ( .A(n192), .B(n13287), .Z(n13286) );
  XNOR U13125 ( .A(n13288), .B(n13289), .Z(n13283) );
  AND U13126 ( .A(n184), .B(n13290), .Z(n13289) );
  XOR U13127 ( .A(p_input[366]), .B(n13288), .Z(n13290) );
  XNOR U13128 ( .A(n13291), .B(n13292), .Z(n13288) );
  AND U13129 ( .A(n188), .B(n13287), .Z(n13292) );
  XNOR U13130 ( .A(n13291), .B(n13285), .Z(n13287) );
  XOR U13131 ( .A(n13293), .B(n13294), .Z(n13285) );
  AND U13132 ( .A(n203), .B(n13295), .Z(n13294) );
  XNOR U13133 ( .A(n13296), .B(n13297), .Z(n13291) );
  AND U13134 ( .A(n195), .B(n13298), .Z(n13297) );
  XOR U13135 ( .A(p_input[398]), .B(n13296), .Z(n13298) );
  XNOR U13136 ( .A(n13299), .B(n13300), .Z(n13296) );
  AND U13137 ( .A(n199), .B(n13295), .Z(n13300) );
  XNOR U13138 ( .A(n13299), .B(n13293), .Z(n13295) );
  XOR U13139 ( .A(n13301), .B(n13302), .Z(n13293) );
  AND U13140 ( .A(n214), .B(n13303), .Z(n13302) );
  XNOR U13141 ( .A(n13304), .B(n13305), .Z(n13299) );
  AND U13142 ( .A(n206), .B(n13306), .Z(n13305) );
  XOR U13143 ( .A(p_input[430]), .B(n13304), .Z(n13306) );
  XNOR U13144 ( .A(n13307), .B(n13308), .Z(n13304) );
  AND U13145 ( .A(n210), .B(n13303), .Z(n13308) );
  XNOR U13146 ( .A(n13307), .B(n13301), .Z(n13303) );
  XOR U13147 ( .A(n13309), .B(n13310), .Z(n13301) );
  AND U13148 ( .A(n225), .B(n13311), .Z(n13310) );
  XNOR U13149 ( .A(n13312), .B(n13313), .Z(n13307) );
  AND U13150 ( .A(n217), .B(n13314), .Z(n13313) );
  XOR U13151 ( .A(p_input[462]), .B(n13312), .Z(n13314) );
  XNOR U13152 ( .A(n13315), .B(n13316), .Z(n13312) );
  AND U13153 ( .A(n221), .B(n13311), .Z(n13316) );
  XNOR U13154 ( .A(n13315), .B(n13309), .Z(n13311) );
  XOR U13155 ( .A(n13317), .B(n13318), .Z(n13309) );
  AND U13156 ( .A(n236), .B(n13319), .Z(n13318) );
  XNOR U13157 ( .A(n13320), .B(n13321), .Z(n13315) );
  AND U13158 ( .A(n228), .B(n13322), .Z(n13321) );
  XOR U13159 ( .A(p_input[494]), .B(n13320), .Z(n13322) );
  XNOR U13160 ( .A(n13323), .B(n13324), .Z(n13320) );
  AND U13161 ( .A(n232), .B(n13319), .Z(n13324) );
  XNOR U13162 ( .A(n13323), .B(n13317), .Z(n13319) );
  XOR U13163 ( .A(n13325), .B(n13326), .Z(n13317) );
  AND U13164 ( .A(n247), .B(n13327), .Z(n13326) );
  XNOR U13165 ( .A(n13328), .B(n13329), .Z(n13323) );
  AND U13166 ( .A(n239), .B(n13330), .Z(n13329) );
  XOR U13167 ( .A(p_input[526]), .B(n13328), .Z(n13330) );
  XNOR U13168 ( .A(n13331), .B(n13332), .Z(n13328) );
  AND U13169 ( .A(n243), .B(n13327), .Z(n13332) );
  XNOR U13170 ( .A(n13331), .B(n13325), .Z(n13327) );
  XOR U13171 ( .A(n13333), .B(n13334), .Z(n13325) );
  AND U13172 ( .A(n258), .B(n13335), .Z(n13334) );
  XNOR U13173 ( .A(n13336), .B(n13337), .Z(n13331) );
  AND U13174 ( .A(n250), .B(n13338), .Z(n13337) );
  XOR U13175 ( .A(p_input[558]), .B(n13336), .Z(n13338) );
  XNOR U13176 ( .A(n13339), .B(n13340), .Z(n13336) );
  AND U13177 ( .A(n254), .B(n13335), .Z(n13340) );
  XNOR U13178 ( .A(n13339), .B(n13333), .Z(n13335) );
  XOR U13179 ( .A(n13341), .B(n13342), .Z(n13333) );
  AND U13180 ( .A(n269), .B(n13343), .Z(n13342) );
  XNOR U13181 ( .A(n13344), .B(n13345), .Z(n13339) );
  AND U13182 ( .A(n261), .B(n13346), .Z(n13345) );
  XOR U13183 ( .A(p_input[590]), .B(n13344), .Z(n13346) );
  XNOR U13184 ( .A(n13347), .B(n13348), .Z(n13344) );
  AND U13185 ( .A(n265), .B(n13343), .Z(n13348) );
  XNOR U13186 ( .A(n13347), .B(n13341), .Z(n13343) );
  XOR U13187 ( .A(n13349), .B(n13350), .Z(n13341) );
  AND U13188 ( .A(n280), .B(n13351), .Z(n13350) );
  XNOR U13189 ( .A(n13352), .B(n13353), .Z(n13347) );
  AND U13190 ( .A(n272), .B(n13354), .Z(n13353) );
  XOR U13191 ( .A(p_input[622]), .B(n13352), .Z(n13354) );
  XNOR U13192 ( .A(n13355), .B(n13356), .Z(n13352) );
  AND U13193 ( .A(n276), .B(n13351), .Z(n13356) );
  XNOR U13194 ( .A(n13355), .B(n13349), .Z(n13351) );
  XOR U13195 ( .A(n13357), .B(n13358), .Z(n13349) );
  AND U13196 ( .A(n291), .B(n13359), .Z(n13358) );
  XNOR U13197 ( .A(n13360), .B(n13361), .Z(n13355) );
  AND U13198 ( .A(n283), .B(n13362), .Z(n13361) );
  XOR U13199 ( .A(p_input[654]), .B(n13360), .Z(n13362) );
  XNOR U13200 ( .A(n13363), .B(n13364), .Z(n13360) );
  AND U13201 ( .A(n287), .B(n13359), .Z(n13364) );
  XNOR U13202 ( .A(n13363), .B(n13357), .Z(n13359) );
  XOR U13203 ( .A(n13365), .B(n13366), .Z(n13357) );
  AND U13204 ( .A(n302), .B(n13367), .Z(n13366) );
  XNOR U13205 ( .A(n13368), .B(n13369), .Z(n13363) );
  AND U13206 ( .A(n294), .B(n13370), .Z(n13369) );
  XOR U13207 ( .A(p_input[686]), .B(n13368), .Z(n13370) );
  XNOR U13208 ( .A(n13371), .B(n13372), .Z(n13368) );
  AND U13209 ( .A(n298), .B(n13367), .Z(n13372) );
  XNOR U13210 ( .A(n13371), .B(n13365), .Z(n13367) );
  XOR U13211 ( .A(n13373), .B(n13374), .Z(n13365) );
  AND U13212 ( .A(n313), .B(n13375), .Z(n13374) );
  XNOR U13213 ( .A(n13376), .B(n13377), .Z(n13371) );
  AND U13214 ( .A(n305), .B(n13378), .Z(n13377) );
  XOR U13215 ( .A(p_input[718]), .B(n13376), .Z(n13378) );
  XNOR U13216 ( .A(n13379), .B(n13380), .Z(n13376) );
  AND U13217 ( .A(n309), .B(n13375), .Z(n13380) );
  XNOR U13218 ( .A(n13379), .B(n13373), .Z(n13375) );
  XOR U13219 ( .A(n13381), .B(n13382), .Z(n13373) );
  AND U13220 ( .A(n324), .B(n13383), .Z(n13382) );
  XNOR U13221 ( .A(n13384), .B(n13385), .Z(n13379) );
  AND U13222 ( .A(n316), .B(n13386), .Z(n13385) );
  XOR U13223 ( .A(p_input[750]), .B(n13384), .Z(n13386) );
  XNOR U13224 ( .A(n13387), .B(n13388), .Z(n13384) );
  AND U13225 ( .A(n320), .B(n13383), .Z(n13388) );
  XNOR U13226 ( .A(n13387), .B(n13381), .Z(n13383) );
  XOR U13227 ( .A(n13389), .B(n13390), .Z(n13381) );
  AND U13228 ( .A(n335), .B(n13391), .Z(n13390) );
  XNOR U13229 ( .A(n13392), .B(n13393), .Z(n13387) );
  AND U13230 ( .A(n327), .B(n13394), .Z(n13393) );
  XOR U13231 ( .A(p_input[782]), .B(n13392), .Z(n13394) );
  XNOR U13232 ( .A(n13395), .B(n13396), .Z(n13392) );
  AND U13233 ( .A(n331), .B(n13391), .Z(n13396) );
  XNOR U13234 ( .A(n13395), .B(n13389), .Z(n13391) );
  XOR U13235 ( .A(n13397), .B(n13398), .Z(n13389) );
  AND U13236 ( .A(n346), .B(n13399), .Z(n13398) );
  XNOR U13237 ( .A(n13400), .B(n13401), .Z(n13395) );
  AND U13238 ( .A(n338), .B(n13402), .Z(n13401) );
  XOR U13239 ( .A(p_input[814]), .B(n13400), .Z(n13402) );
  XNOR U13240 ( .A(n13403), .B(n13404), .Z(n13400) );
  AND U13241 ( .A(n342), .B(n13399), .Z(n13404) );
  XNOR U13242 ( .A(n13403), .B(n13397), .Z(n13399) );
  XOR U13243 ( .A(n13405), .B(n13406), .Z(n13397) );
  AND U13244 ( .A(n357), .B(n13407), .Z(n13406) );
  XNOR U13245 ( .A(n13408), .B(n13409), .Z(n13403) );
  AND U13246 ( .A(n349), .B(n13410), .Z(n13409) );
  XOR U13247 ( .A(p_input[846]), .B(n13408), .Z(n13410) );
  XNOR U13248 ( .A(n13411), .B(n13412), .Z(n13408) );
  AND U13249 ( .A(n353), .B(n13407), .Z(n13412) );
  XNOR U13250 ( .A(n13411), .B(n13405), .Z(n13407) );
  XOR U13251 ( .A(n13413), .B(n13414), .Z(n13405) );
  AND U13252 ( .A(n368), .B(n13415), .Z(n13414) );
  XNOR U13253 ( .A(n13416), .B(n13417), .Z(n13411) );
  AND U13254 ( .A(n360), .B(n13418), .Z(n13417) );
  XOR U13255 ( .A(p_input[878]), .B(n13416), .Z(n13418) );
  XNOR U13256 ( .A(n13419), .B(n13420), .Z(n13416) );
  AND U13257 ( .A(n364), .B(n13415), .Z(n13420) );
  XNOR U13258 ( .A(n13419), .B(n13413), .Z(n13415) );
  XOR U13259 ( .A(n13421), .B(n13422), .Z(n13413) );
  AND U13260 ( .A(n379), .B(n13423), .Z(n13422) );
  XNOR U13261 ( .A(n13424), .B(n13425), .Z(n13419) );
  AND U13262 ( .A(n371), .B(n13426), .Z(n13425) );
  XOR U13263 ( .A(p_input[910]), .B(n13424), .Z(n13426) );
  XNOR U13264 ( .A(n13427), .B(n13428), .Z(n13424) );
  AND U13265 ( .A(n375), .B(n13423), .Z(n13428) );
  XNOR U13266 ( .A(n13427), .B(n13421), .Z(n13423) );
  XOR U13267 ( .A(n13429), .B(n13430), .Z(n13421) );
  AND U13268 ( .A(n390), .B(n13431), .Z(n13430) );
  XNOR U13269 ( .A(n13432), .B(n13433), .Z(n13427) );
  AND U13270 ( .A(n382), .B(n13434), .Z(n13433) );
  XOR U13271 ( .A(p_input[942]), .B(n13432), .Z(n13434) );
  XNOR U13272 ( .A(n13435), .B(n13436), .Z(n13432) );
  AND U13273 ( .A(n386), .B(n13431), .Z(n13436) );
  XNOR U13274 ( .A(n13435), .B(n13429), .Z(n13431) );
  XOR U13275 ( .A(n13437), .B(n13438), .Z(n13429) );
  AND U13276 ( .A(n401), .B(n13439), .Z(n13438) );
  XNOR U13277 ( .A(n13440), .B(n13441), .Z(n13435) );
  AND U13278 ( .A(n393), .B(n13442), .Z(n13441) );
  XOR U13279 ( .A(p_input[974]), .B(n13440), .Z(n13442) );
  XNOR U13280 ( .A(n13443), .B(n13444), .Z(n13440) );
  AND U13281 ( .A(n397), .B(n13439), .Z(n13444) );
  XNOR U13282 ( .A(n13443), .B(n13437), .Z(n13439) );
  XOR U13283 ( .A(n13445), .B(n13446), .Z(n13437) );
  AND U13284 ( .A(n412), .B(n13447), .Z(n13446) );
  XNOR U13285 ( .A(n13448), .B(n13449), .Z(n13443) );
  AND U13286 ( .A(n404), .B(n13450), .Z(n13449) );
  XOR U13287 ( .A(p_input[1006]), .B(n13448), .Z(n13450) );
  XNOR U13288 ( .A(n13451), .B(n13452), .Z(n13448) );
  AND U13289 ( .A(n408), .B(n13447), .Z(n13452) );
  XNOR U13290 ( .A(n13451), .B(n13445), .Z(n13447) );
  XOR U13291 ( .A(n13453), .B(n13454), .Z(n13445) );
  AND U13292 ( .A(n423), .B(n13455), .Z(n13454) );
  XNOR U13293 ( .A(n13456), .B(n13457), .Z(n13451) );
  AND U13294 ( .A(n415), .B(n13458), .Z(n13457) );
  XOR U13295 ( .A(p_input[1038]), .B(n13456), .Z(n13458) );
  XNOR U13296 ( .A(n13459), .B(n13460), .Z(n13456) );
  AND U13297 ( .A(n419), .B(n13455), .Z(n13460) );
  XNOR U13298 ( .A(n13459), .B(n13453), .Z(n13455) );
  XOR U13299 ( .A(n13461), .B(n13462), .Z(n13453) );
  AND U13300 ( .A(n434), .B(n13463), .Z(n13462) );
  XNOR U13301 ( .A(n13464), .B(n13465), .Z(n13459) );
  AND U13302 ( .A(n426), .B(n13466), .Z(n13465) );
  XOR U13303 ( .A(p_input[1070]), .B(n13464), .Z(n13466) );
  XNOR U13304 ( .A(n13467), .B(n13468), .Z(n13464) );
  AND U13305 ( .A(n430), .B(n13463), .Z(n13468) );
  XNOR U13306 ( .A(n13467), .B(n13461), .Z(n13463) );
  XOR U13307 ( .A(n13469), .B(n13470), .Z(n13461) );
  AND U13308 ( .A(n445), .B(n13471), .Z(n13470) );
  XNOR U13309 ( .A(n13472), .B(n13473), .Z(n13467) );
  AND U13310 ( .A(n437), .B(n13474), .Z(n13473) );
  XOR U13311 ( .A(p_input[1102]), .B(n13472), .Z(n13474) );
  XNOR U13312 ( .A(n13475), .B(n13476), .Z(n13472) );
  AND U13313 ( .A(n441), .B(n13471), .Z(n13476) );
  XNOR U13314 ( .A(n13475), .B(n13469), .Z(n13471) );
  XOR U13315 ( .A(n13477), .B(n13478), .Z(n13469) );
  AND U13316 ( .A(n456), .B(n13479), .Z(n13478) );
  XNOR U13317 ( .A(n13480), .B(n13481), .Z(n13475) );
  AND U13318 ( .A(n448), .B(n13482), .Z(n13481) );
  XOR U13319 ( .A(p_input[1134]), .B(n13480), .Z(n13482) );
  XNOR U13320 ( .A(n13483), .B(n13484), .Z(n13480) );
  AND U13321 ( .A(n452), .B(n13479), .Z(n13484) );
  XNOR U13322 ( .A(n13483), .B(n13477), .Z(n13479) );
  XOR U13323 ( .A(n13485), .B(n13486), .Z(n13477) );
  AND U13324 ( .A(n467), .B(n13487), .Z(n13486) );
  XNOR U13325 ( .A(n13488), .B(n13489), .Z(n13483) );
  AND U13326 ( .A(n459), .B(n13490), .Z(n13489) );
  XOR U13327 ( .A(p_input[1166]), .B(n13488), .Z(n13490) );
  XNOR U13328 ( .A(n13491), .B(n13492), .Z(n13488) );
  AND U13329 ( .A(n463), .B(n13487), .Z(n13492) );
  XNOR U13330 ( .A(n13491), .B(n13485), .Z(n13487) );
  XOR U13331 ( .A(n13493), .B(n13494), .Z(n13485) );
  AND U13332 ( .A(n478), .B(n13495), .Z(n13494) );
  XNOR U13333 ( .A(n13496), .B(n13497), .Z(n13491) );
  AND U13334 ( .A(n470), .B(n13498), .Z(n13497) );
  XOR U13335 ( .A(p_input[1198]), .B(n13496), .Z(n13498) );
  XNOR U13336 ( .A(n13499), .B(n13500), .Z(n13496) );
  AND U13337 ( .A(n474), .B(n13495), .Z(n13500) );
  XNOR U13338 ( .A(n13499), .B(n13493), .Z(n13495) );
  XOR U13339 ( .A(n13501), .B(n13502), .Z(n13493) );
  AND U13340 ( .A(n489), .B(n13503), .Z(n13502) );
  XNOR U13341 ( .A(n13504), .B(n13505), .Z(n13499) );
  AND U13342 ( .A(n481), .B(n13506), .Z(n13505) );
  XOR U13343 ( .A(p_input[1230]), .B(n13504), .Z(n13506) );
  XNOR U13344 ( .A(n13507), .B(n13508), .Z(n13504) );
  AND U13345 ( .A(n485), .B(n13503), .Z(n13508) );
  XNOR U13346 ( .A(n13507), .B(n13501), .Z(n13503) );
  XOR U13347 ( .A(n13509), .B(n13510), .Z(n13501) );
  AND U13348 ( .A(n500), .B(n13511), .Z(n13510) );
  XNOR U13349 ( .A(n13512), .B(n13513), .Z(n13507) );
  AND U13350 ( .A(n492), .B(n13514), .Z(n13513) );
  XOR U13351 ( .A(p_input[1262]), .B(n13512), .Z(n13514) );
  XNOR U13352 ( .A(n13515), .B(n13516), .Z(n13512) );
  AND U13353 ( .A(n496), .B(n13511), .Z(n13516) );
  XNOR U13354 ( .A(n13515), .B(n13509), .Z(n13511) );
  XOR U13355 ( .A(n13517), .B(n13518), .Z(n13509) );
  AND U13356 ( .A(n511), .B(n13519), .Z(n13518) );
  XNOR U13357 ( .A(n13520), .B(n13521), .Z(n13515) );
  AND U13358 ( .A(n503), .B(n13522), .Z(n13521) );
  XOR U13359 ( .A(p_input[1294]), .B(n13520), .Z(n13522) );
  XNOR U13360 ( .A(n13523), .B(n13524), .Z(n13520) );
  AND U13361 ( .A(n507), .B(n13519), .Z(n13524) );
  XNOR U13362 ( .A(n13523), .B(n13517), .Z(n13519) );
  XOR U13363 ( .A(n13525), .B(n13526), .Z(n13517) );
  AND U13364 ( .A(n522), .B(n13527), .Z(n13526) );
  XNOR U13365 ( .A(n13528), .B(n13529), .Z(n13523) );
  AND U13366 ( .A(n514), .B(n13530), .Z(n13529) );
  XOR U13367 ( .A(p_input[1326]), .B(n13528), .Z(n13530) );
  XNOR U13368 ( .A(n13531), .B(n13532), .Z(n13528) );
  AND U13369 ( .A(n518), .B(n13527), .Z(n13532) );
  XNOR U13370 ( .A(n13531), .B(n13525), .Z(n13527) );
  XOR U13371 ( .A(n13533), .B(n13534), .Z(n13525) );
  AND U13372 ( .A(n533), .B(n13535), .Z(n13534) );
  XNOR U13373 ( .A(n13536), .B(n13537), .Z(n13531) );
  AND U13374 ( .A(n525), .B(n13538), .Z(n13537) );
  XOR U13375 ( .A(p_input[1358]), .B(n13536), .Z(n13538) );
  XNOR U13376 ( .A(n13539), .B(n13540), .Z(n13536) );
  AND U13377 ( .A(n529), .B(n13535), .Z(n13540) );
  XNOR U13378 ( .A(n13539), .B(n13533), .Z(n13535) );
  XOR U13379 ( .A(n13541), .B(n13542), .Z(n13533) );
  AND U13380 ( .A(n544), .B(n13543), .Z(n13542) );
  XNOR U13381 ( .A(n13544), .B(n13545), .Z(n13539) );
  AND U13382 ( .A(n536), .B(n13546), .Z(n13545) );
  XOR U13383 ( .A(p_input[1390]), .B(n13544), .Z(n13546) );
  XNOR U13384 ( .A(n13547), .B(n13548), .Z(n13544) );
  AND U13385 ( .A(n540), .B(n13543), .Z(n13548) );
  XNOR U13386 ( .A(n13547), .B(n13541), .Z(n13543) );
  XOR U13387 ( .A(n13549), .B(n13550), .Z(n13541) );
  AND U13388 ( .A(n555), .B(n13551), .Z(n13550) );
  XNOR U13389 ( .A(n13552), .B(n13553), .Z(n13547) );
  AND U13390 ( .A(n547), .B(n13554), .Z(n13553) );
  XOR U13391 ( .A(p_input[1422]), .B(n13552), .Z(n13554) );
  XNOR U13392 ( .A(n13555), .B(n13556), .Z(n13552) );
  AND U13393 ( .A(n551), .B(n13551), .Z(n13556) );
  XNOR U13394 ( .A(n13555), .B(n13549), .Z(n13551) );
  XOR U13395 ( .A(n13557), .B(n13558), .Z(n13549) );
  AND U13396 ( .A(n566), .B(n13559), .Z(n13558) );
  XNOR U13397 ( .A(n13560), .B(n13561), .Z(n13555) );
  AND U13398 ( .A(n558), .B(n13562), .Z(n13561) );
  XOR U13399 ( .A(p_input[1454]), .B(n13560), .Z(n13562) );
  XNOR U13400 ( .A(n13563), .B(n13564), .Z(n13560) );
  AND U13401 ( .A(n562), .B(n13559), .Z(n13564) );
  XNOR U13402 ( .A(n13563), .B(n13557), .Z(n13559) );
  XOR U13403 ( .A(n13565), .B(n13566), .Z(n13557) );
  AND U13404 ( .A(n577), .B(n13567), .Z(n13566) );
  XNOR U13405 ( .A(n13568), .B(n13569), .Z(n13563) );
  AND U13406 ( .A(n569), .B(n13570), .Z(n13569) );
  XOR U13407 ( .A(p_input[1486]), .B(n13568), .Z(n13570) );
  XNOR U13408 ( .A(n13571), .B(n13572), .Z(n13568) );
  AND U13409 ( .A(n573), .B(n13567), .Z(n13572) );
  XNOR U13410 ( .A(n13571), .B(n13565), .Z(n13567) );
  XOR U13411 ( .A(n13573), .B(n13574), .Z(n13565) );
  AND U13412 ( .A(n588), .B(n13575), .Z(n13574) );
  XNOR U13413 ( .A(n13576), .B(n13577), .Z(n13571) );
  AND U13414 ( .A(n580), .B(n13578), .Z(n13577) );
  XOR U13415 ( .A(p_input[1518]), .B(n13576), .Z(n13578) );
  XNOR U13416 ( .A(n13579), .B(n13580), .Z(n13576) );
  AND U13417 ( .A(n584), .B(n13575), .Z(n13580) );
  XNOR U13418 ( .A(n13579), .B(n13573), .Z(n13575) );
  XOR U13419 ( .A(n13581), .B(n13582), .Z(n13573) );
  AND U13420 ( .A(n599), .B(n13583), .Z(n13582) );
  XNOR U13421 ( .A(n13584), .B(n13585), .Z(n13579) );
  AND U13422 ( .A(n591), .B(n13586), .Z(n13585) );
  XOR U13423 ( .A(p_input[1550]), .B(n13584), .Z(n13586) );
  XNOR U13424 ( .A(n13587), .B(n13588), .Z(n13584) );
  AND U13425 ( .A(n595), .B(n13583), .Z(n13588) );
  XNOR U13426 ( .A(n13587), .B(n13581), .Z(n13583) );
  XOR U13427 ( .A(n13589), .B(n13590), .Z(n13581) );
  AND U13428 ( .A(n610), .B(n13591), .Z(n13590) );
  XNOR U13429 ( .A(n13592), .B(n13593), .Z(n13587) );
  AND U13430 ( .A(n602), .B(n13594), .Z(n13593) );
  XOR U13431 ( .A(p_input[1582]), .B(n13592), .Z(n13594) );
  XNOR U13432 ( .A(n13595), .B(n13596), .Z(n13592) );
  AND U13433 ( .A(n606), .B(n13591), .Z(n13596) );
  XNOR U13434 ( .A(n13595), .B(n13589), .Z(n13591) );
  XOR U13435 ( .A(n13597), .B(n13598), .Z(n13589) );
  AND U13436 ( .A(n621), .B(n13599), .Z(n13598) );
  XNOR U13437 ( .A(n13600), .B(n13601), .Z(n13595) );
  AND U13438 ( .A(n613), .B(n13602), .Z(n13601) );
  XOR U13439 ( .A(p_input[1614]), .B(n13600), .Z(n13602) );
  XNOR U13440 ( .A(n13603), .B(n13604), .Z(n13600) );
  AND U13441 ( .A(n617), .B(n13599), .Z(n13604) );
  XNOR U13442 ( .A(n13603), .B(n13597), .Z(n13599) );
  XOR U13443 ( .A(n13605), .B(n13606), .Z(n13597) );
  AND U13444 ( .A(n632), .B(n13607), .Z(n13606) );
  XNOR U13445 ( .A(n13608), .B(n13609), .Z(n13603) );
  AND U13446 ( .A(n624), .B(n13610), .Z(n13609) );
  XOR U13447 ( .A(p_input[1646]), .B(n13608), .Z(n13610) );
  XNOR U13448 ( .A(n13611), .B(n13612), .Z(n13608) );
  AND U13449 ( .A(n628), .B(n13607), .Z(n13612) );
  XNOR U13450 ( .A(n13611), .B(n13605), .Z(n13607) );
  XOR U13451 ( .A(n13613), .B(n13614), .Z(n13605) );
  AND U13452 ( .A(n643), .B(n13615), .Z(n13614) );
  XNOR U13453 ( .A(n13616), .B(n13617), .Z(n13611) );
  AND U13454 ( .A(n635), .B(n13618), .Z(n13617) );
  XOR U13455 ( .A(p_input[1678]), .B(n13616), .Z(n13618) );
  XNOR U13456 ( .A(n13619), .B(n13620), .Z(n13616) );
  AND U13457 ( .A(n639), .B(n13615), .Z(n13620) );
  XNOR U13458 ( .A(n13619), .B(n13613), .Z(n13615) );
  XOR U13459 ( .A(n13621), .B(n13622), .Z(n13613) );
  AND U13460 ( .A(n654), .B(n13623), .Z(n13622) );
  XNOR U13461 ( .A(n13624), .B(n13625), .Z(n13619) );
  AND U13462 ( .A(n646), .B(n13626), .Z(n13625) );
  XOR U13463 ( .A(p_input[1710]), .B(n13624), .Z(n13626) );
  XNOR U13464 ( .A(n13627), .B(n13628), .Z(n13624) );
  AND U13465 ( .A(n650), .B(n13623), .Z(n13628) );
  XNOR U13466 ( .A(n13627), .B(n13621), .Z(n13623) );
  XOR U13467 ( .A(n13629), .B(n13630), .Z(n13621) );
  AND U13468 ( .A(n665), .B(n13631), .Z(n13630) );
  XNOR U13469 ( .A(n13632), .B(n13633), .Z(n13627) );
  AND U13470 ( .A(n657), .B(n13634), .Z(n13633) );
  XOR U13471 ( .A(p_input[1742]), .B(n13632), .Z(n13634) );
  XNOR U13472 ( .A(n13635), .B(n13636), .Z(n13632) );
  AND U13473 ( .A(n661), .B(n13631), .Z(n13636) );
  XNOR U13474 ( .A(n13635), .B(n13629), .Z(n13631) );
  XOR U13475 ( .A(n13637), .B(n13638), .Z(n13629) );
  AND U13476 ( .A(n676), .B(n13639), .Z(n13638) );
  XNOR U13477 ( .A(n13640), .B(n13641), .Z(n13635) );
  AND U13478 ( .A(n668), .B(n13642), .Z(n13641) );
  XOR U13479 ( .A(p_input[1774]), .B(n13640), .Z(n13642) );
  XNOR U13480 ( .A(n13643), .B(n13644), .Z(n13640) );
  AND U13481 ( .A(n672), .B(n13639), .Z(n13644) );
  XNOR U13482 ( .A(n13643), .B(n13637), .Z(n13639) );
  XOR U13483 ( .A(n13645), .B(n13646), .Z(n13637) );
  AND U13484 ( .A(n687), .B(n13647), .Z(n13646) );
  XNOR U13485 ( .A(n13648), .B(n13649), .Z(n13643) );
  AND U13486 ( .A(n679), .B(n13650), .Z(n13649) );
  XOR U13487 ( .A(p_input[1806]), .B(n13648), .Z(n13650) );
  XNOR U13488 ( .A(n13651), .B(n13652), .Z(n13648) );
  AND U13489 ( .A(n683), .B(n13647), .Z(n13652) );
  XNOR U13490 ( .A(n13651), .B(n13645), .Z(n13647) );
  XOR U13491 ( .A(n13653), .B(n13654), .Z(n13645) );
  AND U13492 ( .A(n698), .B(n13655), .Z(n13654) );
  XNOR U13493 ( .A(n13656), .B(n13657), .Z(n13651) );
  AND U13494 ( .A(n690), .B(n13658), .Z(n13657) );
  XOR U13495 ( .A(p_input[1838]), .B(n13656), .Z(n13658) );
  XNOR U13496 ( .A(n13659), .B(n13660), .Z(n13656) );
  AND U13497 ( .A(n694), .B(n13655), .Z(n13660) );
  XNOR U13498 ( .A(n13659), .B(n13653), .Z(n13655) );
  XOR U13499 ( .A(n13661), .B(n13662), .Z(n13653) );
  AND U13500 ( .A(n709), .B(n13663), .Z(n13662) );
  XNOR U13501 ( .A(n13664), .B(n13665), .Z(n13659) );
  AND U13502 ( .A(n701), .B(n13666), .Z(n13665) );
  XOR U13503 ( .A(p_input[1870]), .B(n13664), .Z(n13666) );
  XNOR U13504 ( .A(n13667), .B(n13668), .Z(n13664) );
  AND U13505 ( .A(n705), .B(n13663), .Z(n13668) );
  XNOR U13506 ( .A(n13667), .B(n13661), .Z(n13663) );
  XOR U13507 ( .A(n13669), .B(n13670), .Z(n13661) );
  AND U13508 ( .A(n720), .B(n13671), .Z(n13670) );
  XNOR U13509 ( .A(n13672), .B(n13673), .Z(n13667) );
  AND U13510 ( .A(n712), .B(n13674), .Z(n13673) );
  XOR U13511 ( .A(p_input[1902]), .B(n13672), .Z(n13674) );
  XNOR U13512 ( .A(n13675), .B(n13676), .Z(n13672) );
  AND U13513 ( .A(n716), .B(n13671), .Z(n13676) );
  XNOR U13514 ( .A(n13675), .B(n13669), .Z(n13671) );
  XOR U13515 ( .A(n13677), .B(n13678), .Z(n13669) );
  AND U13516 ( .A(n731), .B(n13679), .Z(n13678) );
  XNOR U13517 ( .A(n13680), .B(n13681), .Z(n13675) );
  AND U13518 ( .A(n723), .B(n13682), .Z(n13681) );
  XOR U13519 ( .A(p_input[1934]), .B(n13680), .Z(n13682) );
  XNOR U13520 ( .A(n13683), .B(n13684), .Z(n13680) );
  AND U13521 ( .A(n727), .B(n13679), .Z(n13684) );
  XNOR U13522 ( .A(n13683), .B(n13677), .Z(n13679) );
  XOR U13523 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n13685), .Z(n13677) );
  AND U13524 ( .A(n741), .B(n13686), .Z(n13685) );
  XNOR U13525 ( .A(n13687), .B(n13688), .Z(n13683) );
  AND U13526 ( .A(n734), .B(n13689), .Z(n13688) );
  XOR U13527 ( .A(p_input[1966]), .B(n13687), .Z(n13689) );
  XNOR U13528 ( .A(n13690), .B(n13691), .Z(n13687) );
  AND U13529 ( .A(n738), .B(n13686), .Z(n13691) );
  XOR U13530 ( .A(\knn_comb_/min_val_out[0][14] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n13686) );
  XOR U13531 ( .A(n49), .B(n13692), .Z(o[13]) );
  AND U13532 ( .A(n58), .B(n13693), .Z(n49) );
  XOR U13533 ( .A(n50), .B(n13692), .Z(n13693) );
  XOR U13534 ( .A(n13694), .B(n13695), .Z(n13692) );
  AND U13535 ( .A(n70), .B(n13696), .Z(n13695) );
  XOR U13536 ( .A(n13697), .B(n13698), .Z(n50) );
  AND U13537 ( .A(n62), .B(n13699), .Z(n13698) );
  XOR U13538 ( .A(p_input[13]), .B(n13697), .Z(n13699) );
  XNOR U13539 ( .A(n13700), .B(n13701), .Z(n13697) );
  AND U13540 ( .A(n66), .B(n13696), .Z(n13701) );
  XNOR U13541 ( .A(n13700), .B(n13694), .Z(n13696) );
  XOR U13542 ( .A(n13702), .B(n13703), .Z(n13694) );
  AND U13543 ( .A(n82), .B(n13704), .Z(n13703) );
  XNOR U13544 ( .A(n13705), .B(n13706), .Z(n13700) );
  AND U13545 ( .A(n74), .B(n13707), .Z(n13706) );
  XOR U13546 ( .A(p_input[45]), .B(n13705), .Z(n13707) );
  XNOR U13547 ( .A(n13708), .B(n13709), .Z(n13705) );
  AND U13548 ( .A(n78), .B(n13704), .Z(n13709) );
  XNOR U13549 ( .A(n13708), .B(n13702), .Z(n13704) );
  XOR U13550 ( .A(n13710), .B(n13711), .Z(n13702) );
  AND U13551 ( .A(n93), .B(n13712), .Z(n13711) );
  XNOR U13552 ( .A(n13713), .B(n13714), .Z(n13708) );
  AND U13553 ( .A(n85), .B(n13715), .Z(n13714) );
  XOR U13554 ( .A(p_input[77]), .B(n13713), .Z(n13715) );
  XNOR U13555 ( .A(n13716), .B(n13717), .Z(n13713) );
  AND U13556 ( .A(n89), .B(n13712), .Z(n13717) );
  XNOR U13557 ( .A(n13716), .B(n13710), .Z(n13712) );
  XOR U13558 ( .A(n13718), .B(n13719), .Z(n13710) );
  AND U13559 ( .A(n104), .B(n13720), .Z(n13719) );
  XNOR U13560 ( .A(n13721), .B(n13722), .Z(n13716) );
  AND U13561 ( .A(n96), .B(n13723), .Z(n13722) );
  XOR U13562 ( .A(p_input[109]), .B(n13721), .Z(n13723) );
  XNOR U13563 ( .A(n13724), .B(n13725), .Z(n13721) );
  AND U13564 ( .A(n100), .B(n13720), .Z(n13725) );
  XNOR U13565 ( .A(n13724), .B(n13718), .Z(n13720) );
  XOR U13566 ( .A(n13726), .B(n13727), .Z(n13718) );
  AND U13567 ( .A(n115), .B(n13728), .Z(n13727) );
  XNOR U13568 ( .A(n13729), .B(n13730), .Z(n13724) );
  AND U13569 ( .A(n107), .B(n13731), .Z(n13730) );
  XOR U13570 ( .A(p_input[141]), .B(n13729), .Z(n13731) );
  XNOR U13571 ( .A(n13732), .B(n13733), .Z(n13729) );
  AND U13572 ( .A(n111), .B(n13728), .Z(n13733) );
  XNOR U13573 ( .A(n13732), .B(n13726), .Z(n13728) );
  XOR U13574 ( .A(n13734), .B(n13735), .Z(n13726) );
  AND U13575 ( .A(n126), .B(n13736), .Z(n13735) );
  XNOR U13576 ( .A(n13737), .B(n13738), .Z(n13732) );
  AND U13577 ( .A(n118), .B(n13739), .Z(n13738) );
  XOR U13578 ( .A(p_input[173]), .B(n13737), .Z(n13739) );
  XNOR U13579 ( .A(n13740), .B(n13741), .Z(n13737) );
  AND U13580 ( .A(n122), .B(n13736), .Z(n13741) );
  XNOR U13581 ( .A(n13740), .B(n13734), .Z(n13736) );
  XOR U13582 ( .A(n13742), .B(n13743), .Z(n13734) );
  AND U13583 ( .A(n137), .B(n13744), .Z(n13743) );
  XNOR U13584 ( .A(n13745), .B(n13746), .Z(n13740) );
  AND U13585 ( .A(n129), .B(n13747), .Z(n13746) );
  XOR U13586 ( .A(p_input[205]), .B(n13745), .Z(n13747) );
  XNOR U13587 ( .A(n13748), .B(n13749), .Z(n13745) );
  AND U13588 ( .A(n133), .B(n13744), .Z(n13749) );
  XNOR U13589 ( .A(n13748), .B(n13742), .Z(n13744) );
  XOR U13590 ( .A(n13750), .B(n13751), .Z(n13742) );
  AND U13591 ( .A(n148), .B(n13752), .Z(n13751) );
  XNOR U13592 ( .A(n13753), .B(n13754), .Z(n13748) );
  AND U13593 ( .A(n140), .B(n13755), .Z(n13754) );
  XOR U13594 ( .A(p_input[237]), .B(n13753), .Z(n13755) );
  XNOR U13595 ( .A(n13756), .B(n13757), .Z(n13753) );
  AND U13596 ( .A(n144), .B(n13752), .Z(n13757) );
  XNOR U13597 ( .A(n13756), .B(n13750), .Z(n13752) );
  XOR U13598 ( .A(n13758), .B(n13759), .Z(n13750) );
  AND U13599 ( .A(n159), .B(n13760), .Z(n13759) );
  XNOR U13600 ( .A(n13761), .B(n13762), .Z(n13756) );
  AND U13601 ( .A(n151), .B(n13763), .Z(n13762) );
  XOR U13602 ( .A(p_input[269]), .B(n13761), .Z(n13763) );
  XNOR U13603 ( .A(n13764), .B(n13765), .Z(n13761) );
  AND U13604 ( .A(n155), .B(n13760), .Z(n13765) );
  XNOR U13605 ( .A(n13764), .B(n13758), .Z(n13760) );
  XOR U13606 ( .A(n13766), .B(n13767), .Z(n13758) );
  AND U13607 ( .A(n170), .B(n13768), .Z(n13767) );
  XNOR U13608 ( .A(n13769), .B(n13770), .Z(n13764) );
  AND U13609 ( .A(n162), .B(n13771), .Z(n13770) );
  XOR U13610 ( .A(p_input[301]), .B(n13769), .Z(n13771) );
  XNOR U13611 ( .A(n13772), .B(n13773), .Z(n13769) );
  AND U13612 ( .A(n166), .B(n13768), .Z(n13773) );
  XNOR U13613 ( .A(n13772), .B(n13766), .Z(n13768) );
  XOR U13614 ( .A(n13774), .B(n13775), .Z(n13766) );
  AND U13615 ( .A(n181), .B(n13776), .Z(n13775) );
  XNOR U13616 ( .A(n13777), .B(n13778), .Z(n13772) );
  AND U13617 ( .A(n173), .B(n13779), .Z(n13778) );
  XOR U13618 ( .A(p_input[333]), .B(n13777), .Z(n13779) );
  XNOR U13619 ( .A(n13780), .B(n13781), .Z(n13777) );
  AND U13620 ( .A(n177), .B(n13776), .Z(n13781) );
  XNOR U13621 ( .A(n13780), .B(n13774), .Z(n13776) );
  XOR U13622 ( .A(n13782), .B(n13783), .Z(n13774) );
  AND U13623 ( .A(n192), .B(n13784), .Z(n13783) );
  XNOR U13624 ( .A(n13785), .B(n13786), .Z(n13780) );
  AND U13625 ( .A(n184), .B(n13787), .Z(n13786) );
  XOR U13626 ( .A(p_input[365]), .B(n13785), .Z(n13787) );
  XNOR U13627 ( .A(n13788), .B(n13789), .Z(n13785) );
  AND U13628 ( .A(n188), .B(n13784), .Z(n13789) );
  XNOR U13629 ( .A(n13788), .B(n13782), .Z(n13784) );
  XOR U13630 ( .A(n13790), .B(n13791), .Z(n13782) );
  AND U13631 ( .A(n203), .B(n13792), .Z(n13791) );
  XNOR U13632 ( .A(n13793), .B(n13794), .Z(n13788) );
  AND U13633 ( .A(n195), .B(n13795), .Z(n13794) );
  XOR U13634 ( .A(p_input[397]), .B(n13793), .Z(n13795) );
  XNOR U13635 ( .A(n13796), .B(n13797), .Z(n13793) );
  AND U13636 ( .A(n199), .B(n13792), .Z(n13797) );
  XNOR U13637 ( .A(n13796), .B(n13790), .Z(n13792) );
  XOR U13638 ( .A(n13798), .B(n13799), .Z(n13790) );
  AND U13639 ( .A(n214), .B(n13800), .Z(n13799) );
  XNOR U13640 ( .A(n13801), .B(n13802), .Z(n13796) );
  AND U13641 ( .A(n206), .B(n13803), .Z(n13802) );
  XOR U13642 ( .A(p_input[429]), .B(n13801), .Z(n13803) );
  XNOR U13643 ( .A(n13804), .B(n13805), .Z(n13801) );
  AND U13644 ( .A(n210), .B(n13800), .Z(n13805) );
  XNOR U13645 ( .A(n13804), .B(n13798), .Z(n13800) );
  XOR U13646 ( .A(n13806), .B(n13807), .Z(n13798) );
  AND U13647 ( .A(n225), .B(n13808), .Z(n13807) );
  XNOR U13648 ( .A(n13809), .B(n13810), .Z(n13804) );
  AND U13649 ( .A(n217), .B(n13811), .Z(n13810) );
  XOR U13650 ( .A(p_input[461]), .B(n13809), .Z(n13811) );
  XNOR U13651 ( .A(n13812), .B(n13813), .Z(n13809) );
  AND U13652 ( .A(n221), .B(n13808), .Z(n13813) );
  XNOR U13653 ( .A(n13812), .B(n13806), .Z(n13808) );
  XOR U13654 ( .A(n13814), .B(n13815), .Z(n13806) );
  AND U13655 ( .A(n236), .B(n13816), .Z(n13815) );
  XNOR U13656 ( .A(n13817), .B(n13818), .Z(n13812) );
  AND U13657 ( .A(n228), .B(n13819), .Z(n13818) );
  XOR U13658 ( .A(p_input[493]), .B(n13817), .Z(n13819) );
  XNOR U13659 ( .A(n13820), .B(n13821), .Z(n13817) );
  AND U13660 ( .A(n232), .B(n13816), .Z(n13821) );
  XNOR U13661 ( .A(n13820), .B(n13814), .Z(n13816) );
  XOR U13662 ( .A(n13822), .B(n13823), .Z(n13814) );
  AND U13663 ( .A(n247), .B(n13824), .Z(n13823) );
  XNOR U13664 ( .A(n13825), .B(n13826), .Z(n13820) );
  AND U13665 ( .A(n239), .B(n13827), .Z(n13826) );
  XOR U13666 ( .A(p_input[525]), .B(n13825), .Z(n13827) );
  XNOR U13667 ( .A(n13828), .B(n13829), .Z(n13825) );
  AND U13668 ( .A(n243), .B(n13824), .Z(n13829) );
  XNOR U13669 ( .A(n13828), .B(n13822), .Z(n13824) );
  XOR U13670 ( .A(n13830), .B(n13831), .Z(n13822) );
  AND U13671 ( .A(n258), .B(n13832), .Z(n13831) );
  XNOR U13672 ( .A(n13833), .B(n13834), .Z(n13828) );
  AND U13673 ( .A(n250), .B(n13835), .Z(n13834) );
  XOR U13674 ( .A(p_input[557]), .B(n13833), .Z(n13835) );
  XNOR U13675 ( .A(n13836), .B(n13837), .Z(n13833) );
  AND U13676 ( .A(n254), .B(n13832), .Z(n13837) );
  XNOR U13677 ( .A(n13836), .B(n13830), .Z(n13832) );
  XOR U13678 ( .A(n13838), .B(n13839), .Z(n13830) );
  AND U13679 ( .A(n269), .B(n13840), .Z(n13839) );
  XNOR U13680 ( .A(n13841), .B(n13842), .Z(n13836) );
  AND U13681 ( .A(n261), .B(n13843), .Z(n13842) );
  XOR U13682 ( .A(p_input[589]), .B(n13841), .Z(n13843) );
  XNOR U13683 ( .A(n13844), .B(n13845), .Z(n13841) );
  AND U13684 ( .A(n265), .B(n13840), .Z(n13845) );
  XNOR U13685 ( .A(n13844), .B(n13838), .Z(n13840) );
  XOR U13686 ( .A(n13846), .B(n13847), .Z(n13838) );
  AND U13687 ( .A(n280), .B(n13848), .Z(n13847) );
  XNOR U13688 ( .A(n13849), .B(n13850), .Z(n13844) );
  AND U13689 ( .A(n272), .B(n13851), .Z(n13850) );
  XOR U13690 ( .A(p_input[621]), .B(n13849), .Z(n13851) );
  XNOR U13691 ( .A(n13852), .B(n13853), .Z(n13849) );
  AND U13692 ( .A(n276), .B(n13848), .Z(n13853) );
  XNOR U13693 ( .A(n13852), .B(n13846), .Z(n13848) );
  XOR U13694 ( .A(n13854), .B(n13855), .Z(n13846) );
  AND U13695 ( .A(n291), .B(n13856), .Z(n13855) );
  XNOR U13696 ( .A(n13857), .B(n13858), .Z(n13852) );
  AND U13697 ( .A(n283), .B(n13859), .Z(n13858) );
  XOR U13698 ( .A(p_input[653]), .B(n13857), .Z(n13859) );
  XNOR U13699 ( .A(n13860), .B(n13861), .Z(n13857) );
  AND U13700 ( .A(n287), .B(n13856), .Z(n13861) );
  XNOR U13701 ( .A(n13860), .B(n13854), .Z(n13856) );
  XOR U13702 ( .A(n13862), .B(n13863), .Z(n13854) );
  AND U13703 ( .A(n302), .B(n13864), .Z(n13863) );
  XNOR U13704 ( .A(n13865), .B(n13866), .Z(n13860) );
  AND U13705 ( .A(n294), .B(n13867), .Z(n13866) );
  XOR U13706 ( .A(p_input[685]), .B(n13865), .Z(n13867) );
  XNOR U13707 ( .A(n13868), .B(n13869), .Z(n13865) );
  AND U13708 ( .A(n298), .B(n13864), .Z(n13869) );
  XNOR U13709 ( .A(n13868), .B(n13862), .Z(n13864) );
  XOR U13710 ( .A(n13870), .B(n13871), .Z(n13862) );
  AND U13711 ( .A(n313), .B(n13872), .Z(n13871) );
  XNOR U13712 ( .A(n13873), .B(n13874), .Z(n13868) );
  AND U13713 ( .A(n305), .B(n13875), .Z(n13874) );
  XOR U13714 ( .A(p_input[717]), .B(n13873), .Z(n13875) );
  XNOR U13715 ( .A(n13876), .B(n13877), .Z(n13873) );
  AND U13716 ( .A(n309), .B(n13872), .Z(n13877) );
  XNOR U13717 ( .A(n13876), .B(n13870), .Z(n13872) );
  XOR U13718 ( .A(n13878), .B(n13879), .Z(n13870) );
  AND U13719 ( .A(n324), .B(n13880), .Z(n13879) );
  XNOR U13720 ( .A(n13881), .B(n13882), .Z(n13876) );
  AND U13721 ( .A(n316), .B(n13883), .Z(n13882) );
  XOR U13722 ( .A(p_input[749]), .B(n13881), .Z(n13883) );
  XNOR U13723 ( .A(n13884), .B(n13885), .Z(n13881) );
  AND U13724 ( .A(n320), .B(n13880), .Z(n13885) );
  XNOR U13725 ( .A(n13884), .B(n13878), .Z(n13880) );
  XOR U13726 ( .A(n13886), .B(n13887), .Z(n13878) );
  AND U13727 ( .A(n335), .B(n13888), .Z(n13887) );
  XNOR U13728 ( .A(n13889), .B(n13890), .Z(n13884) );
  AND U13729 ( .A(n327), .B(n13891), .Z(n13890) );
  XOR U13730 ( .A(p_input[781]), .B(n13889), .Z(n13891) );
  XNOR U13731 ( .A(n13892), .B(n13893), .Z(n13889) );
  AND U13732 ( .A(n331), .B(n13888), .Z(n13893) );
  XNOR U13733 ( .A(n13892), .B(n13886), .Z(n13888) );
  XOR U13734 ( .A(n13894), .B(n13895), .Z(n13886) );
  AND U13735 ( .A(n346), .B(n13896), .Z(n13895) );
  XNOR U13736 ( .A(n13897), .B(n13898), .Z(n13892) );
  AND U13737 ( .A(n338), .B(n13899), .Z(n13898) );
  XOR U13738 ( .A(p_input[813]), .B(n13897), .Z(n13899) );
  XNOR U13739 ( .A(n13900), .B(n13901), .Z(n13897) );
  AND U13740 ( .A(n342), .B(n13896), .Z(n13901) );
  XNOR U13741 ( .A(n13900), .B(n13894), .Z(n13896) );
  XOR U13742 ( .A(n13902), .B(n13903), .Z(n13894) );
  AND U13743 ( .A(n357), .B(n13904), .Z(n13903) );
  XNOR U13744 ( .A(n13905), .B(n13906), .Z(n13900) );
  AND U13745 ( .A(n349), .B(n13907), .Z(n13906) );
  XOR U13746 ( .A(p_input[845]), .B(n13905), .Z(n13907) );
  XNOR U13747 ( .A(n13908), .B(n13909), .Z(n13905) );
  AND U13748 ( .A(n353), .B(n13904), .Z(n13909) );
  XNOR U13749 ( .A(n13908), .B(n13902), .Z(n13904) );
  XOR U13750 ( .A(n13910), .B(n13911), .Z(n13902) );
  AND U13751 ( .A(n368), .B(n13912), .Z(n13911) );
  XNOR U13752 ( .A(n13913), .B(n13914), .Z(n13908) );
  AND U13753 ( .A(n360), .B(n13915), .Z(n13914) );
  XOR U13754 ( .A(p_input[877]), .B(n13913), .Z(n13915) );
  XNOR U13755 ( .A(n13916), .B(n13917), .Z(n13913) );
  AND U13756 ( .A(n364), .B(n13912), .Z(n13917) );
  XNOR U13757 ( .A(n13916), .B(n13910), .Z(n13912) );
  XOR U13758 ( .A(n13918), .B(n13919), .Z(n13910) );
  AND U13759 ( .A(n379), .B(n13920), .Z(n13919) );
  XNOR U13760 ( .A(n13921), .B(n13922), .Z(n13916) );
  AND U13761 ( .A(n371), .B(n13923), .Z(n13922) );
  XOR U13762 ( .A(p_input[909]), .B(n13921), .Z(n13923) );
  XNOR U13763 ( .A(n13924), .B(n13925), .Z(n13921) );
  AND U13764 ( .A(n375), .B(n13920), .Z(n13925) );
  XNOR U13765 ( .A(n13924), .B(n13918), .Z(n13920) );
  XOR U13766 ( .A(n13926), .B(n13927), .Z(n13918) );
  AND U13767 ( .A(n390), .B(n13928), .Z(n13927) );
  XNOR U13768 ( .A(n13929), .B(n13930), .Z(n13924) );
  AND U13769 ( .A(n382), .B(n13931), .Z(n13930) );
  XOR U13770 ( .A(p_input[941]), .B(n13929), .Z(n13931) );
  XNOR U13771 ( .A(n13932), .B(n13933), .Z(n13929) );
  AND U13772 ( .A(n386), .B(n13928), .Z(n13933) );
  XNOR U13773 ( .A(n13932), .B(n13926), .Z(n13928) );
  XOR U13774 ( .A(n13934), .B(n13935), .Z(n13926) );
  AND U13775 ( .A(n401), .B(n13936), .Z(n13935) );
  XNOR U13776 ( .A(n13937), .B(n13938), .Z(n13932) );
  AND U13777 ( .A(n393), .B(n13939), .Z(n13938) );
  XOR U13778 ( .A(p_input[973]), .B(n13937), .Z(n13939) );
  XNOR U13779 ( .A(n13940), .B(n13941), .Z(n13937) );
  AND U13780 ( .A(n397), .B(n13936), .Z(n13941) );
  XNOR U13781 ( .A(n13940), .B(n13934), .Z(n13936) );
  XOR U13782 ( .A(n13942), .B(n13943), .Z(n13934) );
  AND U13783 ( .A(n412), .B(n13944), .Z(n13943) );
  XNOR U13784 ( .A(n13945), .B(n13946), .Z(n13940) );
  AND U13785 ( .A(n404), .B(n13947), .Z(n13946) );
  XOR U13786 ( .A(p_input[1005]), .B(n13945), .Z(n13947) );
  XNOR U13787 ( .A(n13948), .B(n13949), .Z(n13945) );
  AND U13788 ( .A(n408), .B(n13944), .Z(n13949) );
  XNOR U13789 ( .A(n13948), .B(n13942), .Z(n13944) );
  XOR U13790 ( .A(n13950), .B(n13951), .Z(n13942) );
  AND U13791 ( .A(n423), .B(n13952), .Z(n13951) );
  XNOR U13792 ( .A(n13953), .B(n13954), .Z(n13948) );
  AND U13793 ( .A(n415), .B(n13955), .Z(n13954) );
  XOR U13794 ( .A(p_input[1037]), .B(n13953), .Z(n13955) );
  XNOR U13795 ( .A(n13956), .B(n13957), .Z(n13953) );
  AND U13796 ( .A(n419), .B(n13952), .Z(n13957) );
  XNOR U13797 ( .A(n13956), .B(n13950), .Z(n13952) );
  XOR U13798 ( .A(n13958), .B(n13959), .Z(n13950) );
  AND U13799 ( .A(n434), .B(n13960), .Z(n13959) );
  XNOR U13800 ( .A(n13961), .B(n13962), .Z(n13956) );
  AND U13801 ( .A(n426), .B(n13963), .Z(n13962) );
  XOR U13802 ( .A(p_input[1069]), .B(n13961), .Z(n13963) );
  XNOR U13803 ( .A(n13964), .B(n13965), .Z(n13961) );
  AND U13804 ( .A(n430), .B(n13960), .Z(n13965) );
  XNOR U13805 ( .A(n13964), .B(n13958), .Z(n13960) );
  XOR U13806 ( .A(n13966), .B(n13967), .Z(n13958) );
  AND U13807 ( .A(n445), .B(n13968), .Z(n13967) );
  XNOR U13808 ( .A(n13969), .B(n13970), .Z(n13964) );
  AND U13809 ( .A(n437), .B(n13971), .Z(n13970) );
  XOR U13810 ( .A(p_input[1101]), .B(n13969), .Z(n13971) );
  XNOR U13811 ( .A(n13972), .B(n13973), .Z(n13969) );
  AND U13812 ( .A(n441), .B(n13968), .Z(n13973) );
  XNOR U13813 ( .A(n13972), .B(n13966), .Z(n13968) );
  XOR U13814 ( .A(n13974), .B(n13975), .Z(n13966) );
  AND U13815 ( .A(n456), .B(n13976), .Z(n13975) );
  XNOR U13816 ( .A(n13977), .B(n13978), .Z(n13972) );
  AND U13817 ( .A(n448), .B(n13979), .Z(n13978) );
  XOR U13818 ( .A(p_input[1133]), .B(n13977), .Z(n13979) );
  XNOR U13819 ( .A(n13980), .B(n13981), .Z(n13977) );
  AND U13820 ( .A(n452), .B(n13976), .Z(n13981) );
  XNOR U13821 ( .A(n13980), .B(n13974), .Z(n13976) );
  XOR U13822 ( .A(n13982), .B(n13983), .Z(n13974) );
  AND U13823 ( .A(n467), .B(n13984), .Z(n13983) );
  XNOR U13824 ( .A(n13985), .B(n13986), .Z(n13980) );
  AND U13825 ( .A(n459), .B(n13987), .Z(n13986) );
  XOR U13826 ( .A(p_input[1165]), .B(n13985), .Z(n13987) );
  XNOR U13827 ( .A(n13988), .B(n13989), .Z(n13985) );
  AND U13828 ( .A(n463), .B(n13984), .Z(n13989) );
  XNOR U13829 ( .A(n13988), .B(n13982), .Z(n13984) );
  XOR U13830 ( .A(n13990), .B(n13991), .Z(n13982) );
  AND U13831 ( .A(n478), .B(n13992), .Z(n13991) );
  XNOR U13832 ( .A(n13993), .B(n13994), .Z(n13988) );
  AND U13833 ( .A(n470), .B(n13995), .Z(n13994) );
  XOR U13834 ( .A(p_input[1197]), .B(n13993), .Z(n13995) );
  XNOR U13835 ( .A(n13996), .B(n13997), .Z(n13993) );
  AND U13836 ( .A(n474), .B(n13992), .Z(n13997) );
  XNOR U13837 ( .A(n13996), .B(n13990), .Z(n13992) );
  XOR U13838 ( .A(n13998), .B(n13999), .Z(n13990) );
  AND U13839 ( .A(n489), .B(n14000), .Z(n13999) );
  XNOR U13840 ( .A(n14001), .B(n14002), .Z(n13996) );
  AND U13841 ( .A(n481), .B(n14003), .Z(n14002) );
  XOR U13842 ( .A(p_input[1229]), .B(n14001), .Z(n14003) );
  XNOR U13843 ( .A(n14004), .B(n14005), .Z(n14001) );
  AND U13844 ( .A(n485), .B(n14000), .Z(n14005) );
  XNOR U13845 ( .A(n14004), .B(n13998), .Z(n14000) );
  XOR U13846 ( .A(n14006), .B(n14007), .Z(n13998) );
  AND U13847 ( .A(n500), .B(n14008), .Z(n14007) );
  XNOR U13848 ( .A(n14009), .B(n14010), .Z(n14004) );
  AND U13849 ( .A(n492), .B(n14011), .Z(n14010) );
  XOR U13850 ( .A(p_input[1261]), .B(n14009), .Z(n14011) );
  XNOR U13851 ( .A(n14012), .B(n14013), .Z(n14009) );
  AND U13852 ( .A(n496), .B(n14008), .Z(n14013) );
  XNOR U13853 ( .A(n14012), .B(n14006), .Z(n14008) );
  XOR U13854 ( .A(n14014), .B(n14015), .Z(n14006) );
  AND U13855 ( .A(n511), .B(n14016), .Z(n14015) );
  XNOR U13856 ( .A(n14017), .B(n14018), .Z(n14012) );
  AND U13857 ( .A(n503), .B(n14019), .Z(n14018) );
  XOR U13858 ( .A(p_input[1293]), .B(n14017), .Z(n14019) );
  XNOR U13859 ( .A(n14020), .B(n14021), .Z(n14017) );
  AND U13860 ( .A(n507), .B(n14016), .Z(n14021) );
  XNOR U13861 ( .A(n14020), .B(n14014), .Z(n14016) );
  XOR U13862 ( .A(n14022), .B(n14023), .Z(n14014) );
  AND U13863 ( .A(n522), .B(n14024), .Z(n14023) );
  XNOR U13864 ( .A(n14025), .B(n14026), .Z(n14020) );
  AND U13865 ( .A(n514), .B(n14027), .Z(n14026) );
  XOR U13866 ( .A(p_input[1325]), .B(n14025), .Z(n14027) );
  XNOR U13867 ( .A(n14028), .B(n14029), .Z(n14025) );
  AND U13868 ( .A(n518), .B(n14024), .Z(n14029) );
  XNOR U13869 ( .A(n14028), .B(n14022), .Z(n14024) );
  XOR U13870 ( .A(n14030), .B(n14031), .Z(n14022) );
  AND U13871 ( .A(n533), .B(n14032), .Z(n14031) );
  XNOR U13872 ( .A(n14033), .B(n14034), .Z(n14028) );
  AND U13873 ( .A(n525), .B(n14035), .Z(n14034) );
  XOR U13874 ( .A(p_input[1357]), .B(n14033), .Z(n14035) );
  XNOR U13875 ( .A(n14036), .B(n14037), .Z(n14033) );
  AND U13876 ( .A(n529), .B(n14032), .Z(n14037) );
  XNOR U13877 ( .A(n14036), .B(n14030), .Z(n14032) );
  XOR U13878 ( .A(n14038), .B(n14039), .Z(n14030) );
  AND U13879 ( .A(n544), .B(n14040), .Z(n14039) );
  XNOR U13880 ( .A(n14041), .B(n14042), .Z(n14036) );
  AND U13881 ( .A(n536), .B(n14043), .Z(n14042) );
  XOR U13882 ( .A(p_input[1389]), .B(n14041), .Z(n14043) );
  XNOR U13883 ( .A(n14044), .B(n14045), .Z(n14041) );
  AND U13884 ( .A(n540), .B(n14040), .Z(n14045) );
  XNOR U13885 ( .A(n14044), .B(n14038), .Z(n14040) );
  XOR U13886 ( .A(n14046), .B(n14047), .Z(n14038) );
  AND U13887 ( .A(n555), .B(n14048), .Z(n14047) );
  XNOR U13888 ( .A(n14049), .B(n14050), .Z(n14044) );
  AND U13889 ( .A(n547), .B(n14051), .Z(n14050) );
  XOR U13890 ( .A(p_input[1421]), .B(n14049), .Z(n14051) );
  XNOR U13891 ( .A(n14052), .B(n14053), .Z(n14049) );
  AND U13892 ( .A(n551), .B(n14048), .Z(n14053) );
  XNOR U13893 ( .A(n14052), .B(n14046), .Z(n14048) );
  XOR U13894 ( .A(n14054), .B(n14055), .Z(n14046) );
  AND U13895 ( .A(n566), .B(n14056), .Z(n14055) );
  XNOR U13896 ( .A(n14057), .B(n14058), .Z(n14052) );
  AND U13897 ( .A(n558), .B(n14059), .Z(n14058) );
  XOR U13898 ( .A(p_input[1453]), .B(n14057), .Z(n14059) );
  XNOR U13899 ( .A(n14060), .B(n14061), .Z(n14057) );
  AND U13900 ( .A(n562), .B(n14056), .Z(n14061) );
  XNOR U13901 ( .A(n14060), .B(n14054), .Z(n14056) );
  XOR U13902 ( .A(n14062), .B(n14063), .Z(n14054) );
  AND U13903 ( .A(n577), .B(n14064), .Z(n14063) );
  XNOR U13904 ( .A(n14065), .B(n14066), .Z(n14060) );
  AND U13905 ( .A(n569), .B(n14067), .Z(n14066) );
  XOR U13906 ( .A(p_input[1485]), .B(n14065), .Z(n14067) );
  XNOR U13907 ( .A(n14068), .B(n14069), .Z(n14065) );
  AND U13908 ( .A(n573), .B(n14064), .Z(n14069) );
  XNOR U13909 ( .A(n14068), .B(n14062), .Z(n14064) );
  XOR U13910 ( .A(n14070), .B(n14071), .Z(n14062) );
  AND U13911 ( .A(n588), .B(n14072), .Z(n14071) );
  XNOR U13912 ( .A(n14073), .B(n14074), .Z(n14068) );
  AND U13913 ( .A(n580), .B(n14075), .Z(n14074) );
  XOR U13914 ( .A(p_input[1517]), .B(n14073), .Z(n14075) );
  XNOR U13915 ( .A(n14076), .B(n14077), .Z(n14073) );
  AND U13916 ( .A(n584), .B(n14072), .Z(n14077) );
  XNOR U13917 ( .A(n14076), .B(n14070), .Z(n14072) );
  XOR U13918 ( .A(n14078), .B(n14079), .Z(n14070) );
  AND U13919 ( .A(n599), .B(n14080), .Z(n14079) );
  XNOR U13920 ( .A(n14081), .B(n14082), .Z(n14076) );
  AND U13921 ( .A(n591), .B(n14083), .Z(n14082) );
  XOR U13922 ( .A(p_input[1549]), .B(n14081), .Z(n14083) );
  XNOR U13923 ( .A(n14084), .B(n14085), .Z(n14081) );
  AND U13924 ( .A(n595), .B(n14080), .Z(n14085) );
  XNOR U13925 ( .A(n14084), .B(n14078), .Z(n14080) );
  XOR U13926 ( .A(n14086), .B(n14087), .Z(n14078) );
  AND U13927 ( .A(n610), .B(n14088), .Z(n14087) );
  XNOR U13928 ( .A(n14089), .B(n14090), .Z(n14084) );
  AND U13929 ( .A(n602), .B(n14091), .Z(n14090) );
  XOR U13930 ( .A(p_input[1581]), .B(n14089), .Z(n14091) );
  XNOR U13931 ( .A(n14092), .B(n14093), .Z(n14089) );
  AND U13932 ( .A(n606), .B(n14088), .Z(n14093) );
  XNOR U13933 ( .A(n14092), .B(n14086), .Z(n14088) );
  XOR U13934 ( .A(n14094), .B(n14095), .Z(n14086) );
  AND U13935 ( .A(n621), .B(n14096), .Z(n14095) );
  XNOR U13936 ( .A(n14097), .B(n14098), .Z(n14092) );
  AND U13937 ( .A(n613), .B(n14099), .Z(n14098) );
  XOR U13938 ( .A(p_input[1613]), .B(n14097), .Z(n14099) );
  XNOR U13939 ( .A(n14100), .B(n14101), .Z(n14097) );
  AND U13940 ( .A(n617), .B(n14096), .Z(n14101) );
  XNOR U13941 ( .A(n14100), .B(n14094), .Z(n14096) );
  XOR U13942 ( .A(n14102), .B(n14103), .Z(n14094) );
  AND U13943 ( .A(n632), .B(n14104), .Z(n14103) );
  XNOR U13944 ( .A(n14105), .B(n14106), .Z(n14100) );
  AND U13945 ( .A(n624), .B(n14107), .Z(n14106) );
  XOR U13946 ( .A(p_input[1645]), .B(n14105), .Z(n14107) );
  XNOR U13947 ( .A(n14108), .B(n14109), .Z(n14105) );
  AND U13948 ( .A(n628), .B(n14104), .Z(n14109) );
  XNOR U13949 ( .A(n14108), .B(n14102), .Z(n14104) );
  XOR U13950 ( .A(n14110), .B(n14111), .Z(n14102) );
  AND U13951 ( .A(n643), .B(n14112), .Z(n14111) );
  XNOR U13952 ( .A(n14113), .B(n14114), .Z(n14108) );
  AND U13953 ( .A(n635), .B(n14115), .Z(n14114) );
  XOR U13954 ( .A(p_input[1677]), .B(n14113), .Z(n14115) );
  XNOR U13955 ( .A(n14116), .B(n14117), .Z(n14113) );
  AND U13956 ( .A(n639), .B(n14112), .Z(n14117) );
  XNOR U13957 ( .A(n14116), .B(n14110), .Z(n14112) );
  XOR U13958 ( .A(n14118), .B(n14119), .Z(n14110) );
  AND U13959 ( .A(n654), .B(n14120), .Z(n14119) );
  XNOR U13960 ( .A(n14121), .B(n14122), .Z(n14116) );
  AND U13961 ( .A(n646), .B(n14123), .Z(n14122) );
  XOR U13962 ( .A(p_input[1709]), .B(n14121), .Z(n14123) );
  XNOR U13963 ( .A(n14124), .B(n14125), .Z(n14121) );
  AND U13964 ( .A(n650), .B(n14120), .Z(n14125) );
  XNOR U13965 ( .A(n14124), .B(n14118), .Z(n14120) );
  XOR U13966 ( .A(n14126), .B(n14127), .Z(n14118) );
  AND U13967 ( .A(n665), .B(n14128), .Z(n14127) );
  XNOR U13968 ( .A(n14129), .B(n14130), .Z(n14124) );
  AND U13969 ( .A(n657), .B(n14131), .Z(n14130) );
  XOR U13970 ( .A(p_input[1741]), .B(n14129), .Z(n14131) );
  XNOR U13971 ( .A(n14132), .B(n14133), .Z(n14129) );
  AND U13972 ( .A(n661), .B(n14128), .Z(n14133) );
  XNOR U13973 ( .A(n14132), .B(n14126), .Z(n14128) );
  XOR U13974 ( .A(n14134), .B(n14135), .Z(n14126) );
  AND U13975 ( .A(n676), .B(n14136), .Z(n14135) );
  XNOR U13976 ( .A(n14137), .B(n14138), .Z(n14132) );
  AND U13977 ( .A(n668), .B(n14139), .Z(n14138) );
  XOR U13978 ( .A(p_input[1773]), .B(n14137), .Z(n14139) );
  XNOR U13979 ( .A(n14140), .B(n14141), .Z(n14137) );
  AND U13980 ( .A(n672), .B(n14136), .Z(n14141) );
  XNOR U13981 ( .A(n14140), .B(n14134), .Z(n14136) );
  XOR U13982 ( .A(n14142), .B(n14143), .Z(n14134) );
  AND U13983 ( .A(n687), .B(n14144), .Z(n14143) );
  XNOR U13984 ( .A(n14145), .B(n14146), .Z(n14140) );
  AND U13985 ( .A(n679), .B(n14147), .Z(n14146) );
  XOR U13986 ( .A(p_input[1805]), .B(n14145), .Z(n14147) );
  XNOR U13987 ( .A(n14148), .B(n14149), .Z(n14145) );
  AND U13988 ( .A(n683), .B(n14144), .Z(n14149) );
  XNOR U13989 ( .A(n14148), .B(n14142), .Z(n14144) );
  XOR U13990 ( .A(n14150), .B(n14151), .Z(n14142) );
  AND U13991 ( .A(n698), .B(n14152), .Z(n14151) );
  XNOR U13992 ( .A(n14153), .B(n14154), .Z(n14148) );
  AND U13993 ( .A(n690), .B(n14155), .Z(n14154) );
  XOR U13994 ( .A(p_input[1837]), .B(n14153), .Z(n14155) );
  XNOR U13995 ( .A(n14156), .B(n14157), .Z(n14153) );
  AND U13996 ( .A(n694), .B(n14152), .Z(n14157) );
  XNOR U13997 ( .A(n14156), .B(n14150), .Z(n14152) );
  XOR U13998 ( .A(n14158), .B(n14159), .Z(n14150) );
  AND U13999 ( .A(n709), .B(n14160), .Z(n14159) );
  XNOR U14000 ( .A(n14161), .B(n14162), .Z(n14156) );
  AND U14001 ( .A(n701), .B(n14163), .Z(n14162) );
  XOR U14002 ( .A(p_input[1869]), .B(n14161), .Z(n14163) );
  XNOR U14003 ( .A(n14164), .B(n14165), .Z(n14161) );
  AND U14004 ( .A(n705), .B(n14160), .Z(n14165) );
  XNOR U14005 ( .A(n14164), .B(n14158), .Z(n14160) );
  XOR U14006 ( .A(n14166), .B(n14167), .Z(n14158) );
  AND U14007 ( .A(n720), .B(n14168), .Z(n14167) );
  XNOR U14008 ( .A(n14169), .B(n14170), .Z(n14164) );
  AND U14009 ( .A(n712), .B(n14171), .Z(n14170) );
  XOR U14010 ( .A(p_input[1901]), .B(n14169), .Z(n14171) );
  XNOR U14011 ( .A(n14172), .B(n14173), .Z(n14169) );
  AND U14012 ( .A(n716), .B(n14168), .Z(n14173) );
  XNOR U14013 ( .A(n14172), .B(n14166), .Z(n14168) );
  XOR U14014 ( .A(n14174), .B(n14175), .Z(n14166) );
  AND U14015 ( .A(n731), .B(n14176), .Z(n14175) );
  XNOR U14016 ( .A(n14177), .B(n14178), .Z(n14172) );
  AND U14017 ( .A(n723), .B(n14179), .Z(n14178) );
  XOR U14018 ( .A(p_input[1933]), .B(n14177), .Z(n14179) );
  XNOR U14019 ( .A(n14180), .B(n14181), .Z(n14177) );
  AND U14020 ( .A(n727), .B(n14176), .Z(n14181) );
  XNOR U14021 ( .A(n14180), .B(n14174), .Z(n14176) );
  XOR U14022 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n14182), .Z(n14174) );
  AND U14023 ( .A(n741), .B(n14183), .Z(n14182) );
  XNOR U14024 ( .A(n14184), .B(n14185), .Z(n14180) );
  AND U14025 ( .A(n734), .B(n14186), .Z(n14185) );
  XOR U14026 ( .A(p_input[1965]), .B(n14184), .Z(n14186) );
  XNOR U14027 ( .A(n14187), .B(n14188), .Z(n14184) );
  AND U14028 ( .A(n738), .B(n14183), .Z(n14188) );
  XOR U14029 ( .A(\knn_comb_/min_val_out[0][13] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n14183) );
  XOR U14030 ( .A(n51), .B(n14189), .Z(o[12]) );
  AND U14031 ( .A(n58), .B(n14190), .Z(n51) );
  XOR U14032 ( .A(n52), .B(n14189), .Z(n14190) );
  XOR U14033 ( .A(n14191), .B(n14192), .Z(n14189) );
  AND U14034 ( .A(n70), .B(n14193), .Z(n14192) );
  XOR U14035 ( .A(n14194), .B(n14195), .Z(n52) );
  AND U14036 ( .A(n62), .B(n14196), .Z(n14195) );
  XOR U14037 ( .A(p_input[12]), .B(n14194), .Z(n14196) );
  XNOR U14038 ( .A(n14197), .B(n14198), .Z(n14194) );
  AND U14039 ( .A(n66), .B(n14193), .Z(n14198) );
  XNOR U14040 ( .A(n14197), .B(n14191), .Z(n14193) );
  XOR U14041 ( .A(n14199), .B(n14200), .Z(n14191) );
  AND U14042 ( .A(n82), .B(n14201), .Z(n14200) );
  XNOR U14043 ( .A(n14202), .B(n14203), .Z(n14197) );
  AND U14044 ( .A(n74), .B(n14204), .Z(n14203) );
  XOR U14045 ( .A(p_input[44]), .B(n14202), .Z(n14204) );
  XNOR U14046 ( .A(n14205), .B(n14206), .Z(n14202) );
  AND U14047 ( .A(n78), .B(n14201), .Z(n14206) );
  XNOR U14048 ( .A(n14205), .B(n14199), .Z(n14201) );
  XOR U14049 ( .A(n14207), .B(n14208), .Z(n14199) );
  AND U14050 ( .A(n93), .B(n14209), .Z(n14208) );
  XNOR U14051 ( .A(n14210), .B(n14211), .Z(n14205) );
  AND U14052 ( .A(n85), .B(n14212), .Z(n14211) );
  XOR U14053 ( .A(p_input[76]), .B(n14210), .Z(n14212) );
  XNOR U14054 ( .A(n14213), .B(n14214), .Z(n14210) );
  AND U14055 ( .A(n89), .B(n14209), .Z(n14214) );
  XNOR U14056 ( .A(n14213), .B(n14207), .Z(n14209) );
  XOR U14057 ( .A(n14215), .B(n14216), .Z(n14207) );
  AND U14058 ( .A(n104), .B(n14217), .Z(n14216) );
  XNOR U14059 ( .A(n14218), .B(n14219), .Z(n14213) );
  AND U14060 ( .A(n96), .B(n14220), .Z(n14219) );
  XOR U14061 ( .A(p_input[108]), .B(n14218), .Z(n14220) );
  XNOR U14062 ( .A(n14221), .B(n14222), .Z(n14218) );
  AND U14063 ( .A(n100), .B(n14217), .Z(n14222) );
  XNOR U14064 ( .A(n14221), .B(n14215), .Z(n14217) );
  XOR U14065 ( .A(n14223), .B(n14224), .Z(n14215) );
  AND U14066 ( .A(n115), .B(n14225), .Z(n14224) );
  XNOR U14067 ( .A(n14226), .B(n14227), .Z(n14221) );
  AND U14068 ( .A(n107), .B(n14228), .Z(n14227) );
  XOR U14069 ( .A(p_input[140]), .B(n14226), .Z(n14228) );
  XNOR U14070 ( .A(n14229), .B(n14230), .Z(n14226) );
  AND U14071 ( .A(n111), .B(n14225), .Z(n14230) );
  XNOR U14072 ( .A(n14229), .B(n14223), .Z(n14225) );
  XOR U14073 ( .A(n14231), .B(n14232), .Z(n14223) );
  AND U14074 ( .A(n126), .B(n14233), .Z(n14232) );
  XNOR U14075 ( .A(n14234), .B(n14235), .Z(n14229) );
  AND U14076 ( .A(n118), .B(n14236), .Z(n14235) );
  XOR U14077 ( .A(p_input[172]), .B(n14234), .Z(n14236) );
  XNOR U14078 ( .A(n14237), .B(n14238), .Z(n14234) );
  AND U14079 ( .A(n122), .B(n14233), .Z(n14238) );
  XNOR U14080 ( .A(n14237), .B(n14231), .Z(n14233) );
  XOR U14081 ( .A(n14239), .B(n14240), .Z(n14231) );
  AND U14082 ( .A(n137), .B(n14241), .Z(n14240) );
  XNOR U14083 ( .A(n14242), .B(n14243), .Z(n14237) );
  AND U14084 ( .A(n129), .B(n14244), .Z(n14243) );
  XOR U14085 ( .A(p_input[204]), .B(n14242), .Z(n14244) );
  XNOR U14086 ( .A(n14245), .B(n14246), .Z(n14242) );
  AND U14087 ( .A(n133), .B(n14241), .Z(n14246) );
  XNOR U14088 ( .A(n14245), .B(n14239), .Z(n14241) );
  XOR U14089 ( .A(n14247), .B(n14248), .Z(n14239) );
  AND U14090 ( .A(n148), .B(n14249), .Z(n14248) );
  XNOR U14091 ( .A(n14250), .B(n14251), .Z(n14245) );
  AND U14092 ( .A(n140), .B(n14252), .Z(n14251) );
  XOR U14093 ( .A(p_input[236]), .B(n14250), .Z(n14252) );
  XNOR U14094 ( .A(n14253), .B(n14254), .Z(n14250) );
  AND U14095 ( .A(n144), .B(n14249), .Z(n14254) );
  XNOR U14096 ( .A(n14253), .B(n14247), .Z(n14249) );
  XOR U14097 ( .A(n14255), .B(n14256), .Z(n14247) );
  AND U14098 ( .A(n159), .B(n14257), .Z(n14256) );
  XNOR U14099 ( .A(n14258), .B(n14259), .Z(n14253) );
  AND U14100 ( .A(n151), .B(n14260), .Z(n14259) );
  XOR U14101 ( .A(p_input[268]), .B(n14258), .Z(n14260) );
  XNOR U14102 ( .A(n14261), .B(n14262), .Z(n14258) );
  AND U14103 ( .A(n155), .B(n14257), .Z(n14262) );
  XNOR U14104 ( .A(n14261), .B(n14255), .Z(n14257) );
  XOR U14105 ( .A(n14263), .B(n14264), .Z(n14255) );
  AND U14106 ( .A(n170), .B(n14265), .Z(n14264) );
  XNOR U14107 ( .A(n14266), .B(n14267), .Z(n14261) );
  AND U14108 ( .A(n162), .B(n14268), .Z(n14267) );
  XOR U14109 ( .A(p_input[300]), .B(n14266), .Z(n14268) );
  XNOR U14110 ( .A(n14269), .B(n14270), .Z(n14266) );
  AND U14111 ( .A(n166), .B(n14265), .Z(n14270) );
  XNOR U14112 ( .A(n14269), .B(n14263), .Z(n14265) );
  XOR U14113 ( .A(n14271), .B(n14272), .Z(n14263) );
  AND U14114 ( .A(n181), .B(n14273), .Z(n14272) );
  XNOR U14115 ( .A(n14274), .B(n14275), .Z(n14269) );
  AND U14116 ( .A(n173), .B(n14276), .Z(n14275) );
  XOR U14117 ( .A(p_input[332]), .B(n14274), .Z(n14276) );
  XNOR U14118 ( .A(n14277), .B(n14278), .Z(n14274) );
  AND U14119 ( .A(n177), .B(n14273), .Z(n14278) );
  XNOR U14120 ( .A(n14277), .B(n14271), .Z(n14273) );
  XOR U14121 ( .A(n14279), .B(n14280), .Z(n14271) );
  AND U14122 ( .A(n192), .B(n14281), .Z(n14280) );
  XNOR U14123 ( .A(n14282), .B(n14283), .Z(n14277) );
  AND U14124 ( .A(n184), .B(n14284), .Z(n14283) );
  XOR U14125 ( .A(p_input[364]), .B(n14282), .Z(n14284) );
  XNOR U14126 ( .A(n14285), .B(n14286), .Z(n14282) );
  AND U14127 ( .A(n188), .B(n14281), .Z(n14286) );
  XNOR U14128 ( .A(n14285), .B(n14279), .Z(n14281) );
  XOR U14129 ( .A(n14287), .B(n14288), .Z(n14279) );
  AND U14130 ( .A(n203), .B(n14289), .Z(n14288) );
  XNOR U14131 ( .A(n14290), .B(n14291), .Z(n14285) );
  AND U14132 ( .A(n195), .B(n14292), .Z(n14291) );
  XOR U14133 ( .A(p_input[396]), .B(n14290), .Z(n14292) );
  XNOR U14134 ( .A(n14293), .B(n14294), .Z(n14290) );
  AND U14135 ( .A(n199), .B(n14289), .Z(n14294) );
  XNOR U14136 ( .A(n14293), .B(n14287), .Z(n14289) );
  XOR U14137 ( .A(n14295), .B(n14296), .Z(n14287) );
  AND U14138 ( .A(n214), .B(n14297), .Z(n14296) );
  XNOR U14139 ( .A(n14298), .B(n14299), .Z(n14293) );
  AND U14140 ( .A(n206), .B(n14300), .Z(n14299) );
  XOR U14141 ( .A(p_input[428]), .B(n14298), .Z(n14300) );
  XNOR U14142 ( .A(n14301), .B(n14302), .Z(n14298) );
  AND U14143 ( .A(n210), .B(n14297), .Z(n14302) );
  XNOR U14144 ( .A(n14301), .B(n14295), .Z(n14297) );
  XOR U14145 ( .A(n14303), .B(n14304), .Z(n14295) );
  AND U14146 ( .A(n225), .B(n14305), .Z(n14304) );
  XNOR U14147 ( .A(n14306), .B(n14307), .Z(n14301) );
  AND U14148 ( .A(n217), .B(n14308), .Z(n14307) );
  XOR U14149 ( .A(p_input[460]), .B(n14306), .Z(n14308) );
  XNOR U14150 ( .A(n14309), .B(n14310), .Z(n14306) );
  AND U14151 ( .A(n221), .B(n14305), .Z(n14310) );
  XNOR U14152 ( .A(n14309), .B(n14303), .Z(n14305) );
  XOR U14153 ( .A(n14311), .B(n14312), .Z(n14303) );
  AND U14154 ( .A(n236), .B(n14313), .Z(n14312) );
  XNOR U14155 ( .A(n14314), .B(n14315), .Z(n14309) );
  AND U14156 ( .A(n228), .B(n14316), .Z(n14315) );
  XOR U14157 ( .A(p_input[492]), .B(n14314), .Z(n14316) );
  XNOR U14158 ( .A(n14317), .B(n14318), .Z(n14314) );
  AND U14159 ( .A(n232), .B(n14313), .Z(n14318) );
  XNOR U14160 ( .A(n14317), .B(n14311), .Z(n14313) );
  XOR U14161 ( .A(n14319), .B(n14320), .Z(n14311) );
  AND U14162 ( .A(n247), .B(n14321), .Z(n14320) );
  XNOR U14163 ( .A(n14322), .B(n14323), .Z(n14317) );
  AND U14164 ( .A(n239), .B(n14324), .Z(n14323) );
  XOR U14165 ( .A(p_input[524]), .B(n14322), .Z(n14324) );
  XNOR U14166 ( .A(n14325), .B(n14326), .Z(n14322) );
  AND U14167 ( .A(n243), .B(n14321), .Z(n14326) );
  XNOR U14168 ( .A(n14325), .B(n14319), .Z(n14321) );
  XOR U14169 ( .A(n14327), .B(n14328), .Z(n14319) );
  AND U14170 ( .A(n258), .B(n14329), .Z(n14328) );
  XNOR U14171 ( .A(n14330), .B(n14331), .Z(n14325) );
  AND U14172 ( .A(n250), .B(n14332), .Z(n14331) );
  XOR U14173 ( .A(p_input[556]), .B(n14330), .Z(n14332) );
  XNOR U14174 ( .A(n14333), .B(n14334), .Z(n14330) );
  AND U14175 ( .A(n254), .B(n14329), .Z(n14334) );
  XNOR U14176 ( .A(n14333), .B(n14327), .Z(n14329) );
  XOR U14177 ( .A(n14335), .B(n14336), .Z(n14327) );
  AND U14178 ( .A(n269), .B(n14337), .Z(n14336) );
  XNOR U14179 ( .A(n14338), .B(n14339), .Z(n14333) );
  AND U14180 ( .A(n261), .B(n14340), .Z(n14339) );
  XOR U14181 ( .A(p_input[588]), .B(n14338), .Z(n14340) );
  XNOR U14182 ( .A(n14341), .B(n14342), .Z(n14338) );
  AND U14183 ( .A(n265), .B(n14337), .Z(n14342) );
  XNOR U14184 ( .A(n14341), .B(n14335), .Z(n14337) );
  XOR U14185 ( .A(n14343), .B(n14344), .Z(n14335) );
  AND U14186 ( .A(n280), .B(n14345), .Z(n14344) );
  XNOR U14187 ( .A(n14346), .B(n14347), .Z(n14341) );
  AND U14188 ( .A(n272), .B(n14348), .Z(n14347) );
  XOR U14189 ( .A(p_input[620]), .B(n14346), .Z(n14348) );
  XNOR U14190 ( .A(n14349), .B(n14350), .Z(n14346) );
  AND U14191 ( .A(n276), .B(n14345), .Z(n14350) );
  XNOR U14192 ( .A(n14349), .B(n14343), .Z(n14345) );
  XOR U14193 ( .A(n14351), .B(n14352), .Z(n14343) );
  AND U14194 ( .A(n291), .B(n14353), .Z(n14352) );
  XNOR U14195 ( .A(n14354), .B(n14355), .Z(n14349) );
  AND U14196 ( .A(n283), .B(n14356), .Z(n14355) );
  XOR U14197 ( .A(p_input[652]), .B(n14354), .Z(n14356) );
  XNOR U14198 ( .A(n14357), .B(n14358), .Z(n14354) );
  AND U14199 ( .A(n287), .B(n14353), .Z(n14358) );
  XNOR U14200 ( .A(n14357), .B(n14351), .Z(n14353) );
  XOR U14201 ( .A(n14359), .B(n14360), .Z(n14351) );
  AND U14202 ( .A(n302), .B(n14361), .Z(n14360) );
  XNOR U14203 ( .A(n14362), .B(n14363), .Z(n14357) );
  AND U14204 ( .A(n294), .B(n14364), .Z(n14363) );
  XOR U14205 ( .A(p_input[684]), .B(n14362), .Z(n14364) );
  XNOR U14206 ( .A(n14365), .B(n14366), .Z(n14362) );
  AND U14207 ( .A(n298), .B(n14361), .Z(n14366) );
  XNOR U14208 ( .A(n14365), .B(n14359), .Z(n14361) );
  XOR U14209 ( .A(n14367), .B(n14368), .Z(n14359) );
  AND U14210 ( .A(n313), .B(n14369), .Z(n14368) );
  XNOR U14211 ( .A(n14370), .B(n14371), .Z(n14365) );
  AND U14212 ( .A(n305), .B(n14372), .Z(n14371) );
  XOR U14213 ( .A(p_input[716]), .B(n14370), .Z(n14372) );
  XNOR U14214 ( .A(n14373), .B(n14374), .Z(n14370) );
  AND U14215 ( .A(n309), .B(n14369), .Z(n14374) );
  XNOR U14216 ( .A(n14373), .B(n14367), .Z(n14369) );
  XOR U14217 ( .A(n14375), .B(n14376), .Z(n14367) );
  AND U14218 ( .A(n324), .B(n14377), .Z(n14376) );
  XNOR U14219 ( .A(n14378), .B(n14379), .Z(n14373) );
  AND U14220 ( .A(n316), .B(n14380), .Z(n14379) );
  XOR U14221 ( .A(p_input[748]), .B(n14378), .Z(n14380) );
  XNOR U14222 ( .A(n14381), .B(n14382), .Z(n14378) );
  AND U14223 ( .A(n320), .B(n14377), .Z(n14382) );
  XNOR U14224 ( .A(n14381), .B(n14375), .Z(n14377) );
  XOR U14225 ( .A(n14383), .B(n14384), .Z(n14375) );
  AND U14226 ( .A(n335), .B(n14385), .Z(n14384) );
  XNOR U14227 ( .A(n14386), .B(n14387), .Z(n14381) );
  AND U14228 ( .A(n327), .B(n14388), .Z(n14387) );
  XOR U14229 ( .A(p_input[780]), .B(n14386), .Z(n14388) );
  XNOR U14230 ( .A(n14389), .B(n14390), .Z(n14386) );
  AND U14231 ( .A(n331), .B(n14385), .Z(n14390) );
  XNOR U14232 ( .A(n14389), .B(n14383), .Z(n14385) );
  XOR U14233 ( .A(n14391), .B(n14392), .Z(n14383) );
  AND U14234 ( .A(n346), .B(n14393), .Z(n14392) );
  XNOR U14235 ( .A(n14394), .B(n14395), .Z(n14389) );
  AND U14236 ( .A(n338), .B(n14396), .Z(n14395) );
  XOR U14237 ( .A(p_input[812]), .B(n14394), .Z(n14396) );
  XNOR U14238 ( .A(n14397), .B(n14398), .Z(n14394) );
  AND U14239 ( .A(n342), .B(n14393), .Z(n14398) );
  XNOR U14240 ( .A(n14397), .B(n14391), .Z(n14393) );
  XOR U14241 ( .A(n14399), .B(n14400), .Z(n14391) );
  AND U14242 ( .A(n357), .B(n14401), .Z(n14400) );
  XNOR U14243 ( .A(n14402), .B(n14403), .Z(n14397) );
  AND U14244 ( .A(n349), .B(n14404), .Z(n14403) );
  XOR U14245 ( .A(p_input[844]), .B(n14402), .Z(n14404) );
  XNOR U14246 ( .A(n14405), .B(n14406), .Z(n14402) );
  AND U14247 ( .A(n353), .B(n14401), .Z(n14406) );
  XNOR U14248 ( .A(n14405), .B(n14399), .Z(n14401) );
  XOR U14249 ( .A(n14407), .B(n14408), .Z(n14399) );
  AND U14250 ( .A(n368), .B(n14409), .Z(n14408) );
  XNOR U14251 ( .A(n14410), .B(n14411), .Z(n14405) );
  AND U14252 ( .A(n360), .B(n14412), .Z(n14411) );
  XOR U14253 ( .A(p_input[876]), .B(n14410), .Z(n14412) );
  XNOR U14254 ( .A(n14413), .B(n14414), .Z(n14410) );
  AND U14255 ( .A(n364), .B(n14409), .Z(n14414) );
  XNOR U14256 ( .A(n14413), .B(n14407), .Z(n14409) );
  XOR U14257 ( .A(n14415), .B(n14416), .Z(n14407) );
  AND U14258 ( .A(n379), .B(n14417), .Z(n14416) );
  XNOR U14259 ( .A(n14418), .B(n14419), .Z(n14413) );
  AND U14260 ( .A(n371), .B(n14420), .Z(n14419) );
  XOR U14261 ( .A(p_input[908]), .B(n14418), .Z(n14420) );
  XNOR U14262 ( .A(n14421), .B(n14422), .Z(n14418) );
  AND U14263 ( .A(n375), .B(n14417), .Z(n14422) );
  XNOR U14264 ( .A(n14421), .B(n14415), .Z(n14417) );
  XOR U14265 ( .A(n14423), .B(n14424), .Z(n14415) );
  AND U14266 ( .A(n390), .B(n14425), .Z(n14424) );
  XNOR U14267 ( .A(n14426), .B(n14427), .Z(n14421) );
  AND U14268 ( .A(n382), .B(n14428), .Z(n14427) );
  XOR U14269 ( .A(p_input[940]), .B(n14426), .Z(n14428) );
  XNOR U14270 ( .A(n14429), .B(n14430), .Z(n14426) );
  AND U14271 ( .A(n386), .B(n14425), .Z(n14430) );
  XNOR U14272 ( .A(n14429), .B(n14423), .Z(n14425) );
  XOR U14273 ( .A(n14431), .B(n14432), .Z(n14423) );
  AND U14274 ( .A(n401), .B(n14433), .Z(n14432) );
  XNOR U14275 ( .A(n14434), .B(n14435), .Z(n14429) );
  AND U14276 ( .A(n393), .B(n14436), .Z(n14435) );
  XOR U14277 ( .A(p_input[972]), .B(n14434), .Z(n14436) );
  XNOR U14278 ( .A(n14437), .B(n14438), .Z(n14434) );
  AND U14279 ( .A(n397), .B(n14433), .Z(n14438) );
  XNOR U14280 ( .A(n14437), .B(n14431), .Z(n14433) );
  XOR U14281 ( .A(n14439), .B(n14440), .Z(n14431) );
  AND U14282 ( .A(n412), .B(n14441), .Z(n14440) );
  XNOR U14283 ( .A(n14442), .B(n14443), .Z(n14437) );
  AND U14284 ( .A(n404), .B(n14444), .Z(n14443) );
  XOR U14285 ( .A(p_input[1004]), .B(n14442), .Z(n14444) );
  XNOR U14286 ( .A(n14445), .B(n14446), .Z(n14442) );
  AND U14287 ( .A(n408), .B(n14441), .Z(n14446) );
  XNOR U14288 ( .A(n14445), .B(n14439), .Z(n14441) );
  XOR U14289 ( .A(n14447), .B(n14448), .Z(n14439) );
  AND U14290 ( .A(n423), .B(n14449), .Z(n14448) );
  XNOR U14291 ( .A(n14450), .B(n14451), .Z(n14445) );
  AND U14292 ( .A(n415), .B(n14452), .Z(n14451) );
  XOR U14293 ( .A(p_input[1036]), .B(n14450), .Z(n14452) );
  XNOR U14294 ( .A(n14453), .B(n14454), .Z(n14450) );
  AND U14295 ( .A(n419), .B(n14449), .Z(n14454) );
  XNOR U14296 ( .A(n14453), .B(n14447), .Z(n14449) );
  XOR U14297 ( .A(n14455), .B(n14456), .Z(n14447) );
  AND U14298 ( .A(n434), .B(n14457), .Z(n14456) );
  XNOR U14299 ( .A(n14458), .B(n14459), .Z(n14453) );
  AND U14300 ( .A(n426), .B(n14460), .Z(n14459) );
  XOR U14301 ( .A(p_input[1068]), .B(n14458), .Z(n14460) );
  XNOR U14302 ( .A(n14461), .B(n14462), .Z(n14458) );
  AND U14303 ( .A(n430), .B(n14457), .Z(n14462) );
  XNOR U14304 ( .A(n14461), .B(n14455), .Z(n14457) );
  XOR U14305 ( .A(n14463), .B(n14464), .Z(n14455) );
  AND U14306 ( .A(n445), .B(n14465), .Z(n14464) );
  XNOR U14307 ( .A(n14466), .B(n14467), .Z(n14461) );
  AND U14308 ( .A(n437), .B(n14468), .Z(n14467) );
  XOR U14309 ( .A(p_input[1100]), .B(n14466), .Z(n14468) );
  XNOR U14310 ( .A(n14469), .B(n14470), .Z(n14466) );
  AND U14311 ( .A(n441), .B(n14465), .Z(n14470) );
  XNOR U14312 ( .A(n14469), .B(n14463), .Z(n14465) );
  XOR U14313 ( .A(n14471), .B(n14472), .Z(n14463) );
  AND U14314 ( .A(n456), .B(n14473), .Z(n14472) );
  XNOR U14315 ( .A(n14474), .B(n14475), .Z(n14469) );
  AND U14316 ( .A(n448), .B(n14476), .Z(n14475) );
  XOR U14317 ( .A(p_input[1132]), .B(n14474), .Z(n14476) );
  XNOR U14318 ( .A(n14477), .B(n14478), .Z(n14474) );
  AND U14319 ( .A(n452), .B(n14473), .Z(n14478) );
  XNOR U14320 ( .A(n14477), .B(n14471), .Z(n14473) );
  XOR U14321 ( .A(n14479), .B(n14480), .Z(n14471) );
  AND U14322 ( .A(n467), .B(n14481), .Z(n14480) );
  XNOR U14323 ( .A(n14482), .B(n14483), .Z(n14477) );
  AND U14324 ( .A(n459), .B(n14484), .Z(n14483) );
  XOR U14325 ( .A(p_input[1164]), .B(n14482), .Z(n14484) );
  XNOR U14326 ( .A(n14485), .B(n14486), .Z(n14482) );
  AND U14327 ( .A(n463), .B(n14481), .Z(n14486) );
  XNOR U14328 ( .A(n14485), .B(n14479), .Z(n14481) );
  XOR U14329 ( .A(n14487), .B(n14488), .Z(n14479) );
  AND U14330 ( .A(n478), .B(n14489), .Z(n14488) );
  XNOR U14331 ( .A(n14490), .B(n14491), .Z(n14485) );
  AND U14332 ( .A(n470), .B(n14492), .Z(n14491) );
  XOR U14333 ( .A(p_input[1196]), .B(n14490), .Z(n14492) );
  XNOR U14334 ( .A(n14493), .B(n14494), .Z(n14490) );
  AND U14335 ( .A(n474), .B(n14489), .Z(n14494) );
  XNOR U14336 ( .A(n14493), .B(n14487), .Z(n14489) );
  XOR U14337 ( .A(n14495), .B(n14496), .Z(n14487) );
  AND U14338 ( .A(n489), .B(n14497), .Z(n14496) );
  XNOR U14339 ( .A(n14498), .B(n14499), .Z(n14493) );
  AND U14340 ( .A(n481), .B(n14500), .Z(n14499) );
  XOR U14341 ( .A(p_input[1228]), .B(n14498), .Z(n14500) );
  XNOR U14342 ( .A(n14501), .B(n14502), .Z(n14498) );
  AND U14343 ( .A(n485), .B(n14497), .Z(n14502) );
  XNOR U14344 ( .A(n14501), .B(n14495), .Z(n14497) );
  XOR U14345 ( .A(n14503), .B(n14504), .Z(n14495) );
  AND U14346 ( .A(n500), .B(n14505), .Z(n14504) );
  XNOR U14347 ( .A(n14506), .B(n14507), .Z(n14501) );
  AND U14348 ( .A(n492), .B(n14508), .Z(n14507) );
  XOR U14349 ( .A(p_input[1260]), .B(n14506), .Z(n14508) );
  XNOR U14350 ( .A(n14509), .B(n14510), .Z(n14506) );
  AND U14351 ( .A(n496), .B(n14505), .Z(n14510) );
  XNOR U14352 ( .A(n14509), .B(n14503), .Z(n14505) );
  XOR U14353 ( .A(n14511), .B(n14512), .Z(n14503) );
  AND U14354 ( .A(n511), .B(n14513), .Z(n14512) );
  XNOR U14355 ( .A(n14514), .B(n14515), .Z(n14509) );
  AND U14356 ( .A(n503), .B(n14516), .Z(n14515) );
  XOR U14357 ( .A(p_input[1292]), .B(n14514), .Z(n14516) );
  XNOR U14358 ( .A(n14517), .B(n14518), .Z(n14514) );
  AND U14359 ( .A(n507), .B(n14513), .Z(n14518) );
  XNOR U14360 ( .A(n14517), .B(n14511), .Z(n14513) );
  XOR U14361 ( .A(n14519), .B(n14520), .Z(n14511) );
  AND U14362 ( .A(n522), .B(n14521), .Z(n14520) );
  XNOR U14363 ( .A(n14522), .B(n14523), .Z(n14517) );
  AND U14364 ( .A(n514), .B(n14524), .Z(n14523) );
  XOR U14365 ( .A(p_input[1324]), .B(n14522), .Z(n14524) );
  XNOR U14366 ( .A(n14525), .B(n14526), .Z(n14522) );
  AND U14367 ( .A(n518), .B(n14521), .Z(n14526) );
  XNOR U14368 ( .A(n14525), .B(n14519), .Z(n14521) );
  XOR U14369 ( .A(n14527), .B(n14528), .Z(n14519) );
  AND U14370 ( .A(n533), .B(n14529), .Z(n14528) );
  XNOR U14371 ( .A(n14530), .B(n14531), .Z(n14525) );
  AND U14372 ( .A(n525), .B(n14532), .Z(n14531) );
  XOR U14373 ( .A(p_input[1356]), .B(n14530), .Z(n14532) );
  XNOR U14374 ( .A(n14533), .B(n14534), .Z(n14530) );
  AND U14375 ( .A(n529), .B(n14529), .Z(n14534) );
  XNOR U14376 ( .A(n14533), .B(n14527), .Z(n14529) );
  XOR U14377 ( .A(n14535), .B(n14536), .Z(n14527) );
  AND U14378 ( .A(n544), .B(n14537), .Z(n14536) );
  XNOR U14379 ( .A(n14538), .B(n14539), .Z(n14533) );
  AND U14380 ( .A(n536), .B(n14540), .Z(n14539) );
  XOR U14381 ( .A(p_input[1388]), .B(n14538), .Z(n14540) );
  XNOR U14382 ( .A(n14541), .B(n14542), .Z(n14538) );
  AND U14383 ( .A(n540), .B(n14537), .Z(n14542) );
  XNOR U14384 ( .A(n14541), .B(n14535), .Z(n14537) );
  XOR U14385 ( .A(n14543), .B(n14544), .Z(n14535) );
  AND U14386 ( .A(n555), .B(n14545), .Z(n14544) );
  XNOR U14387 ( .A(n14546), .B(n14547), .Z(n14541) );
  AND U14388 ( .A(n547), .B(n14548), .Z(n14547) );
  XOR U14389 ( .A(p_input[1420]), .B(n14546), .Z(n14548) );
  XNOR U14390 ( .A(n14549), .B(n14550), .Z(n14546) );
  AND U14391 ( .A(n551), .B(n14545), .Z(n14550) );
  XNOR U14392 ( .A(n14549), .B(n14543), .Z(n14545) );
  XOR U14393 ( .A(n14551), .B(n14552), .Z(n14543) );
  AND U14394 ( .A(n566), .B(n14553), .Z(n14552) );
  XNOR U14395 ( .A(n14554), .B(n14555), .Z(n14549) );
  AND U14396 ( .A(n558), .B(n14556), .Z(n14555) );
  XOR U14397 ( .A(p_input[1452]), .B(n14554), .Z(n14556) );
  XNOR U14398 ( .A(n14557), .B(n14558), .Z(n14554) );
  AND U14399 ( .A(n562), .B(n14553), .Z(n14558) );
  XNOR U14400 ( .A(n14557), .B(n14551), .Z(n14553) );
  XOR U14401 ( .A(n14559), .B(n14560), .Z(n14551) );
  AND U14402 ( .A(n577), .B(n14561), .Z(n14560) );
  XNOR U14403 ( .A(n14562), .B(n14563), .Z(n14557) );
  AND U14404 ( .A(n569), .B(n14564), .Z(n14563) );
  XOR U14405 ( .A(p_input[1484]), .B(n14562), .Z(n14564) );
  XNOR U14406 ( .A(n14565), .B(n14566), .Z(n14562) );
  AND U14407 ( .A(n573), .B(n14561), .Z(n14566) );
  XNOR U14408 ( .A(n14565), .B(n14559), .Z(n14561) );
  XOR U14409 ( .A(n14567), .B(n14568), .Z(n14559) );
  AND U14410 ( .A(n588), .B(n14569), .Z(n14568) );
  XNOR U14411 ( .A(n14570), .B(n14571), .Z(n14565) );
  AND U14412 ( .A(n580), .B(n14572), .Z(n14571) );
  XOR U14413 ( .A(p_input[1516]), .B(n14570), .Z(n14572) );
  XNOR U14414 ( .A(n14573), .B(n14574), .Z(n14570) );
  AND U14415 ( .A(n584), .B(n14569), .Z(n14574) );
  XNOR U14416 ( .A(n14573), .B(n14567), .Z(n14569) );
  XOR U14417 ( .A(n14575), .B(n14576), .Z(n14567) );
  AND U14418 ( .A(n599), .B(n14577), .Z(n14576) );
  XNOR U14419 ( .A(n14578), .B(n14579), .Z(n14573) );
  AND U14420 ( .A(n591), .B(n14580), .Z(n14579) );
  XOR U14421 ( .A(p_input[1548]), .B(n14578), .Z(n14580) );
  XNOR U14422 ( .A(n14581), .B(n14582), .Z(n14578) );
  AND U14423 ( .A(n595), .B(n14577), .Z(n14582) );
  XNOR U14424 ( .A(n14581), .B(n14575), .Z(n14577) );
  XOR U14425 ( .A(n14583), .B(n14584), .Z(n14575) );
  AND U14426 ( .A(n610), .B(n14585), .Z(n14584) );
  XNOR U14427 ( .A(n14586), .B(n14587), .Z(n14581) );
  AND U14428 ( .A(n602), .B(n14588), .Z(n14587) );
  XOR U14429 ( .A(p_input[1580]), .B(n14586), .Z(n14588) );
  XNOR U14430 ( .A(n14589), .B(n14590), .Z(n14586) );
  AND U14431 ( .A(n606), .B(n14585), .Z(n14590) );
  XNOR U14432 ( .A(n14589), .B(n14583), .Z(n14585) );
  XOR U14433 ( .A(n14591), .B(n14592), .Z(n14583) );
  AND U14434 ( .A(n621), .B(n14593), .Z(n14592) );
  XNOR U14435 ( .A(n14594), .B(n14595), .Z(n14589) );
  AND U14436 ( .A(n613), .B(n14596), .Z(n14595) );
  XOR U14437 ( .A(p_input[1612]), .B(n14594), .Z(n14596) );
  XNOR U14438 ( .A(n14597), .B(n14598), .Z(n14594) );
  AND U14439 ( .A(n617), .B(n14593), .Z(n14598) );
  XNOR U14440 ( .A(n14597), .B(n14591), .Z(n14593) );
  XOR U14441 ( .A(n14599), .B(n14600), .Z(n14591) );
  AND U14442 ( .A(n632), .B(n14601), .Z(n14600) );
  XNOR U14443 ( .A(n14602), .B(n14603), .Z(n14597) );
  AND U14444 ( .A(n624), .B(n14604), .Z(n14603) );
  XOR U14445 ( .A(p_input[1644]), .B(n14602), .Z(n14604) );
  XNOR U14446 ( .A(n14605), .B(n14606), .Z(n14602) );
  AND U14447 ( .A(n628), .B(n14601), .Z(n14606) );
  XNOR U14448 ( .A(n14605), .B(n14599), .Z(n14601) );
  XOR U14449 ( .A(n14607), .B(n14608), .Z(n14599) );
  AND U14450 ( .A(n643), .B(n14609), .Z(n14608) );
  XNOR U14451 ( .A(n14610), .B(n14611), .Z(n14605) );
  AND U14452 ( .A(n635), .B(n14612), .Z(n14611) );
  XOR U14453 ( .A(p_input[1676]), .B(n14610), .Z(n14612) );
  XNOR U14454 ( .A(n14613), .B(n14614), .Z(n14610) );
  AND U14455 ( .A(n639), .B(n14609), .Z(n14614) );
  XNOR U14456 ( .A(n14613), .B(n14607), .Z(n14609) );
  XOR U14457 ( .A(n14615), .B(n14616), .Z(n14607) );
  AND U14458 ( .A(n654), .B(n14617), .Z(n14616) );
  XNOR U14459 ( .A(n14618), .B(n14619), .Z(n14613) );
  AND U14460 ( .A(n646), .B(n14620), .Z(n14619) );
  XOR U14461 ( .A(p_input[1708]), .B(n14618), .Z(n14620) );
  XNOR U14462 ( .A(n14621), .B(n14622), .Z(n14618) );
  AND U14463 ( .A(n650), .B(n14617), .Z(n14622) );
  XNOR U14464 ( .A(n14621), .B(n14615), .Z(n14617) );
  XOR U14465 ( .A(n14623), .B(n14624), .Z(n14615) );
  AND U14466 ( .A(n665), .B(n14625), .Z(n14624) );
  XNOR U14467 ( .A(n14626), .B(n14627), .Z(n14621) );
  AND U14468 ( .A(n657), .B(n14628), .Z(n14627) );
  XOR U14469 ( .A(p_input[1740]), .B(n14626), .Z(n14628) );
  XNOR U14470 ( .A(n14629), .B(n14630), .Z(n14626) );
  AND U14471 ( .A(n661), .B(n14625), .Z(n14630) );
  XNOR U14472 ( .A(n14629), .B(n14623), .Z(n14625) );
  XOR U14473 ( .A(n14631), .B(n14632), .Z(n14623) );
  AND U14474 ( .A(n676), .B(n14633), .Z(n14632) );
  XNOR U14475 ( .A(n14634), .B(n14635), .Z(n14629) );
  AND U14476 ( .A(n668), .B(n14636), .Z(n14635) );
  XOR U14477 ( .A(p_input[1772]), .B(n14634), .Z(n14636) );
  XNOR U14478 ( .A(n14637), .B(n14638), .Z(n14634) );
  AND U14479 ( .A(n672), .B(n14633), .Z(n14638) );
  XNOR U14480 ( .A(n14637), .B(n14631), .Z(n14633) );
  XOR U14481 ( .A(n14639), .B(n14640), .Z(n14631) );
  AND U14482 ( .A(n687), .B(n14641), .Z(n14640) );
  XNOR U14483 ( .A(n14642), .B(n14643), .Z(n14637) );
  AND U14484 ( .A(n679), .B(n14644), .Z(n14643) );
  XOR U14485 ( .A(p_input[1804]), .B(n14642), .Z(n14644) );
  XNOR U14486 ( .A(n14645), .B(n14646), .Z(n14642) );
  AND U14487 ( .A(n683), .B(n14641), .Z(n14646) );
  XNOR U14488 ( .A(n14645), .B(n14639), .Z(n14641) );
  XOR U14489 ( .A(n14647), .B(n14648), .Z(n14639) );
  AND U14490 ( .A(n698), .B(n14649), .Z(n14648) );
  XNOR U14491 ( .A(n14650), .B(n14651), .Z(n14645) );
  AND U14492 ( .A(n690), .B(n14652), .Z(n14651) );
  XOR U14493 ( .A(p_input[1836]), .B(n14650), .Z(n14652) );
  XNOR U14494 ( .A(n14653), .B(n14654), .Z(n14650) );
  AND U14495 ( .A(n694), .B(n14649), .Z(n14654) );
  XNOR U14496 ( .A(n14653), .B(n14647), .Z(n14649) );
  XOR U14497 ( .A(n14655), .B(n14656), .Z(n14647) );
  AND U14498 ( .A(n709), .B(n14657), .Z(n14656) );
  XNOR U14499 ( .A(n14658), .B(n14659), .Z(n14653) );
  AND U14500 ( .A(n701), .B(n14660), .Z(n14659) );
  XOR U14501 ( .A(p_input[1868]), .B(n14658), .Z(n14660) );
  XNOR U14502 ( .A(n14661), .B(n14662), .Z(n14658) );
  AND U14503 ( .A(n705), .B(n14657), .Z(n14662) );
  XNOR U14504 ( .A(n14661), .B(n14655), .Z(n14657) );
  XOR U14505 ( .A(n14663), .B(n14664), .Z(n14655) );
  AND U14506 ( .A(n720), .B(n14665), .Z(n14664) );
  XNOR U14507 ( .A(n14666), .B(n14667), .Z(n14661) );
  AND U14508 ( .A(n712), .B(n14668), .Z(n14667) );
  XOR U14509 ( .A(p_input[1900]), .B(n14666), .Z(n14668) );
  XNOR U14510 ( .A(n14669), .B(n14670), .Z(n14666) );
  AND U14511 ( .A(n716), .B(n14665), .Z(n14670) );
  XNOR U14512 ( .A(n14669), .B(n14663), .Z(n14665) );
  XOR U14513 ( .A(n14671), .B(n14672), .Z(n14663) );
  AND U14514 ( .A(n731), .B(n14673), .Z(n14672) );
  XNOR U14515 ( .A(n14674), .B(n14675), .Z(n14669) );
  AND U14516 ( .A(n723), .B(n14676), .Z(n14675) );
  XOR U14517 ( .A(p_input[1932]), .B(n14674), .Z(n14676) );
  XNOR U14518 ( .A(n14677), .B(n14678), .Z(n14674) );
  AND U14519 ( .A(n727), .B(n14673), .Z(n14678) );
  XNOR U14520 ( .A(n14677), .B(n14671), .Z(n14673) );
  XOR U14521 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n14679), .Z(n14671) );
  AND U14522 ( .A(n741), .B(n14680), .Z(n14679) );
  XNOR U14523 ( .A(n14681), .B(n14682), .Z(n14677) );
  AND U14524 ( .A(n734), .B(n14683), .Z(n14682) );
  XOR U14525 ( .A(p_input[1964]), .B(n14681), .Z(n14683) );
  XNOR U14526 ( .A(n14684), .B(n14685), .Z(n14681) );
  AND U14527 ( .A(n738), .B(n14680), .Z(n14685) );
  XOR U14528 ( .A(n14686), .B(n14684), .Z(n14680) );
  IV U14529 ( .A(\knn_comb_/min_val_out[0][12] ), .Z(n14686) );
  IV U14530 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n14684)
         );
  XOR U14531 ( .A(n53), .B(n14687), .Z(o[11]) );
  AND U14532 ( .A(n58), .B(n14688), .Z(n53) );
  XOR U14533 ( .A(n54), .B(n14687), .Z(n14688) );
  XOR U14534 ( .A(n14689), .B(n14690), .Z(n14687) );
  AND U14535 ( .A(n70), .B(n14691), .Z(n14690) );
  XOR U14536 ( .A(n14692), .B(n14693), .Z(n54) );
  AND U14537 ( .A(n62), .B(n14694), .Z(n14693) );
  XOR U14538 ( .A(p_input[11]), .B(n14692), .Z(n14694) );
  XNOR U14539 ( .A(n14695), .B(n14696), .Z(n14692) );
  AND U14540 ( .A(n66), .B(n14691), .Z(n14696) );
  XNOR U14541 ( .A(n14695), .B(n14689), .Z(n14691) );
  XOR U14542 ( .A(n14697), .B(n14698), .Z(n14689) );
  AND U14543 ( .A(n82), .B(n14699), .Z(n14698) );
  XNOR U14544 ( .A(n14700), .B(n14701), .Z(n14695) );
  AND U14545 ( .A(n74), .B(n14702), .Z(n14701) );
  XOR U14546 ( .A(p_input[43]), .B(n14700), .Z(n14702) );
  XNOR U14547 ( .A(n14703), .B(n14704), .Z(n14700) );
  AND U14548 ( .A(n78), .B(n14699), .Z(n14704) );
  XNOR U14549 ( .A(n14703), .B(n14697), .Z(n14699) );
  XOR U14550 ( .A(n14705), .B(n14706), .Z(n14697) );
  AND U14551 ( .A(n93), .B(n14707), .Z(n14706) );
  XNOR U14552 ( .A(n14708), .B(n14709), .Z(n14703) );
  AND U14553 ( .A(n85), .B(n14710), .Z(n14709) );
  XOR U14554 ( .A(p_input[75]), .B(n14708), .Z(n14710) );
  XNOR U14555 ( .A(n14711), .B(n14712), .Z(n14708) );
  AND U14556 ( .A(n89), .B(n14707), .Z(n14712) );
  XNOR U14557 ( .A(n14711), .B(n14705), .Z(n14707) );
  XOR U14558 ( .A(n14713), .B(n14714), .Z(n14705) );
  AND U14559 ( .A(n104), .B(n14715), .Z(n14714) );
  XNOR U14560 ( .A(n14716), .B(n14717), .Z(n14711) );
  AND U14561 ( .A(n96), .B(n14718), .Z(n14717) );
  XOR U14562 ( .A(p_input[107]), .B(n14716), .Z(n14718) );
  XNOR U14563 ( .A(n14719), .B(n14720), .Z(n14716) );
  AND U14564 ( .A(n100), .B(n14715), .Z(n14720) );
  XNOR U14565 ( .A(n14719), .B(n14713), .Z(n14715) );
  XOR U14566 ( .A(n14721), .B(n14722), .Z(n14713) );
  AND U14567 ( .A(n115), .B(n14723), .Z(n14722) );
  XNOR U14568 ( .A(n14724), .B(n14725), .Z(n14719) );
  AND U14569 ( .A(n107), .B(n14726), .Z(n14725) );
  XOR U14570 ( .A(p_input[139]), .B(n14724), .Z(n14726) );
  XNOR U14571 ( .A(n14727), .B(n14728), .Z(n14724) );
  AND U14572 ( .A(n111), .B(n14723), .Z(n14728) );
  XNOR U14573 ( .A(n14727), .B(n14721), .Z(n14723) );
  XOR U14574 ( .A(n14729), .B(n14730), .Z(n14721) );
  AND U14575 ( .A(n126), .B(n14731), .Z(n14730) );
  XNOR U14576 ( .A(n14732), .B(n14733), .Z(n14727) );
  AND U14577 ( .A(n118), .B(n14734), .Z(n14733) );
  XOR U14578 ( .A(p_input[171]), .B(n14732), .Z(n14734) );
  XNOR U14579 ( .A(n14735), .B(n14736), .Z(n14732) );
  AND U14580 ( .A(n122), .B(n14731), .Z(n14736) );
  XNOR U14581 ( .A(n14735), .B(n14729), .Z(n14731) );
  XOR U14582 ( .A(n14737), .B(n14738), .Z(n14729) );
  AND U14583 ( .A(n137), .B(n14739), .Z(n14738) );
  XNOR U14584 ( .A(n14740), .B(n14741), .Z(n14735) );
  AND U14585 ( .A(n129), .B(n14742), .Z(n14741) );
  XOR U14586 ( .A(p_input[203]), .B(n14740), .Z(n14742) );
  XNOR U14587 ( .A(n14743), .B(n14744), .Z(n14740) );
  AND U14588 ( .A(n133), .B(n14739), .Z(n14744) );
  XNOR U14589 ( .A(n14743), .B(n14737), .Z(n14739) );
  XOR U14590 ( .A(n14745), .B(n14746), .Z(n14737) );
  AND U14591 ( .A(n148), .B(n14747), .Z(n14746) );
  XNOR U14592 ( .A(n14748), .B(n14749), .Z(n14743) );
  AND U14593 ( .A(n140), .B(n14750), .Z(n14749) );
  XOR U14594 ( .A(p_input[235]), .B(n14748), .Z(n14750) );
  XNOR U14595 ( .A(n14751), .B(n14752), .Z(n14748) );
  AND U14596 ( .A(n144), .B(n14747), .Z(n14752) );
  XNOR U14597 ( .A(n14751), .B(n14745), .Z(n14747) );
  XOR U14598 ( .A(n14753), .B(n14754), .Z(n14745) );
  AND U14599 ( .A(n159), .B(n14755), .Z(n14754) );
  XNOR U14600 ( .A(n14756), .B(n14757), .Z(n14751) );
  AND U14601 ( .A(n151), .B(n14758), .Z(n14757) );
  XOR U14602 ( .A(p_input[267]), .B(n14756), .Z(n14758) );
  XNOR U14603 ( .A(n14759), .B(n14760), .Z(n14756) );
  AND U14604 ( .A(n155), .B(n14755), .Z(n14760) );
  XNOR U14605 ( .A(n14759), .B(n14753), .Z(n14755) );
  XOR U14606 ( .A(n14761), .B(n14762), .Z(n14753) );
  AND U14607 ( .A(n170), .B(n14763), .Z(n14762) );
  XNOR U14608 ( .A(n14764), .B(n14765), .Z(n14759) );
  AND U14609 ( .A(n162), .B(n14766), .Z(n14765) );
  XOR U14610 ( .A(p_input[299]), .B(n14764), .Z(n14766) );
  XNOR U14611 ( .A(n14767), .B(n14768), .Z(n14764) );
  AND U14612 ( .A(n166), .B(n14763), .Z(n14768) );
  XNOR U14613 ( .A(n14767), .B(n14761), .Z(n14763) );
  XOR U14614 ( .A(n14769), .B(n14770), .Z(n14761) );
  AND U14615 ( .A(n181), .B(n14771), .Z(n14770) );
  XNOR U14616 ( .A(n14772), .B(n14773), .Z(n14767) );
  AND U14617 ( .A(n173), .B(n14774), .Z(n14773) );
  XOR U14618 ( .A(p_input[331]), .B(n14772), .Z(n14774) );
  XNOR U14619 ( .A(n14775), .B(n14776), .Z(n14772) );
  AND U14620 ( .A(n177), .B(n14771), .Z(n14776) );
  XNOR U14621 ( .A(n14775), .B(n14769), .Z(n14771) );
  XOR U14622 ( .A(n14777), .B(n14778), .Z(n14769) );
  AND U14623 ( .A(n192), .B(n14779), .Z(n14778) );
  XNOR U14624 ( .A(n14780), .B(n14781), .Z(n14775) );
  AND U14625 ( .A(n184), .B(n14782), .Z(n14781) );
  XOR U14626 ( .A(p_input[363]), .B(n14780), .Z(n14782) );
  XNOR U14627 ( .A(n14783), .B(n14784), .Z(n14780) );
  AND U14628 ( .A(n188), .B(n14779), .Z(n14784) );
  XNOR U14629 ( .A(n14783), .B(n14777), .Z(n14779) );
  XOR U14630 ( .A(n14785), .B(n14786), .Z(n14777) );
  AND U14631 ( .A(n203), .B(n14787), .Z(n14786) );
  XNOR U14632 ( .A(n14788), .B(n14789), .Z(n14783) );
  AND U14633 ( .A(n195), .B(n14790), .Z(n14789) );
  XOR U14634 ( .A(p_input[395]), .B(n14788), .Z(n14790) );
  XNOR U14635 ( .A(n14791), .B(n14792), .Z(n14788) );
  AND U14636 ( .A(n199), .B(n14787), .Z(n14792) );
  XNOR U14637 ( .A(n14791), .B(n14785), .Z(n14787) );
  XOR U14638 ( .A(n14793), .B(n14794), .Z(n14785) );
  AND U14639 ( .A(n214), .B(n14795), .Z(n14794) );
  XNOR U14640 ( .A(n14796), .B(n14797), .Z(n14791) );
  AND U14641 ( .A(n206), .B(n14798), .Z(n14797) );
  XOR U14642 ( .A(p_input[427]), .B(n14796), .Z(n14798) );
  XNOR U14643 ( .A(n14799), .B(n14800), .Z(n14796) );
  AND U14644 ( .A(n210), .B(n14795), .Z(n14800) );
  XNOR U14645 ( .A(n14799), .B(n14793), .Z(n14795) );
  XOR U14646 ( .A(n14801), .B(n14802), .Z(n14793) );
  AND U14647 ( .A(n225), .B(n14803), .Z(n14802) );
  XNOR U14648 ( .A(n14804), .B(n14805), .Z(n14799) );
  AND U14649 ( .A(n217), .B(n14806), .Z(n14805) );
  XOR U14650 ( .A(p_input[459]), .B(n14804), .Z(n14806) );
  XNOR U14651 ( .A(n14807), .B(n14808), .Z(n14804) );
  AND U14652 ( .A(n221), .B(n14803), .Z(n14808) );
  XNOR U14653 ( .A(n14807), .B(n14801), .Z(n14803) );
  XOR U14654 ( .A(n14809), .B(n14810), .Z(n14801) );
  AND U14655 ( .A(n236), .B(n14811), .Z(n14810) );
  XNOR U14656 ( .A(n14812), .B(n14813), .Z(n14807) );
  AND U14657 ( .A(n228), .B(n14814), .Z(n14813) );
  XOR U14658 ( .A(p_input[491]), .B(n14812), .Z(n14814) );
  XNOR U14659 ( .A(n14815), .B(n14816), .Z(n14812) );
  AND U14660 ( .A(n232), .B(n14811), .Z(n14816) );
  XNOR U14661 ( .A(n14815), .B(n14809), .Z(n14811) );
  XOR U14662 ( .A(n14817), .B(n14818), .Z(n14809) );
  AND U14663 ( .A(n247), .B(n14819), .Z(n14818) );
  XNOR U14664 ( .A(n14820), .B(n14821), .Z(n14815) );
  AND U14665 ( .A(n239), .B(n14822), .Z(n14821) );
  XOR U14666 ( .A(p_input[523]), .B(n14820), .Z(n14822) );
  XNOR U14667 ( .A(n14823), .B(n14824), .Z(n14820) );
  AND U14668 ( .A(n243), .B(n14819), .Z(n14824) );
  XNOR U14669 ( .A(n14823), .B(n14817), .Z(n14819) );
  XOR U14670 ( .A(n14825), .B(n14826), .Z(n14817) );
  AND U14671 ( .A(n258), .B(n14827), .Z(n14826) );
  XNOR U14672 ( .A(n14828), .B(n14829), .Z(n14823) );
  AND U14673 ( .A(n250), .B(n14830), .Z(n14829) );
  XOR U14674 ( .A(p_input[555]), .B(n14828), .Z(n14830) );
  XNOR U14675 ( .A(n14831), .B(n14832), .Z(n14828) );
  AND U14676 ( .A(n254), .B(n14827), .Z(n14832) );
  XNOR U14677 ( .A(n14831), .B(n14825), .Z(n14827) );
  XOR U14678 ( .A(n14833), .B(n14834), .Z(n14825) );
  AND U14679 ( .A(n269), .B(n14835), .Z(n14834) );
  XNOR U14680 ( .A(n14836), .B(n14837), .Z(n14831) );
  AND U14681 ( .A(n261), .B(n14838), .Z(n14837) );
  XOR U14682 ( .A(p_input[587]), .B(n14836), .Z(n14838) );
  XNOR U14683 ( .A(n14839), .B(n14840), .Z(n14836) );
  AND U14684 ( .A(n265), .B(n14835), .Z(n14840) );
  XNOR U14685 ( .A(n14839), .B(n14833), .Z(n14835) );
  XOR U14686 ( .A(n14841), .B(n14842), .Z(n14833) );
  AND U14687 ( .A(n280), .B(n14843), .Z(n14842) );
  XNOR U14688 ( .A(n14844), .B(n14845), .Z(n14839) );
  AND U14689 ( .A(n272), .B(n14846), .Z(n14845) );
  XOR U14690 ( .A(p_input[619]), .B(n14844), .Z(n14846) );
  XNOR U14691 ( .A(n14847), .B(n14848), .Z(n14844) );
  AND U14692 ( .A(n276), .B(n14843), .Z(n14848) );
  XNOR U14693 ( .A(n14847), .B(n14841), .Z(n14843) );
  XOR U14694 ( .A(n14849), .B(n14850), .Z(n14841) );
  AND U14695 ( .A(n291), .B(n14851), .Z(n14850) );
  XNOR U14696 ( .A(n14852), .B(n14853), .Z(n14847) );
  AND U14697 ( .A(n283), .B(n14854), .Z(n14853) );
  XOR U14698 ( .A(p_input[651]), .B(n14852), .Z(n14854) );
  XNOR U14699 ( .A(n14855), .B(n14856), .Z(n14852) );
  AND U14700 ( .A(n287), .B(n14851), .Z(n14856) );
  XNOR U14701 ( .A(n14855), .B(n14849), .Z(n14851) );
  XOR U14702 ( .A(n14857), .B(n14858), .Z(n14849) );
  AND U14703 ( .A(n302), .B(n14859), .Z(n14858) );
  XNOR U14704 ( .A(n14860), .B(n14861), .Z(n14855) );
  AND U14705 ( .A(n294), .B(n14862), .Z(n14861) );
  XOR U14706 ( .A(p_input[683]), .B(n14860), .Z(n14862) );
  XNOR U14707 ( .A(n14863), .B(n14864), .Z(n14860) );
  AND U14708 ( .A(n298), .B(n14859), .Z(n14864) );
  XNOR U14709 ( .A(n14863), .B(n14857), .Z(n14859) );
  XOR U14710 ( .A(n14865), .B(n14866), .Z(n14857) );
  AND U14711 ( .A(n313), .B(n14867), .Z(n14866) );
  XNOR U14712 ( .A(n14868), .B(n14869), .Z(n14863) );
  AND U14713 ( .A(n305), .B(n14870), .Z(n14869) );
  XOR U14714 ( .A(p_input[715]), .B(n14868), .Z(n14870) );
  XNOR U14715 ( .A(n14871), .B(n14872), .Z(n14868) );
  AND U14716 ( .A(n309), .B(n14867), .Z(n14872) );
  XNOR U14717 ( .A(n14871), .B(n14865), .Z(n14867) );
  XOR U14718 ( .A(n14873), .B(n14874), .Z(n14865) );
  AND U14719 ( .A(n324), .B(n14875), .Z(n14874) );
  XNOR U14720 ( .A(n14876), .B(n14877), .Z(n14871) );
  AND U14721 ( .A(n316), .B(n14878), .Z(n14877) );
  XOR U14722 ( .A(p_input[747]), .B(n14876), .Z(n14878) );
  XNOR U14723 ( .A(n14879), .B(n14880), .Z(n14876) );
  AND U14724 ( .A(n320), .B(n14875), .Z(n14880) );
  XNOR U14725 ( .A(n14879), .B(n14873), .Z(n14875) );
  XOR U14726 ( .A(n14881), .B(n14882), .Z(n14873) );
  AND U14727 ( .A(n335), .B(n14883), .Z(n14882) );
  XNOR U14728 ( .A(n14884), .B(n14885), .Z(n14879) );
  AND U14729 ( .A(n327), .B(n14886), .Z(n14885) );
  XOR U14730 ( .A(p_input[779]), .B(n14884), .Z(n14886) );
  XNOR U14731 ( .A(n14887), .B(n14888), .Z(n14884) );
  AND U14732 ( .A(n331), .B(n14883), .Z(n14888) );
  XNOR U14733 ( .A(n14887), .B(n14881), .Z(n14883) );
  XOR U14734 ( .A(n14889), .B(n14890), .Z(n14881) );
  AND U14735 ( .A(n346), .B(n14891), .Z(n14890) );
  XNOR U14736 ( .A(n14892), .B(n14893), .Z(n14887) );
  AND U14737 ( .A(n338), .B(n14894), .Z(n14893) );
  XOR U14738 ( .A(p_input[811]), .B(n14892), .Z(n14894) );
  XNOR U14739 ( .A(n14895), .B(n14896), .Z(n14892) );
  AND U14740 ( .A(n342), .B(n14891), .Z(n14896) );
  XNOR U14741 ( .A(n14895), .B(n14889), .Z(n14891) );
  XOR U14742 ( .A(n14897), .B(n14898), .Z(n14889) );
  AND U14743 ( .A(n357), .B(n14899), .Z(n14898) );
  XNOR U14744 ( .A(n14900), .B(n14901), .Z(n14895) );
  AND U14745 ( .A(n349), .B(n14902), .Z(n14901) );
  XOR U14746 ( .A(p_input[843]), .B(n14900), .Z(n14902) );
  XNOR U14747 ( .A(n14903), .B(n14904), .Z(n14900) );
  AND U14748 ( .A(n353), .B(n14899), .Z(n14904) );
  XNOR U14749 ( .A(n14903), .B(n14897), .Z(n14899) );
  XOR U14750 ( .A(n14905), .B(n14906), .Z(n14897) );
  AND U14751 ( .A(n368), .B(n14907), .Z(n14906) );
  XNOR U14752 ( .A(n14908), .B(n14909), .Z(n14903) );
  AND U14753 ( .A(n360), .B(n14910), .Z(n14909) );
  XOR U14754 ( .A(p_input[875]), .B(n14908), .Z(n14910) );
  XNOR U14755 ( .A(n14911), .B(n14912), .Z(n14908) );
  AND U14756 ( .A(n364), .B(n14907), .Z(n14912) );
  XNOR U14757 ( .A(n14911), .B(n14905), .Z(n14907) );
  XOR U14758 ( .A(n14913), .B(n14914), .Z(n14905) );
  AND U14759 ( .A(n379), .B(n14915), .Z(n14914) );
  XNOR U14760 ( .A(n14916), .B(n14917), .Z(n14911) );
  AND U14761 ( .A(n371), .B(n14918), .Z(n14917) );
  XOR U14762 ( .A(p_input[907]), .B(n14916), .Z(n14918) );
  XNOR U14763 ( .A(n14919), .B(n14920), .Z(n14916) );
  AND U14764 ( .A(n375), .B(n14915), .Z(n14920) );
  XNOR U14765 ( .A(n14919), .B(n14913), .Z(n14915) );
  XOR U14766 ( .A(n14921), .B(n14922), .Z(n14913) );
  AND U14767 ( .A(n390), .B(n14923), .Z(n14922) );
  XNOR U14768 ( .A(n14924), .B(n14925), .Z(n14919) );
  AND U14769 ( .A(n382), .B(n14926), .Z(n14925) );
  XOR U14770 ( .A(p_input[939]), .B(n14924), .Z(n14926) );
  XNOR U14771 ( .A(n14927), .B(n14928), .Z(n14924) );
  AND U14772 ( .A(n386), .B(n14923), .Z(n14928) );
  XNOR U14773 ( .A(n14927), .B(n14921), .Z(n14923) );
  XOR U14774 ( .A(n14929), .B(n14930), .Z(n14921) );
  AND U14775 ( .A(n401), .B(n14931), .Z(n14930) );
  XNOR U14776 ( .A(n14932), .B(n14933), .Z(n14927) );
  AND U14777 ( .A(n393), .B(n14934), .Z(n14933) );
  XOR U14778 ( .A(p_input[971]), .B(n14932), .Z(n14934) );
  XNOR U14779 ( .A(n14935), .B(n14936), .Z(n14932) );
  AND U14780 ( .A(n397), .B(n14931), .Z(n14936) );
  XNOR U14781 ( .A(n14935), .B(n14929), .Z(n14931) );
  XOR U14782 ( .A(n14937), .B(n14938), .Z(n14929) );
  AND U14783 ( .A(n412), .B(n14939), .Z(n14938) );
  XNOR U14784 ( .A(n14940), .B(n14941), .Z(n14935) );
  AND U14785 ( .A(n404), .B(n14942), .Z(n14941) );
  XOR U14786 ( .A(p_input[1003]), .B(n14940), .Z(n14942) );
  XNOR U14787 ( .A(n14943), .B(n14944), .Z(n14940) );
  AND U14788 ( .A(n408), .B(n14939), .Z(n14944) );
  XNOR U14789 ( .A(n14943), .B(n14937), .Z(n14939) );
  XOR U14790 ( .A(n14945), .B(n14946), .Z(n14937) );
  AND U14791 ( .A(n423), .B(n14947), .Z(n14946) );
  XNOR U14792 ( .A(n14948), .B(n14949), .Z(n14943) );
  AND U14793 ( .A(n415), .B(n14950), .Z(n14949) );
  XOR U14794 ( .A(p_input[1035]), .B(n14948), .Z(n14950) );
  XNOR U14795 ( .A(n14951), .B(n14952), .Z(n14948) );
  AND U14796 ( .A(n419), .B(n14947), .Z(n14952) );
  XNOR U14797 ( .A(n14951), .B(n14945), .Z(n14947) );
  XOR U14798 ( .A(n14953), .B(n14954), .Z(n14945) );
  AND U14799 ( .A(n434), .B(n14955), .Z(n14954) );
  XNOR U14800 ( .A(n14956), .B(n14957), .Z(n14951) );
  AND U14801 ( .A(n426), .B(n14958), .Z(n14957) );
  XOR U14802 ( .A(p_input[1067]), .B(n14956), .Z(n14958) );
  XNOR U14803 ( .A(n14959), .B(n14960), .Z(n14956) );
  AND U14804 ( .A(n430), .B(n14955), .Z(n14960) );
  XNOR U14805 ( .A(n14959), .B(n14953), .Z(n14955) );
  XOR U14806 ( .A(n14961), .B(n14962), .Z(n14953) );
  AND U14807 ( .A(n445), .B(n14963), .Z(n14962) );
  XNOR U14808 ( .A(n14964), .B(n14965), .Z(n14959) );
  AND U14809 ( .A(n437), .B(n14966), .Z(n14965) );
  XOR U14810 ( .A(p_input[1099]), .B(n14964), .Z(n14966) );
  XNOR U14811 ( .A(n14967), .B(n14968), .Z(n14964) );
  AND U14812 ( .A(n441), .B(n14963), .Z(n14968) );
  XNOR U14813 ( .A(n14967), .B(n14961), .Z(n14963) );
  XOR U14814 ( .A(n14969), .B(n14970), .Z(n14961) );
  AND U14815 ( .A(n456), .B(n14971), .Z(n14970) );
  XNOR U14816 ( .A(n14972), .B(n14973), .Z(n14967) );
  AND U14817 ( .A(n448), .B(n14974), .Z(n14973) );
  XOR U14818 ( .A(p_input[1131]), .B(n14972), .Z(n14974) );
  XNOR U14819 ( .A(n14975), .B(n14976), .Z(n14972) );
  AND U14820 ( .A(n452), .B(n14971), .Z(n14976) );
  XNOR U14821 ( .A(n14975), .B(n14969), .Z(n14971) );
  XOR U14822 ( .A(n14977), .B(n14978), .Z(n14969) );
  AND U14823 ( .A(n467), .B(n14979), .Z(n14978) );
  XNOR U14824 ( .A(n14980), .B(n14981), .Z(n14975) );
  AND U14825 ( .A(n459), .B(n14982), .Z(n14981) );
  XOR U14826 ( .A(p_input[1163]), .B(n14980), .Z(n14982) );
  XNOR U14827 ( .A(n14983), .B(n14984), .Z(n14980) );
  AND U14828 ( .A(n463), .B(n14979), .Z(n14984) );
  XNOR U14829 ( .A(n14983), .B(n14977), .Z(n14979) );
  XOR U14830 ( .A(n14985), .B(n14986), .Z(n14977) );
  AND U14831 ( .A(n478), .B(n14987), .Z(n14986) );
  XNOR U14832 ( .A(n14988), .B(n14989), .Z(n14983) );
  AND U14833 ( .A(n470), .B(n14990), .Z(n14989) );
  XOR U14834 ( .A(p_input[1195]), .B(n14988), .Z(n14990) );
  XNOR U14835 ( .A(n14991), .B(n14992), .Z(n14988) );
  AND U14836 ( .A(n474), .B(n14987), .Z(n14992) );
  XNOR U14837 ( .A(n14991), .B(n14985), .Z(n14987) );
  XOR U14838 ( .A(n14993), .B(n14994), .Z(n14985) );
  AND U14839 ( .A(n489), .B(n14995), .Z(n14994) );
  XNOR U14840 ( .A(n14996), .B(n14997), .Z(n14991) );
  AND U14841 ( .A(n481), .B(n14998), .Z(n14997) );
  XOR U14842 ( .A(p_input[1227]), .B(n14996), .Z(n14998) );
  XNOR U14843 ( .A(n14999), .B(n15000), .Z(n14996) );
  AND U14844 ( .A(n485), .B(n14995), .Z(n15000) );
  XNOR U14845 ( .A(n14999), .B(n14993), .Z(n14995) );
  XOR U14846 ( .A(n15001), .B(n15002), .Z(n14993) );
  AND U14847 ( .A(n500), .B(n15003), .Z(n15002) );
  XNOR U14848 ( .A(n15004), .B(n15005), .Z(n14999) );
  AND U14849 ( .A(n492), .B(n15006), .Z(n15005) );
  XOR U14850 ( .A(p_input[1259]), .B(n15004), .Z(n15006) );
  XNOR U14851 ( .A(n15007), .B(n15008), .Z(n15004) );
  AND U14852 ( .A(n496), .B(n15003), .Z(n15008) );
  XNOR U14853 ( .A(n15007), .B(n15001), .Z(n15003) );
  XOR U14854 ( .A(n15009), .B(n15010), .Z(n15001) );
  AND U14855 ( .A(n511), .B(n15011), .Z(n15010) );
  XNOR U14856 ( .A(n15012), .B(n15013), .Z(n15007) );
  AND U14857 ( .A(n503), .B(n15014), .Z(n15013) );
  XOR U14858 ( .A(p_input[1291]), .B(n15012), .Z(n15014) );
  XNOR U14859 ( .A(n15015), .B(n15016), .Z(n15012) );
  AND U14860 ( .A(n507), .B(n15011), .Z(n15016) );
  XNOR U14861 ( .A(n15015), .B(n15009), .Z(n15011) );
  XOR U14862 ( .A(n15017), .B(n15018), .Z(n15009) );
  AND U14863 ( .A(n522), .B(n15019), .Z(n15018) );
  XNOR U14864 ( .A(n15020), .B(n15021), .Z(n15015) );
  AND U14865 ( .A(n514), .B(n15022), .Z(n15021) );
  XOR U14866 ( .A(p_input[1323]), .B(n15020), .Z(n15022) );
  XNOR U14867 ( .A(n15023), .B(n15024), .Z(n15020) );
  AND U14868 ( .A(n518), .B(n15019), .Z(n15024) );
  XNOR U14869 ( .A(n15023), .B(n15017), .Z(n15019) );
  XOR U14870 ( .A(n15025), .B(n15026), .Z(n15017) );
  AND U14871 ( .A(n533), .B(n15027), .Z(n15026) );
  XNOR U14872 ( .A(n15028), .B(n15029), .Z(n15023) );
  AND U14873 ( .A(n525), .B(n15030), .Z(n15029) );
  XOR U14874 ( .A(p_input[1355]), .B(n15028), .Z(n15030) );
  XNOR U14875 ( .A(n15031), .B(n15032), .Z(n15028) );
  AND U14876 ( .A(n529), .B(n15027), .Z(n15032) );
  XNOR U14877 ( .A(n15031), .B(n15025), .Z(n15027) );
  XOR U14878 ( .A(n15033), .B(n15034), .Z(n15025) );
  AND U14879 ( .A(n544), .B(n15035), .Z(n15034) );
  XNOR U14880 ( .A(n15036), .B(n15037), .Z(n15031) );
  AND U14881 ( .A(n536), .B(n15038), .Z(n15037) );
  XOR U14882 ( .A(p_input[1387]), .B(n15036), .Z(n15038) );
  XNOR U14883 ( .A(n15039), .B(n15040), .Z(n15036) );
  AND U14884 ( .A(n540), .B(n15035), .Z(n15040) );
  XNOR U14885 ( .A(n15039), .B(n15033), .Z(n15035) );
  XOR U14886 ( .A(n15041), .B(n15042), .Z(n15033) );
  AND U14887 ( .A(n555), .B(n15043), .Z(n15042) );
  XNOR U14888 ( .A(n15044), .B(n15045), .Z(n15039) );
  AND U14889 ( .A(n547), .B(n15046), .Z(n15045) );
  XOR U14890 ( .A(p_input[1419]), .B(n15044), .Z(n15046) );
  XNOR U14891 ( .A(n15047), .B(n15048), .Z(n15044) );
  AND U14892 ( .A(n551), .B(n15043), .Z(n15048) );
  XNOR U14893 ( .A(n15047), .B(n15041), .Z(n15043) );
  XOR U14894 ( .A(n15049), .B(n15050), .Z(n15041) );
  AND U14895 ( .A(n566), .B(n15051), .Z(n15050) );
  XNOR U14896 ( .A(n15052), .B(n15053), .Z(n15047) );
  AND U14897 ( .A(n558), .B(n15054), .Z(n15053) );
  XOR U14898 ( .A(p_input[1451]), .B(n15052), .Z(n15054) );
  XNOR U14899 ( .A(n15055), .B(n15056), .Z(n15052) );
  AND U14900 ( .A(n562), .B(n15051), .Z(n15056) );
  XNOR U14901 ( .A(n15055), .B(n15049), .Z(n15051) );
  XOR U14902 ( .A(n15057), .B(n15058), .Z(n15049) );
  AND U14903 ( .A(n577), .B(n15059), .Z(n15058) );
  XNOR U14904 ( .A(n15060), .B(n15061), .Z(n15055) );
  AND U14905 ( .A(n569), .B(n15062), .Z(n15061) );
  XOR U14906 ( .A(p_input[1483]), .B(n15060), .Z(n15062) );
  XNOR U14907 ( .A(n15063), .B(n15064), .Z(n15060) );
  AND U14908 ( .A(n573), .B(n15059), .Z(n15064) );
  XNOR U14909 ( .A(n15063), .B(n15057), .Z(n15059) );
  XOR U14910 ( .A(n15065), .B(n15066), .Z(n15057) );
  AND U14911 ( .A(n588), .B(n15067), .Z(n15066) );
  XNOR U14912 ( .A(n15068), .B(n15069), .Z(n15063) );
  AND U14913 ( .A(n580), .B(n15070), .Z(n15069) );
  XOR U14914 ( .A(p_input[1515]), .B(n15068), .Z(n15070) );
  XNOR U14915 ( .A(n15071), .B(n15072), .Z(n15068) );
  AND U14916 ( .A(n584), .B(n15067), .Z(n15072) );
  XNOR U14917 ( .A(n15071), .B(n15065), .Z(n15067) );
  XOR U14918 ( .A(n15073), .B(n15074), .Z(n15065) );
  AND U14919 ( .A(n599), .B(n15075), .Z(n15074) );
  XNOR U14920 ( .A(n15076), .B(n15077), .Z(n15071) );
  AND U14921 ( .A(n591), .B(n15078), .Z(n15077) );
  XOR U14922 ( .A(p_input[1547]), .B(n15076), .Z(n15078) );
  XNOR U14923 ( .A(n15079), .B(n15080), .Z(n15076) );
  AND U14924 ( .A(n595), .B(n15075), .Z(n15080) );
  XNOR U14925 ( .A(n15079), .B(n15073), .Z(n15075) );
  XOR U14926 ( .A(n15081), .B(n15082), .Z(n15073) );
  AND U14927 ( .A(n610), .B(n15083), .Z(n15082) );
  XNOR U14928 ( .A(n15084), .B(n15085), .Z(n15079) );
  AND U14929 ( .A(n602), .B(n15086), .Z(n15085) );
  XOR U14930 ( .A(p_input[1579]), .B(n15084), .Z(n15086) );
  XNOR U14931 ( .A(n15087), .B(n15088), .Z(n15084) );
  AND U14932 ( .A(n606), .B(n15083), .Z(n15088) );
  XNOR U14933 ( .A(n15087), .B(n15081), .Z(n15083) );
  XOR U14934 ( .A(n15089), .B(n15090), .Z(n15081) );
  AND U14935 ( .A(n621), .B(n15091), .Z(n15090) );
  XNOR U14936 ( .A(n15092), .B(n15093), .Z(n15087) );
  AND U14937 ( .A(n613), .B(n15094), .Z(n15093) );
  XOR U14938 ( .A(p_input[1611]), .B(n15092), .Z(n15094) );
  XNOR U14939 ( .A(n15095), .B(n15096), .Z(n15092) );
  AND U14940 ( .A(n617), .B(n15091), .Z(n15096) );
  XNOR U14941 ( .A(n15095), .B(n15089), .Z(n15091) );
  XOR U14942 ( .A(n15097), .B(n15098), .Z(n15089) );
  AND U14943 ( .A(n632), .B(n15099), .Z(n15098) );
  XNOR U14944 ( .A(n15100), .B(n15101), .Z(n15095) );
  AND U14945 ( .A(n624), .B(n15102), .Z(n15101) );
  XOR U14946 ( .A(p_input[1643]), .B(n15100), .Z(n15102) );
  XNOR U14947 ( .A(n15103), .B(n15104), .Z(n15100) );
  AND U14948 ( .A(n628), .B(n15099), .Z(n15104) );
  XNOR U14949 ( .A(n15103), .B(n15097), .Z(n15099) );
  XOR U14950 ( .A(n15105), .B(n15106), .Z(n15097) );
  AND U14951 ( .A(n643), .B(n15107), .Z(n15106) );
  XNOR U14952 ( .A(n15108), .B(n15109), .Z(n15103) );
  AND U14953 ( .A(n635), .B(n15110), .Z(n15109) );
  XOR U14954 ( .A(p_input[1675]), .B(n15108), .Z(n15110) );
  XNOR U14955 ( .A(n15111), .B(n15112), .Z(n15108) );
  AND U14956 ( .A(n639), .B(n15107), .Z(n15112) );
  XNOR U14957 ( .A(n15111), .B(n15105), .Z(n15107) );
  XOR U14958 ( .A(n15113), .B(n15114), .Z(n15105) );
  AND U14959 ( .A(n654), .B(n15115), .Z(n15114) );
  XNOR U14960 ( .A(n15116), .B(n15117), .Z(n15111) );
  AND U14961 ( .A(n646), .B(n15118), .Z(n15117) );
  XOR U14962 ( .A(p_input[1707]), .B(n15116), .Z(n15118) );
  XNOR U14963 ( .A(n15119), .B(n15120), .Z(n15116) );
  AND U14964 ( .A(n650), .B(n15115), .Z(n15120) );
  XNOR U14965 ( .A(n15119), .B(n15113), .Z(n15115) );
  XOR U14966 ( .A(n15121), .B(n15122), .Z(n15113) );
  AND U14967 ( .A(n665), .B(n15123), .Z(n15122) );
  XNOR U14968 ( .A(n15124), .B(n15125), .Z(n15119) );
  AND U14969 ( .A(n657), .B(n15126), .Z(n15125) );
  XOR U14970 ( .A(p_input[1739]), .B(n15124), .Z(n15126) );
  XNOR U14971 ( .A(n15127), .B(n15128), .Z(n15124) );
  AND U14972 ( .A(n661), .B(n15123), .Z(n15128) );
  XNOR U14973 ( .A(n15127), .B(n15121), .Z(n15123) );
  XOR U14974 ( .A(n15129), .B(n15130), .Z(n15121) );
  AND U14975 ( .A(n676), .B(n15131), .Z(n15130) );
  XNOR U14976 ( .A(n15132), .B(n15133), .Z(n15127) );
  AND U14977 ( .A(n668), .B(n15134), .Z(n15133) );
  XOR U14978 ( .A(p_input[1771]), .B(n15132), .Z(n15134) );
  XNOR U14979 ( .A(n15135), .B(n15136), .Z(n15132) );
  AND U14980 ( .A(n672), .B(n15131), .Z(n15136) );
  XNOR U14981 ( .A(n15135), .B(n15129), .Z(n15131) );
  XOR U14982 ( .A(n15137), .B(n15138), .Z(n15129) );
  AND U14983 ( .A(n687), .B(n15139), .Z(n15138) );
  XNOR U14984 ( .A(n15140), .B(n15141), .Z(n15135) );
  AND U14985 ( .A(n679), .B(n15142), .Z(n15141) );
  XOR U14986 ( .A(p_input[1803]), .B(n15140), .Z(n15142) );
  XNOR U14987 ( .A(n15143), .B(n15144), .Z(n15140) );
  AND U14988 ( .A(n683), .B(n15139), .Z(n15144) );
  XNOR U14989 ( .A(n15143), .B(n15137), .Z(n15139) );
  XOR U14990 ( .A(n15145), .B(n15146), .Z(n15137) );
  AND U14991 ( .A(n698), .B(n15147), .Z(n15146) );
  XNOR U14992 ( .A(n15148), .B(n15149), .Z(n15143) );
  AND U14993 ( .A(n690), .B(n15150), .Z(n15149) );
  XOR U14994 ( .A(p_input[1835]), .B(n15148), .Z(n15150) );
  XNOR U14995 ( .A(n15151), .B(n15152), .Z(n15148) );
  AND U14996 ( .A(n694), .B(n15147), .Z(n15152) );
  XNOR U14997 ( .A(n15151), .B(n15145), .Z(n15147) );
  XOR U14998 ( .A(n15153), .B(n15154), .Z(n15145) );
  AND U14999 ( .A(n709), .B(n15155), .Z(n15154) );
  XNOR U15000 ( .A(n15156), .B(n15157), .Z(n15151) );
  AND U15001 ( .A(n701), .B(n15158), .Z(n15157) );
  XOR U15002 ( .A(p_input[1867]), .B(n15156), .Z(n15158) );
  XNOR U15003 ( .A(n15159), .B(n15160), .Z(n15156) );
  AND U15004 ( .A(n705), .B(n15155), .Z(n15160) );
  XNOR U15005 ( .A(n15159), .B(n15153), .Z(n15155) );
  XOR U15006 ( .A(n15161), .B(n15162), .Z(n15153) );
  AND U15007 ( .A(n720), .B(n15163), .Z(n15162) );
  XNOR U15008 ( .A(n15164), .B(n15165), .Z(n15159) );
  AND U15009 ( .A(n712), .B(n15166), .Z(n15165) );
  XOR U15010 ( .A(p_input[1899]), .B(n15164), .Z(n15166) );
  XNOR U15011 ( .A(n15167), .B(n15168), .Z(n15164) );
  AND U15012 ( .A(n716), .B(n15163), .Z(n15168) );
  XNOR U15013 ( .A(n15167), .B(n15161), .Z(n15163) );
  XOR U15014 ( .A(n15169), .B(n15170), .Z(n15161) );
  AND U15015 ( .A(n731), .B(n15171), .Z(n15170) );
  XNOR U15016 ( .A(n15172), .B(n15173), .Z(n15167) );
  AND U15017 ( .A(n723), .B(n15174), .Z(n15173) );
  XOR U15018 ( .A(p_input[1931]), .B(n15172), .Z(n15174) );
  XNOR U15019 ( .A(n15175), .B(n15176), .Z(n15172) );
  AND U15020 ( .A(n727), .B(n15171), .Z(n15176) );
  XNOR U15021 ( .A(n15175), .B(n15169), .Z(n15171) );
  XOR U15022 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n15177), .Z(n15169) );
  AND U15023 ( .A(n741), .B(n15178), .Z(n15177) );
  XNOR U15024 ( .A(n15179), .B(n15180), .Z(n15175) );
  AND U15025 ( .A(n734), .B(n15181), .Z(n15180) );
  XOR U15026 ( .A(p_input[1963]), .B(n15179), .Z(n15181) );
  XNOR U15027 ( .A(n15182), .B(n15183), .Z(n15179) );
  AND U15028 ( .A(n738), .B(n15178), .Z(n15183) );
  XOR U15029 ( .A(\knn_comb_/min_val_out[0][11] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n15178) );
  XOR U15030 ( .A(n55), .B(n15184), .Z(o[10]) );
  AND U15031 ( .A(n58), .B(n15185), .Z(n55) );
  XOR U15032 ( .A(n56), .B(n15184), .Z(n15185) );
  XOR U15033 ( .A(n15186), .B(n15187), .Z(n15184) );
  AND U15034 ( .A(n70), .B(n15188), .Z(n15187) );
  XOR U15035 ( .A(n15189), .B(n15190), .Z(n56) );
  AND U15036 ( .A(n62), .B(n15191), .Z(n15190) );
  XOR U15037 ( .A(p_input[10]), .B(n15189), .Z(n15191) );
  XNOR U15038 ( .A(n15192), .B(n15193), .Z(n15189) );
  AND U15039 ( .A(n66), .B(n15188), .Z(n15193) );
  XNOR U15040 ( .A(n15192), .B(n15186), .Z(n15188) );
  XOR U15041 ( .A(n15194), .B(n15195), .Z(n15186) );
  AND U15042 ( .A(n82), .B(n15196), .Z(n15195) );
  XNOR U15043 ( .A(n15197), .B(n15198), .Z(n15192) );
  AND U15044 ( .A(n74), .B(n15199), .Z(n15198) );
  XOR U15045 ( .A(p_input[42]), .B(n15197), .Z(n15199) );
  XNOR U15046 ( .A(n15200), .B(n15201), .Z(n15197) );
  AND U15047 ( .A(n78), .B(n15196), .Z(n15201) );
  XNOR U15048 ( .A(n15200), .B(n15194), .Z(n15196) );
  XOR U15049 ( .A(n15202), .B(n15203), .Z(n15194) );
  AND U15050 ( .A(n93), .B(n15204), .Z(n15203) );
  XNOR U15051 ( .A(n15205), .B(n15206), .Z(n15200) );
  AND U15052 ( .A(n85), .B(n15207), .Z(n15206) );
  XOR U15053 ( .A(p_input[74]), .B(n15205), .Z(n15207) );
  XNOR U15054 ( .A(n15208), .B(n15209), .Z(n15205) );
  AND U15055 ( .A(n89), .B(n15204), .Z(n15209) );
  XNOR U15056 ( .A(n15208), .B(n15202), .Z(n15204) );
  XOR U15057 ( .A(n15210), .B(n15211), .Z(n15202) );
  AND U15058 ( .A(n104), .B(n15212), .Z(n15211) );
  XNOR U15059 ( .A(n15213), .B(n15214), .Z(n15208) );
  AND U15060 ( .A(n96), .B(n15215), .Z(n15214) );
  XOR U15061 ( .A(p_input[106]), .B(n15213), .Z(n15215) );
  XNOR U15062 ( .A(n15216), .B(n15217), .Z(n15213) );
  AND U15063 ( .A(n100), .B(n15212), .Z(n15217) );
  XNOR U15064 ( .A(n15216), .B(n15210), .Z(n15212) );
  XOR U15065 ( .A(n15218), .B(n15219), .Z(n15210) );
  AND U15066 ( .A(n115), .B(n15220), .Z(n15219) );
  XNOR U15067 ( .A(n15221), .B(n15222), .Z(n15216) );
  AND U15068 ( .A(n107), .B(n15223), .Z(n15222) );
  XOR U15069 ( .A(p_input[138]), .B(n15221), .Z(n15223) );
  XNOR U15070 ( .A(n15224), .B(n15225), .Z(n15221) );
  AND U15071 ( .A(n111), .B(n15220), .Z(n15225) );
  XNOR U15072 ( .A(n15224), .B(n15218), .Z(n15220) );
  XOR U15073 ( .A(n15226), .B(n15227), .Z(n15218) );
  AND U15074 ( .A(n126), .B(n15228), .Z(n15227) );
  XNOR U15075 ( .A(n15229), .B(n15230), .Z(n15224) );
  AND U15076 ( .A(n118), .B(n15231), .Z(n15230) );
  XOR U15077 ( .A(p_input[170]), .B(n15229), .Z(n15231) );
  XNOR U15078 ( .A(n15232), .B(n15233), .Z(n15229) );
  AND U15079 ( .A(n122), .B(n15228), .Z(n15233) );
  XNOR U15080 ( .A(n15232), .B(n15226), .Z(n15228) );
  XOR U15081 ( .A(n15234), .B(n15235), .Z(n15226) );
  AND U15082 ( .A(n137), .B(n15236), .Z(n15235) );
  XNOR U15083 ( .A(n15237), .B(n15238), .Z(n15232) );
  AND U15084 ( .A(n129), .B(n15239), .Z(n15238) );
  XOR U15085 ( .A(p_input[202]), .B(n15237), .Z(n15239) );
  XNOR U15086 ( .A(n15240), .B(n15241), .Z(n15237) );
  AND U15087 ( .A(n133), .B(n15236), .Z(n15241) );
  XNOR U15088 ( .A(n15240), .B(n15234), .Z(n15236) );
  XOR U15089 ( .A(n15242), .B(n15243), .Z(n15234) );
  AND U15090 ( .A(n148), .B(n15244), .Z(n15243) );
  XNOR U15091 ( .A(n15245), .B(n15246), .Z(n15240) );
  AND U15092 ( .A(n140), .B(n15247), .Z(n15246) );
  XOR U15093 ( .A(p_input[234]), .B(n15245), .Z(n15247) );
  XNOR U15094 ( .A(n15248), .B(n15249), .Z(n15245) );
  AND U15095 ( .A(n144), .B(n15244), .Z(n15249) );
  XNOR U15096 ( .A(n15248), .B(n15242), .Z(n15244) );
  XOR U15097 ( .A(n15250), .B(n15251), .Z(n15242) );
  AND U15098 ( .A(n159), .B(n15252), .Z(n15251) );
  XNOR U15099 ( .A(n15253), .B(n15254), .Z(n15248) );
  AND U15100 ( .A(n151), .B(n15255), .Z(n15254) );
  XOR U15101 ( .A(p_input[266]), .B(n15253), .Z(n15255) );
  XNOR U15102 ( .A(n15256), .B(n15257), .Z(n15253) );
  AND U15103 ( .A(n155), .B(n15252), .Z(n15257) );
  XNOR U15104 ( .A(n15256), .B(n15250), .Z(n15252) );
  XOR U15105 ( .A(n15258), .B(n15259), .Z(n15250) );
  AND U15106 ( .A(n170), .B(n15260), .Z(n15259) );
  XNOR U15107 ( .A(n15261), .B(n15262), .Z(n15256) );
  AND U15108 ( .A(n162), .B(n15263), .Z(n15262) );
  XOR U15109 ( .A(p_input[298]), .B(n15261), .Z(n15263) );
  XNOR U15110 ( .A(n15264), .B(n15265), .Z(n15261) );
  AND U15111 ( .A(n166), .B(n15260), .Z(n15265) );
  XNOR U15112 ( .A(n15264), .B(n15258), .Z(n15260) );
  XOR U15113 ( .A(n15266), .B(n15267), .Z(n15258) );
  AND U15114 ( .A(n181), .B(n15268), .Z(n15267) );
  XNOR U15115 ( .A(n15269), .B(n15270), .Z(n15264) );
  AND U15116 ( .A(n173), .B(n15271), .Z(n15270) );
  XOR U15117 ( .A(p_input[330]), .B(n15269), .Z(n15271) );
  XNOR U15118 ( .A(n15272), .B(n15273), .Z(n15269) );
  AND U15119 ( .A(n177), .B(n15268), .Z(n15273) );
  XNOR U15120 ( .A(n15272), .B(n15266), .Z(n15268) );
  XOR U15121 ( .A(n15274), .B(n15275), .Z(n15266) );
  AND U15122 ( .A(n192), .B(n15276), .Z(n15275) );
  XNOR U15123 ( .A(n15277), .B(n15278), .Z(n15272) );
  AND U15124 ( .A(n184), .B(n15279), .Z(n15278) );
  XOR U15125 ( .A(p_input[362]), .B(n15277), .Z(n15279) );
  XNOR U15126 ( .A(n15280), .B(n15281), .Z(n15277) );
  AND U15127 ( .A(n188), .B(n15276), .Z(n15281) );
  XNOR U15128 ( .A(n15280), .B(n15274), .Z(n15276) );
  XOR U15129 ( .A(n15282), .B(n15283), .Z(n15274) );
  AND U15130 ( .A(n203), .B(n15284), .Z(n15283) );
  XNOR U15131 ( .A(n15285), .B(n15286), .Z(n15280) );
  AND U15132 ( .A(n195), .B(n15287), .Z(n15286) );
  XOR U15133 ( .A(p_input[394]), .B(n15285), .Z(n15287) );
  XNOR U15134 ( .A(n15288), .B(n15289), .Z(n15285) );
  AND U15135 ( .A(n199), .B(n15284), .Z(n15289) );
  XNOR U15136 ( .A(n15288), .B(n15282), .Z(n15284) );
  XOR U15137 ( .A(n15290), .B(n15291), .Z(n15282) );
  AND U15138 ( .A(n214), .B(n15292), .Z(n15291) );
  XNOR U15139 ( .A(n15293), .B(n15294), .Z(n15288) );
  AND U15140 ( .A(n206), .B(n15295), .Z(n15294) );
  XOR U15141 ( .A(p_input[426]), .B(n15293), .Z(n15295) );
  XNOR U15142 ( .A(n15296), .B(n15297), .Z(n15293) );
  AND U15143 ( .A(n210), .B(n15292), .Z(n15297) );
  XNOR U15144 ( .A(n15296), .B(n15290), .Z(n15292) );
  XOR U15145 ( .A(n15298), .B(n15299), .Z(n15290) );
  AND U15146 ( .A(n225), .B(n15300), .Z(n15299) );
  XNOR U15147 ( .A(n15301), .B(n15302), .Z(n15296) );
  AND U15148 ( .A(n217), .B(n15303), .Z(n15302) );
  XOR U15149 ( .A(p_input[458]), .B(n15301), .Z(n15303) );
  XNOR U15150 ( .A(n15304), .B(n15305), .Z(n15301) );
  AND U15151 ( .A(n221), .B(n15300), .Z(n15305) );
  XNOR U15152 ( .A(n15304), .B(n15298), .Z(n15300) );
  XOR U15153 ( .A(n15306), .B(n15307), .Z(n15298) );
  AND U15154 ( .A(n236), .B(n15308), .Z(n15307) );
  XNOR U15155 ( .A(n15309), .B(n15310), .Z(n15304) );
  AND U15156 ( .A(n228), .B(n15311), .Z(n15310) );
  XOR U15157 ( .A(p_input[490]), .B(n15309), .Z(n15311) );
  XNOR U15158 ( .A(n15312), .B(n15313), .Z(n15309) );
  AND U15159 ( .A(n232), .B(n15308), .Z(n15313) );
  XNOR U15160 ( .A(n15312), .B(n15306), .Z(n15308) );
  XOR U15161 ( .A(n15314), .B(n15315), .Z(n15306) );
  AND U15162 ( .A(n247), .B(n15316), .Z(n15315) );
  XNOR U15163 ( .A(n15317), .B(n15318), .Z(n15312) );
  AND U15164 ( .A(n239), .B(n15319), .Z(n15318) );
  XOR U15165 ( .A(p_input[522]), .B(n15317), .Z(n15319) );
  XNOR U15166 ( .A(n15320), .B(n15321), .Z(n15317) );
  AND U15167 ( .A(n243), .B(n15316), .Z(n15321) );
  XNOR U15168 ( .A(n15320), .B(n15314), .Z(n15316) );
  XOR U15169 ( .A(n15322), .B(n15323), .Z(n15314) );
  AND U15170 ( .A(n258), .B(n15324), .Z(n15323) );
  XNOR U15171 ( .A(n15325), .B(n15326), .Z(n15320) );
  AND U15172 ( .A(n250), .B(n15327), .Z(n15326) );
  XOR U15173 ( .A(p_input[554]), .B(n15325), .Z(n15327) );
  XNOR U15174 ( .A(n15328), .B(n15329), .Z(n15325) );
  AND U15175 ( .A(n254), .B(n15324), .Z(n15329) );
  XNOR U15176 ( .A(n15328), .B(n15322), .Z(n15324) );
  XOR U15177 ( .A(n15330), .B(n15331), .Z(n15322) );
  AND U15178 ( .A(n269), .B(n15332), .Z(n15331) );
  XNOR U15179 ( .A(n15333), .B(n15334), .Z(n15328) );
  AND U15180 ( .A(n261), .B(n15335), .Z(n15334) );
  XOR U15181 ( .A(p_input[586]), .B(n15333), .Z(n15335) );
  XNOR U15182 ( .A(n15336), .B(n15337), .Z(n15333) );
  AND U15183 ( .A(n265), .B(n15332), .Z(n15337) );
  XNOR U15184 ( .A(n15336), .B(n15330), .Z(n15332) );
  XOR U15185 ( .A(n15338), .B(n15339), .Z(n15330) );
  AND U15186 ( .A(n280), .B(n15340), .Z(n15339) );
  XNOR U15187 ( .A(n15341), .B(n15342), .Z(n15336) );
  AND U15188 ( .A(n272), .B(n15343), .Z(n15342) );
  XOR U15189 ( .A(p_input[618]), .B(n15341), .Z(n15343) );
  XNOR U15190 ( .A(n15344), .B(n15345), .Z(n15341) );
  AND U15191 ( .A(n276), .B(n15340), .Z(n15345) );
  XNOR U15192 ( .A(n15344), .B(n15338), .Z(n15340) );
  XOR U15193 ( .A(n15346), .B(n15347), .Z(n15338) );
  AND U15194 ( .A(n291), .B(n15348), .Z(n15347) );
  XNOR U15195 ( .A(n15349), .B(n15350), .Z(n15344) );
  AND U15196 ( .A(n283), .B(n15351), .Z(n15350) );
  XOR U15197 ( .A(p_input[650]), .B(n15349), .Z(n15351) );
  XNOR U15198 ( .A(n15352), .B(n15353), .Z(n15349) );
  AND U15199 ( .A(n287), .B(n15348), .Z(n15353) );
  XNOR U15200 ( .A(n15352), .B(n15346), .Z(n15348) );
  XOR U15201 ( .A(n15354), .B(n15355), .Z(n15346) );
  AND U15202 ( .A(n302), .B(n15356), .Z(n15355) );
  XNOR U15203 ( .A(n15357), .B(n15358), .Z(n15352) );
  AND U15204 ( .A(n294), .B(n15359), .Z(n15358) );
  XOR U15205 ( .A(p_input[682]), .B(n15357), .Z(n15359) );
  XNOR U15206 ( .A(n15360), .B(n15361), .Z(n15357) );
  AND U15207 ( .A(n298), .B(n15356), .Z(n15361) );
  XNOR U15208 ( .A(n15360), .B(n15354), .Z(n15356) );
  XOR U15209 ( .A(n15362), .B(n15363), .Z(n15354) );
  AND U15210 ( .A(n313), .B(n15364), .Z(n15363) );
  XNOR U15211 ( .A(n15365), .B(n15366), .Z(n15360) );
  AND U15212 ( .A(n305), .B(n15367), .Z(n15366) );
  XOR U15213 ( .A(p_input[714]), .B(n15365), .Z(n15367) );
  XNOR U15214 ( .A(n15368), .B(n15369), .Z(n15365) );
  AND U15215 ( .A(n309), .B(n15364), .Z(n15369) );
  XNOR U15216 ( .A(n15368), .B(n15362), .Z(n15364) );
  XOR U15217 ( .A(n15370), .B(n15371), .Z(n15362) );
  AND U15218 ( .A(n324), .B(n15372), .Z(n15371) );
  XNOR U15219 ( .A(n15373), .B(n15374), .Z(n15368) );
  AND U15220 ( .A(n316), .B(n15375), .Z(n15374) );
  XOR U15221 ( .A(p_input[746]), .B(n15373), .Z(n15375) );
  XNOR U15222 ( .A(n15376), .B(n15377), .Z(n15373) );
  AND U15223 ( .A(n320), .B(n15372), .Z(n15377) );
  XNOR U15224 ( .A(n15376), .B(n15370), .Z(n15372) );
  XOR U15225 ( .A(n15378), .B(n15379), .Z(n15370) );
  AND U15226 ( .A(n335), .B(n15380), .Z(n15379) );
  XNOR U15227 ( .A(n15381), .B(n15382), .Z(n15376) );
  AND U15228 ( .A(n327), .B(n15383), .Z(n15382) );
  XOR U15229 ( .A(p_input[778]), .B(n15381), .Z(n15383) );
  XNOR U15230 ( .A(n15384), .B(n15385), .Z(n15381) );
  AND U15231 ( .A(n331), .B(n15380), .Z(n15385) );
  XNOR U15232 ( .A(n15384), .B(n15378), .Z(n15380) );
  XOR U15233 ( .A(n15386), .B(n15387), .Z(n15378) );
  AND U15234 ( .A(n346), .B(n15388), .Z(n15387) );
  XNOR U15235 ( .A(n15389), .B(n15390), .Z(n15384) );
  AND U15236 ( .A(n338), .B(n15391), .Z(n15390) );
  XOR U15237 ( .A(p_input[810]), .B(n15389), .Z(n15391) );
  XNOR U15238 ( .A(n15392), .B(n15393), .Z(n15389) );
  AND U15239 ( .A(n342), .B(n15388), .Z(n15393) );
  XNOR U15240 ( .A(n15392), .B(n15386), .Z(n15388) );
  XOR U15241 ( .A(n15394), .B(n15395), .Z(n15386) );
  AND U15242 ( .A(n357), .B(n15396), .Z(n15395) );
  XNOR U15243 ( .A(n15397), .B(n15398), .Z(n15392) );
  AND U15244 ( .A(n349), .B(n15399), .Z(n15398) );
  XOR U15245 ( .A(p_input[842]), .B(n15397), .Z(n15399) );
  XNOR U15246 ( .A(n15400), .B(n15401), .Z(n15397) );
  AND U15247 ( .A(n353), .B(n15396), .Z(n15401) );
  XNOR U15248 ( .A(n15400), .B(n15394), .Z(n15396) );
  XOR U15249 ( .A(n15402), .B(n15403), .Z(n15394) );
  AND U15250 ( .A(n368), .B(n15404), .Z(n15403) );
  XNOR U15251 ( .A(n15405), .B(n15406), .Z(n15400) );
  AND U15252 ( .A(n360), .B(n15407), .Z(n15406) );
  XOR U15253 ( .A(p_input[874]), .B(n15405), .Z(n15407) );
  XNOR U15254 ( .A(n15408), .B(n15409), .Z(n15405) );
  AND U15255 ( .A(n364), .B(n15404), .Z(n15409) );
  XNOR U15256 ( .A(n15408), .B(n15402), .Z(n15404) );
  XOR U15257 ( .A(n15410), .B(n15411), .Z(n15402) );
  AND U15258 ( .A(n379), .B(n15412), .Z(n15411) );
  XNOR U15259 ( .A(n15413), .B(n15414), .Z(n15408) );
  AND U15260 ( .A(n371), .B(n15415), .Z(n15414) );
  XOR U15261 ( .A(p_input[906]), .B(n15413), .Z(n15415) );
  XNOR U15262 ( .A(n15416), .B(n15417), .Z(n15413) );
  AND U15263 ( .A(n375), .B(n15412), .Z(n15417) );
  XNOR U15264 ( .A(n15416), .B(n15410), .Z(n15412) );
  XOR U15265 ( .A(n15418), .B(n15419), .Z(n15410) );
  AND U15266 ( .A(n390), .B(n15420), .Z(n15419) );
  XNOR U15267 ( .A(n15421), .B(n15422), .Z(n15416) );
  AND U15268 ( .A(n382), .B(n15423), .Z(n15422) );
  XOR U15269 ( .A(p_input[938]), .B(n15421), .Z(n15423) );
  XNOR U15270 ( .A(n15424), .B(n15425), .Z(n15421) );
  AND U15271 ( .A(n386), .B(n15420), .Z(n15425) );
  XNOR U15272 ( .A(n15424), .B(n15418), .Z(n15420) );
  XOR U15273 ( .A(n15426), .B(n15427), .Z(n15418) );
  AND U15274 ( .A(n401), .B(n15428), .Z(n15427) );
  XNOR U15275 ( .A(n15429), .B(n15430), .Z(n15424) );
  AND U15276 ( .A(n393), .B(n15431), .Z(n15430) );
  XOR U15277 ( .A(p_input[970]), .B(n15429), .Z(n15431) );
  XNOR U15278 ( .A(n15432), .B(n15433), .Z(n15429) );
  AND U15279 ( .A(n397), .B(n15428), .Z(n15433) );
  XNOR U15280 ( .A(n15432), .B(n15426), .Z(n15428) );
  XOR U15281 ( .A(n15434), .B(n15435), .Z(n15426) );
  AND U15282 ( .A(n412), .B(n15436), .Z(n15435) );
  XNOR U15283 ( .A(n15437), .B(n15438), .Z(n15432) );
  AND U15284 ( .A(n404), .B(n15439), .Z(n15438) );
  XOR U15285 ( .A(p_input[1002]), .B(n15437), .Z(n15439) );
  XNOR U15286 ( .A(n15440), .B(n15441), .Z(n15437) );
  AND U15287 ( .A(n408), .B(n15436), .Z(n15441) );
  XNOR U15288 ( .A(n15440), .B(n15434), .Z(n15436) );
  XOR U15289 ( .A(n15442), .B(n15443), .Z(n15434) );
  AND U15290 ( .A(n423), .B(n15444), .Z(n15443) );
  XNOR U15291 ( .A(n15445), .B(n15446), .Z(n15440) );
  AND U15292 ( .A(n415), .B(n15447), .Z(n15446) );
  XOR U15293 ( .A(p_input[1034]), .B(n15445), .Z(n15447) );
  XNOR U15294 ( .A(n15448), .B(n15449), .Z(n15445) );
  AND U15295 ( .A(n419), .B(n15444), .Z(n15449) );
  XNOR U15296 ( .A(n15448), .B(n15442), .Z(n15444) );
  XOR U15297 ( .A(n15450), .B(n15451), .Z(n15442) );
  AND U15298 ( .A(n434), .B(n15452), .Z(n15451) );
  XNOR U15299 ( .A(n15453), .B(n15454), .Z(n15448) );
  AND U15300 ( .A(n426), .B(n15455), .Z(n15454) );
  XOR U15301 ( .A(p_input[1066]), .B(n15453), .Z(n15455) );
  XNOR U15302 ( .A(n15456), .B(n15457), .Z(n15453) );
  AND U15303 ( .A(n430), .B(n15452), .Z(n15457) );
  XNOR U15304 ( .A(n15456), .B(n15450), .Z(n15452) );
  XOR U15305 ( .A(n15458), .B(n15459), .Z(n15450) );
  AND U15306 ( .A(n445), .B(n15460), .Z(n15459) );
  XNOR U15307 ( .A(n15461), .B(n15462), .Z(n15456) );
  AND U15308 ( .A(n437), .B(n15463), .Z(n15462) );
  XOR U15309 ( .A(p_input[1098]), .B(n15461), .Z(n15463) );
  XNOR U15310 ( .A(n15464), .B(n15465), .Z(n15461) );
  AND U15311 ( .A(n441), .B(n15460), .Z(n15465) );
  XNOR U15312 ( .A(n15464), .B(n15458), .Z(n15460) );
  XOR U15313 ( .A(n15466), .B(n15467), .Z(n15458) );
  AND U15314 ( .A(n456), .B(n15468), .Z(n15467) );
  XNOR U15315 ( .A(n15469), .B(n15470), .Z(n15464) );
  AND U15316 ( .A(n448), .B(n15471), .Z(n15470) );
  XOR U15317 ( .A(p_input[1130]), .B(n15469), .Z(n15471) );
  XNOR U15318 ( .A(n15472), .B(n15473), .Z(n15469) );
  AND U15319 ( .A(n452), .B(n15468), .Z(n15473) );
  XNOR U15320 ( .A(n15472), .B(n15466), .Z(n15468) );
  XOR U15321 ( .A(n15474), .B(n15475), .Z(n15466) );
  AND U15322 ( .A(n467), .B(n15476), .Z(n15475) );
  XNOR U15323 ( .A(n15477), .B(n15478), .Z(n15472) );
  AND U15324 ( .A(n459), .B(n15479), .Z(n15478) );
  XOR U15325 ( .A(p_input[1162]), .B(n15477), .Z(n15479) );
  XNOR U15326 ( .A(n15480), .B(n15481), .Z(n15477) );
  AND U15327 ( .A(n463), .B(n15476), .Z(n15481) );
  XNOR U15328 ( .A(n15480), .B(n15474), .Z(n15476) );
  XOR U15329 ( .A(n15482), .B(n15483), .Z(n15474) );
  AND U15330 ( .A(n478), .B(n15484), .Z(n15483) );
  XNOR U15331 ( .A(n15485), .B(n15486), .Z(n15480) );
  AND U15332 ( .A(n470), .B(n15487), .Z(n15486) );
  XOR U15333 ( .A(p_input[1194]), .B(n15485), .Z(n15487) );
  XNOR U15334 ( .A(n15488), .B(n15489), .Z(n15485) );
  AND U15335 ( .A(n474), .B(n15484), .Z(n15489) );
  XNOR U15336 ( .A(n15488), .B(n15482), .Z(n15484) );
  XOR U15337 ( .A(n15490), .B(n15491), .Z(n15482) );
  AND U15338 ( .A(n489), .B(n15492), .Z(n15491) );
  XNOR U15339 ( .A(n15493), .B(n15494), .Z(n15488) );
  AND U15340 ( .A(n481), .B(n15495), .Z(n15494) );
  XOR U15341 ( .A(p_input[1226]), .B(n15493), .Z(n15495) );
  XNOR U15342 ( .A(n15496), .B(n15497), .Z(n15493) );
  AND U15343 ( .A(n485), .B(n15492), .Z(n15497) );
  XNOR U15344 ( .A(n15496), .B(n15490), .Z(n15492) );
  XOR U15345 ( .A(n15498), .B(n15499), .Z(n15490) );
  AND U15346 ( .A(n500), .B(n15500), .Z(n15499) );
  XNOR U15347 ( .A(n15501), .B(n15502), .Z(n15496) );
  AND U15348 ( .A(n492), .B(n15503), .Z(n15502) );
  XOR U15349 ( .A(p_input[1258]), .B(n15501), .Z(n15503) );
  XNOR U15350 ( .A(n15504), .B(n15505), .Z(n15501) );
  AND U15351 ( .A(n496), .B(n15500), .Z(n15505) );
  XNOR U15352 ( .A(n15504), .B(n15498), .Z(n15500) );
  XOR U15353 ( .A(n15506), .B(n15507), .Z(n15498) );
  AND U15354 ( .A(n511), .B(n15508), .Z(n15507) );
  XNOR U15355 ( .A(n15509), .B(n15510), .Z(n15504) );
  AND U15356 ( .A(n503), .B(n15511), .Z(n15510) );
  XOR U15357 ( .A(p_input[1290]), .B(n15509), .Z(n15511) );
  XNOR U15358 ( .A(n15512), .B(n15513), .Z(n15509) );
  AND U15359 ( .A(n507), .B(n15508), .Z(n15513) );
  XNOR U15360 ( .A(n15512), .B(n15506), .Z(n15508) );
  XOR U15361 ( .A(n15514), .B(n15515), .Z(n15506) );
  AND U15362 ( .A(n522), .B(n15516), .Z(n15515) );
  XNOR U15363 ( .A(n15517), .B(n15518), .Z(n15512) );
  AND U15364 ( .A(n514), .B(n15519), .Z(n15518) );
  XOR U15365 ( .A(p_input[1322]), .B(n15517), .Z(n15519) );
  XNOR U15366 ( .A(n15520), .B(n15521), .Z(n15517) );
  AND U15367 ( .A(n518), .B(n15516), .Z(n15521) );
  XNOR U15368 ( .A(n15520), .B(n15514), .Z(n15516) );
  XOR U15369 ( .A(n15522), .B(n15523), .Z(n15514) );
  AND U15370 ( .A(n533), .B(n15524), .Z(n15523) );
  XNOR U15371 ( .A(n15525), .B(n15526), .Z(n15520) );
  AND U15372 ( .A(n525), .B(n15527), .Z(n15526) );
  XOR U15373 ( .A(p_input[1354]), .B(n15525), .Z(n15527) );
  XNOR U15374 ( .A(n15528), .B(n15529), .Z(n15525) );
  AND U15375 ( .A(n529), .B(n15524), .Z(n15529) );
  XNOR U15376 ( .A(n15528), .B(n15522), .Z(n15524) );
  XOR U15377 ( .A(n15530), .B(n15531), .Z(n15522) );
  AND U15378 ( .A(n544), .B(n15532), .Z(n15531) );
  XNOR U15379 ( .A(n15533), .B(n15534), .Z(n15528) );
  AND U15380 ( .A(n536), .B(n15535), .Z(n15534) );
  XOR U15381 ( .A(p_input[1386]), .B(n15533), .Z(n15535) );
  XNOR U15382 ( .A(n15536), .B(n15537), .Z(n15533) );
  AND U15383 ( .A(n540), .B(n15532), .Z(n15537) );
  XNOR U15384 ( .A(n15536), .B(n15530), .Z(n15532) );
  XOR U15385 ( .A(n15538), .B(n15539), .Z(n15530) );
  AND U15386 ( .A(n555), .B(n15540), .Z(n15539) );
  XNOR U15387 ( .A(n15541), .B(n15542), .Z(n15536) );
  AND U15388 ( .A(n547), .B(n15543), .Z(n15542) );
  XOR U15389 ( .A(p_input[1418]), .B(n15541), .Z(n15543) );
  XNOR U15390 ( .A(n15544), .B(n15545), .Z(n15541) );
  AND U15391 ( .A(n551), .B(n15540), .Z(n15545) );
  XNOR U15392 ( .A(n15544), .B(n15538), .Z(n15540) );
  XOR U15393 ( .A(n15546), .B(n15547), .Z(n15538) );
  AND U15394 ( .A(n566), .B(n15548), .Z(n15547) );
  XNOR U15395 ( .A(n15549), .B(n15550), .Z(n15544) );
  AND U15396 ( .A(n558), .B(n15551), .Z(n15550) );
  XOR U15397 ( .A(p_input[1450]), .B(n15549), .Z(n15551) );
  XNOR U15398 ( .A(n15552), .B(n15553), .Z(n15549) );
  AND U15399 ( .A(n562), .B(n15548), .Z(n15553) );
  XNOR U15400 ( .A(n15552), .B(n15546), .Z(n15548) );
  XOR U15401 ( .A(n15554), .B(n15555), .Z(n15546) );
  AND U15402 ( .A(n577), .B(n15556), .Z(n15555) );
  XNOR U15403 ( .A(n15557), .B(n15558), .Z(n15552) );
  AND U15404 ( .A(n569), .B(n15559), .Z(n15558) );
  XOR U15405 ( .A(p_input[1482]), .B(n15557), .Z(n15559) );
  XNOR U15406 ( .A(n15560), .B(n15561), .Z(n15557) );
  AND U15407 ( .A(n573), .B(n15556), .Z(n15561) );
  XNOR U15408 ( .A(n15560), .B(n15554), .Z(n15556) );
  XOR U15409 ( .A(n15562), .B(n15563), .Z(n15554) );
  AND U15410 ( .A(n588), .B(n15564), .Z(n15563) );
  XNOR U15411 ( .A(n15565), .B(n15566), .Z(n15560) );
  AND U15412 ( .A(n580), .B(n15567), .Z(n15566) );
  XOR U15413 ( .A(p_input[1514]), .B(n15565), .Z(n15567) );
  XNOR U15414 ( .A(n15568), .B(n15569), .Z(n15565) );
  AND U15415 ( .A(n584), .B(n15564), .Z(n15569) );
  XNOR U15416 ( .A(n15568), .B(n15562), .Z(n15564) );
  XOR U15417 ( .A(n15570), .B(n15571), .Z(n15562) );
  AND U15418 ( .A(n599), .B(n15572), .Z(n15571) );
  XNOR U15419 ( .A(n15573), .B(n15574), .Z(n15568) );
  AND U15420 ( .A(n591), .B(n15575), .Z(n15574) );
  XOR U15421 ( .A(p_input[1546]), .B(n15573), .Z(n15575) );
  XNOR U15422 ( .A(n15576), .B(n15577), .Z(n15573) );
  AND U15423 ( .A(n595), .B(n15572), .Z(n15577) );
  XNOR U15424 ( .A(n15576), .B(n15570), .Z(n15572) );
  XOR U15425 ( .A(n15578), .B(n15579), .Z(n15570) );
  AND U15426 ( .A(n610), .B(n15580), .Z(n15579) );
  XNOR U15427 ( .A(n15581), .B(n15582), .Z(n15576) );
  AND U15428 ( .A(n602), .B(n15583), .Z(n15582) );
  XOR U15429 ( .A(p_input[1578]), .B(n15581), .Z(n15583) );
  XNOR U15430 ( .A(n15584), .B(n15585), .Z(n15581) );
  AND U15431 ( .A(n606), .B(n15580), .Z(n15585) );
  XNOR U15432 ( .A(n15584), .B(n15578), .Z(n15580) );
  XOR U15433 ( .A(n15586), .B(n15587), .Z(n15578) );
  AND U15434 ( .A(n621), .B(n15588), .Z(n15587) );
  XNOR U15435 ( .A(n15589), .B(n15590), .Z(n15584) );
  AND U15436 ( .A(n613), .B(n15591), .Z(n15590) );
  XOR U15437 ( .A(p_input[1610]), .B(n15589), .Z(n15591) );
  XNOR U15438 ( .A(n15592), .B(n15593), .Z(n15589) );
  AND U15439 ( .A(n617), .B(n15588), .Z(n15593) );
  XNOR U15440 ( .A(n15592), .B(n15586), .Z(n15588) );
  XOR U15441 ( .A(n15594), .B(n15595), .Z(n15586) );
  AND U15442 ( .A(n632), .B(n15596), .Z(n15595) );
  XNOR U15443 ( .A(n15597), .B(n15598), .Z(n15592) );
  AND U15444 ( .A(n624), .B(n15599), .Z(n15598) );
  XOR U15445 ( .A(p_input[1642]), .B(n15597), .Z(n15599) );
  XNOR U15446 ( .A(n15600), .B(n15601), .Z(n15597) );
  AND U15447 ( .A(n628), .B(n15596), .Z(n15601) );
  XNOR U15448 ( .A(n15600), .B(n15594), .Z(n15596) );
  XOR U15449 ( .A(n15602), .B(n15603), .Z(n15594) );
  AND U15450 ( .A(n643), .B(n15604), .Z(n15603) );
  XNOR U15451 ( .A(n15605), .B(n15606), .Z(n15600) );
  AND U15452 ( .A(n635), .B(n15607), .Z(n15606) );
  XOR U15453 ( .A(p_input[1674]), .B(n15605), .Z(n15607) );
  XNOR U15454 ( .A(n15608), .B(n15609), .Z(n15605) );
  AND U15455 ( .A(n639), .B(n15604), .Z(n15609) );
  XNOR U15456 ( .A(n15608), .B(n15602), .Z(n15604) );
  XOR U15457 ( .A(n15610), .B(n15611), .Z(n15602) );
  AND U15458 ( .A(n654), .B(n15612), .Z(n15611) );
  XNOR U15459 ( .A(n15613), .B(n15614), .Z(n15608) );
  AND U15460 ( .A(n646), .B(n15615), .Z(n15614) );
  XOR U15461 ( .A(p_input[1706]), .B(n15613), .Z(n15615) );
  XNOR U15462 ( .A(n15616), .B(n15617), .Z(n15613) );
  AND U15463 ( .A(n650), .B(n15612), .Z(n15617) );
  XNOR U15464 ( .A(n15616), .B(n15610), .Z(n15612) );
  XOR U15465 ( .A(n15618), .B(n15619), .Z(n15610) );
  AND U15466 ( .A(n665), .B(n15620), .Z(n15619) );
  XNOR U15467 ( .A(n15621), .B(n15622), .Z(n15616) );
  AND U15468 ( .A(n657), .B(n15623), .Z(n15622) );
  XOR U15469 ( .A(p_input[1738]), .B(n15621), .Z(n15623) );
  XNOR U15470 ( .A(n15624), .B(n15625), .Z(n15621) );
  AND U15471 ( .A(n661), .B(n15620), .Z(n15625) );
  XNOR U15472 ( .A(n15624), .B(n15618), .Z(n15620) );
  XOR U15473 ( .A(n15626), .B(n15627), .Z(n15618) );
  AND U15474 ( .A(n676), .B(n15628), .Z(n15627) );
  XNOR U15475 ( .A(n15629), .B(n15630), .Z(n15624) );
  AND U15476 ( .A(n668), .B(n15631), .Z(n15630) );
  XOR U15477 ( .A(p_input[1770]), .B(n15629), .Z(n15631) );
  XNOR U15478 ( .A(n15632), .B(n15633), .Z(n15629) );
  AND U15479 ( .A(n672), .B(n15628), .Z(n15633) );
  XNOR U15480 ( .A(n15632), .B(n15626), .Z(n15628) );
  XOR U15481 ( .A(n15634), .B(n15635), .Z(n15626) );
  AND U15482 ( .A(n687), .B(n15636), .Z(n15635) );
  XNOR U15483 ( .A(n15637), .B(n15638), .Z(n15632) );
  AND U15484 ( .A(n679), .B(n15639), .Z(n15638) );
  XOR U15485 ( .A(p_input[1802]), .B(n15637), .Z(n15639) );
  XNOR U15486 ( .A(n15640), .B(n15641), .Z(n15637) );
  AND U15487 ( .A(n683), .B(n15636), .Z(n15641) );
  XNOR U15488 ( .A(n15640), .B(n15634), .Z(n15636) );
  XOR U15489 ( .A(n15642), .B(n15643), .Z(n15634) );
  AND U15490 ( .A(n698), .B(n15644), .Z(n15643) );
  XNOR U15491 ( .A(n15645), .B(n15646), .Z(n15640) );
  AND U15492 ( .A(n690), .B(n15647), .Z(n15646) );
  XOR U15493 ( .A(p_input[1834]), .B(n15645), .Z(n15647) );
  XNOR U15494 ( .A(n15648), .B(n15649), .Z(n15645) );
  AND U15495 ( .A(n694), .B(n15644), .Z(n15649) );
  XNOR U15496 ( .A(n15648), .B(n15642), .Z(n15644) );
  XOR U15497 ( .A(n15650), .B(n15651), .Z(n15642) );
  AND U15498 ( .A(n709), .B(n15652), .Z(n15651) );
  XNOR U15499 ( .A(n15653), .B(n15654), .Z(n15648) );
  AND U15500 ( .A(n701), .B(n15655), .Z(n15654) );
  XOR U15501 ( .A(p_input[1866]), .B(n15653), .Z(n15655) );
  XNOR U15502 ( .A(n15656), .B(n15657), .Z(n15653) );
  AND U15503 ( .A(n705), .B(n15652), .Z(n15657) );
  XNOR U15504 ( .A(n15656), .B(n15650), .Z(n15652) );
  XOR U15505 ( .A(n15658), .B(n15659), .Z(n15650) );
  AND U15506 ( .A(n720), .B(n15660), .Z(n15659) );
  XNOR U15507 ( .A(n15661), .B(n15662), .Z(n15656) );
  AND U15508 ( .A(n712), .B(n15663), .Z(n15662) );
  XOR U15509 ( .A(p_input[1898]), .B(n15661), .Z(n15663) );
  XNOR U15510 ( .A(n15664), .B(n15665), .Z(n15661) );
  AND U15511 ( .A(n716), .B(n15660), .Z(n15665) );
  XNOR U15512 ( .A(n15664), .B(n15658), .Z(n15660) );
  XOR U15513 ( .A(n15666), .B(n15667), .Z(n15658) );
  AND U15514 ( .A(n731), .B(n15668), .Z(n15667) );
  XNOR U15515 ( .A(n15669), .B(n15670), .Z(n15664) );
  AND U15516 ( .A(n723), .B(n15671), .Z(n15670) );
  XOR U15517 ( .A(p_input[1930]), .B(n15669), .Z(n15671) );
  XNOR U15518 ( .A(n15672), .B(n15673), .Z(n15669) );
  AND U15519 ( .A(n727), .B(n15668), .Z(n15673) );
  XNOR U15520 ( .A(n15672), .B(n15666), .Z(n15668) );
  XOR U15521 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n15674), .Z(n15666) );
  AND U15522 ( .A(n741), .B(n15675), .Z(n15674) );
  XNOR U15523 ( .A(n15676), .B(n15677), .Z(n15672) );
  AND U15524 ( .A(n734), .B(n15678), .Z(n15677) );
  XOR U15525 ( .A(p_input[1962]), .B(n15676), .Z(n15678) );
  XNOR U15526 ( .A(n15679), .B(n15680), .Z(n15676) );
  AND U15527 ( .A(n738), .B(n15675), .Z(n15680) );
  XOR U15528 ( .A(\knn_comb_/min_val_out[0][10] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n15675) );
  XOR U15529 ( .A(n3743), .B(n15681), .Z(o[0]) );
  AND U15530 ( .A(n58), .B(n15682), .Z(n3743) );
  XOR U15531 ( .A(n3744), .B(n15681), .Z(n15682) );
  XOR U15532 ( .A(n15683), .B(n15684), .Z(n15681) );
  AND U15533 ( .A(n70), .B(n15685), .Z(n15684) );
  XOR U15534 ( .A(n15686), .B(n15687), .Z(n3744) );
  AND U15535 ( .A(n62), .B(n15688), .Z(n15687) );
  XOR U15536 ( .A(p_input[0]), .B(n15686), .Z(n15688) );
  XNOR U15537 ( .A(n15689), .B(n15690), .Z(n15686) );
  AND U15538 ( .A(n66), .B(n15685), .Z(n15690) );
  XNOR U15539 ( .A(n15689), .B(n15683), .Z(n15685) );
  XOR U15540 ( .A(n15691), .B(n15692), .Z(n15683) );
  AND U15541 ( .A(n82), .B(n15693), .Z(n15692) );
  XNOR U15542 ( .A(n15694), .B(n15695), .Z(n15689) );
  AND U15543 ( .A(n74), .B(n15696), .Z(n15695) );
  XOR U15544 ( .A(p_input[32]), .B(n15694), .Z(n15696) );
  XNOR U15545 ( .A(n15697), .B(n15698), .Z(n15694) );
  AND U15546 ( .A(n78), .B(n15693), .Z(n15698) );
  XNOR U15547 ( .A(n15697), .B(n15691), .Z(n15693) );
  XOR U15548 ( .A(n15699), .B(n15700), .Z(n15691) );
  AND U15549 ( .A(n93), .B(n15701), .Z(n15700) );
  XNOR U15550 ( .A(n15702), .B(n15703), .Z(n15697) );
  AND U15551 ( .A(n85), .B(n15704), .Z(n15703) );
  XOR U15552 ( .A(p_input[64]), .B(n15702), .Z(n15704) );
  XNOR U15553 ( .A(n15705), .B(n15706), .Z(n15702) );
  AND U15554 ( .A(n89), .B(n15701), .Z(n15706) );
  XNOR U15555 ( .A(n15705), .B(n15699), .Z(n15701) );
  XOR U15556 ( .A(n15707), .B(n15708), .Z(n15699) );
  AND U15557 ( .A(n104), .B(n15709), .Z(n15708) );
  XNOR U15558 ( .A(n15710), .B(n15711), .Z(n15705) );
  AND U15559 ( .A(n96), .B(n15712), .Z(n15711) );
  XOR U15560 ( .A(p_input[96]), .B(n15710), .Z(n15712) );
  XNOR U15561 ( .A(n15713), .B(n15714), .Z(n15710) );
  AND U15562 ( .A(n100), .B(n15709), .Z(n15714) );
  XNOR U15563 ( .A(n15713), .B(n15707), .Z(n15709) );
  XOR U15564 ( .A(n15715), .B(n15716), .Z(n15707) );
  AND U15565 ( .A(n115), .B(n15717), .Z(n15716) );
  XNOR U15566 ( .A(n15718), .B(n15719), .Z(n15713) );
  AND U15567 ( .A(n107), .B(n15720), .Z(n15719) );
  XOR U15568 ( .A(p_input[128]), .B(n15718), .Z(n15720) );
  XNOR U15569 ( .A(n15721), .B(n15722), .Z(n15718) );
  AND U15570 ( .A(n111), .B(n15717), .Z(n15722) );
  XNOR U15571 ( .A(n15721), .B(n15715), .Z(n15717) );
  XOR U15572 ( .A(n15723), .B(n15724), .Z(n15715) );
  AND U15573 ( .A(n126), .B(n15725), .Z(n15724) );
  XNOR U15574 ( .A(n15726), .B(n15727), .Z(n15721) );
  AND U15575 ( .A(n118), .B(n15728), .Z(n15727) );
  XOR U15576 ( .A(p_input[160]), .B(n15726), .Z(n15728) );
  XNOR U15577 ( .A(n15729), .B(n15730), .Z(n15726) );
  AND U15578 ( .A(n122), .B(n15725), .Z(n15730) );
  XNOR U15579 ( .A(n15729), .B(n15723), .Z(n15725) );
  XOR U15580 ( .A(n15731), .B(n15732), .Z(n15723) );
  AND U15581 ( .A(n137), .B(n15733), .Z(n15732) );
  XNOR U15582 ( .A(n15734), .B(n15735), .Z(n15729) );
  AND U15583 ( .A(n129), .B(n15736), .Z(n15735) );
  XOR U15584 ( .A(p_input[192]), .B(n15734), .Z(n15736) );
  XNOR U15585 ( .A(n15737), .B(n15738), .Z(n15734) );
  AND U15586 ( .A(n133), .B(n15733), .Z(n15738) );
  XNOR U15587 ( .A(n15737), .B(n15731), .Z(n15733) );
  XOR U15588 ( .A(n15739), .B(n15740), .Z(n15731) );
  AND U15589 ( .A(n148), .B(n15741), .Z(n15740) );
  XNOR U15590 ( .A(n15742), .B(n15743), .Z(n15737) );
  AND U15591 ( .A(n140), .B(n15744), .Z(n15743) );
  XOR U15592 ( .A(p_input[224]), .B(n15742), .Z(n15744) );
  XNOR U15593 ( .A(n15745), .B(n15746), .Z(n15742) );
  AND U15594 ( .A(n144), .B(n15741), .Z(n15746) );
  XNOR U15595 ( .A(n15745), .B(n15739), .Z(n15741) );
  XOR U15596 ( .A(n15747), .B(n15748), .Z(n15739) );
  AND U15597 ( .A(n159), .B(n15749), .Z(n15748) );
  XNOR U15598 ( .A(n15750), .B(n15751), .Z(n15745) );
  AND U15599 ( .A(n151), .B(n15752), .Z(n15751) );
  XOR U15600 ( .A(p_input[256]), .B(n15750), .Z(n15752) );
  XNOR U15601 ( .A(n15753), .B(n15754), .Z(n15750) );
  AND U15602 ( .A(n155), .B(n15749), .Z(n15754) );
  XNOR U15603 ( .A(n15753), .B(n15747), .Z(n15749) );
  XOR U15604 ( .A(n15755), .B(n15756), .Z(n15747) );
  AND U15605 ( .A(n170), .B(n15757), .Z(n15756) );
  XNOR U15606 ( .A(n15758), .B(n15759), .Z(n15753) );
  AND U15607 ( .A(n162), .B(n15760), .Z(n15759) );
  XOR U15608 ( .A(p_input[288]), .B(n15758), .Z(n15760) );
  XNOR U15609 ( .A(n15761), .B(n15762), .Z(n15758) );
  AND U15610 ( .A(n166), .B(n15757), .Z(n15762) );
  XNOR U15611 ( .A(n15761), .B(n15755), .Z(n15757) );
  XOR U15612 ( .A(n15763), .B(n15764), .Z(n15755) );
  AND U15613 ( .A(n181), .B(n15765), .Z(n15764) );
  XNOR U15614 ( .A(n15766), .B(n15767), .Z(n15761) );
  AND U15615 ( .A(n173), .B(n15768), .Z(n15767) );
  XOR U15616 ( .A(p_input[320]), .B(n15766), .Z(n15768) );
  XNOR U15617 ( .A(n15769), .B(n15770), .Z(n15766) );
  AND U15618 ( .A(n177), .B(n15765), .Z(n15770) );
  XNOR U15619 ( .A(n15769), .B(n15763), .Z(n15765) );
  XOR U15620 ( .A(n15771), .B(n15772), .Z(n15763) );
  AND U15621 ( .A(n192), .B(n15773), .Z(n15772) );
  XNOR U15622 ( .A(n15774), .B(n15775), .Z(n15769) );
  AND U15623 ( .A(n184), .B(n15776), .Z(n15775) );
  XOR U15624 ( .A(p_input[352]), .B(n15774), .Z(n15776) );
  XNOR U15625 ( .A(n15777), .B(n15778), .Z(n15774) );
  AND U15626 ( .A(n188), .B(n15773), .Z(n15778) );
  XNOR U15627 ( .A(n15777), .B(n15771), .Z(n15773) );
  XOR U15628 ( .A(n15779), .B(n15780), .Z(n15771) );
  AND U15629 ( .A(n203), .B(n15781), .Z(n15780) );
  XNOR U15630 ( .A(n15782), .B(n15783), .Z(n15777) );
  AND U15631 ( .A(n195), .B(n15784), .Z(n15783) );
  XOR U15632 ( .A(p_input[384]), .B(n15782), .Z(n15784) );
  XNOR U15633 ( .A(n15785), .B(n15786), .Z(n15782) );
  AND U15634 ( .A(n199), .B(n15781), .Z(n15786) );
  XNOR U15635 ( .A(n15785), .B(n15779), .Z(n15781) );
  XOR U15636 ( .A(n15787), .B(n15788), .Z(n15779) );
  AND U15637 ( .A(n214), .B(n15789), .Z(n15788) );
  XNOR U15638 ( .A(n15790), .B(n15791), .Z(n15785) );
  AND U15639 ( .A(n206), .B(n15792), .Z(n15791) );
  XOR U15640 ( .A(p_input[416]), .B(n15790), .Z(n15792) );
  XNOR U15641 ( .A(n15793), .B(n15794), .Z(n15790) );
  AND U15642 ( .A(n210), .B(n15789), .Z(n15794) );
  XNOR U15643 ( .A(n15793), .B(n15787), .Z(n15789) );
  XOR U15644 ( .A(n15795), .B(n15796), .Z(n15787) );
  AND U15645 ( .A(n225), .B(n15797), .Z(n15796) );
  XNOR U15646 ( .A(n15798), .B(n15799), .Z(n15793) );
  AND U15647 ( .A(n217), .B(n15800), .Z(n15799) );
  XOR U15648 ( .A(p_input[448]), .B(n15798), .Z(n15800) );
  XNOR U15649 ( .A(n15801), .B(n15802), .Z(n15798) );
  AND U15650 ( .A(n221), .B(n15797), .Z(n15802) );
  XNOR U15651 ( .A(n15801), .B(n15795), .Z(n15797) );
  XOR U15652 ( .A(n15803), .B(n15804), .Z(n15795) );
  AND U15653 ( .A(n236), .B(n15805), .Z(n15804) );
  XNOR U15654 ( .A(n15806), .B(n15807), .Z(n15801) );
  AND U15655 ( .A(n228), .B(n15808), .Z(n15807) );
  XOR U15656 ( .A(p_input[480]), .B(n15806), .Z(n15808) );
  XNOR U15657 ( .A(n15809), .B(n15810), .Z(n15806) );
  AND U15658 ( .A(n232), .B(n15805), .Z(n15810) );
  XNOR U15659 ( .A(n15809), .B(n15803), .Z(n15805) );
  XOR U15660 ( .A(n15811), .B(n15812), .Z(n15803) );
  AND U15661 ( .A(n247), .B(n15813), .Z(n15812) );
  XNOR U15662 ( .A(n15814), .B(n15815), .Z(n15809) );
  AND U15663 ( .A(n239), .B(n15816), .Z(n15815) );
  XOR U15664 ( .A(p_input[512]), .B(n15814), .Z(n15816) );
  XNOR U15665 ( .A(n15817), .B(n15818), .Z(n15814) );
  AND U15666 ( .A(n243), .B(n15813), .Z(n15818) );
  XNOR U15667 ( .A(n15817), .B(n15811), .Z(n15813) );
  XOR U15668 ( .A(n15819), .B(n15820), .Z(n15811) );
  AND U15669 ( .A(n258), .B(n15821), .Z(n15820) );
  XNOR U15670 ( .A(n15822), .B(n15823), .Z(n15817) );
  AND U15671 ( .A(n250), .B(n15824), .Z(n15823) );
  XOR U15672 ( .A(p_input[544]), .B(n15822), .Z(n15824) );
  XNOR U15673 ( .A(n15825), .B(n15826), .Z(n15822) );
  AND U15674 ( .A(n254), .B(n15821), .Z(n15826) );
  XNOR U15675 ( .A(n15825), .B(n15819), .Z(n15821) );
  XOR U15676 ( .A(n15827), .B(n15828), .Z(n15819) );
  AND U15677 ( .A(n269), .B(n15829), .Z(n15828) );
  XNOR U15678 ( .A(n15830), .B(n15831), .Z(n15825) );
  AND U15679 ( .A(n261), .B(n15832), .Z(n15831) );
  XOR U15680 ( .A(p_input[576]), .B(n15830), .Z(n15832) );
  XNOR U15681 ( .A(n15833), .B(n15834), .Z(n15830) );
  AND U15682 ( .A(n265), .B(n15829), .Z(n15834) );
  XNOR U15683 ( .A(n15833), .B(n15827), .Z(n15829) );
  XOR U15684 ( .A(n15835), .B(n15836), .Z(n15827) );
  AND U15685 ( .A(n280), .B(n15837), .Z(n15836) );
  XNOR U15686 ( .A(n15838), .B(n15839), .Z(n15833) );
  AND U15687 ( .A(n272), .B(n15840), .Z(n15839) );
  XOR U15688 ( .A(p_input[608]), .B(n15838), .Z(n15840) );
  XNOR U15689 ( .A(n15841), .B(n15842), .Z(n15838) );
  AND U15690 ( .A(n276), .B(n15837), .Z(n15842) );
  XNOR U15691 ( .A(n15841), .B(n15835), .Z(n15837) );
  XOR U15692 ( .A(n15843), .B(n15844), .Z(n15835) );
  AND U15693 ( .A(n291), .B(n15845), .Z(n15844) );
  XNOR U15694 ( .A(n15846), .B(n15847), .Z(n15841) );
  AND U15695 ( .A(n283), .B(n15848), .Z(n15847) );
  XOR U15696 ( .A(p_input[640]), .B(n15846), .Z(n15848) );
  XNOR U15697 ( .A(n15849), .B(n15850), .Z(n15846) );
  AND U15698 ( .A(n287), .B(n15845), .Z(n15850) );
  XNOR U15699 ( .A(n15849), .B(n15843), .Z(n15845) );
  XOR U15700 ( .A(n15851), .B(n15852), .Z(n15843) );
  AND U15701 ( .A(n302), .B(n15853), .Z(n15852) );
  XNOR U15702 ( .A(n15854), .B(n15855), .Z(n15849) );
  AND U15703 ( .A(n294), .B(n15856), .Z(n15855) );
  XOR U15704 ( .A(p_input[672]), .B(n15854), .Z(n15856) );
  XNOR U15705 ( .A(n15857), .B(n15858), .Z(n15854) );
  AND U15706 ( .A(n298), .B(n15853), .Z(n15858) );
  XNOR U15707 ( .A(n15857), .B(n15851), .Z(n15853) );
  XOR U15708 ( .A(n15859), .B(n15860), .Z(n15851) );
  AND U15709 ( .A(n313), .B(n15861), .Z(n15860) );
  XNOR U15710 ( .A(n15862), .B(n15863), .Z(n15857) );
  AND U15711 ( .A(n305), .B(n15864), .Z(n15863) );
  XOR U15712 ( .A(p_input[704]), .B(n15862), .Z(n15864) );
  XNOR U15713 ( .A(n15865), .B(n15866), .Z(n15862) );
  AND U15714 ( .A(n309), .B(n15861), .Z(n15866) );
  XNOR U15715 ( .A(n15865), .B(n15859), .Z(n15861) );
  XOR U15716 ( .A(n15867), .B(n15868), .Z(n15859) );
  AND U15717 ( .A(n324), .B(n15869), .Z(n15868) );
  XNOR U15718 ( .A(n15870), .B(n15871), .Z(n15865) );
  AND U15719 ( .A(n316), .B(n15872), .Z(n15871) );
  XOR U15720 ( .A(p_input[736]), .B(n15870), .Z(n15872) );
  XNOR U15721 ( .A(n15873), .B(n15874), .Z(n15870) );
  AND U15722 ( .A(n320), .B(n15869), .Z(n15874) );
  XNOR U15723 ( .A(n15873), .B(n15867), .Z(n15869) );
  XOR U15724 ( .A(n15875), .B(n15876), .Z(n15867) );
  AND U15725 ( .A(n335), .B(n15877), .Z(n15876) );
  XNOR U15726 ( .A(n15878), .B(n15879), .Z(n15873) );
  AND U15727 ( .A(n327), .B(n15880), .Z(n15879) );
  XOR U15728 ( .A(p_input[768]), .B(n15878), .Z(n15880) );
  XNOR U15729 ( .A(n15881), .B(n15882), .Z(n15878) );
  AND U15730 ( .A(n331), .B(n15877), .Z(n15882) );
  XNOR U15731 ( .A(n15881), .B(n15875), .Z(n15877) );
  XOR U15732 ( .A(n15883), .B(n15884), .Z(n15875) );
  AND U15733 ( .A(n346), .B(n15885), .Z(n15884) );
  XNOR U15734 ( .A(n15886), .B(n15887), .Z(n15881) );
  AND U15735 ( .A(n338), .B(n15888), .Z(n15887) );
  XOR U15736 ( .A(p_input[800]), .B(n15886), .Z(n15888) );
  XNOR U15737 ( .A(n15889), .B(n15890), .Z(n15886) );
  AND U15738 ( .A(n342), .B(n15885), .Z(n15890) );
  XNOR U15739 ( .A(n15889), .B(n15883), .Z(n15885) );
  XOR U15740 ( .A(n15891), .B(n15892), .Z(n15883) );
  AND U15741 ( .A(n357), .B(n15893), .Z(n15892) );
  XNOR U15742 ( .A(n15894), .B(n15895), .Z(n15889) );
  AND U15743 ( .A(n349), .B(n15896), .Z(n15895) );
  XOR U15744 ( .A(p_input[832]), .B(n15894), .Z(n15896) );
  XNOR U15745 ( .A(n15897), .B(n15898), .Z(n15894) );
  AND U15746 ( .A(n353), .B(n15893), .Z(n15898) );
  XNOR U15747 ( .A(n15897), .B(n15891), .Z(n15893) );
  XOR U15748 ( .A(n15899), .B(n15900), .Z(n15891) );
  AND U15749 ( .A(n368), .B(n15901), .Z(n15900) );
  XNOR U15750 ( .A(n15902), .B(n15903), .Z(n15897) );
  AND U15751 ( .A(n360), .B(n15904), .Z(n15903) );
  XOR U15752 ( .A(p_input[864]), .B(n15902), .Z(n15904) );
  XNOR U15753 ( .A(n15905), .B(n15906), .Z(n15902) );
  AND U15754 ( .A(n364), .B(n15901), .Z(n15906) );
  XNOR U15755 ( .A(n15905), .B(n15899), .Z(n15901) );
  XOR U15756 ( .A(n15907), .B(n15908), .Z(n15899) );
  AND U15757 ( .A(n379), .B(n15909), .Z(n15908) );
  XNOR U15758 ( .A(n15910), .B(n15911), .Z(n15905) );
  AND U15759 ( .A(n371), .B(n15912), .Z(n15911) );
  XOR U15760 ( .A(p_input[896]), .B(n15910), .Z(n15912) );
  XNOR U15761 ( .A(n15913), .B(n15914), .Z(n15910) );
  AND U15762 ( .A(n375), .B(n15909), .Z(n15914) );
  XNOR U15763 ( .A(n15913), .B(n15907), .Z(n15909) );
  XOR U15764 ( .A(n15915), .B(n15916), .Z(n15907) );
  AND U15765 ( .A(n390), .B(n15917), .Z(n15916) );
  XNOR U15766 ( .A(n15918), .B(n15919), .Z(n15913) );
  AND U15767 ( .A(n382), .B(n15920), .Z(n15919) );
  XOR U15768 ( .A(p_input[928]), .B(n15918), .Z(n15920) );
  XNOR U15769 ( .A(n15921), .B(n15922), .Z(n15918) );
  AND U15770 ( .A(n386), .B(n15917), .Z(n15922) );
  XNOR U15771 ( .A(n15921), .B(n15915), .Z(n15917) );
  XOR U15772 ( .A(n15923), .B(n15924), .Z(n15915) );
  AND U15773 ( .A(n401), .B(n15925), .Z(n15924) );
  XNOR U15774 ( .A(n15926), .B(n15927), .Z(n15921) );
  AND U15775 ( .A(n393), .B(n15928), .Z(n15927) );
  XOR U15776 ( .A(p_input[960]), .B(n15926), .Z(n15928) );
  XNOR U15777 ( .A(n15929), .B(n15930), .Z(n15926) );
  AND U15778 ( .A(n397), .B(n15925), .Z(n15930) );
  XNOR U15779 ( .A(n15929), .B(n15923), .Z(n15925) );
  XOR U15780 ( .A(n15931), .B(n15932), .Z(n15923) );
  AND U15781 ( .A(n412), .B(n15933), .Z(n15932) );
  XNOR U15782 ( .A(n15934), .B(n15935), .Z(n15929) );
  AND U15783 ( .A(n404), .B(n15936), .Z(n15935) );
  XOR U15784 ( .A(p_input[992]), .B(n15934), .Z(n15936) );
  XNOR U15785 ( .A(n15937), .B(n15938), .Z(n15934) );
  AND U15786 ( .A(n408), .B(n15933), .Z(n15938) );
  XNOR U15787 ( .A(n15937), .B(n15931), .Z(n15933) );
  XOR U15788 ( .A(n15939), .B(n15940), .Z(n15931) );
  AND U15789 ( .A(n423), .B(n15941), .Z(n15940) );
  XNOR U15790 ( .A(n15942), .B(n15943), .Z(n15937) );
  AND U15791 ( .A(n415), .B(n15944), .Z(n15943) );
  XOR U15792 ( .A(p_input[1024]), .B(n15942), .Z(n15944) );
  XNOR U15793 ( .A(n15945), .B(n15946), .Z(n15942) );
  AND U15794 ( .A(n419), .B(n15941), .Z(n15946) );
  XNOR U15795 ( .A(n15945), .B(n15939), .Z(n15941) );
  XOR U15796 ( .A(n15947), .B(n15948), .Z(n15939) );
  AND U15797 ( .A(n434), .B(n15949), .Z(n15948) );
  XNOR U15798 ( .A(n15950), .B(n15951), .Z(n15945) );
  AND U15799 ( .A(n426), .B(n15952), .Z(n15951) );
  XOR U15800 ( .A(p_input[1056]), .B(n15950), .Z(n15952) );
  XNOR U15801 ( .A(n15953), .B(n15954), .Z(n15950) );
  AND U15802 ( .A(n430), .B(n15949), .Z(n15954) );
  XNOR U15803 ( .A(n15953), .B(n15947), .Z(n15949) );
  XOR U15804 ( .A(n15955), .B(n15956), .Z(n15947) );
  AND U15805 ( .A(n445), .B(n15957), .Z(n15956) );
  XNOR U15806 ( .A(n15958), .B(n15959), .Z(n15953) );
  AND U15807 ( .A(n437), .B(n15960), .Z(n15959) );
  XOR U15808 ( .A(p_input[1088]), .B(n15958), .Z(n15960) );
  XNOR U15809 ( .A(n15961), .B(n15962), .Z(n15958) );
  AND U15810 ( .A(n441), .B(n15957), .Z(n15962) );
  XNOR U15811 ( .A(n15961), .B(n15955), .Z(n15957) );
  XOR U15812 ( .A(n15963), .B(n15964), .Z(n15955) );
  AND U15813 ( .A(n456), .B(n15965), .Z(n15964) );
  XNOR U15814 ( .A(n15966), .B(n15967), .Z(n15961) );
  AND U15815 ( .A(n448), .B(n15968), .Z(n15967) );
  XOR U15816 ( .A(p_input[1120]), .B(n15966), .Z(n15968) );
  XNOR U15817 ( .A(n15969), .B(n15970), .Z(n15966) );
  AND U15818 ( .A(n452), .B(n15965), .Z(n15970) );
  XNOR U15819 ( .A(n15969), .B(n15963), .Z(n15965) );
  XOR U15820 ( .A(n15971), .B(n15972), .Z(n15963) );
  AND U15821 ( .A(n467), .B(n15973), .Z(n15972) );
  XNOR U15822 ( .A(n15974), .B(n15975), .Z(n15969) );
  AND U15823 ( .A(n459), .B(n15976), .Z(n15975) );
  XOR U15824 ( .A(p_input[1152]), .B(n15974), .Z(n15976) );
  XNOR U15825 ( .A(n15977), .B(n15978), .Z(n15974) );
  AND U15826 ( .A(n463), .B(n15973), .Z(n15978) );
  XNOR U15827 ( .A(n15977), .B(n15971), .Z(n15973) );
  XOR U15828 ( .A(n15979), .B(n15980), .Z(n15971) );
  AND U15829 ( .A(n478), .B(n15981), .Z(n15980) );
  XNOR U15830 ( .A(n15982), .B(n15983), .Z(n15977) );
  AND U15831 ( .A(n470), .B(n15984), .Z(n15983) );
  XOR U15832 ( .A(p_input[1184]), .B(n15982), .Z(n15984) );
  XNOR U15833 ( .A(n15985), .B(n15986), .Z(n15982) );
  AND U15834 ( .A(n474), .B(n15981), .Z(n15986) );
  XNOR U15835 ( .A(n15985), .B(n15979), .Z(n15981) );
  XOR U15836 ( .A(n15987), .B(n15988), .Z(n15979) );
  AND U15837 ( .A(n489), .B(n15989), .Z(n15988) );
  XNOR U15838 ( .A(n15990), .B(n15991), .Z(n15985) );
  AND U15839 ( .A(n481), .B(n15992), .Z(n15991) );
  XOR U15840 ( .A(p_input[1216]), .B(n15990), .Z(n15992) );
  XNOR U15841 ( .A(n15993), .B(n15994), .Z(n15990) );
  AND U15842 ( .A(n485), .B(n15989), .Z(n15994) );
  XNOR U15843 ( .A(n15993), .B(n15987), .Z(n15989) );
  XOR U15844 ( .A(n15995), .B(n15996), .Z(n15987) );
  AND U15845 ( .A(n500), .B(n15997), .Z(n15996) );
  XNOR U15846 ( .A(n15998), .B(n15999), .Z(n15993) );
  AND U15847 ( .A(n492), .B(n16000), .Z(n15999) );
  XOR U15848 ( .A(p_input[1248]), .B(n15998), .Z(n16000) );
  XNOR U15849 ( .A(n16001), .B(n16002), .Z(n15998) );
  AND U15850 ( .A(n496), .B(n15997), .Z(n16002) );
  XNOR U15851 ( .A(n16001), .B(n15995), .Z(n15997) );
  XOR U15852 ( .A(n16003), .B(n16004), .Z(n15995) );
  AND U15853 ( .A(n511), .B(n16005), .Z(n16004) );
  XNOR U15854 ( .A(n16006), .B(n16007), .Z(n16001) );
  AND U15855 ( .A(n503), .B(n16008), .Z(n16007) );
  XOR U15856 ( .A(p_input[1280]), .B(n16006), .Z(n16008) );
  XNOR U15857 ( .A(n16009), .B(n16010), .Z(n16006) );
  AND U15858 ( .A(n507), .B(n16005), .Z(n16010) );
  XNOR U15859 ( .A(n16009), .B(n16003), .Z(n16005) );
  XOR U15860 ( .A(n16011), .B(n16012), .Z(n16003) );
  AND U15861 ( .A(n522), .B(n16013), .Z(n16012) );
  XNOR U15862 ( .A(n16014), .B(n16015), .Z(n16009) );
  AND U15863 ( .A(n514), .B(n16016), .Z(n16015) );
  XOR U15864 ( .A(p_input[1312]), .B(n16014), .Z(n16016) );
  XNOR U15865 ( .A(n16017), .B(n16018), .Z(n16014) );
  AND U15866 ( .A(n518), .B(n16013), .Z(n16018) );
  XNOR U15867 ( .A(n16017), .B(n16011), .Z(n16013) );
  XOR U15868 ( .A(n16019), .B(n16020), .Z(n16011) );
  AND U15869 ( .A(n533), .B(n16021), .Z(n16020) );
  XNOR U15870 ( .A(n16022), .B(n16023), .Z(n16017) );
  AND U15871 ( .A(n525), .B(n16024), .Z(n16023) );
  XOR U15872 ( .A(p_input[1344]), .B(n16022), .Z(n16024) );
  XNOR U15873 ( .A(n16025), .B(n16026), .Z(n16022) );
  AND U15874 ( .A(n529), .B(n16021), .Z(n16026) );
  XNOR U15875 ( .A(n16025), .B(n16019), .Z(n16021) );
  XOR U15876 ( .A(n16027), .B(n16028), .Z(n16019) );
  AND U15877 ( .A(n544), .B(n16029), .Z(n16028) );
  XNOR U15878 ( .A(n16030), .B(n16031), .Z(n16025) );
  AND U15879 ( .A(n536), .B(n16032), .Z(n16031) );
  XOR U15880 ( .A(p_input[1376]), .B(n16030), .Z(n16032) );
  XNOR U15881 ( .A(n16033), .B(n16034), .Z(n16030) );
  AND U15882 ( .A(n540), .B(n16029), .Z(n16034) );
  XNOR U15883 ( .A(n16033), .B(n16027), .Z(n16029) );
  XOR U15884 ( .A(n16035), .B(n16036), .Z(n16027) );
  AND U15885 ( .A(n555), .B(n16037), .Z(n16036) );
  XNOR U15886 ( .A(n16038), .B(n16039), .Z(n16033) );
  AND U15887 ( .A(n547), .B(n16040), .Z(n16039) );
  XOR U15888 ( .A(p_input[1408]), .B(n16038), .Z(n16040) );
  XNOR U15889 ( .A(n16041), .B(n16042), .Z(n16038) );
  AND U15890 ( .A(n551), .B(n16037), .Z(n16042) );
  XNOR U15891 ( .A(n16041), .B(n16035), .Z(n16037) );
  XOR U15892 ( .A(n16043), .B(n16044), .Z(n16035) );
  AND U15893 ( .A(n566), .B(n16045), .Z(n16044) );
  XNOR U15894 ( .A(n16046), .B(n16047), .Z(n16041) );
  AND U15895 ( .A(n558), .B(n16048), .Z(n16047) );
  XOR U15896 ( .A(p_input[1440]), .B(n16046), .Z(n16048) );
  XNOR U15897 ( .A(n16049), .B(n16050), .Z(n16046) );
  AND U15898 ( .A(n562), .B(n16045), .Z(n16050) );
  XNOR U15899 ( .A(n16049), .B(n16043), .Z(n16045) );
  XOR U15900 ( .A(n16051), .B(n16052), .Z(n16043) );
  AND U15901 ( .A(n577), .B(n16053), .Z(n16052) );
  XNOR U15902 ( .A(n16054), .B(n16055), .Z(n16049) );
  AND U15903 ( .A(n569), .B(n16056), .Z(n16055) );
  XOR U15904 ( .A(p_input[1472]), .B(n16054), .Z(n16056) );
  XNOR U15905 ( .A(n16057), .B(n16058), .Z(n16054) );
  AND U15906 ( .A(n573), .B(n16053), .Z(n16058) );
  XNOR U15907 ( .A(n16057), .B(n16051), .Z(n16053) );
  XOR U15908 ( .A(n16059), .B(n16060), .Z(n16051) );
  AND U15909 ( .A(n588), .B(n16061), .Z(n16060) );
  XNOR U15910 ( .A(n16062), .B(n16063), .Z(n16057) );
  AND U15911 ( .A(n580), .B(n16064), .Z(n16063) );
  XOR U15912 ( .A(p_input[1504]), .B(n16062), .Z(n16064) );
  XNOR U15913 ( .A(n16065), .B(n16066), .Z(n16062) );
  AND U15914 ( .A(n584), .B(n16061), .Z(n16066) );
  XNOR U15915 ( .A(n16065), .B(n16059), .Z(n16061) );
  XOR U15916 ( .A(n16067), .B(n16068), .Z(n16059) );
  AND U15917 ( .A(n599), .B(n16069), .Z(n16068) );
  XNOR U15918 ( .A(n16070), .B(n16071), .Z(n16065) );
  AND U15919 ( .A(n591), .B(n16072), .Z(n16071) );
  XOR U15920 ( .A(p_input[1536]), .B(n16070), .Z(n16072) );
  XNOR U15921 ( .A(n16073), .B(n16074), .Z(n16070) );
  AND U15922 ( .A(n595), .B(n16069), .Z(n16074) );
  XNOR U15923 ( .A(n16073), .B(n16067), .Z(n16069) );
  XOR U15924 ( .A(n16075), .B(n16076), .Z(n16067) );
  AND U15925 ( .A(n610), .B(n16077), .Z(n16076) );
  XNOR U15926 ( .A(n16078), .B(n16079), .Z(n16073) );
  AND U15927 ( .A(n602), .B(n16080), .Z(n16079) );
  XOR U15928 ( .A(p_input[1568]), .B(n16078), .Z(n16080) );
  XNOR U15929 ( .A(n16081), .B(n16082), .Z(n16078) );
  AND U15930 ( .A(n606), .B(n16077), .Z(n16082) );
  XNOR U15931 ( .A(n16081), .B(n16075), .Z(n16077) );
  XOR U15932 ( .A(n16083), .B(n16084), .Z(n16075) );
  AND U15933 ( .A(n621), .B(n16085), .Z(n16084) );
  XNOR U15934 ( .A(n16086), .B(n16087), .Z(n16081) );
  AND U15935 ( .A(n613), .B(n16088), .Z(n16087) );
  XOR U15936 ( .A(p_input[1600]), .B(n16086), .Z(n16088) );
  XNOR U15937 ( .A(n16089), .B(n16090), .Z(n16086) );
  AND U15938 ( .A(n617), .B(n16085), .Z(n16090) );
  XNOR U15939 ( .A(n16089), .B(n16083), .Z(n16085) );
  XOR U15940 ( .A(n16091), .B(n16092), .Z(n16083) );
  AND U15941 ( .A(n632), .B(n16093), .Z(n16092) );
  XNOR U15942 ( .A(n16094), .B(n16095), .Z(n16089) );
  AND U15943 ( .A(n624), .B(n16096), .Z(n16095) );
  XOR U15944 ( .A(p_input[1632]), .B(n16094), .Z(n16096) );
  XNOR U15945 ( .A(n16097), .B(n16098), .Z(n16094) );
  AND U15946 ( .A(n628), .B(n16093), .Z(n16098) );
  XNOR U15947 ( .A(n16097), .B(n16091), .Z(n16093) );
  XOR U15948 ( .A(n16099), .B(n16100), .Z(n16091) );
  AND U15949 ( .A(n643), .B(n16101), .Z(n16100) );
  XNOR U15950 ( .A(n16102), .B(n16103), .Z(n16097) );
  AND U15951 ( .A(n635), .B(n16104), .Z(n16103) );
  XOR U15952 ( .A(p_input[1664]), .B(n16102), .Z(n16104) );
  XNOR U15953 ( .A(n16105), .B(n16106), .Z(n16102) );
  AND U15954 ( .A(n639), .B(n16101), .Z(n16106) );
  XNOR U15955 ( .A(n16105), .B(n16099), .Z(n16101) );
  XOR U15956 ( .A(n16107), .B(n16108), .Z(n16099) );
  AND U15957 ( .A(n654), .B(n16109), .Z(n16108) );
  XNOR U15958 ( .A(n16110), .B(n16111), .Z(n16105) );
  AND U15959 ( .A(n646), .B(n16112), .Z(n16111) );
  XOR U15960 ( .A(p_input[1696]), .B(n16110), .Z(n16112) );
  XNOR U15961 ( .A(n16113), .B(n16114), .Z(n16110) );
  AND U15962 ( .A(n650), .B(n16109), .Z(n16114) );
  XNOR U15963 ( .A(n16113), .B(n16107), .Z(n16109) );
  XOR U15964 ( .A(n16115), .B(n16116), .Z(n16107) );
  AND U15965 ( .A(n665), .B(n16117), .Z(n16116) );
  XNOR U15966 ( .A(n16118), .B(n16119), .Z(n16113) );
  AND U15967 ( .A(n657), .B(n16120), .Z(n16119) );
  XOR U15968 ( .A(p_input[1728]), .B(n16118), .Z(n16120) );
  XNOR U15969 ( .A(n16121), .B(n16122), .Z(n16118) );
  AND U15970 ( .A(n661), .B(n16117), .Z(n16122) );
  XNOR U15971 ( .A(n16121), .B(n16115), .Z(n16117) );
  XOR U15972 ( .A(n16123), .B(n16124), .Z(n16115) );
  AND U15973 ( .A(n676), .B(n16125), .Z(n16124) );
  XNOR U15974 ( .A(n16126), .B(n16127), .Z(n16121) );
  AND U15975 ( .A(n668), .B(n16128), .Z(n16127) );
  XOR U15976 ( .A(p_input[1760]), .B(n16126), .Z(n16128) );
  XNOR U15977 ( .A(n16129), .B(n16130), .Z(n16126) );
  AND U15978 ( .A(n672), .B(n16125), .Z(n16130) );
  XNOR U15979 ( .A(n16129), .B(n16123), .Z(n16125) );
  XOR U15980 ( .A(n16131), .B(n16132), .Z(n16123) );
  AND U15981 ( .A(n687), .B(n16133), .Z(n16132) );
  XNOR U15982 ( .A(n16134), .B(n16135), .Z(n16129) );
  AND U15983 ( .A(n679), .B(n16136), .Z(n16135) );
  XOR U15984 ( .A(p_input[1792]), .B(n16134), .Z(n16136) );
  XNOR U15985 ( .A(n16137), .B(n16138), .Z(n16134) );
  AND U15986 ( .A(n683), .B(n16133), .Z(n16138) );
  XNOR U15987 ( .A(n16137), .B(n16131), .Z(n16133) );
  XOR U15988 ( .A(n16139), .B(n16140), .Z(n16131) );
  AND U15989 ( .A(n698), .B(n16141), .Z(n16140) );
  XNOR U15990 ( .A(n16142), .B(n16143), .Z(n16137) );
  AND U15991 ( .A(n690), .B(n16144), .Z(n16143) );
  XOR U15992 ( .A(p_input[1824]), .B(n16142), .Z(n16144) );
  XNOR U15993 ( .A(n16145), .B(n16146), .Z(n16142) );
  AND U15994 ( .A(n694), .B(n16141), .Z(n16146) );
  XNOR U15995 ( .A(n16145), .B(n16139), .Z(n16141) );
  XOR U15996 ( .A(n16147), .B(n16148), .Z(n16139) );
  AND U15997 ( .A(n709), .B(n16149), .Z(n16148) );
  XNOR U15998 ( .A(n16150), .B(n16151), .Z(n16145) );
  AND U15999 ( .A(n701), .B(n16152), .Z(n16151) );
  XOR U16000 ( .A(p_input[1856]), .B(n16150), .Z(n16152) );
  XNOR U16001 ( .A(n16153), .B(n16154), .Z(n16150) );
  AND U16002 ( .A(n705), .B(n16149), .Z(n16154) );
  XNOR U16003 ( .A(n16153), .B(n16147), .Z(n16149) );
  XOR U16004 ( .A(n16155), .B(n16156), .Z(n16147) );
  AND U16005 ( .A(n720), .B(n16157), .Z(n16156) );
  XNOR U16006 ( .A(n16158), .B(n16159), .Z(n16153) );
  AND U16007 ( .A(n712), .B(n16160), .Z(n16159) );
  XOR U16008 ( .A(p_input[1888]), .B(n16158), .Z(n16160) );
  XNOR U16009 ( .A(n16161), .B(n16162), .Z(n16158) );
  AND U16010 ( .A(n716), .B(n16157), .Z(n16162) );
  XNOR U16011 ( .A(n16161), .B(n16155), .Z(n16157) );
  XOR U16012 ( .A(n16163), .B(n16164), .Z(n16155) );
  AND U16013 ( .A(n731), .B(n16165), .Z(n16164) );
  XNOR U16014 ( .A(n16166), .B(n16167), .Z(n16161) );
  AND U16015 ( .A(n723), .B(n16168), .Z(n16167) );
  XOR U16016 ( .A(p_input[1920]), .B(n16166), .Z(n16168) );
  XNOR U16017 ( .A(n16169), .B(n16170), .Z(n16166) );
  AND U16018 ( .A(n727), .B(n16165), .Z(n16170) );
  XNOR U16019 ( .A(n16169), .B(n16163), .Z(n16165) );
  XOR U16020 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n16171), .Z(n16163) );
  AND U16021 ( .A(n741), .B(n16172), .Z(n16171) );
  XNOR U16022 ( .A(n16173), .B(n16174), .Z(n16169) );
  AND U16023 ( .A(n734), .B(n16175), .Z(n16174) );
  XOR U16024 ( .A(p_input[1952]), .B(n16173), .Z(n16175) );
  XNOR U16025 ( .A(n16176), .B(n16177), .Z(n16173) );
  AND U16026 ( .A(n738), .B(n16172), .Z(n16177) );
  XOR U16027 ( .A(\knn_comb_/min_val_out[0][0] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n16172) );
  IV U16028 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n16176) );
  XNOR U16029 ( .A(n16178), .B(n16179), .Z(n58) );
  AND U16030 ( .A(n16180), .B(n16181), .Z(n16179) );
  XNOR U16031 ( .A(n16178), .B(n16182), .Z(n16181) );
  XOR U16032 ( .A(n16183), .B(n16184), .Z(n16182) );
  AND U16033 ( .A(n62), .B(n16185), .Z(n16184) );
  XNOR U16034 ( .A(n16183), .B(n16186), .Z(n16185) );
  XNOR U16035 ( .A(n16178), .B(n16187), .Z(n16180) );
  XOR U16036 ( .A(n16188), .B(n16189), .Z(n16187) );
  AND U16037 ( .A(n70), .B(n16190), .Z(n16189) );
  XOR U16038 ( .A(n16191), .B(n16192), .Z(n16178) );
  AND U16039 ( .A(n16193), .B(n16194), .Z(n16192) );
  XOR U16040 ( .A(n16195), .B(n16191), .Z(n16194) );
  XOR U16041 ( .A(n16196), .B(n16197), .Z(n16195) );
  AND U16042 ( .A(n62), .B(n16198), .Z(n16197) );
  XOR U16043 ( .A(n16199), .B(n16196), .Z(n16198) );
  XNOR U16044 ( .A(n16191), .B(n16200), .Z(n16193) );
  XOR U16045 ( .A(n16201), .B(n16202), .Z(n16200) );
  AND U16046 ( .A(n70), .B(n16203), .Z(n16202) );
  XOR U16047 ( .A(n16204), .B(n16205), .Z(n16191) );
  AND U16048 ( .A(n16206), .B(n16207), .Z(n16205) );
  XOR U16049 ( .A(n16208), .B(n16204), .Z(n16207) );
  XOR U16050 ( .A(n16209), .B(n16210), .Z(n16208) );
  AND U16051 ( .A(n62), .B(n16211), .Z(n16210) );
  XNOR U16052 ( .A(n16212), .B(n16209), .Z(n16211) );
  XNOR U16053 ( .A(n16204), .B(n16213), .Z(n16206) );
  XOR U16054 ( .A(n16214), .B(n16215), .Z(n16213) );
  AND U16055 ( .A(n70), .B(n16216), .Z(n16215) );
  XOR U16056 ( .A(n16217), .B(n16218), .Z(n16204) );
  AND U16057 ( .A(n16219), .B(n16220), .Z(n16218) );
  XOR U16058 ( .A(n16221), .B(n16217), .Z(n16220) );
  XOR U16059 ( .A(n16222), .B(n16223), .Z(n16221) );
  AND U16060 ( .A(n62), .B(n16224), .Z(n16223) );
  XOR U16061 ( .A(n16225), .B(n16222), .Z(n16224) );
  XNOR U16062 ( .A(n16217), .B(n16226), .Z(n16219) );
  XOR U16063 ( .A(n16227), .B(n16228), .Z(n16226) );
  AND U16064 ( .A(n70), .B(n16229), .Z(n16228) );
  XOR U16065 ( .A(n16230), .B(n16231), .Z(n16217) );
  AND U16066 ( .A(n16232), .B(n16233), .Z(n16231) );
  XOR U16067 ( .A(n16230), .B(n16234), .Z(n16233) );
  XOR U16068 ( .A(n16235), .B(n16236), .Z(n16234) );
  AND U16069 ( .A(n62), .B(n16237), .Z(n16236) );
  XNOR U16070 ( .A(n16238), .B(n16235), .Z(n16237) );
  XNOR U16071 ( .A(n16239), .B(n16230), .Z(n16232) );
  XNOR U16072 ( .A(n16240), .B(n16241), .Z(n16239) );
  AND U16073 ( .A(n70), .B(n16242), .Z(n16241) );
  AND U16074 ( .A(n16243), .B(n16244), .Z(n16230) );
  XNOR U16075 ( .A(n16245), .B(n16246), .Z(n16244) );
  AND U16076 ( .A(n62), .B(n16247), .Z(n16246) );
  XNOR U16077 ( .A(n16248), .B(n16245), .Z(n16247) );
  XNOR U16078 ( .A(n16249), .B(n16250), .Z(n62) );
  AND U16079 ( .A(n16251), .B(n16252), .Z(n16250) );
  XOR U16080 ( .A(n16186), .B(n16249), .Z(n16252) );
  AND U16081 ( .A(n16253), .B(n16254), .Z(n16186) );
  XOR U16082 ( .A(n16249), .B(n16183), .Z(n16251) );
  XNOR U16083 ( .A(n16255), .B(n16256), .Z(n16183) );
  AND U16084 ( .A(n66), .B(n16190), .Z(n16256) );
  XOR U16085 ( .A(n16188), .B(n16255), .Z(n16190) );
  XOR U16086 ( .A(n16257), .B(n16258), .Z(n16249) );
  AND U16087 ( .A(n16259), .B(n16260), .Z(n16258) );
  XNOR U16088 ( .A(n16257), .B(n16253), .Z(n16260) );
  IV U16089 ( .A(n16199), .Z(n16253) );
  XOR U16090 ( .A(n16261), .B(n16262), .Z(n16199) );
  XOR U16091 ( .A(n16263), .B(n16254), .Z(n16262) );
  AND U16092 ( .A(n16212), .B(n16264), .Z(n16254) );
  AND U16093 ( .A(n16265), .B(n16266), .Z(n16263) );
  XOR U16094 ( .A(n16267), .B(n16261), .Z(n16265) );
  XNOR U16095 ( .A(n16196), .B(n16257), .Z(n16259) );
  XNOR U16096 ( .A(n16268), .B(n16269), .Z(n16196) );
  AND U16097 ( .A(n66), .B(n16203), .Z(n16269) );
  XOR U16098 ( .A(n16268), .B(n16270), .Z(n16203) );
  XOR U16099 ( .A(n16271), .B(n16272), .Z(n16257) );
  AND U16100 ( .A(n16273), .B(n16274), .Z(n16272) );
  XNOR U16101 ( .A(n16271), .B(n16212), .Z(n16274) );
  XOR U16102 ( .A(n16275), .B(n16266), .Z(n16212) );
  XNOR U16103 ( .A(n16276), .B(n16261), .Z(n16266) );
  XOR U16104 ( .A(n16277), .B(n16278), .Z(n16261) );
  AND U16105 ( .A(n16279), .B(n16280), .Z(n16278) );
  XOR U16106 ( .A(n16281), .B(n16277), .Z(n16279) );
  XNOR U16107 ( .A(n16282), .B(n16283), .Z(n16276) );
  AND U16108 ( .A(n16284), .B(n16285), .Z(n16283) );
  XOR U16109 ( .A(n16282), .B(n16286), .Z(n16284) );
  XNOR U16110 ( .A(n16267), .B(n16264), .Z(n16275) );
  AND U16111 ( .A(n16287), .B(n16288), .Z(n16264) );
  XOR U16112 ( .A(n16289), .B(n16290), .Z(n16267) );
  AND U16113 ( .A(n16291), .B(n16292), .Z(n16290) );
  XOR U16114 ( .A(n16289), .B(n16293), .Z(n16291) );
  XNOR U16115 ( .A(n16209), .B(n16271), .Z(n16273) );
  XNOR U16116 ( .A(n16294), .B(n16295), .Z(n16209) );
  AND U16117 ( .A(n66), .B(n16216), .Z(n16295) );
  XOR U16118 ( .A(n16294), .B(n16296), .Z(n16216) );
  XOR U16119 ( .A(n16297), .B(n16298), .Z(n16271) );
  AND U16120 ( .A(n16299), .B(n16300), .Z(n16298) );
  XNOR U16121 ( .A(n16297), .B(n16287), .Z(n16300) );
  IV U16122 ( .A(n16225), .Z(n16287) );
  XNOR U16123 ( .A(n16301), .B(n16280), .Z(n16225) );
  XNOR U16124 ( .A(n16302), .B(n16286), .Z(n16280) );
  XOR U16125 ( .A(n16303), .B(n16304), .Z(n16286) );
  AND U16126 ( .A(n16305), .B(n16306), .Z(n16304) );
  XOR U16127 ( .A(n16303), .B(n16307), .Z(n16305) );
  XNOR U16128 ( .A(n16285), .B(n16277), .Z(n16302) );
  XOR U16129 ( .A(n16308), .B(n16309), .Z(n16277) );
  AND U16130 ( .A(n16310), .B(n16311), .Z(n16309) );
  XNOR U16131 ( .A(n16312), .B(n16308), .Z(n16310) );
  XNOR U16132 ( .A(n16313), .B(n16282), .Z(n16285) );
  XOR U16133 ( .A(n16314), .B(n16315), .Z(n16282) );
  AND U16134 ( .A(n16316), .B(n16317), .Z(n16315) );
  XOR U16135 ( .A(n16314), .B(n16318), .Z(n16316) );
  XNOR U16136 ( .A(n16319), .B(n16320), .Z(n16313) );
  AND U16137 ( .A(n16321), .B(n16322), .Z(n16320) );
  XNOR U16138 ( .A(n16319), .B(n16323), .Z(n16321) );
  XNOR U16139 ( .A(n16281), .B(n16288), .Z(n16301) );
  AND U16140 ( .A(n16238), .B(n16324), .Z(n16288) );
  XOR U16141 ( .A(n16293), .B(n16292), .Z(n16281) );
  XNOR U16142 ( .A(n16325), .B(n16289), .Z(n16292) );
  XOR U16143 ( .A(n16326), .B(n16327), .Z(n16289) );
  AND U16144 ( .A(n16328), .B(n16329), .Z(n16327) );
  XOR U16145 ( .A(n16326), .B(n16330), .Z(n16328) );
  XNOR U16146 ( .A(n16331), .B(n16332), .Z(n16325) );
  AND U16147 ( .A(n16333), .B(n16334), .Z(n16332) );
  XOR U16148 ( .A(n16331), .B(n16335), .Z(n16333) );
  XOR U16149 ( .A(n16336), .B(n16337), .Z(n16293) );
  AND U16150 ( .A(n16338), .B(n16339), .Z(n16337) );
  XOR U16151 ( .A(n16336), .B(n16340), .Z(n16338) );
  XNOR U16152 ( .A(n16222), .B(n16297), .Z(n16299) );
  XNOR U16153 ( .A(n16341), .B(n16342), .Z(n16222) );
  AND U16154 ( .A(n66), .B(n16229), .Z(n16342) );
  XOR U16155 ( .A(n16341), .B(n16343), .Z(n16229) );
  XOR U16156 ( .A(n16344), .B(n16345), .Z(n16297) );
  AND U16157 ( .A(n16346), .B(n16347), .Z(n16345) );
  XNOR U16158 ( .A(n16344), .B(n16238), .Z(n16347) );
  XOR U16159 ( .A(n16348), .B(n16311), .Z(n16238) );
  XNOR U16160 ( .A(n16349), .B(n16318), .Z(n16311) );
  XOR U16161 ( .A(n16307), .B(n16306), .Z(n16318) );
  XNOR U16162 ( .A(n16350), .B(n16303), .Z(n16306) );
  XOR U16163 ( .A(n16351), .B(n16352), .Z(n16303) );
  AND U16164 ( .A(n16353), .B(n16354), .Z(n16352) );
  XNOR U16165 ( .A(n16355), .B(n16356), .Z(n16353) );
  IV U16166 ( .A(n16351), .Z(n16355) );
  XNOR U16167 ( .A(n16357), .B(n16358), .Z(n16350) );
  NOR U16168 ( .A(n16359), .B(n16360), .Z(n16358) );
  XNOR U16169 ( .A(n16357), .B(n16361), .Z(n16359) );
  XOR U16170 ( .A(n16362), .B(n16363), .Z(n16307) );
  NOR U16171 ( .A(n16364), .B(n16365), .Z(n16363) );
  XNOR U16172 ( .A(n16362), .B(n16366), .Z(n16364) );
  XNOR U16173 ( .A(n16317), .B(n16308), .Z(n16349) );
  XOR U16174 ( .A(n16367), .B(n16368), .Z(n16308) );
  NOR U16175 ( .A(n16369), .B(n16370), .Z(n16368) );
  XOR U16176 ( .A(n16371), .B(n16372), .Z(n16369) );
  XOR U16177 ( .A(n16373), .B(n16323), .Z(n16317) );
  XNOR U16178 ( .A(n16374), .B(n16375), .Z(n16323) );
  NOR U16179 ( .A(n16376), .B(n16377), .Z(n16375) );
  XNOR U16180 ( .A(n16374), .B(n16378), .Z(n16376) );
  XNOR U16181 ( .A(n16322), .B(n16314), .Z(n16373) );
  XOR U16182 ( .A(n16379), .B(n16380), .Z(n16314) );
  AND U16183 ( .A(n16381), .B(n16382), .Z(n16380) );
  XOR U16184 ( .A(n16379), .B(n16383), .Z(n16381) );
  XNOR U16185 ( .A(n16384), .B(n16319), .Z(n16322) );
  XOR U16186 ( .A(n16385), .B(n16386), .Z(n16319) );
  AND U16187 ( .A(n16387), .B(n16388), .Z(n16386) );
  XOR U16188 ( .A(n16385), .B(n16389), .Z(n16387) );
  XNOR U16189 ( .A(n16390), .B(n16391), .Z(n16384) );
  NOR U16190 ( .A(n16392), .B(n16393), .Z(n16391) );
  XOR U16191 ( .A(n16390), .B(n16394), .Z(n16392) );
  XOR U16192 ( .A(n16312), .B(n16324), .Z(n16348) );
  NOR U16193 ( .A(n16248), .B(n16395), .Z(n16324) );
  XNOR U16194 ( .A(n16330), .B(n16329), .Z(n16312) );
  XNOR U16195 ( .A(n16396), .B(n16335), .Z(n16329) );
  XNOR U16196 ( .A(n16397), .B(n16398), .Z(n16335) );
  NOR U16197 ( .A(n16399), .B(n16400), .Z(n16398) );
  XOR U16198 ( .A(n16397), .B(n16401), .Z(n16399) );
  XNOR U16199 ( .A(n16334), .B(n16326), .Z(n16396) );
  XOR U16200 ( .A(n16402), .B(n16403), .Z(n16326) );
  AND U16201 ( .A(n16404), .B(n16405), .Z(n16403) );
  XNOR U16202 ( .A(n16402), .B(n16406), .Z(n16404) );
  XNOR U16203 ( .A(n16407), .B(n16331), .Z(n16334) );
  XOR U16204 ( .A(n16408), .B(n16409), .Z(n16331) );
  AND U16205 ( .A(n16410), .B(n16411), .Z(n16409) );
  XNOR U16206 ( .A(n16412), .B(n16413), .Z(n16410) );
  IV U16207 ( .A(n16408), .Z(n16412) );
  XNOR U16208 ( .A(n16414), .B(n16415), .Z(n16407) );
  NOR U16209 ( .A(n16416), .B(n16417), .Z(n16415) );
  XNOR U16210 ( .A(n16414), .B(n16418), .Z(n16416) );
  XOR U16211 ( .A(n16340), .B(n16339), .Z(n16330) );
  XNOR U16212 ( .A(n16419), .B(n16336), .Z(n16339) );
  XOR U16213 ( .A(n16420), .B(n16421), .Z(n16336) );
  AND U16214 ( .A(n16422), .B(n16423), .Z(n16421) );
  XOR U16215 ( .A(n16420), .B(n16424), .Z(n16422) );
  XNOR U16216 ( .A(n16425), .B(n16426), .Z(n16419) );
  NOR U16217 ( .A(n16427), .B(n16428), .Z(n16426) );
  XNOR U16218 ( .A(n16425), .B(n16429), .Z(n16427) );
  XOR U16219 ( .A(n16430), .B(n16431), .Z(n16340) );
  NOR U16220 ( .A(n16432), .B(n16433), .Z(n16431) );
  XNOR U16221 ( .A(n16430), .B(n16434), .Z(n16432) );
  XNOR U16222 ( .A(n16235), .B(n16344), .Z(n16346) );
  XNOR U16223 ( .A(n16435), .B(n16436), .Z(n16235) );
  AND U16224 ( .A(n66), .B(n16242), .Z(n16436) );
  XOR U16225 ( .A(n16435), .B(n16240), .Z(n16242) );
  AND U16226 ( .A(n16245), .B(n16248), .Z(n16344) );
  XOR U16227 ( .A(n16437), .B(n16395), .Z(n16248) );
  XNOR U16228 ( .A(p_input[0]), .B(p_input[2048]), .Z(n16395) );
  XOR U16229 ( .A(n16372), .B(n16370), .Z(n16437) );
  XOR U16230 ( .A(n16438), .B(n16383), .Z(n16370) );
  XOR U16231 ( .A(n16356), .B(n16354), .Z(n16383) );
  XNOR U16232 ( .A(n16439), .B(n16361), .Z(n16354) );
  XOR U16233 ( .A(p_input[2072]), .B(p_input[24]), .Z(n16361) );
  XOR U16234 ( .A(n16351), .B(n16360), .Z(n16439) );
  XOR U16235 ( .A(n16440), .B(n16357), .Z(n16360) );
  XOR U16236 ( .A(p_input[2070]), .B(p_input[22]), .Z(n16357) );
  XNOR U16237 ( .A(p_input[2071]), .B(p_input[23]), .Z(n16440) );
  XOR U16238 ( .A(p_input[18]), .B(p_input[2066]), .Z(n16351) );
  XNOR U16239 ( .A(n16366), .B(n16365), .Z(n16356) );
  XOR U16240 ( .A(n16441), .B(n16362), .Z(n16365) );
  XOR U16241 ( .A(p_input[19]), .B(p_input[2067]), .Z(n16362) );
  XNOR U16242 ( .A(p_input[2068]), .B(p_input[20]), .Z(n16441) );
  XOR U16243 ( .A(p_input[2069]), .B(p_input[21]), .Z(n16366) );
  XOR U16244 ( .A(n16382), .B(n16371), .Z(n16438) );
  IV U16245 ( .A(n16367), .Z(n16371) );
  XOR U16246 ( .A(p_input[1]), .B(p_input[2049]), .Z(n16367) );
  XNOR U16247 ( .A(n16442), .B(n16389), .Z(n16382) );
  XNOR U16248 ( .A(n16378), .B(n16377), .Z(n16389) );
  XOR U16249 ( .A(n16443), .B(n16374), .Z(n16377) );
  XNOR U16250 ( .A(n16444), .B(p_input[26]), .Z(n16374) );
  XNOR U16251 ( .A(p_input[2075]), .B(p_input[27]), .Z(n16443) );
  XOR U16252 ( .A(p_input[2076]), .B(p_input[28]), .Z(n16378) );
  XOR U16253 ( .A(n16388), .B(n16445), .Z(n16442) );
  IV U16254 ( .A(n16379), .Z(n16445) );
  XOR U16255 ( .A(p_input[17]), .B(p_input[2065]), .Z(n16379) );
  XOR U16256 ( .A(n16446), .B(n16394), .Z(n16388) );
  XNOR U16257 ( .A(p_input[2079]), .B(p_input[31]), .Z(n16394) );
  XOR U16258 ( .A(n16385), .B(n16393), .Z(n16446) );
  XOR U16259 ( .A(n16447), .B(n16390), .Z(n16393) );
  XOR U16260 ( .A(p_input[2077]), .B(p_input[29]), .Z(n16390) );
  XNOR U16261 ( .A(p_input[2078]), .B(p_input[30]), .Z(n16447) );
  XNOR U16262 ( .A(n16448), .B(p_input[25]), .Z(n16385) );
  XNOR U16263 ( .A(n16406), .B(n16405), .Z(n16372) );
  XNOR U16264 ( .A(n16449), .B(n16413), .Z(n16405) );
  XNOR U16265 ( .A(n16401), .B(n16400), .Z(n16413) );
  XNOR U16266 ( .A(n16450), .B(n16397), .Z(n16400) );
  XNOR U16267 ( .A(p_input[11]), .B(p_input[2059]), .Z(n16397) );
  XOR U16268 ( .A(p_input[12]), .B(n16451), .Z(n16450) );
  XOR U16269 ( .A(p_input[13]), .B(p_input[2061]), .Z(n16401) );
  XNOR U16270 ( .A(n16411), .B(n16402), .Z(n16449) );
  XNOR U16271 ( .A(n16452), .B(p_input[2]), .Z(n16402) );
  XNOR U16272 ( .A(n16453), .B(n16418), .Z(n16411) );
  XNOR U16273 ( .A(p_input[16]), .B(n16454), .Z(n16418) );
  XOR U16274 ( .A(n16408), .B(n16417), .Z(n16453) );
  XOR U16275 ( .A(n16455), .B(n16414), .Z(n16417) );
  XOR U16276 ( .A(p_input[14]), .B(p_input[2062]), .Z(n16414) );
  XOR U16277 ( .A(p_input[15]), .B(n16456), .Z(n16455) );
  XOR U16278 ( .A(p_input[10]), .B(p_input[2058]), .Z(n16408) );
  XNOR U16279 ( .A(n16424), .B(n16423), .Z(n16406) );
  XNOR U16280 ( .A(n16457), .B(n16429), .Z(n16423) );
  XOR U16281 ( .A(p_input[2057]), .B(p_input[9]), .Z(n16429) );
  XOR U16282 ( .A(n16420), .B(n16428), .Z(n16457) );
  XOR U16283 ( .A(n16458), .B(n16425), .Z(n16428) );
  XOR U16284 ( .A(p_input[2055]), .B(p_input[7]), .Z(n16425) );
  XNOR U16285 ( .A(p_input[2056]), .B(p_input[8]), .Z(n16458) );
  XNOR U16286 ( .A(n16459), .B(p_input[3]), .Z(n16420) );
  XNOR U16287 ( .A(n16434), .B(n16433), .Z(n16424) );
  XOR U16288 ( .A(n16460), .B(n16430), .Z(n16433) );
  XOR U16289 ( .A(p_input[2052]), .B(p_input[4]), .Z(n16430) );
  XNOR U16290 ( .A(p_input[2053]), .B(p_input[5]), .Z(n16460) );
  XOR U16291 ( .A(p_input[2054]), .B(p_input[6]), .Z(n16434) );
  XNOR U16292 ( .A(n16461), .B(n16462), .Z(n16245) );
  AND U16293 ( .A(n66), .B(n16463), .Z(n16462) );
  XNOR U16294 ( .A(n16464), .B(n16465), .Z(n66) );
  AND U16295 ( .A(n16466), .B(n16467), .Z(n16465) );
  XOR U16296 ( .A(n16464), .B(n16255), .Z(n16467) );
  XNOR U16297 ( .A(n16464), .B(n16188), .Z(n16466) );
  XOR U16298 ( .A(n16468), .B(n16469), .Z(n16464) );
  AND U16299 ( .A(n16470), .B(n16471), .Z(n16469) );
  XNOR U16300 ( .A(n16268), .B(n16468), .Z(n16471) );
  XOR U16301 ( .A(n16468), .B(n16270), .Z(n16470) );
  XOR U16302 ( .A(n16472), .B(n16473), .Z(n16468) );
  AND U16303 ( .A(n16474), .B(n16475), .Z(n16473) );
  XNOR U16304 ( .A(n16294), .B(n16472), .Z(n16475) );
  XOR U16305 ( .A(n16472), .B(n16296), .Z(n16474) );
  IV U16306 ( .A(n16214), .Z(n16296) );
  XOR U16307 ( .A(n16476), .B(n16477), .Z(n16472) );
  AND U16308 ( .A(n16478), .B(n16479), .Z(n16477) );
  XOR U16309 ( .A(n16476), .B(n16343), .Z(n16478) );
  XOR U16310 ( .A(n16480), .B(n16481), .Z(n16243) );
  AND U16311 ( .A(n70), .B(n16463), .Z(n16481) );
  XNOR U16312 ( .A(n16461), .B(n16480), .Z(n16463) );
  XNOR U16313 ( .A(n16482), .B(n16483), .Z(n70) );
  AND U16314 ( .A(n16484), .B(n16485), .Z(n16483) );
  XNOR U16315 ( .A(n16486), .B(n16482), .Z(n16485) );
  IV U16316 ( .A(n16255), .Z(n16486) );
  XNOR U16317 ( .A(n16487), .B(n16488), .Z(n16255) );
  AND U16318 ( .A(n74), .B(n16489), .Z(n16488) );
  XNOR U16319 ( .A(n16487), .B(n16490), .Z(n16489) );
  XNOR U16320 ( .A(n16188), .B(n16482), .Z(n16484) );
  XOR U16321 ( .A(n16491), .B(n16492), .Z(n16188) );
  AND U16322 ( .A(n82), .B(n16493), .Z(n16492) );
  XOR U16323 ( .A(n16494), .B(n16495), .Z(n16482) );
  AND U16324 ( .A(n16496), .B(n16497), .Z(n16495) );
  XNOR U16325 ( .A(n16494), .B(n16268), .Z(n16497) );
  XNOR U16326 ( .A(n16498), .B(n16499), .Z(n16268) );
  AND U16327 ( .A(n74), .B(n16500), .Z(n16499) );
  XOR U16328 ( .A(n16501), .B(n16498), .Z(n16500) );
  XNOR U16329 ( .A(n16201), .B(n16494), .Z(n16496) );
  IV U16330 ( .A(n16270), .Z(n16201) );
  XOR U16331 ( .A(n16502), .B(n16503), .Z(n16270) );
  AND U16332 ( .A(n82), .B(n16504), .Z(n16503) );
  XOR U16333 ( .A(n16505), .B(n16506), .Z(n16494) );
  AND U16334 ( .A(n16507), .B(n16508), .Z(n16506) );
  XNOR U16335 ( .A(n16505), .B(n16294), .Z(n16508) );
  XNOR U16336 ( .A(n16509), .B(n16510), .Z(n16294) );
  AND U16337 ( .A(n74), .B(n16511), .Z(n16510) );
  XNOR U16338 ( .A(n16512), .B(n16509), .Z(n16511) );
  XNOR U16339 ( .A(n16214), .B(n16505), .Z(n16507) );
  XNOR U16340 ( .A(n16513), .B(n16514), .Z(n16214) );
  AND U16341 ( .A(n82), .B(n16515), .Z(n16514) );
  XOR U16342 ( .A(n16476), .B(n16516), .Z(n16505) );
  AND U16343 ( .A(n16517), .B(n16479), .Z(n16516) );
  XNOR U16344 ( .A(n16341), .B(n16476), .Z(n16479) );
  XNOR U16345 ( .A(n16518), .B(n16519), .Z(n16341) );
  AND U16346 ( .A(n74), .B(n16520), .Z(n16519) );
  XOR U16347 ( .A(n16521), .B(n16518), .Z(n16520) );
  XNOR U16348 ( .A(n16227), .B(n16476), .Z(n16517) );
  IV U16349 ( .A(n16343), .Z(n16227) );
  XOR U16350 ( .A(n16522), .B(n16523), .Z(n16343) );
  AND U16351 ( .A(n82), .B(n16524), .Z(n16523) );
  XOR U16352 ( .A(n16525), .B(n16526), .Z(n16476) );
  AND U16353 ( .A(n16527), .B(n16528), .Z(n16526) );
  XNOR U16354 ( .A(n16525), .B(n16435), .Z(n16528) );
  XNOR U16355 ( .A(n16529), .B(n16530), .Z(n16435) );
  AND U16356 ( .A(n74), .B(n16531), .Z(n16530) );
  XNOR U16357 ( .A(n16532), .B(n16529), .Z(n16531) );
  XNOR U16358 ( .A(n16533), .B(n16525), .Z(n16527) );
  IV U16359 ( .A(n16240), .Z(n16533) );
  XOR U16360 ( .A(n16534), .B(n16535), .Z(n16240) );
  AND U16361 ( .A(n82), .B(n16536), .Z(n16535) );
  AND U16362 ( .A(n16480), .B(n16461), .Z(n16525) );
  XNOR U16363 ( .A(n16537), .B(n16538), .Z(n16461) );
  AND U16364 ( .A(n74), .B(n16539), .Z(n16538) );
  XNOR U16365 ( .A(n16540), .B(n16537), .Z(n16539) );
  XNOR U16366 ( .A(n16541), .B(n16542), .Z(n74) );
  AND U16367 ( .A(n16543), .B(n16544), .Z(n16542) );
  XOR U16368 ( .A(n16490), .B(n16541), .Z(n16544) );
  AND U16369 ( .A(n16545), .B(n16546), .Z(n16490) );
  XOR U16370 ( .A(n16541), .B(n16487), .Z(n16543) );
  XNOR U16371 ( .A(n16547), .B(n16548), .Z(n16487) );
  AND U16372 ( .A(n78), .B(n16493), .Z(n16548) );
  XOR U16373 ( .A(n16491), .B(n16547), .Z(n16493) );
  XOR U16374 ( .A(n16549), .B(n16550), .Z(n16541) );
  AND U16375 ( .A(n16551), .B(n16552), .Z(n16550) );
  XNOR U16376 ( .A(n16549), .B(n16545), .Z(n16552) );
  IV U16377 ( .A(n16501), .Z(n16545) );
  XOR U16378 ( .A(n16553), .B(n16554), .Z(n16501) );
  XOR U16379 ( .A(n16555), .B(n16546), .Z(n16554) );
  AND U16380 ( .A(n16512), .B(n16556), .Z(n16546) );
  AND U16381 ( .A(n16557), .B(n16558), .Z(n16555) );
  XOR U16382 ( .A(n16559), .B(n16553), .Z(n16557) );
  XNOR U16383 ( .A(n16498), .B(n16549), .Z(n16551) );
  XNOR U16384 ( .A(n16560), .B(n16561), .Z(n16498) );
  AND U16385 ( .A(n78), .B(n16504), .Z(n16561) );
  XOR U16386 ( .A(n16560), .B(n16502), .Z(n16504) );
  XOR U16387 ( .A(n16562), .B(n16563), .Z(n16549) );
  AND U16388 ( .A(n16564), .B(n16565), .Z(n16563) );
  XNOR U16389 ( .A(n16562), .B(n16512), .Z(n16565) );
  XOR U16390 ( .A(n16566), .B(n16558), .Z(n16512) );
  XNOR U16391 ( .A(n16567), .B(n16553), .Z(n16558) );
  XOR U16392 ( .A(n16568), .B(n16569), .Z(n16553) );
  AND U16393 ( .A(n16570), .B(n16571), .Z(n16569) );
  XOR U16394 ( .A(n16572), .B(n16568), .Z(n16570) );
  XNOR U16395 ( .A(n16573), .B(n16574), .Z(n16567) );
  AND U16396 ( .A(n16575), .B(n16576), .Z(n16574) );
  XOR U16397 ( .A(n16573), .B(n16577), .Z(n16575) );
  XNOR U16398 ( .A(n16559), .B(n16556), .Z(n16566) );
  AND U16399 ( .A(n16578), .B(n16579), .Z(n16556) );
  XOR U16400 ( .A(n16580), .B(n16581), .Z(n16559) );
  AND U16401 ( .A(n16582), .B(n16583), .Z(n16581) );
  XOR U16402 ( .A(n16580), .B(n16584), .Z(n16582) );
  XNOR U16403 ( .A(n16509), .B(n16562), .Z(n16564) );
  XNOR U16404 ( .A(n16585), .B(n16586), .Z(n16509) );
  AND U16405 ( .A(n78), .B(n16515), .Z(n16586) );
  XOR U16406 ( .A(n16585), .B(n16513), .Z(n16515) );
  XOR U16407 ( .A(n16587), .B(n16588), .Z(n16562) );
  AND U16408 ( .A(n16589), .B(n16590), .Z(n16588) );
  XNOR U16409 ( .A(n16587), .B(n16578), .Z(n16590) );
  IV U16410 ( .A(n16521), .Z(n16578) );
  XNOR U16411 ( .A(n16591), .B(n16571), .Z(n16521) );
  XNOR U16412 ( .A(n16592), .B(n16577), .Z(n16571) );
  XOR U16413 ( .A(n16593), .B(n16594), .Z(n16577) );
  AND U16414 ( .A(n16595), .B(n16596), .Z(n16594) );
  XOR U16415 ( .A(n16593), .B(n16597), .Z(n16595) );
  XNOR U16416 ( .A(n16576), .B(n16568), .Z(n16592) );
  XOR U16417 ( .A(n16598), .B(n16599), .Z(n16568) );
  AND U16418 ( .A(n16600), .B(n16601), .Z(n16599) );
  XNOR U16419 ( .A(n16602), .B(n16598), .Z(n16600) );
  XNOR U16420 ( .A(n16603), .B(n16573), .Z(n16576) );
  XOR U16421 ( .A(n16604), .B(n16605), .Z(n16573) );
  AND U16422 ( .A(n16606), .B(n16607), .Z(n16605) );
  XOR U16423 ( .A(n16604), .B(n16608), .Z(n16606) );
  XNOR U16424 ( .A(n16609), .B(n16610), .Z(n16603) );
  AND U16425 ( .A(n16611), .B(n16612), .Z(n16610) );
  XNOR U16426 ( .A(n16609), .B(n16613), .Z(n16611) );
  XNOR U16427 ( .A(n16572), .B(n16579), .Z(n16591) );
  AND U16428 ( .A(n16532), .B(n16614), .Z(n16579) );
  XOR U16429 ( .A(n16584), .B(n16583), .Z(n16572) );
  XNOR U16430 ( .A(n16615), .B(n16580), .Z(n16583) );
  XOR U16431 ( .A(n16616), .B(n16617), .Z(n16580) );
  AND U16432 ( .A(n16618), .B(n16619), .Z(n16617) );
  XOR U16433 ( .A(n16616), .B(n16620), .Z(n16618) );
  XNOR U16434 ( .A(n16621), .B(n16622), .Z(n16615) );
  AND U16435 ( .A(n16623), .B(n16624), .Z(n16622) );
  XOR U16436 ( .A(n16621), .B(n16625), .Z(n16623) );
  XOR U16437 ( .A(n16626), .B(n16627), .Z(n16584) );
  AND U16438 ( .A(n16628), .B(n16629), .Z(n16627) );
  XOR U16439 ( .A(n16626), .B(n16630), .Z(n16628) );
  XNOR U16440 ( .A(n16518), .B(n16587), .Z(n16589) );
  XNOR U16441 ( .A(n16631), .B(n16632), .Z(n16518) );
  AND U16442 ( .A(n78), .B(n16524), .Z(n16632) );
  XOR U16443 ( .A(n16631), .B(n16522), .Z(n16524) );
  XOR U16444 ( .A(n16633), .B(n16634), .Z(n16587) );
  AND U16445 ( .A(n16635), .B(n16636), .Z(n16634) );
  XNOR U16446 ( .A(n16633), .B(n16532), .Z(n16636) );
  XOR U16447 ( .A(n16637), .B(n16601), .Z(n16532) );
  XNOR U16448 ( .A(n16638), .B(n16608), .Z(n16601) );
  XOR U16449 ( .A(n16597), .B(n16596), .Z(n16608) );
  XNOR U16450 ( .A(n16639), .B(n16593), .Z(n16596) );
  XOR U16451 ( .A(n16640), .B(n16641), .Z(n16593) );
  AND U16452 ( .A(n16642), .B(n16643), .Z(n16641) );
  XOR U16453 ( .A(n16640), .B(n16644), .Z(n16642) );
  XNOR U16454 ( .A(n16645), .B(n16646), .Z(n16639) );
  NOR U16455 ( .A(n16647), .B(n16648), .Z(n16646) );
  XNOR U16456 ( .A(n16645), .B(n16649), .Z(n16647) );
  XOR U16457 ( .A(n16650), .B(n16651), .Z(n16597) );
  NOR U16458 ( .A(n16652), .B(n16653), .Z(n16651) );
  XNOR U16459 ( .A(n16650), .B(n16654), .Z(n16652) );
  XNOR U16460 ( .A(n16607), .B(n16598), .Z(n16638) );
  XOR U16461 ( .A(n16655), .B(n16656), .Z(n16598) );
  NOR U16462 ( .A(n16657), .B(n16658), .Z(n16656) );
  XNOR U16463 ( .A(n16655), .B(n16659), .Z(n16657) );
  XOR U16464 ( .A(n16660), .B(n16613), .Z(n16607) );
  XNOR U16465 ( .A(n16661), .B(n16662), .Z(n16613) );
  NOR U16466 ( .A(n16663), .B(n16664), .Z(n16662) );
  XNOR U16467 ( .A(n16661), .B(n16665), .Z(n16663) );
  XNOR U16468 ( .A(n16612), .B(n16604), .Z(n16660) );
  XOR U16469 ( .A(n16666), .B(n16667), .Z(n16604) );
  AND U16470 ( .A(n16668), .B(n16669), .Z(n16667) );
  XOR U16471 ( .A(n16666), .B(n16670), .Z(n16668) );
  XNOR U16472 ( .A(n16671), .B(n16609), .Z(n16612) );
  XOR U16473 ( .A(n16672), .B(n16673), .Z(n16609) );
  AND U16474 ( .A(n16674), .B(n16675), .Z(n16673) );
  XOR U16475 ( .A(n16672), .B(n16676), .Z(n16674) );
  XNOR U16476 ( .A(n16677), .B(n16678), .Z(n16671) );
  NOR U16477 ( .A(n16679), .B(n16680), .Z(n16678) );
  XOR U16478 ( .A(n16677), .B(n16681), .Z(n16679) );
  XOR U16479 ( .A(n16602), .B(n16614), .Z(n16637) );
  NOR U16480 ( .A(n16540), .B(n16682), .Z(n16614) );
  XNOR U16481 ( .A(n16620), .B(n16619), .Z(n16602) );
  XNOR U16482 ( .A(n16683), .B(n16625), .Z(n16619) );
  XOR U16483 ( .A(n16684), .B(n16685), .Z(n16625) );
  NOR U16484 ( .A(n16686), .B(n16687), .Z(n16685) );
  XNOR U16485 ( .A(n16684), .B(n16688), .Z(n16686) );
  XNOR U16486 ( .A(n16624), .B(n16616), .Z(n16683) );
  XOR U16487 ( .A(n16689), .B(n16690), .Z(n16616) );
  AND U16488 ( .A(n16691), .B(n16692), .Z(n16690) );
  XNOR U16489 ( .A(n16689), .B(n16693), .Z(n16691) );
  XNOR U16490 ( .A(n16694), .B(n16621), .Z(n16624) );
  XOR U16491 ( .A(n16695), .B(n16696), .Z(n16621) );
  AND U16492 ( .A(n16697), .B(n16698), .Z(n16696) );
  XOR U16493 ( .A(n16695), .B(n16699), .Z(n16697) );
  XNOR U16494 ( .A(n16700), .B(n16701), .Z(n16694) );
  NOR U16495 ( .A(n16702), .B(n16703), .Z(n16701) );
  XOR U16496 ( .A(n16700), .B(n16704), .Z(n16702) );
  XOR U16497 ( .A(n16630), .B(n16629), .Z(n16620) );
  XNOR U16498 ( .A(n16705), .B(n16626), .Z(n16629) );
  XOR U16499 ( .A(n16706), .B(n16707), .Z(n16626) );
  AND U16500 ( .A(n16708), .B(n16709), .Z(n16707) );
  XOR U16501 ( .A(n16706), .B(n16710), .Z(n16708) );
  XNOR U16502 ( .A(n16711), .B(n16712), .Z(n16705) );
  NOR U16503 ( .A(n16713), .B(n16714), .Z(n16712) );
  XNOR U16504 ( .A(n16711), .B(n16715), .Z(n16713) );
  XOR U16505 ( .A(n16716), .B(n16717), .Z(n16630) );
  NOR U16506 ( .A(n16718), .B(n16719), .Z(n16717) );
  XNOR U16507 ( .A(n16716), .B(n16720), .Z(n16718) );
  XNOR U16508 ( .A(n16529), .B(n16633), .Z(n16635) );
  XNOR U16509 ( .A(n16721), .B(n16722), .Z(n16529) );
  AND U16510 ( .A(n78), .B(n16536), .Z(n16722) );
  XOR U16511 ( .A(n16721), .B(n16534), .Z(n16536) );
  AND U16512 ( .A(n16537), .B(n16540), .Z(n16633) );
  XOR U16513 ( .A(n16723), .B(n16682), .Z(n16540) );
  XNOR U16514 ( .A(p_input[2048]), .B(p_input[32]), .Z(n16682) );
  XOR U16515 ( .A(n16659), .B(n16658), .Z(n16723) );
  XOR U16516 ( .A(n16724), .B(n16670), .Z(n16658) );
  XOR U16517 ( .A(n16644), .B(n16643), .Z(n16670) );
  XNOR U16518 ( .A(n16725), .B(n16649), .Z(n16643) );
  XOR U16519 ( .A(p_input[2072]), .B(p_input[56]), .Z(n16649) );
  XOR U16520 ( .A(n16640), .B(n16648), .Z(n16725) );
  XOR U16521 ( .A(n16726), .B(n16645), .Z(n16648) );
  XOR U16522 ( .A(p_input[2070]), .B(p_input[54]), .Z(n16645) );
  XNOR U16523 ( .A(p_input[2071]), .B(p_input[55]), .Z(n16726) );
  XNOR U16524 ( .A(n16727), .B(p_input[50]), .Z(n16640) );
  XNOR U16525 ( .A(n16654), .B(n16653), .Z(n16644) );
  XOR U16526 ( .A(n16728), .B(n16650), .Z(n16653) );
  XOR U16527 ( .A(p_input[2067]), .B(p_input[51]), .Z(n16650) );
  XNOR U16528 ( .A(p_input[2068]), .B(p_input[52]), .Z(n16728) );
  XOR U16529 ( .A(p_input[2069]), .B(p_input[53]), .Z(n16654) );
  XNOR U16530 ( .A(n16669), .B(n16655), .Z(n16724) );
  XNOR U16531 ( .A(n16729), .B(p_input[33]), .Z(n16655) );
  XNOR U16532 ( .A(n16730), .B(n16676), .Z(n16669) );
  XNOR U16533 ( .A(n16665), .B(n16664), .Z(n16676) );
  XOR U16534 ( .A(n16731), .B(n16661), .Z(n16664) );
  XNOR U16535 ( .A(n16444), .B(p_input[58]), .Z(n16661) );
  XNOR U16536 ( .A(p_input[2075]), .B(p_input[59]), .Z(n16731) );
  XOR U16537 ( .A(p_input[2076]), .B(p_input[60]), .Z(n16665) );
  XNOR U16538 ( .A(n16675), .B(n16666), .Z(n16730) );
  XNOR U16539 ( .A(n16732), .B(p_input[49]), .Z(n16666) );
  XOR U16540 ( .A(n16733), .B(n16681), .Z(n16675) );
  XNOR U16541 ( .A(p_input[2079]), .B(p_input[63]), .Z(n16681) );
  XOR U16542 ( .A(n16672), .B(n16680), .Z(n16733) );
  XOR U16543 ( .A(n16734), .B(n16677), .Z(n16680) );
  XOR U16544 ( .A(p_input[2077]), .B(p_input[61]), .Z(n16677) );
  XNOR U16545 ( .A(p_input[2078]), .B(p_input[62]), .Z(n16734) );
  XNOR U16546 ( .A(n16448), .B(p_input[57]), .Z(n16672) );
  XNOR U16547 ( .A(n16693), .B(n16692), .Z(n16659) );
  XNOR U16548 ( .A(n16735), .B(n16699), .Z(n16692) );
  XNOR U16549 ( .A(n16688), .B(n16687), .Z(n16699) );
  XOR U16550 ( .A(n16736), .B(n16684), .Z(n16687) );
  XNOR U16551 ( .A(n16737), .B(p_input[43]), .Z(n16684) );
  XNOR U16552 ( .A(p_input[2060]), .B(p_input[44]), .Z(n16736) );
  XOR U16553 ( .A(p_input[2061]), .B(p_input[45]), .Z(n16688) );
  XNOR U16554 ( .A(n16698), .B(n16689), .Z(n16735) );
  XNOR U16555 ( .A(n16452), .B(p_input[34]), .Z(n16689) );
  XOR U16556 ( .A(n16738), .B(n16704), .Z(n16698) );
  XNOR U16557 ( .A(p_input[2064]), .B(p_input[48]), .Z(n16704) );
  XOR U16558 ( .A(n16695), .B(n16703), .Z(n16738) );
  XOR U16559 ( .A(n16739), .B(n16700), .Z(n16703) );
  XOR U16560 ( .A(p_input[2062]), .B(p_input[46]), .Z(n16700) );
  XNOR U16561 ( .A(p_input[2063]), .B(p_input[47]), .Z(n16739) );
  XNOR U16562 ( .A(n16740), .B(p_input[42]), .Z(n16695) );
  XNOR U16563 ( .A(n16710), .B(n16709), .Z(n16693) );
  XNOR U16564 ( .A(n16741), .B(n16715), .Z(n16709) );
  XOR U16565 ( .A(p_input[2057]), .B(p_input[41]), .Z(n16715) );
  XOR U16566 ( .A(n16706), .B(n16714), .Z(n16741) );
  XOR U16567 ( .A(n16742), .B(n16711), .Z(n16714) );
  XOR U16568 ( .A(p_input[2055]), .B(p_input[39]), .Z(n16711) );
  XNOR U16569 ( .A(p_input[2056]), .B(p_input[40]), .Z(n16742) );
  XNOR U16570 ( .A(n16459), .B(p_input[35]), .Z(n16706) );
  XNOR U16571 ( .A(n16720), .B(n16719), .Z(n16710) );
  XOR U16572 ( .A(n16743), .B(n16716), .Z(n16719) );
  XOR U16573 ( .A(p_input[2052]), .B(p_input[36]), .Z(n16716) );
  XNOR U16574 ( .A(p_input[2053]), .B(p_input[37]), .Z(n16743) );
  XOR U16575 ( .A(p_input[2054]), .B(p_input[38]), .Z(n16720) );
  XNOR U16576 ( .A(n16744), .B(n16745), .Z(n16537) );
  AND U16577 ( .A(n78), .B(n16746), .Z(n16745) );
  XNOR U16578 ( .A(n16747), .B(n16748), .Z(n78) );
  AND U16579 ( .A(n16749), .B(n16750), .Z(n16748) );
  XOR U16580 ( .A(n16747), .B(n16547), .Z(n16750) );
  XNOR U16581 ( .A(n16747), .B(n16491), .Z(n16749) );
  XOR U16582 ( .A(n16751), .B(n16752), .Z(n16747) );
  AND U16583 ( .A(n16753), .B(n16754), .Z(n16752) );
  XNOR U16584 ( .A(n16560), .B(n16751), .Z(n16754) );
  XOR U16585 ( .A(n16751), .B(n16502), .Z(n16753) );
  XOR U16586 ( .A(n16755), .B(n16756), .Z(n16751) );
  AND U16587 ( .A(n16757), .B(n16758), .Z(n16756) );
  XNOR U16588 ( .A(n16585), .B(n16755), .Z(n16758) );
  XOR U16589 ( .A(n16755), .B(n16513), .Z(n16757) );
  XOR U16590 ( .A(n16759), .B(n16760), .Z(n16755) );
  AND U16591 ( .A(n16761), .B(n16762), .Z(n16760) );
  XOR U16592 ( .A(n16759), .B(n16522), .Z(n16761) );
  XOR U16593 ( .A(n16763), .B(n16764), .Z(n16480) );
  AND U16594 ( .A(n82), .B(n16746), .Z(n16764) );
  XNOR U16595 ( .A(n16744), .B(n16763), .Z(n16746) );
  XNOR U16596 ( .A(n16765), .B(n16766), .Z(n82) );
  AND U16597 ( .A(n16767), .B(n16768), .Z(n16766) );
  XNOR U16598 ( .A(n16769), .B(n16765), .Z(n16768) );
  IV U16599 ( .A(n16547), .Z(n16769) );
  XNOR U16600 ( .A(n16770), .B(n16771), .Z(n16547) );
  AND U16601 ( .A(n85), .B(n16772), .Z(n16771) );
  XNOR U16602 ( .A(n16770), .B(n16773), .Z(n16772) );
  XNOR U16603 ( .A(n16491), .B(n16765), .Z(n16767) );
  XOR U16604 ( .A(n16774), .B(n16775), .Z(n16491) );
  AND U16605 ( .A(n93), .B(n16776), .Z(n16775) );
  XOR U16606 ( .A(n16777), .B(n16778), .Z(n16765) );
  AND U16607 ( .A(n16779), .B(n16780), .Z(n16778) );
  XNOR U16608 ( .A(n16777), .B(n16560), .Z(n16780) );
  XNOR U16609 ( .A(n16781), .B(n16782), .Z(n16560) );
  AND U16610 ( .A(n85), .B(n16783), .Z(n16782) );
  XOR U16611 ( .A(n16784), .B(n16781), .Z(n16783) );
  XNOR U16612 ( .A(n16785), .B(n16777), .Z(n16779) );
  IV U16613 ( .A(n16502), .Z(n16785) );
  XOR U16614 ( .A(n16786), .B(n16787), .Z(n16502) );
  AND U16615 ( .A(n93), .B(n16788), .Z(n16787) );
  XOR U16616 ( .A(n16789), .B(n16790), .Z(n16777) );
  AND U16617 ( .A(n16791), .B(n16792), .Z(n16790) );
  XNOR U16618 ( .A(n16789), .B(n16585), .Z(n16792) );
  XNOR U16619 ( .A(n16793), .B(n16794), .Z(n16585) );
  AND U16620 ( .A(n85), .B(n16795), .Z(n16794) );
  XNOR U16621 ( .A(n16796), .B(n16793), .Z(n16795) );
  XOR U16622 ( .A(n16513), .B(n16789), .Z(n16791) );
  XOR U16623 ( .A(n16797), .B(n16798), .Z(n16513) );
  AND U16624 ( .A(n93), .B(n16799), .Z(n16798) );
  XOR U16625 ( .A(n16759), .B(n16800), .Z(n16789) );
  AND U16626 ( .A(n16801), .B(n16762), .Z(n16800) );
  XNOR U16627 ( .A(n16631), .B(n16759), .Z(n16762) );
  XNOR U16628 ( .A(n16802), .B(n16803), .Z(n16631) );
  AND U16629 ( .A(n85), .B(n16804), .Z(n16803) );
  XOR U16630 ( .A(n16805), .B(n16802), .Z(n16804) );
  XNOR U16631 ( .A(n16806), .B(n16759), .Z(n16801) );
  IV U16632 ( .A(n16522), .Z(n16806) );
  XOR U16633 ( .A(n16807), .B(n16808), .Z(n16522) );
  AND U16634 ( .A(n93), .B(n16809), .Z(n16808) );
  XOR U16635 ( .A(n16810), .B(n16811), .Z(n16759) );
  AND U16636 ( .A(n16812), .B(n16813), .Z(n16811) );
  XNOR U16637 ( .A(n16810), .B(n16721), .Z(n16813) );
  XNOR U16638 ( .A(n16814), .B(n16815), .Z(n16721) );
  AND U16639 ( .A(n85), .B(n16816), .Z(n16815) );
  XNOR U16640 ( .A(n16817), .B(n16814), .Z(n16816) );
  XNOR U16641 ( .A(n16818), .B(n16810), .Z(n16812) );
  IV U16642 ( .A(n16534), .Z(n16818) );
  XOR U16643 ( .A(n16819), .B(n16820), .Z(n16534) );
  AND U16644 ( .A(n93), .B(n16821), .Z(n16820) );
  AND U16645 ( .A(n16763), .B(n16744), .Z(n16810) );
  XNOR U16646 ( .A(n16822), .B(n16823), .Z(n16744) );
  AND U16647 ( .A(n85), .B(n16824), .Z(n16823) );
  XNOR U16648 ( .A(n16825), .B(n16822), .Z(n16824) );
  XNOR U16649 ( .A(n16826), .B(n16827), .Z(n85) );
  AND U16650 ( .A(n16828), .B(n16829), .Z(n16827) );
  XOR U16651 ( .A(n16773), .B(n16826), .Z(n16829) );
  AND U16652 ( .A(n16830), .B(n16831), .Z(n16773) );
  XOR U16653 ( .A(n16826), .B(n16770), .Z(n16828) );
  XNOR U16654 ( .A(n16832), .B(n16833), .Z(n16770) );
  AND U16655 ( .A(n89), .B(n16776), .Z(n16833) );
  XOR U16656 ( .A(n16774), .B(n16832), .Z(n16776) );
  XOR U16657 ( .A(n16834), .B(n16835), .Z(n16826) );
  AND U16658 ( .A(n16836), .B(n16837), .Z(n16835) );
  XNOR U16659 ( .A(n16834), .B(n16830), .Z(n16837) );
  IV U16660 ( .A(n16784), .Z(n16830) );
  XOR U16661 ( .A(n16838), .B(n16839), .Z(n16784) );
  XOR U16662 ( .A(n16840), .B(n16831), .Z(n16839) );
  AND U16663 ( .A(n16796), .B(n16841), .Z(n16831) );
  AND U16664 ( .A(n16842), .B(n16843), .Z(n16840) );
  XOR U16665 ( .A(n16844), .B(n16838), .Z(n16842) );
  XNOR U16666 ( .A(n16781), .B(n16834), .Z(n16836) );
  XNOR U16667 ( .A(n16845), .B(n16846), .Z(n16781) );
  AND U16668 ( .A(n89), .B(n16788), .Z(n16846) );
  XOR U16669 ( .A(n16845), .B(n16786), .Z(n16788) );
  XOR U16670 ( .A(n16847), .B(n16848), .Z(n16834) );
  AND U16671 ( .A(n16849), .B(n16850), .Z(n16848) );
  XNOR U16672 ( .A(n16847), .B(n16796), .Z(n16850) );
  XOR U16673 ( .A(n16851), .B(n16843), .Z(n16796) );
  XNOR U16674 ( .A(n16852), .B(n16838), .Z(n16843) );
  XOR U16675 ( .A(n16853), .B(n16854), .Z(n16838) );
  AND U16676 ( .A(n16855), .B(n16856), .Z(n16854) );
  XOR U16677 ( .A(n16857), .B(n16853), .Z(n16855) );
  XNOR U16678 ( .A(n16858), .B(n16859), .Z(n16852) );
  AND U16679 ( .A(n16860), .B(n16861), .Z(n16859) );
  XOR U16680 ( .A(n16858), .B(n16862), .Z(n16860) );
  XNOR U16681 ( .A(n16844), .B(n16841), .Z(n16851) );
  AND U16682 ( .A(n16863), .B(n16864), .Z(n16841) );
  XOR U16683 ( .A(n16865), .B(n16866), .Z(n16844) );
  AND U16684 ( .A(n16867), .B(n16868), .Z(n16866) );
  XOR U16685 ( .A(n16865), .B(n16869), .Z(n16867) );
  XNOR U16686 ( .A(n16793), .B(n16847), .Z(n16849) );
  XNOR U16687 ( .A(n16870), .B(n16871), .Z(n16793) );
  AND U16688 ( .A(n89), .B(n16799), .Z(n16871) );
  XOR U16689 ( .A(n16870), .B(n16797), .Z(n16799) );
  XOR U16690 ( .A(n16872), .B(n16873), .Z(n16847) );
  AND U16691 ( .A(n16874), .B(n16875), .Z(n16873) );
  XNOR U16692 ( .A(n16872), .B(n16863), .Z(n16875) );
  IV U16693 ( .A(n16805), .Z(n16863) );
  XNOR U16694 ( .A(n16876), .B(n16856), .Z(n16805) );
  XNOR U16695 ( .A(n16877), .B(n16862), .Z(n16856) );
  XOR U16696 ( .A(n16878), .B(n16879), .Z(n16862) );
  AND U16697 ( .A(n16880), .B(n16881), .Z(n16879) );
  XOR U16698 ( .A(n16878), .B(n16882), .Z(n16880) );
  XNOR U16699 ( .A(n16861), .B(n16853), .Z(n16877) );
  XOR U16700 ( .A(n16883), .B(n16884), .Z(n16853) );
  AND U16701 ( .A(n16885), .B(n16886), .Z(n16884) );
  XNOR U16702 ( .A(n16887), .B(n16883), .Z(n16885) );
  XNOR U16703 ( .A(n16888), .B(n16858), .Z(n16861) );
  XOR U16704 ( .A(n16889), .B(n16890), .Z(n16858) );
  AND U16705 ( .A(n16891), .B(n16892), .Z(n16890) );
  XOR U16706 ( .A(n16889), .B(n16893), .Z(n16891) );
  XNOR U16707 ( .A(n16894), .B(n16895), .Z(n16888) );
  AND U16708 ( .A(n16896), .B(n16897), .Z(n16895) );
  XNOR U16709 ( .A(n16894), .B(n16898), .Z(n16896) );
  XNOR U16710 ( .A(n16857), .B(n16864), .Z(n16876) );
  AND U16711 ( .A(n16817), .B(n16899), .Z(n16864) );
  XOR U16712 ( .A(n16869), .B(n16868), .Z(n16857) );
  XNOR U16713 ( .A(n16900), .B(n16865), .Z(n16868) );
  XOR U16714 ( .A(n16901), .B(n16902), .Z(n16865) );
  AND U16715 ( .A(n16903), .B(n16904), .Z(n16902) );
  XOR U16716 ( .A(n16901), .B(n16905), .Z(n16903) );
  XNOR U16717 ( .A(n16906), .B(n16907), .Z(n16900) );
  AND U16718 ( .A(n16908), .B(n16909), .Z(n16907) );
  XOR U16719 ( .A(n16906), .B(n16910), .Z(n16908) );
  XOR U16720 ( .A(n16911), .B(n16912), .Z(n16869) );
  AND U16721 ( .A(n16913), .B(n16914), .Z(n16912) );
  XOR U16722 ( .A(n16911), .B(n16915), .Z(n16913) );
  XNOR U16723 ( .A(n16802), .B(n16872), .Z(n16874) );
  XNOR U16724 ( .A(n16916), .B(n16917), .Z(n16802) );
  AND U16725 ( .A(n89), .B(n16809), .Z(n16917) );
  XOR U16726 ( .A(n16916), .B(n16807), .Z(n16809) );
  XOR U16727 ( .A(n16918), .B(n16919), .Z(n16872) );
  AND U16728 ( .A(n16920), .B(n16921), .Z(n16919) );
  XNOR U16729 ( .A(n16918), .B(n16817), .Z(n16921) );
  XOR U16730 ( .A(n16922), .B(n16886), .Z(n16817) );
  XNOR U16731 ( .A(n16923), .B(n16893), .Z(n16886) );
  XOR U16732 ( .A(n16882), .B(n16881), .Z(n16893) );
  XNOR U16733 ( .A(n16924), .B(n16878), .Z(n16881) );
  XOR U16734 ( .A(n16925), .B(n16926), .Z(n16878) );
  AND U16735 ( .A(n16927), .B(n16928), .Z(n16926) );
  XOR U16736 ( .A(n16925), .B(n16929), .Z(n16927) );
  XNOR U16737 ( .A(n16930), .B(n16931), .Z(n16924) );
  NOR U16738 ( .A(n16932), .B(n16933), .Z(n16931) );
  XNOR U16739 ( .A(n16930), .B(n16934), .Z(n16932) );
  XOR U16740 ( .A(n16935), .B(n16936), .Z(n16882) );
  NOR U16741 ( .A(n16937), .B(n16938), .Z(n16936) );
  XNOR U16742 ( .A(n16935), .B(n16939), .Z(n16937) );
  XNOR U16743 ( .A(n16892), .B(n16883), .Z(n16923) );
  XOR U16744 ( .A(n16940), .B(n16941), .Z(n16883) );
  NOR U16745 ( .A(n16942), .B(n16943), .Z(n16941) );
  XNOR U16746 ( .A(n16940), .B(n16944), .Z(n16942) );
  XOR U16747 ( .A(n16945), .B(n16898), .Z(n16892) );
  XNOR U16748 ( .A(n16946), .B(n16947), .Z(n16898) );
  NOR U16749 ( .A(n16948), .B(n16949), .Z(n16947) );
  XNOR U16750 ( .A(n16946), .B(n16950), .Z(n16948) );
  XNOR U16751 ( .A(n16897), .B(n16889), .Z(n16945) );
  XOR U16752 ( .A(n16951), .B(n16952), .Z(n16889) );
  AND U16753 ( .A(n16953), .B(n16954), .Z(n16952) );
  XOR U16754 ( .A(n16951), .B(n16955), .Z(n16953) );
  XNOR U16755 ( .A(n16956), .B(n16894), .Z(n16897) );
  XOR U16756 ( .A(n16957), .B(n16958), .Z(n16894) );
  AND U16757 ( .A(n16959), .B(n16960), .Z(n16958) );
  XOR U16758 ( .A(n16957), .B(n16961), .Z(n16959) );
  XNOR U16759 ( .A(n16962), .B(n16963), .Z(n16956) );
  NOR U16760 ( .A(n16964), .B(n16965), .Z(n16963) );
  XOR U16761 ( .A(n16962), .B(n16966), .Z(n16964) );
  XOR U16762 ( .A(n16887), .B(n16899), .Z(n16922) );
  NOR U16763 ( .A(n16825), .B(n16967), .Z(n16899) );
  XNOR U16764 ( .A(n16905), .B(n16904), .Z(n16887) );
  XNOR U16765 ( .A(n16968), .B(n16910), .Z(n16904) );
  XOR U16766 ( .A(n16969), .B(n16970), .Z(n16910) );
  NOR U16767 ( .A(n16971), .B(n16972), .Z(n16970) );
  XNOR U16768 ( .A(n16969), .B(n16973), .Z(n16971) );
  XNOR U16769 ( .A(n16909), .B(n16901), .Z(n16968) );
  XOR U16770 ( .A(n16974), .B(n16975), .Z(n16901) );
  AND U16771 ( .A(n16976), .B(n16977), .Z(n16975) );
  XNOR U16772 ( .A(n16974), .B(n16978), .Z(n16976) );
  XNOR U16773 ( .A(n16979), .B(n16906), .Z(n16909) );
  XOR U16774 ( .A(n16980), .B(n16981), .Z(n16906) );
  AND U16775 ( .A(n16982), .B(n16983), .Z(n16981) );
  XOR U16776 ( .A(n16980), .B(n16984), .Z(n16982) );
  XNOR U16777 ( .A(n16985), .B(n16986), .Z(n16979) );
  NOR U16778 ( .A(n16987), .B(n16988), .Z(n16986) );
  XOR U16779 ( .A(n16985), .B(n16989), .Z(n16987) );
  XOR U16780 ( .A(n16915), .B(n16914), .Z(n16905) );
  XNOR U16781 ( .A(n16990), .B(n16911), .Z(n16914) );
  XOR U16782 ( .A(n16991), .B(n16992), .Z(n16911) );
  AND U16783 ( .A(n16993), .B(n16994), .Z(n16992) );
  XOR U16784 ( .A(n16991), .B(n16995), .Z(n16993) );
  XNOR U16785 ( .A(n16996), .B(n16997), .Z(n16990) );
  NOR U16786 ( .A(n16998), .B(n16999), .Z(n16997) );
  XNOR U16787 ( .A(n16996), .B(n17000), .Z(n16998) );
  XOR U16788 ( .A(n17001), .B(n17002), .Z(n16915) );
  NOR U16789 ( .A(n17003), .B(n17004), .Z(n17002) );
  XNOR U16790 ( .A(n17001), .B(n17005), .Z(n17003) );
  XNOR U16791 ( .A(n16814), .B(n16918), .Z(n16920) );
  XNOR U16792 ( .A(n17006), .B(n17007), .Z(n16814) );
  AND U16793 ( .A(n89), .B(n16821), .Z(n17007) );
  XOR U16794 ( .A(n17006), .B(n16819), .Z(n16821) );
  AND U16795 ( .A(n16822), .B(n16825), .Z(n16918) );
  XOR U16796 ( .A(n17008), .B(n16967), .Z(n16825) );
  XNOR U16797 ( .A(p_input[2048]), .B(p_input[64]), .Z(n16967) );
  XOR U16798 ( .A(n16944), .B(n16943), .Z(n17008) );
  XOR U16799 ( .A(n17009), .B(n16955), .Z(n16943) );
  XOR U16800 ( .A(n16929), .B(n16928), .Z(n16955) );
  XNOR U16801 ( .A(n17010), .B(n16934), .Z(n16928) );
  XOR U16802 ( .A(p_input[2072]), .B(p_input[88]), .Z(n16934) );
  XOR U16803 ( .A(n16925), .B(n16933), .Z(n17010) );
  XOR U16804 ( .A(n17011), .B(n16930), .Z(n16933) );
  XOR U16805 ( .A(p_input[2070]), .B(p_input[86]), .Z(n16930) );
  XNOR U16806 ( .A(p_input[2071]), .B(p_input[87]), .Z(n17011) );
  XNOR U16807 ( .A(n16727), .B(p_input[82]), .Z(n16925) );
  XNOR U16808 ( .A(n16939), .B(n16938), .Z(n16929) );
  XOR U16809 ( .A(n17012), .B(n16935), .Z(n16938) );
  XOR U16810 ( .A(p_input[2067]), .B(p_input[83]), .Z(n16935) );
  XNOR U16811 ( .A(p_input[2068]), .B(p_input[84]), .Z(n17012) );
  XOR U16812 ( .A(p_input[2069]), .B(p_input[85]), .Z(n16939) );
  XNOR U16813 ( .A(n16954), .B(n16940), .Z(n17009) );
  XNOR U16814 ( .A(n16729), .B(p_input[65]), .Z(n16940) );
  XNOR U16815 ( .A(n17013), .B(n16961), .Z(n16954) );
  XNOR U16816 ( .A(n16950), .B(n16949), .Z(n16961) );
  XOR U16817 ( .A(n17014), .B(n16946), .Z(n16949) );
  XNOR U16818 ( .A(n16444), .B(p_input[90]), .Z(n16946) );
  XNOR U16819 ( .A(p_input[2075]), .B(p_input[91]), .Z(n17014) );
  XOR U16820 ( .A(p_input[2076]), .B(p_input[92]), .Z(n16950) );
  XNOR U16821 ( .A(n16960), .B(n16951), .Z(n17013) );
  XNOR U16822 ( .A(n16732), .B(p_input[81]), .Z(n16951) );
  XOR U16823 ( .A(n17015), .B(n16966), .Z(n16960) );
  XNOR U16824 ( .A(p_input[2079]), .B(p_input[95]), .Z(n16966) );
  XOR U16825 ( .A(n16957), .B(n16965), .Z(n17015) );
  XOR U16826 ( .A(n17016), .B(n16962), .Z(n16965) );
  XOR U16827 ( .A(p_input[2077]), .B(p_input[93]), .Z(n16962) );
  XNOR U16828 ( .A(p_input[2078]), .B(p_input[94]), .Z(n17016) );
  XNOR U16829 ( .A(n16448), .B(p_input[89]), .Z(n16957) );
  XNOR U16830 ( .A(n16978), .B(n16977), .Z(n16944) );
  XNOR U16831 ( .A(n17017), .B(n16984), .Z(n16977) );
  XNOR U16832 ( .A(n16973), .B(n16972), .Z(n16984) );
  XOR U16833 ( .A(n17018), .B(n16969), .Z(n16972) );
  XNOR U16834 ( .A(n16737), .B(p_input[75]), .Z(n16969) );
  XNOR U16835 ( .A(p_input[2060]), .B(p_input[76]), .Z(n17018) );
  XOR U16836 ( .A(p_input[2061]), .B(p_input[77]), .Z(n16973) );
  XNOR U16837 ( .A(n16983), .B(n16974), .Z(n17017) );
  XNOR U16838 ( .A(n16452), .B(p_input[66]), .Z(n16974) );
  XOR U16839 ( .A(n17019), .B(n16989), .Z(n16983) );
  XNOR U16840 ( .A(p_input[2064]), .B(p_input[80]), .Z(n16989) );
  XOR U16841 ( .A(n16980), .B(n16988), .Z(n17019) );
  XOR U16842 ( .A(n17020), .B(n16985), .Z(n16988) );
  XOR U16843 ( .A(p_input[2062]), .B(p_input[78]), .Z(n16985) );
  XNOR U16844 ( .A(p_input[2063]), .B(p_input[79]), .Z(n17020) );
  XNOR U16845 ( .A(n16740), .B(p_input[74]), .Z(n16980) );
  XNOR U16846 ( .A(n16995), .B(n16994), .Z(n16978) );
  XNOR U16847 ( .A(n17021), .B(n17000), .Z(n16994) );
  XOR U16848 ( .A(p_input[2057]), .B(p_input[73]), .Z(n17000) );
  XOR U16849 ( .A(n16991), .B(n16999), .Z(n17021) );
  XOR U16850 ( .A(n17022), .B(n16996), .Z(n16999) );
  XOR U16851 ( .A(p_input[2055]), .B(p_input[71]), .Z(n16996) );
  XNOR U16852 ( .A(p_input[2056]), .B(p_input[72]), .Z(n17022) );
  XNOR U16853 ( .A(n16459), .B(p_input[67]), .Z(n16991) );
  XNOR U16854 ( .A(n17005), .B(n17004), .Z(n16995) );
  XOR U16855 ( .A(n17023), .B(n17001), .Z(n17004) );
  XOR U16856 ( .A(p_input[2052]), .B(p_input[68]), .Z(n17001) );
  XNOR U16857 ( .A(p_input[2053]), .B(p_input[69]), .Z(n17023) );
  XOR U16858 ( .A(p_input[2054]), .B(p_input[70]), .Z(n17005) );
  XNOR U16859 ( .A(n17024), .B(n17025), .Z(n16822) );
  AND U16860 ( .A(n89), .B(n17026), .Z(n17025) );
  XNOR U16861 ( .A(n17027), .B(n17028), .Z(n89) );
  AND U16862 ( .A(n17029), .B(n17030), .Z(n17028) );
  XOR U16863 ( .A(n17027), .B(n16832), .Z(n17030) );
  XNOR U16864 ( .A(n17027), .B(n16774), .Z(n17029) );
  XOR U16865 ( .A(n17031), .B(n17032), .Z(n17027) );
  AND U16866 ( .A(n17033), .B(n17034), .Z(n17032) );
  XNOR U16867 ( .A(n16845), .B(n17031), .Z(n17034) );
  XOR U16868 ( .A(n17031), .B(n16786), .Z(n17033) );
  XOR U16869 ( .A(n17035), .B(n17036), .Z(n17031) );
  AND U16870 ( .A(n17037), .B(n17038), .Z(n17036) );
  XNOR U16871 ( .A(n16870), .B(n17035), .Z(n17038) );
  XOR U16872 ( .A(n17035), .B(n16797), .Z(n17037) );
  XOR U16873 ( .A(n17039), .B(n17040), .Z(n17035) );
  AND U16874 ( .A(n17041), .B(n17042), .Z(n17040) );
  XOR U16875 ( .A(n17039), .B(n16807), .Z(n17041) );
  XOR U16876 ( .A(n17043), .B(n17044), .Z(n16763) );
  AND U16877 ( .A(n93), .B(n17026), .Z(n17044) );
  XNOR U16878 ( .A(n17024), .B(n17043), .Z(n17026) );
  XNOR U16879 ( .A(n17045), .B(n17046), .Z(n93) );
  AND U16880 ( .A(n17047), .B(n17048), .Z(n17046) );
  XNOR U16881 ( .A(n17049), .B(n17045), .Z(n17048) );
  IV U16882 ( .A(n16832), .Z(n17049) );
  XNOR U16883 ( .A(n17050), .B(n17051), .Z(n16832) );
  AND U16884 ( .A(n96), .B(n17052), .Z(n17051) );
  XNOR U16885 ( .A(n17050), .B(n17053), .Z(n17052) );
  XNOR U16886 ( .A(n16774), .B(n17045), .Z(n17047) );
  XOR U16887 ( .A(n17054), .B(n17055), .Z(n16774) );
  AND U16888 ( .A(n104), .B(n17056), .Z(n17055) );
  XOR U16889 ( .A(n17057), .B(n17058), .Z(n17045) );
  AND U16890 ( .A(n17059), .B(n17060), .Z(n17058) );
  XNOR U16891 ( .A(n17057), .B(n16845), .Z(n17060) );
  XNOR U16892 ( .A(n17061), .B(n17062), .Z(n16845) );
  AND U16893 ( .A(n96), .B(n17063), .Z(n17062) );
  XOR U16894 ( .A(n17064), .B(n17061), .Z(n17063) );
  XNOR U16895 ( .A(n17065), .B(n17057), .Z(n17059) );
  IV U16896 ( .A(n16786), .Z(n17065) );
  XOR U16897 ( .A(n17066), .B(n17067), .Z(n16786) );
  AND U16898 ( .A(n104), .B(n17068), .Z(n17067) );
  XOR U16899 ( .A(n17069), .B(n17070), .Z(n17057) );
  AND U16900 ( .A(n17071), .B(n17072), .Z(n17070) );
  XNOR U16901 ( .A(n17069), .B(n16870), .Z(n17072) );
  XNOR U16902 ( .A(n17073), .B(n17074), .Z(n16870) );
  AND U16903 ( .A(n96), .B(n17075), .Z(n17074) );
  XNOR U16904 ( .A(n17076), .B(n17073), .Z(n17075) );
  XOR U16905 ( .A(n16797), .B(n17069), .Z(n17071) );
  XOR U16906 ( .A(n17077), .B(n17078), .Z(n16797) );
  AND U16907 ( .A(n104), .B(n17079), .Z(n17078) );
  XOR U16908 ( .A(n17039), .B(n17080), .Z(n17069) );
  AND U16909 ( .A(n17081), .B(n17042), .Z(n17080) );
  XNOR U16910 ( .A(n16916), .B(n17039), .Z(n17042) );
  XNOR U16911 ( .A(n17082), .B(n17083), .Z(n16916) );
  AND U16912 ( .A(n96), .B(n17084), .Z(n17083) );
  XOR U16913 ( .A(n17085), .B(n17082), .Z(n17084) );
  XNOR U16914 ( .A(n17086), .B(n17039), .Z(n17081) );
  IV U16915 ( .A(n16807), .Z(n17086) );
  XOR U16916 ( .A(n17087), .B(n17088), .Z(n16807) );
  AND U16917 ( .A(n104), .B(n17089), .Z(n17088) );
  XOR U16918 ( .A(n17090), .B(n17091), .Z(n17039) );
  AND U16919 ( .A(n17092), .B(n17093), .Z(n17091) );
  XNOR U16920 ( .A(n17090), .B(n17006), .Z(n17093) );
  XNOR U16921 ( .A(n17094), .B(n17095), .Z(n17006) );
  AND U16922 ( .A(n96), .B(n17096), .Z(n17095) );
  XNOR U16923 ( .A(n17097), .B(n17094), .Z(n17096) );
  XNOR U16924 ( .A(n17098), .B(n17090), .Z(n17092) );
  IV U16925 ( .A(n16819), .Z(n17098) );
  XOR U16926 ( .A(n17099), .B(n17100), .Z(n16819) );
  AND U16927 ( .A(n104), .B(n17101), .Z(n17100) );
  AND U16928 ( .A(n17043), .B(n17024), .Z(n17090) );
  XNOR U16929 ( .A(n17102), .B(n17103), .Z(n17024) );
  AND U16930 ( .A(n96), .B(n17104), .Z(n17103) );
  XNOR U16931 ( .A(n17105), .B(n17102), .Z(n17104) );
  XNOR U16932 ( .A(n17106), .B(n17107), .Z(n96) );
  AND U16933 ( .A(n17108), .B(n17109), .Z(n17107) );
  XOR U16934 ( .A(n17053), .B(n17106), .Z(n17109) );
  AND U16935 ( .A(n17110), .B(n17111), .Z(n17053) );
  XOR U16936 ( .A(n17106), .B(n17050), .Z(n17108) );
  XNOR U16937 ( .A(n17112), .B(n17113), .Z(n17050) );
  AND U16938 ( .A(n100), .B(n17056), .Z(n17113) );
  XOR U16939 ( .A(n17054), .B(n17112), .Z(n17056) );
  XOR U16940 ( .A(n17114), .B(n17115), .Z(n17106) );
  AND U16941 ( .A(n17116), .B(n17117), .Z(n17115) );
  XNOR U16942 ( .A(n17114), .B(n17110), .Z(n17117) );
  IV U16943 ( .A(n17064), .Z(n17110) );
  XOR U16944 ( .A(n17118), .B(n17119), .Z(n17064) );
  XOR U16945 ( .A(n17120), .B(n17111), .Z(n17119) );
  AND U16946 ( .A(n17076), .B(n17121), .Z(n17111) );
  AND U16947 ( .A(n17122), .B(n17123), .Z(n17120) );
  XOR U16948 ( .A(n17124), .B(n17118), .Z(n17122) );
  XNOR U16949 ( .A(n17061), .B(n17114), .Z(n17116) );
  XNOR U16950 ( .A(n17125), .B(n17126), .Z(n17061) );
  AND U16951 ( .A(n100), .B(n17068), .Z(n17126) );
  XOR U16952 ( .A(n17125), .B(n17066), .Z(n17068) );
  XOR U16953 ( .A(n17127), .B(n17128), .Z(n17114) );
  AND U16954 ( .A(n17129), .B(n17130), .Z(n17128) );
  XNOR U16955 ( .A(n17127), .B(n17076), .Z(n17130) );
  XOR U16956 ( .A(n17131), .B(n17123), .Z(n17076) );
  XNOR U16957 ( .A(n17132), .B(n17118), .Z(n17123) );
  XOR U16958 ( .A(n17133), .B(n17134), .Z(n17118) );
  AND U16959 ( .A(n17135), .B(n17136), .Z(n17134) );
  XOR U16960 ( .A(n17137), .B(n17133), .Z(n17135) );
  XNOR U16961 ( .A(n17138), .B(n17139), .Z(n17132) );
  AND U16962 ( .A(n17140), .B(n17141), .Z(n17139) );
  XOR U16963 ( .A(n17138), .B(n17142), .Z(n17140) );
  XNOR U16964 ( .A(n17124), .B(n17121), .Z(n17131) );
  AND U16965 ( .A(n17143), .B(n17144), .Z(n17121) );
  XOR U16966 ( .A(n17145), .B(n17146), .Z(n17124) );
  AND U16967 ( .A(n17147), .B(n17148), .Z(n17146) );
  XOR U16968 ( .A(n17145), .B(n17149), .Z(n17147) );
  XNOR U16969 ( .A(n17073), .B(n17127), .Z(n17129) );
  XNOR U16970 ( .A(n17150), .B(n17151), .Z(n17073) );
  AND U16971 ( .A(n100), .B(n17079), .Z(n17151) );
  XOR U16972 ( .A(n17150), .B(n17077), .Z(n17079) );
  XOR U16973 ( .A(n17152), .B(n17153), .Z(n17127) );
  AND U16974 ( .A(n17154), .B(n17155), .Z(n17153) );
  XNOR U16975 ( .A(n17152), .B(n17143), .Z(n17155) );
  IV U16976 ( .A(n17085), .Z(n17143) );
  XNOR U16977 ( .A(n17156), .B(n17136), .Z(n17085) );
  XNOR U16978 ( .A(n17157), .B(n17142), .Z(n17136) );
  XOR U16979 ( .A(n17158), .B(n17159), .Z(n17142) );
  AND U16980 ( .A(n17160), .B(n17161), .Z(n17159) );
  XOR U16981 ( .A(n17158), .B(n17162), .Z(n17160) );
  XNOR U16982 ( .A(n17141), .B(n17133), .Z(n17157) );
  XOR U16983 ( .A(n17163), .B(n17164), .Z(n17133) );
  AND U16984 ( .A(n17165), .B(n17166), .Z(n17164) );
  XNOR U16985 ( .A(n17167), .B(n17163), .Z(n17165) );
  XNOR U16986 ( .A(n17168), .B(n17138), .Z(n17141) );
  XOR U16987 ( .A(n17169), .B(n17170), .Z(n17138) );
  AND U16988 ( .A(n17171), .B(n17172), .Z(n17170) );
  XOR U16989 ( .A(n17169), .B(n17173), .Z(n17171) );
  XNOR U16990 ( .A(n17174), .B(n17175), .Z(n17168) );
  AND U16991 ( .A(n17176), .B(n17177), .Z(n17175) );
  XNOR U16992 ( .A(n17174), .B(n17178), .Z(n17176) );
  XNOR U16993 ( .A(n17137), .B(n17144), .Z(n17156) );
  AND U16994 ( .A(n17097), .B(n17179), .Z(n17144) );
  XOR U16995 ( .A(n17149), .B(n17148), .Z(n17137) );
  XNOR U16996 ( .A(n17180), .B(n17145), .Z(n17148) );
  XOR U16997 ( .A(n17181), .B(n17182), .Z(n17145) );
  AND U16998 ( .A(n17183), .B(n17184), .Z(n17182) );
  XOR U16999 ( .A(n17181), .B(n17185), .Z(n17183) );
  XNOR U17000 ( .A(n17186), .B(n17187), .Z(n17180) );
  AND U17001 ( .A(n17188), .B(n17189), .Z(n17187) );
  XOR U17002 ( .A(n17186), .B(n17190), .Z(n17188) );
  XOR U17003 ( .A(n17191), .B(n17192), .Z(n17149) );
  AND U17004 ( .A(n17193), .B(n17194), .Z(n17192) );
  XOR U17005 ( .A(n17191), .B(n17195), .Z(n17193) );
  XNOR U17006 ( .A(n17082), .B(n17152), .Z(n17154) );
  XNOR U17007 ( .A(n17196), .B(n17197), .Z(n17082) );
  AND U17008 ( .A(n100), .B(n17089), .Z(n17197) );
  XOR U17009 ( .A(n17196), .B(n17087), .Z(n17089) );
  XOR U17010 ( .A(n17198), .B(n17199), .Z(n17152) );
  AND U17011 ( .A(n17200), .B(n17201), .Z(n17199) );
  XNOR U17012 ( .A(n17198), .B(n17097), .Z(n17201) );
  XOR U17013 ( .A(n17202), .B(n17166), .Z(n17097) );
  XNOR U17014 ( .A(n17203), .B(n17173), .Z(n17166) );
  XOR U17015 ( .A(n17162), .B(n17161), .Z(n17173) );
  XNOR U17016 ( .A(n17204), .B(n17158), .Z(n17161) );
  XOR U17017 ( .A(n17205), .B(n17206), .Z(n17158) );
  AND U17018 ( .A(n17207), .B(n17208), .Z(n17206) );
  XNOR U17019 ( .A(n17209), .B(n17210), .Z(n17207) );
  IV U17020 ( .A(n17205), .Z(n17209) );
  XNOR U17021 ( .A(n17211), .B(n17212), .Z(n17204) );
  NOR U17022 ( .A(n17213), .B(n17214), .Z(n17212) );
  XNOR U17023 ( .A(n17211), .B(n17215), .Z(n17213) );
  XOR U17024 ( .A(n17216), .B(n17217), .Z(n17162) );
  NOR U17025 ( .A(n17218), .B(n17219), .Z(n17217) );
  XNOR U17026 ( .A(n17216), .B(n17220), .Z(n17218) );
  XNOR U17027 ( .A(n17172), .B(n17163), .Z(n17203) );
  XOR U17028 ( .A(n17221), .B(n17222), .Z(n17163) );
  AND U17029 ( .A(n17223), .B(n17224), .Z(n17222) );
  XOR U17030 ( .A(n17221), .B(n17225), .Z(n17223) );
  XOR U17031 ( .A(n17226), .B(n17178), .Z(n17172) );
  XOR U17032 ( .A(n17227), .B(n17228), .Z(n17178) );
  NOR U17033 ( .A(n17229), .B(n17230), .Z(n17228) );
  XOR U17034 ( .A(n17227), .B(n17231), .Z(n17229) );
  XNOR U17035 ( .A(n17177), .B(n17169), .Z(n17226) );
  XOR U17036 ( .A(n17232), .B(n17233), .Z(n17169) );
  AND U17037 ( .A(n17234), .B(n17235), .Z(n17233) );
  XOR U17038 ( .A(n17232), .B(n17236), .Z(n17234) );
  XNOR U17039 ( .A(n17237), .B(n17174), .Z(n17177) );
  XOR U17040 ( .A(n17238), .B(n17239), .Z(n17174) );
  AND U17041 ( .A(n17240), .B(n17241), .Z(n17239) );
  XNOR U17042 ( .A(n17242), .B(n17243), .Z(n17240) );
  IV U17043 ( .A(n17238), .Z(n17242) );
  XNOR U17044 ( .A(n17244), .B(n17245), .Z(n17237) );
  NOR U17045 ( .A(n17246), .B(n17247), .Z(n17245) );
  XNOR U17046 ( .A(n17244), .B(n17248), .Z(n17246) );
  XOR U17047 ( .A(n17167), .B(n17179), .Z(n17202) );
  NOR U17048 ( .A(n17105), .B(n17249), .Z(n17179) );
  XNOR U17049 ( .A(n17185), .B(n17184), .Z(n17167) );
  XNOR U17050 ( .A(n17250), .B(n17190), .Z(n17184) );
  XNOR U17051 ( .A(n17251), .B(n17252), .Z(n17190) );
  NOR U17052 ( .A(n17253), .B(n17254), .Z(n17252) );
  XOR U17053 ( .A(n17251), .B(n17255), .Z(n17253) );
  XNOR U17054 ( .A(n17189), .B(n17181), .Z(n17250) );
  XOR U17055 ( .A(n17256), .B(n17257), .Z(n17181) );
  AND U17056 ( .A(n17258), .B(n17259), .Z(n17257) );
  XOR U17057 ( .A(n17256), .B(n17260), .Z(n17258) );
  XNOR U17058 ( .A(n17261), .B(n17186), .Z(n17189) );
  XOR U17059 ( .A(n17262), .B(n17263), .Z(n17186) );
  AND U17060 ( .A(n17264), .B(n17265), .Z(n17263) );
  XNOR U17061 ( .A(n17266), .B(n17267), .Z(n17264) );
  IV U17062 ( .A(n17262), .Z(n17266) );
  XNOR U17063 ( .A(n17268), .B(n17269), .Z(n17261) );
  NOR U17064 ( .A(n17270), .B(n17271), .Z(n17269) );
  XNOR U17065 ( .A(n17268), .B(n17272), .Z(n17270) );
  XOR U17066 ( .A(n17195), .B(n17194), .Z(n17185) );
  XNOR U17067 ( .A(n17273), .B(n17191), .Z(n17194) );
  XOR U17068 ( .A(n17274), .B(n17275), .Z(n17191) );
  AND U17069 ( .A(n17276), .B(n17277), .Z(n17275) );
  XOR U17070 ( .A(n17274), .B(n17278), .Z(n17276) );
  XNOR U17071 ( .A(n17279), .B(n17280), .Z(n17273) );
  NOR U17072 ( .A(n17281), .B(n17282), .Z(n17280) );
  XNOR U17073 ( .A(n17279), .B(n17283), .Z(n17281) );
  XOR U17074 ( .A(n17284), .B(n17285), .Z(n17195) );
  NOR U17075 ( .A(n17286), .B(n17287), .Z(n17285) );
  XNOR U17076 ( .A(n17284), .B(n17288), .Z(n17286) );
  XNOR U17077 ( .A(n17094), .B(n17198), .Z(n17200) );
  XNOR U17078 ( .A(n17289), .B(n17290), .Z(n17094) );
  AND U17079 ( .A(n100), .B(n17101), .Z(n17290) );
  XOR U17080 ( .A(n17289), .B(n17099), .Z(n17101) );
  AND U17081 ( .A(n17102), .B(n17105), .Z(n17198) );
  XOR U17082 ( .A(n17291), .B(n17249), .Z(n17105) );
  XNOR U17083 ( .A(p_input[2048]), .B(p_input[96]), .Z(n17249) );
  XNOR U17084 ( .A(n17225), .B(n17224), .Z(n17291) );
  XNOR U17085 ( .A(n17292), .B(n17236), .Z(n17224) );
  XOR U17086 ( .A(n17210), .B(n17208), .Z(n17236) );
  XNOR U17087 ( .A(n17293), .B(n17215), .Z(n17208) );
  XOR U17088 ( .A(p_input[120]), .B(p_input[2072]), .Z(n17215) );
  XOR U17089 ( .A(n17205), .B(n17214), .Z(n17293) );
  XOR U17090 ( .A(n17294), .B(n17211), .Z(n17214) );
  XOR U17091 ( .A(p_input[118]), .B(p_input[2070]), .Z(n17211) );
  XOR U17092 ( .A(p_input[119]), .B(n17295), .Z(n17294) );
  XOR U17093 ( .A(p_input[114]), .B(p_input[2066]), .Z(n17205) );
  XNOR U17094 ( .A(n17220), .B(n17219), .Z(n17210) );
  XOR U17095 ( .A(n17296), .B(n17216), .Z(n17219) );
  XOR U17096 ( .A(p_input[115]), .B(p_input[2067]), .Z(n17216) );
  XOR U17097 ( .A(p_input[116]), .B(n17297), .Z(n17296) );
  XOR U17098 ( .A(p_input[117]), .B(p_input[2069]), .Z(n17220) );
  XNOR U17099 ( .A(n17235), .B(n17221), .Z(n17292) );
  XNOR U17100 ( .A(n16729), .B(p_input[97]), .Z(n17221) );
  XNOR U17101 ( .A(n17298), .B(n17243), .Z(n17235) );
  XNOR U17102 ( .A(n17231), .B(n17230), .Z(n17243) );
  XNOR U17103 ( .A(n17299), .B(n17227), .Z(n17230) );
  XNOR U17104 ( .A(p_input[122]), .B(p_input[2074]), .Z(n17227) );
  XOR U17105 ( .A(p_input[123]), .B(n17300), .Z(n17299) );
  XOR U17106 ( .A(p_input[124]), .B(p_input[2076]), .Z(n17231) );
  XOR U17107 ( .A(n17241), .B(n17301), .Z(n17298) );
  IV U17108 ( .A(n17232), .Z(n17301) );
  XOR U17109 ( .A(p_input[113]), .B(p_input[2065]), .Z(n17232) );
  XNOR U17110 ( .A(n17302), .B(n17248), .Z(n17241) );
  XNOR U17111 ( .A(p_input[127]), .B(n17303), .Z(n17248) );
  XOR U17112 ( .A(n17238), .B(n17247), .Z(n17302) );
  XOR U17113 ( .A(n17304), .B(n17244), .Z(n17247) );
  XOR U17114 ( .A(p_input[125]), .B(p_input[2077]), .Z(n17244) );
  XOR U17115 ( .A(p_input[126]), .B(n17305), .Z(n17304) );
  XOR U17116 ( .A(p_input[121]), .B(p_input[2073]), .Z(n17238) );
  XOR U17117 ( .A(n17260), .B(n17259), .Z(n17225) );
  XNOR U17118 ( .A(n17306), .B(n17267), .Z(n17259) );
  XNOR U17119 ( .A(n17255), .B(n17254), .Z(n17267) );
  XNOR U17120 ( .A(n17307), .B(n17251), .Z(n17254) );
  XNOR U17121 ( .A(p_input[107]), .B(p_input[2059]), .Z(n17251) );
  XOR U17122 ( .A(p_input[108]), .B(n16451), .Z(n17307) );
  XOR U17123 ( .A(p_input[109]), .B(p_input[2061]), .Z(n17255) );
  XNOR U17124 ( .A(n17265), .B(n17256), .Z(n17306) );
  XNOR U17125 ( .A(n16452), .B(p_input[98]), .Z(n17256) );
  XNOR U17126 ( .A(n17308), .B(n17272), .Z(n17265) );
  XNOR U17127 ( .A(p_input[112]), .B(n16454), .Z(n17272) );
  XOR U17128 ( .A(n17262), .B(n17271), .Z(n17308) );
  XOR U17129 ( .A(n17309), .B(n17268), .Z(n17271) );
  XOR U17130 ( .A(p_input[110]), .B(p_input[2062]), .Z(n17268) );
  XOR U17131 ( .A(p_input[111]), .B(n16456), .Z(n17309) );
  XOR U17132 ( .A(p_input[106]), .B(p_input[2058]), .Z(n17262) );
  XOR U17133 ( .A(n17278), .B(n17277), .Z(n17260) );
  XNOR U17134 ( .A(n17310), .B(n17283), .Z(n17277) );
  XOR U17135 ( .A(p_input[105]), .B(p_input[2057]), .Z(n17283) );
  XOR U17136 ( .A(n17274), .B(n17282), .Z(n17310) );
  XOR U17137 ( .A(n17311), .B(n17279), .Z(n17282) );
  XOR U17138 ( .A(p_input[103]), .B(p_input[2055]), .Z(n17279) );
  XOR U17139 ( .A(p_input[104]), .B(n17312), .Z(n17311) );
  XNOR U17140 ( .A(n16459), .B(p_input[99]), .Z(n17274) );
  XNOR U17141 ( .A(n17288), .B(n17287), .Z(n17278) );
  XOR U17142 ( .A(n17313), .B(n17284), .Z(n17287) );
  XOR U17143 ( .A(p_input[100]), .B(p_input[2052]), .Z(n17284) );
  XOR U17144 ( .A(p_input[101]), .B(n17314), .Z(n17313) );
  XOR U17145 ( .A(p_input[102]), .B(p_input[2054]), .Z(n17288) );
  XNOR U17146 ( .A(n17315), .B(n17316), .Z(n17102) );
  AND U17147 ( .A(n100), .B(n17317), .Z(n17316) );
  XNOR U17148 ( .A(n17318), .B(n17319), .Z(n100) );
  AND U17149 ( .A(n17320), .B(n17321), .Z(n17319) );
  XOR U17150 ( .A(n17318), .B(n17112), .Z(n17321) );
  XNOR U17151 ( .A(n17318), .B(n17054), .Z(n17320) );
  XOR U17152 ( .A(n17322), .B(n17323), .Z(n17318) );
  AND U17153 ( .A(n17324), .B(n17325), .Z(n17323) );
  XNOR U17154 ( .A(n17125), .B(n17322), .Z(n17325) );
  XOR U17155 ( .A(n17322), .B(n17066), .Z(n17324) );
  XOR U17156 ( .A(n17326), .B(n17327), .Z(n17322) );
  AND U17157 ( .A(n17328), .B(n17329), .Z(n17327) );
  XNOR U17158 ( .A(n17150), .B(n17326), .Z(n17329) );
  XOR U17159 ( .A(n17326), .B(n17077), .Z(n17328) );
  XOR U17160 ( .A(n17330), .B(n17331), .Z(n17326) );
  AND U17161 ( .A(n17332), .B(n17333), .Z(n17331) );
  XOR U17162 ( .A(n17330), .B(n17087), .Z(n17332) );
  XOR U17163 ( .A(n17334), .B(n17335), .Z(n17043) );
  AND U17164 ( .A(n104), .B(n17317), .Z(n17335) );
  XNOR U17165 ( .A(n17315), .B(n17334), .Z(n17317) );
  XNOR U17166 ( .A(n17336), .B(n17337), .Z(n104) );
  AND U17167 ( .A(n17338), .B(n17339), .Z(n17337) );
  XNOR U17168 ( .A(n17340), .B(n17336), .Z(n17339) );
  IV U17169 ( .A(n17112), .Z(n17340) );
  XNOR U17170 ( .A(n17341), .B(n17342), .Z(n17112) );
  AND U17171 ( .A(n107), .B(n17343), .Z(n17342) );
  XNOR U17172 ( .A(n17341), .B(n17344), .Z(n17343) );
  XNOR U17173 ( .A(n17054), .B(n17336), .Z(n17338) );
  XOR U17174 ( .A(n17345), .B(n17346), .Z(n17054) );
  AND U17175 ( .A(n115), .B(n17347), .Z(n17346) );
  XOR U17176 ( .A(n17348), .B(n17349), .Z(n17336) );
  AND U17177 ( .A(n17350), .B(n17351), .Z(n17349) );
  XNOR U17178 ( .A(n17348), .B(n17125), .Z(n17351) );
  XNOR U17179 ( .A(n17352), .B(n17353), .Z(n17125) );
  AND U17180 ( .A(n107), .B(n17354), .Z(n17353) );
  XOR U17181 ( .A(n17355), .B(n17352), .Z(n17354) );
  XNOR U17182 ( .A(n17356), .B(n17348), .Z(n17350) );
  IV U17183 ( .A(n17066), .Z(n17356) );
  XOR U17184 ( .A(n17357), .B(n17358), .Z(n17066) );
  AND U17185 ( .A(n115), .B(n17359), .Z(n17358) );
  XOR U17186 ( .A(n17360), .B(n17361), .Z(n17348) );
  AND U17187 ( .A(n17362), .B(n17363), .Z(n17361) );
  XNOR U17188 ( .A(n17360), .B(n17150), .Z(n17363) );
  XNOR U17189 ( .A(n17364), .B(n17365), .Z(n17150) );
  AND U17190 ( .A(n107), .B(n17366), .Z(n17365) );
  XNOR U17191 ( .A(n17367), .B(n17364), .Z(n17366) );
  XOR U17192 ( .A(n17077), .B(n17360), .Z(n17362) );
  XOR U17193 ( .A(n17368), .B(n17369), .Z(n17077) );
  AND U17194 ( .A(n115), .B(n17370), .Z(n17369) );
  XOR U17195 ( .A(n17330), .B(n17371), .Z(n17360) );
  AND U17196 ( .A(n17372), .B(n17333), .Z(n17371) );
  XNOR U17197 ( .A(n17196), .B(n17330), .Z(n17333) );
  XNOR U17198 ( .A(n17373), .B(n17374), .Z(n17196) );
  AND U17199 ( .A(n107), .B(n17375), .Z(n17374) );
  XOR U17200 ( .A(n17376), .B(n17373), .Z(n17375) );
  XNOR U17201 ( .A(n17377), .B(n17330), .Z(n17372) );
  IV U17202 ( .A(n17087), .Z(n17377) );
  XOR U17203 ( .A(n17378), .B(n17379), .Z(n17087) );
  AND U17204 ( .A(n115), .B(n17380), .Z(n17379) );
  XOR U17205 ( .A(n17381), .B(n17382), .Z(n17330) );
  AND U17206 ( .A(n17383), .B(n17384), .Z(n17382) );
  XNOR U17207 ( .A(n17381), .B(n17289), .Z(n17384) );
  XNOR U17208 ( .A(n17385), .B(n17386), .Z(n17289) );
  AND U17209 ( .A(n107), .B(n17387), .Z(n17386) );
  XNOR U17210 ( .A(n17388), .B(n17385), .Z(n17387) );
  XNOR U17211 ( .A(n17389), .B(n17381), .Z(n17383) );
  IV U17212 ( .A(n17099), .Z(n17389) );
  XOR U17213 ( .A(n17390), .B(n17391), .Z(n17099) );
  AND U17214 ( .A(n115), .B(n17392), .Z(n17391) );
  AND U17215 ( .A(n17334), .B(n17315), .Z(n17381) );
  XNOR U17216 ( .A(n17393), .B(n17394), .Z(n17315) );
  AND U17217 ( .A(n107), .B(n17395), .Z(n17394) );
  XNOR U17218 ( .A(n17396), .B(n17393), .Z(n17395) );
  XNOR U17219 ( .A(n17397), .B(n17398), .Z(n107) );
  AND U17220 ( .A(n17399), .B(n17400), .Z(n17398) );
  XOR U17221 ( .A(n17344), .B(n17397), .Z(n17400) );
  AND U17222 ( .A(n17401), .B(n17402), .Z(n17344) );
  XOR U17223 ( .A(n17397), .B(n17341), .Z(n17399) );
  XNOR U17224 ( .A(n17403), .B(n17404), .Z(n17341) );
  AND U17225 ( .A(n111), .B(n17347), .Z(n17404) );
  XOR U17226 ( .A(n17345), .B(n17403), .Z(n17347) );
  XOR U17227 ( .A(n17405), .B(n17406), .Z(n17397) );
  AND U17228 ( .A(n17407), .B(n17408), .Z(n17406) );
  XNOR U17229 ( .A(n17405), .B(n17401), .Z(n17408) );
  IV U17230 ( .A(n17355), .Z(n17401) );
  XOR U17231 ( .A(n17409), .B(n17410), .Z(n17355) );
  XOR U17232 ( .A(n17411), .B(n17402), .Z(n17410) );
  AND U17233 ( .A(n17367), .B(n17412), .Z(n17402) );
  AND U17234 ( .A(n17413), .B(n17414), .Z(n17411) );
  XOR U17235 ( .A(n17415), .B(n17409), .Z(n17413) );
  XNOR U17236 ( .A(n17352), .B(n17405), .Z(n17407) );
  XNOR U17237 ( .A(n17416), .B(n17417), .Z(n17352) );
  AND U17238 ( .A(n111), .B(n17359), .Z(n17417) );
  XOR U17239 ( .A(n17416), .B(n17357), .Z(n17359) );
  XOR U17240 ( .A(n17418), .B(n17419), .Z(n17405) );
  AND U17241 ( .A(n17420), .B(n17421), .Z(n17419) );
  XNOR U17242 ( .A(n17418), .B(n17367), .Z(n17421) );
  XOR U17243 ( .A(n17422), .B(n17414), .Z(n17367) );
  XNOR U17244 ( .A(n17423), .B(n17409), .Z(n17414) );
  XOR U17245 ( .A(n17424), .B(n17425), .Z(n17409) );
  AND U17246 ( .A(n17426), .B(n17427), .Z(n17425) );
  XOR U17247 ( .A(n17428), .B(n17424), .Z(n17426) );
  XNOR U17248 ( .A(n17429), .B(n17430), .Z(n17423) );
  AND U17249 ( .A(n17431), .B(n17432), .Z(n17430) );
  XOR U17250 ( .A(n17429), .B(n17433), .Z(n17431) );
  XNOR U17251 ( .A(n17415), .B(n17412), .Z(n17422) );
  AND U17252 ( .A(n17434), .B(n17435), .Z(n17412) );
  XOR U17253 ( .A(n17436), .B(n17437), .Z(n17415) );
  AND U17254 ( .A(n17438), .B(n17439), .Z(n17437) );
  XOR U17255 ( .A(n17436), .B(n17440), .Z(n17438) );
  XNOR U17256 ( .A(n17364), .B(n17418), .Z(n17420) );
  XNOR U17257 ( .A(n17441), .B(n17442), .Z(n17364) );
  AND U17258 ( .A(n111), .B(n17370), .Z(n17442) );
  XOR U17259 ( .A(n17441), .B(n17368), .Z(n17370) );
  XOR U17260 ( .A(n17443), .B(n17444), .Z(n17418) );
  AND U17261 ( .A(n17445), .B(n17446), .Z(n17444) );
  XNOR U17262 ( .A(n17443), .B(n17434), .Z(n17446) );
  IV U17263 ( .A(n17376), .Z(n17434) );
  XNOR U17264 ( .A(n17447), .B(n17427), .Z(n17376) );
  XNOR U17265 ( .A(n17448), .B(n17433), .Z(n17427) );
  XOR U17266 ( .A(n17449), .B(n17450), .Z(n17433) );
  AND U17267 ( .A(n17451), .B(n17452), .Z(n17450) );
  XOR U17268 ( .A(n17449), .B(n17453), .Z(n17451) );
  XNOR U17269 ( .A(n17432), .B(n17424), .Z(n17448) );
  XOR U17270 ( .A(n17454), .B(n17455), .Z(n17424) );
  AND U17271 ( .A(n17456), .B(n17457), .Z(n17455) );
  XNOR U17272 ( .A(n17458), .B(n17454), .Z(n17456) );
  XNOR U17273 ( .A(n17459), .B(n17429), .Z(n17432) );
  XOR U17274 ( .A(n17460), .B(n17461), .Z(n17429) );
  AND U17275 ( .A(n17462), .B(n17463), .Z(n17461) );
  XOR U17276 ( .A(n17460), .B(n17464), .Z(n17462) );
  XNOR U17277 ( .A(n17465), .B(n17466), .Z(n17459) );
  AND U17278 ( .A(n17467), .B(n17468), .Z(n17466) );
  XNOR U17279 ( .A(n17465), .B(n17469), .Z(n17467) );
  XNOR U17280 ( .A(n17428), .B(n17435), .Z(n17447) );
  AND U17281 ( .A(n17388), .B(n17470), .Z(n17435) );
  XOR U17282 ( .A(n17440), .B(n17439), .Z(n17428) );
  XNOR U17283 ( .A(n17471), .B(n17436), .Z(n17439) );
  XOR U17284 ( .A(n17472), .B(n17473), .Z(n17436) );
  AND U17285 ( .A(n17474), .B(n17475), .Z(n17473) );
  XOR U17286 ( .A(n17472), .B(n17476), .Z(n17474) );
  XNOR U17287 ( .A(n17477), .B(n17478), .Z(n17471) );
  AND U17288 ( .A(n17479), .B(n17480), .Z(n17478) );
  XOR U17289 ( .A(n17477), .B(n17481), .Z(n17479) );
  XOR U17290 ( .A(n17482), .B(n17483), .Z(n17440) );
  AND U17291 ( .A(n17484), .B(n17485), .Z(n17483) );
  XOR U17292 ( .A(n17482), .B(n17486), .Z(n17484) );
  XNOR U17293 ( .A(n17373), .B(n17443), .Z(n17445) );
  XNOR U17294 ( .A(n17487), .B(n17488), .Z(n17373) );
  AND U17295 ( .A(n111), .B(n17380), .Z(n17488) );
  XOR U17296 ( .A(n17487), .B(n17378), .Z(n17380) );
  XOR U17297 ( .A(n17489), .B(n17490), .Z(n17443) );
  AND U17298 ( .A(n17491), .B(n17492), .Z(n17490) );
  XNOR U17299 ( .A(n17489), .B(n17388), .Z(n17492) );
  XOR U17300 ( .A(n17493), .B(n17457), .Z(n17388) );
  XNOR U17301 ( .A(n17494), .B(n17464), .Z(n17457) );
  XOR U17302 ( .A(n17453), .B(n17452), .Z(n17464) );
  XNOR U17303 ( .A(n17495), .B(n17449), .Z(n17452) );
  XOR U17304 ( .A(n17496), .B(n17497), .Z(n17449) );
  AND U17305 ( .A(n17498), .B(n17499), .Z(n17497) );
  XNOR U17306 ( .A(n17500), .B(n17501), .Z(n17498) );
  IV U17307 ( .A(n17496), .Z(n17500) );
  XNOR U17308 ( .A(n17502), .B(n17503), .Z(n17495) );
  NOR U17309 ( .A(n17504), .B(n17505), .Z(n17503) );
  XNOR U17310 ( .A(n17502), .B(n17506), .Z(n17504) );
  XOR U17311 ( .A(n17507), .B(n17508), .Z(n17453) );
  NOR U17312 ( .A(n17509), .B(n17510), .Z(n17508) );
  XNOR U17313 ( .A(n17507), .B(n17511), .Z(n17509) );
  XNOR U17314 ( .A(n17463), .B(n17454), .Z(n17494) );
  XOR U17315 ( .A(n17512), .B(n17513), .Z(n17454) );
  AND U17316 ( .A(n17514), .B(n17515), .Z(n17513) );
  XOR U17317 ( .A(n17512), .B(n17516), .Z(n17514) );
  XOR U17318 ( .A(n17517), .B(n17469), .Z(n17463) );
  XOR U17319 ( .A(n17518), .B(n17519), .Z(n17469) );
  NOR U17320 ( .A(n17520), .B(n17521), .Z(n17519) );
  XOR U17321 ( .A(n17518), .B(n17522), .Z(n17520) );
  XNOR U17322 ( .A(n17468), .B(n17460), .Z(n17517) );
  XOR U17323 ( .A(n17523), .B(n17524), .Z(n17460) );
  AND U17324 ( .A(n17525), .B(n17526), .Z(n17524) );
  XOR U17325 ( .A(n17523), .B(n17527), .Z(n17525) );
  XNOR U17326 ( .A(n17528), .B(n17465), .Z(n17468) );
  XOR U17327 ( .A(n17529), .B(n17530), .Z(n17465) );
  AND U17328 ( .A(n17531), .B(n17532), .Z(n17530) );
  XNOR U17329 ( .A(n17533), .B(n17534), .Z(n17531) );
  IV U17330 ( .A(n17529), .Z(n17533) );
  XNOR U17331 ( .A(n17535), .B(n17536), .Z(n17528) );
  NOR U17332 ( .A(n17537), .B(n17538), .Z(n17536) );
  XNOR U17333 ( .A(n17535), .B(n17539), .Z(n17537) );
  XOR U17334 ( .A(n17458), .B(n17470), .Z(n17493) );
  NOR U17335 ( .A(n17396), .B(n17540), .Z(n17470) );
  XNOR U17336 ( .A(n17476), .B(n17475), .Z(n17458) );
  XNOR U17337 ( .A(n17541), .B(n17481), .Z(n17475) );
  XNOR U17338 ( .A(n17542), .B(n17543), .Z(n17481) );
  NOR U17339 ( .A(n17544), .B(n17545), .Z(n17543) );
  XOR U17340 ( .A(n17542), .B(n17546), .Z(n17544) );
  XNOR U17341 ( .A(n17480), .B(n17472), .Z(n17541) );
  XOR U17342 ( .A(n17547), .B(n17548), .Z(n17472) );
  AND U17343 ( .A(n17549), .B(n17550), .Z(n17548) );
  XOR U17344 ( .A(n17547), .B(n17551), .Z(n17549) );
  XNOR U17345 ( .A(n17552), .B(n17477), .Z(n17480) );
  XOR U17346 ( .A(n17553), .B(n17554), .Z(n17477) );
  AND U17347 ( .A(n17555), .B(n17556), .Z(n17554) );
  XNOR U17348 ( .A(n17557), .B(n17558), .Z(n17555) );
  IV U17349 ( .A(n17553), .Z(n17557) );
  XNOR U17350 ( .A(n17559), .B(n17560), .Z(n17552) );
  NOR U17351 ( .A(n17561), .B(n17562), .Z(n17560) );
  XNOR U17352 ( .A(n17559), .B(n17563), .Z(n17561) );
  XOR U17353 ( .A(n17486), .B(n17485), .Z(n17476) );
  XNOR U17354 ( .A(n17564), .B(n17482), .Z(n17485) );
  XOR U17355 ( .A(n17565), .B(n17566), .Z(n17482) );
  AND U17356 ( .A(n17567), .B(n17568), .Z(n17566) );
  XNOR U17357 ( .A(n17569), .B(n17570), .Z(n17567) );
  IV U17358 ( .A(n17565), .Z(n17569) );
  XNOR U17359 ( .A(n17571), .B(n17572), .Z(n17564) );
  NOR U17360 ( .A(n17573), .B(n17574), .Z(n17572) );
  XNOR U17361 ( .A(n17571), .B(n17575), .Z(n17573) );
  XOR U17362 ( .A(n17576), .B(n17577), .Z(n17486) );
  NOR U17363 ( .A(n17578), .B(n17579), .Z(n17577) );
  XNOR U17364 ( .A(n17576), .B(n17580), .Z(n17578) );
  XNOR U17365 ( .A(n17385), .B(n17489), .Z(n17491) );
  XNOR U17366 ( .A(n17581), .B(n17582), .Z(n17385) );
  AND U17367 ( .A(n111), .B(n17392), .Z(n17582) );
  XOR U17368 ( .A(n17581), .B(n17390), .Z(n17392) );
  AND U17369 ( .A(n17393), .B(n17396), .Z(n17489) );
  XOR U17370 ( .A(n17583), .B(n17540), .Z(n17396) );
  XNOR U17371 ( .A(p_input[128]), .B(p_input[2048]), .Z(n17540) );
  XNOR U17372 ( .A(n17516), .B(n17515), .Z(n17583) );
  XNOR U17373 ( .A(n17584), .B(n17527), .Z(n17515) );
  XOR U17374 ( .A(n17501), .B(n17499), .Z(n17527) );
  XNOR U17375 ( .A(n17585), .B(n17506), .Z(n17499) );
  XOR U17376 ( .A(p_input[152]), .B(p_input[2072]), .Z(n17506) );
  XOR U17377 ( .A(n17496), .B(n17505), .Z(n17585) );
  XOR U17378 ( .A(n17586), .B(n17502), .Z(n17505) );
  XOR U17379 ( .A(p_input[150]), .B(p_input[2070]), .Z(n17502) );
  XOR U17380 ( .A(p_input[151]), .B(n17295), .Z(n17586) );
  XOR U17381 ( .A(p_input[146]), .B(p_input[2066]), .Z(n17496) );
  XNOR U17382 ( .A(n17511), .B(n17510), .Z(n17501) );
  XOR U17383 ( .A(n17587), .B(n17507), .Z(n17510) );
  XOR U17384 ( .A(p_input[147]), .B(p_input[2067]), .Z(n17507) );
  XOR U17385 ( .A(p_input[148]), .B(n17297), .Z(n17587) );
  XOR U17386 ( .A(p_input[149]), .B(p_input[2069]), .Z(n17511) );
  XOR U17387 ( .A(n17526), .B(n17588), .Z(n17584) );
  IV U17388 ( .A(n17512), .Z(n17588) );
  XOR U17389 ( .A(p_input[129]), .B(p_input[2049]), .Z(n17512) );
  XNOR U17390 ( .A(n17589), .B(n17534), .Z(n17526) );
  XNOR U17391 ( .A(n17522), .B(n17521), .Z(n17534) );
  XNOR U17392 ( .A(n17590), .B(n17518), .Z(n17521) );
  XNOR U17393 ( .A(p_input[154]), .B(p_input[2074]), .Z(n17518) );
  XOR U17394 ( .A(p_input[155]), .B(n17300), .Z(n17590) );
  XOR U17395 ( .A(p_input[156]), .B(p_input[2076]), .Z(n17522) );
  XOR U17396 ( .A(n17532), .B(n17591), .Z(n17589) );
  IV U17397 ( .A(n17523), .Z(n17591) );
  XOR U17398 ( .A(p_input[145]), .B(p_input[2065]), .Z(n17523) );
  XNOR U17399 ( .A(n17592), .B(n17539), .Z(n17532) );
  XNOR U17400 ( .A(p_input[159]), .B(n17303), .Z(n17539) );
  XOR U17401 ( .A(n17529), .B(n17538), .Z(n17592) );
  XOR U17402 ( .A(n17593), .B(n17535), .Z(n17538) );
  XOR U17403 ( .A(p_input[157]), .B(p_input[2077]), .Z(n17535) );
  XOR U17404 ( .A(p_input[158]), .B(n17305), .Z(n17593) );
  XOR U17405 ( .A(p_input[153]), .B(p_input[2073]), .Z(n17529) );
  XOR U17406 ( .A(n17551), .B(n17550), .Z(n17516) );
  XNOR U17407 ( .A(n17594), .B(n17558), .Z(n17550) );
  XNOR U17408 ( .A(n17546), .B(n17545), .Z(n17558) );
  XNOR U17409 ( .A(n17595), .B(n17542), .Z(n17545) );
  XNOR U17410 ( .A(p_input[139]), .B(p_input[2059]), .Z(n17542) );
  XOR U17411 ( .A(p_input[140]), .B(n16451), .Z(n17595) );
  XOR U17412 ( .A(p_input[141]), .B(p_input[2061]), .Z(n17546) );
  XOR U17413 ( .A(n17556), .B(n17596), .Z(n17594) );
  IV U17414 ( .A(n17547), .Z(n17596) );
  XOR U17415 ( .A(p_input[130]), .B(p_input[2050]), .Z(n17547) );
  XNOR U17416 ( .A(n17597), .B(n17563), .Z(n17556) );
  XNOR U17417 ( .A(p_input[144]), .B(n16454), .Z(n17563) );
  XOR U17418 ( .A(n17553), .B(n17562), .Z(n17597) );
  XOR U17419 ( .A(n17598), .B(n17559), .Z(n17562) );
  XOR U17420 ( .A(p_input[142]), .B(p_input[2062]), .Z(n17559) );
  XOR U17421 ( .A(p_input[143]), .B(n16456), .Z(n17598) );
  XOR U17422 ( .A(p_input[138]), .B(p_input[2058]), .Z(n17553) );
  XOR U17423 ( .A(n17570), .B(n17568), .Z(n17551) );
  XNOR U17424 ( .A(n17599), .B(n17575), .Z(n17568) );
  XOR U17425 ( .A(p_input[137]), .B(p_input[2057]), .Z(n17575) );
  XOR U17426 ( .A(n17565), .B(n17574), .Z(n17599) );
  XOR U17427 ( .A(n17600), .B(n17571), .Z(n17574) );
  XOR U17428 ( .A(p_input[135]), .B(p_input[2055]), .Z(n17571) );
  XOR U17429 ( .A(p_input[136]), .B(n17312), .Z(n17600) );
  XOR U17430 ( .A(p_input[131]), .B(p_input[2051]), .Z(n17565) );
  XNOR U17431 ( .A(n17580), .B(n17579), .Z(n17570) );
  XOR U17432 ( .A(n17601), .B(n17576), .Z(n17579) );
  XOR U17433 ( .A(p_input[132]), .B(p_input[2052]), .Z(n17576) );
  XOR U17434 ( .A(p_input[133]), .B(n17314), .Z(n17601) );
  XOR U17435 ( .A(p_input[134]), .B(p_input[2054]), .Z(n17580) );
  XNOR U17436 ( .A(n17602), .B(n17603), .Z(n17393) );
  AND U17437 ( .A(n111), .B(n17604), .Z(n17603) );
  XNOR U17438 ( .A(n17605), .B(n17606), .Z(n111) );
  AND U17439 ( .A(n17607), .B(n17608), .Z(n17606) );
  XOR U17440 ( .A(n17605), .B(n17403), .Z(n17608) );
  XNOR U17441 ( .A(n17605), .B(n17345), .Z(n17607) );
  XOR U17442 ( .A(n17609), .B(n17610), .Z(n17605) );
  AND U17443 ( .A(n17611), .B(n17612), .Z(n17610) );
  XNOR U17444 ( .A(n17416), .B(n17609), .Z(n17612) );
  XOR U17445 ( .A(n17609), .B(n17357), .Z(n17611) );
  XOR U17446 ( .A(n17613), .B(n17614), .Z(n17609) );
  AND U17447 ( .A(n17615), .B(n17616), .Z(n17614) );
  XNOR U17448 ( .A(n17441), .B(n17613), .Z(n17616) );
  XOR U17449 ( .A(n17613), .B(n17368), .Z(n17615) );
  XOR U17450 ( .A(n17617), .B(n17618), .Z(n17613) );
  AND U17451 ( .A(n17619), .B(n17620), .Z(n17618) );
  XOR U17452 ( .A(n17617), .B(n17378), .Z(n17619) );
  XOR U17453 ( .A(n17621), .B(n17622), .Z(n17334) );
  AND U17454 ( .A(n115), .B(n17604), .Z(n17622) );
  XNOR U17455 ( .A(n17602), .B(n17621), .Z(n17604) );
  XNOR U17456 ( .A(n17623), .B(n17624), .Z(n115) );
  AND U17457 ( .A(n17625), .B(n17626), .Z(n17624) );
  XNOR U17458 ( .A(n17627), .B(n17623), .Z(n17626) );
  IV U17459 ( .A(n17403), .Z(n17627) );
  XNOR U17460 ( .A(n17628), .B(n17629), .Z(n17403) );
  AND U17461 ( .A(n118), .B(n17630), .Z(n17629) );
  XNOR U17462 ( .A(n17628), .B(n17631), .Z(n17630) );
  XNOR U17463 ( .A(n17345), .B(n17623), .Z(n17625) );
  XOR U17464 ( .A(n17632), .B(n17633), .Z(n17345) );
  AND U17465 ( .A(n126), .B(n17634), .Z(n17633) );
  XOR U17466 ( .A(n17635), .B(n17636), .Z(n17623) );
  AND U17467 ( .A(n17637), .B(n17638), .Z(n17636) );
  XNOR U17468 ( .A(n17635), .B(n17416), .Z(n17638) );
  XNOR U17469 ( .A(n17639), .B(n17640), .Z(n17416) );
  AND U17470 ( .A(n118), .B(n17641), .Z(n17640) );
  XOR U17471 ( .A(n17642), .B(n17639), .Z(n17641) );
  XNOR U17472 ( .A(n17643), .B(n17635), .Z(n17637) );
  IV U17473 ( .A(n17357), .Z(n17643) );
  XOR U17474 ( .A(n17644), .B(n17645), .Z(n17357) );
  AND U17475 ( .A(n126), .B(n17646), .Z(n17645) );
  XOR U17476 ( .A(n17647), .B(n17648), .Z(n17635) );
  AND U17477 ( .A(n17649), .B(n17650), .Z(n17648) );
  XNOR U17478 ( .A(n17647), .B(n17441), .Z(n17650) );
  XNOR U17479 ( .A(n17651), .B(n17652), .Z(n17441) );
  AND U17480 ( .A(n118), .B(n17653), .Z(n17652) );
  XNOR U17481 ( .A(n17654), .B(n17651), .Z(n17653) );
  XOR U17482 ( .A(n17368), .B(n17647), .Z(n17649) );
  XOR U17483 ( .A(n17655), .B(n17656), .Z(n17368) );
  AND U17484 ( .A(n126), .B(n17657), .Z(n17656) );
  XOR U17485 ( .A(n17617), .B(n17658), .Z(n17647) );
  AND U17486 ( .A(n17659), .B(n17620), .Z(n17658) );
  XNOR U17487 ( .A(n17487), .B(n17617), .Z(n17620) );
  XNOR U17488 ( .A(n17660), .B(n17661), .Z(n17487) );
  AND U17489 ( .A(n118), .B(n17662), .Z(n17661) );
  XOR U17490 ( .A(n17663), .B(n17660), .Z(n17662) );
  XNOR U17491 ( .A(n17664), .B(n17617), .Z(n17659) );
  IV U17492 ( .A(n17378), .Z(n17664) );
  XOR U17493 ( .A(n17665), .B(n17666), .Z(n17378) );
  AND U17494 ( .A(n126), .B(n17667), .Z(n17666) );
  XOR U17495 ( .A(n17668), .B(n17669), .Z(n17617) );
  AND U17496 ( .A(n17670), .B(n17671), .Z(n17669) );
  XNOR U17497 ( .A(n17668), .B(n17581), .Z(n17671) );
  XNOR U17498 ( .A(n17672), .B(n17673), .Z(n17581) );
  AND U17499 ( .A(n118), .B(n17674), .Z(n17673) );
  XNOR U17500 ( .A(n17675), .B(n17672), .Z(n17674) );
  XNOR U17501 ( .A(n17676), .B(n17668), .Z(n17670) );
  IV U17502 ( .A(n17390), .Z(n17676) );
  XOR U17503 ( .A(n17677), .B(n17678), .Z(n17390) );
  AND U17504 ( .A(n126), .B(n17679), .Z(n17678) );
  AND U17505 ( .A(n17621), .B(n17602), .Z(n17668) );
  XNOR U17506 ( .A(n17680), .B(n17681), .Z(n17602) );
  AND U17507 ( .A(n118), .B(n17682), .Z(n17681) );
  XNOR U17508 ( .A(n17683), .B(n17680), .Z(n17682) );
  XNOR U17509 ( .A(n17684), .B(n17685), .Z(n118) );
  AND U17510 ( .A(n17686), .B(n17687), .Z(n17685) );
  XOR U17511 ( .A(n17631), .B(n17684), .Z(n17687) );
  AND U17512 ( .A(n17688), .B(n17689), .Z(n17631) );
  XOR U17513 ( .A(n17684), .B(n17628), .Z(n17686) );
  XNOR U17514 ( .A(n17690), .B(n17691), .Z(n17628) );
  AND U17515 ( .A(n122), .B(n17634), .Z(n17691) );
  XOR U17516 ( .A(n17632), .B(n17690), .Z(n17634) );
  XOR U17517 ( .A(n17692), .B(n17693), .Z(n17684) );
  AND U17518 ( .A(n17694), .B(n17695), .Z(n17693) );
  XNOR U17519 ( .A(n17692), .B(n17688), .Z(n17695) );
  IV U17520 ( .A(n17642), .Z(n17688) );
  XOR U17521 ( .A(n17696), .B(n17697), .Z(n17642) );
  XOR U17522 ( .A(n17698), .B(n17689), .Z(n17697) );
  AND U17523 ( .A(n17654), .B(n17699), .Z(n17689) );
  AND U17524 ( .A(n17700), .B(n17701), .Z(n17698) );
  XOR U17525 ( .A(n17702), .B(n17696), .Z(n17700) );
  XNOR U17526 ( .A(n17639), .B(n17692), .Z(n17694) );
  XNOR U17527 ( .A(n17703), .B(n17704), .Z(n17639) );
  AND U17528 ( .A(n122), .B(n17646), .Z(n17704) );
  XOR U17529 ( .A(n17703), .B(n17644), .Z(n17646) );
  XOR U17530 ( .A(n17705), .B(n17706), .Z(n17692) );
  AND U17531 ( .A(n17707), .B(n17708), .Z(n17706) );
  XNOR U17532 ( .A(n17705), .B(n17654), .Z(n17708) );
  XOR U17533 ( .A(n17709), .B(n17701), .Z(n17654) );
  XNOR U17534 ( .A(n17710), .B(n17696), .Z(n17701) );
  XOR U17535 ( .A(n17711), .B(n17712), .Z(n17696) );
  AND U17536 ( .A(n17713), .B(n17714), .Z(n17712) );
  XOR U17537 ( .A(n17715), .B(n17711), .Z(n17713) );
  XNOR U17538 ( .A(n17716), .B(n17717), .Z(n17710) );
  AND U17539 ( .A(n17718), .B(n17719), .Z(n17717) );
  XOR U17540 ( .A(n17716), .B(n17720), .Z(n17718) );
  XNOR U17541 ( .A(n17702), .B(n17699), .Z(n17709) );
  AND U17542 ( .A(n17721), .B(n17722), .Z(n17699) );
  XOR U17543 ( .A(n17723), .B(n17724), .Z(n17702) );
  AND U17544 ( .A(n17725), .B(n17726), .Z(n17724) );
  XOR U17545 ( .A(n17723), .B(n17727), .Z(n17725) );
  XNOR U17546 ( .A(n17651), .B(n17705), .Z(n17707) );
  XNOR U17547 ( .A(n17728), .B(n17729), .Z(n17651) );
  AND U17548 ( .A(n122), .B(n17657), .Z(n17729) );
  XOR U17549 ( .A(n17728), .B(n17655), .Z(n17657) );
  XOR U17550 ( .A(n17730), .B(n17731), .Z(n17705) );
  AND U17551 ( .A(n17732), .B(n17733), .Z(n17731) );
  XNOR U17552 ( .A(n17730), .B(n17721), .Z(n17733) );
  IV U17553 ( .A(n17663), .Z(n17721) );
  XNOR U17554 ( .A(n17734), .B(n17714), .Z(n17663) );
  XNOR U17555 ( .A(n17735), .B(n17720), .Z(n17714) );
  XOR U17556 ( .A(n17736), .B(n17737), .Z(n17720) );
  AND U17557 ( .A(n17738), .B(n17739), .Z(n17737) );
  XOR U17558 ( .A(n17736), .B(n17740), .Z(n17738) );
  XNOR U17559 ( .A(n17719), .B(n17711), .Z(n17735) );
  XOR U17560 ( .A(n17741), .B(n17742), .Z(n17711) );
  AND U17561 ( .A(n17743), .B(n17744), .Z(n17742) );
  XNOR U17562 ( .A(n17745), .B(n17741), .Z(n17743) );
  XNOR U17563 ( .A(n17746), .B(n17716), .Z(n17719) );
  XOR U17564 ( .A(n17747), .B(n17748), .Z(n17716) );
  AND U17565 ( .A(n17749), .B(n17750), .Z(n17748) );
  XOR U17566 ( .A(n17747), .B(n17751), .Z(n17749) );
  XNOR U17567 ( .A(n17752), .B(n17753), .Z(n17746) );
  AND U17568 ( .A(n17754), .B(n17755), .Z(n17753) );
  XNOR U17569 ( .A(n17752), .B(n17756), .Z(n17754) );
  XNOR U17570 ( .A(n17715), .B(n17722), .Z(n17734) );
  AND U17571 ( .A(n17675), .B(n17757), .Z(n17722) );
  XOR U17572 ( .A(n17727), .B(n17726), .Z(n17715) );
  XNOR U17573 ( .A(n17758), .B(n17723), .Z(n17726) );
  XOR U17574 ( .A(n17759), .B(n17760), .Z(n17723) );
  AND U17575 ( .A(n17761), .B(n17762), .Z(n17760) );
  XOR U17576 ( .A(n17759), .B(n17763), .Z(n17761) );
  XNOR U17577 ( .A(n17764), .B(n17765), .Z(n17758) );
  AND U17578 ( .A(n17766), .B(n17767), .Z(n17765) );
  XOR U17579 ( .A(n17764), .B(n17768), .Z(n17766) );
  XOR U17580 ( .A(n17769), .B(n17770), .Z(n17727) );
  AND U17581 ( .A(n17771), .B(n17772), .Z(n17770) );
  XOR U17582 ( .A(n17769), .B(n17773), .Z(n17771) );
  XNOR U17583 ( .A(n17660), .B(n17730), .Z(n17732) );
  XNOR U17584 ( .A(n17774), .B(n17775), .Z(n17660) );
  AND U17585 ( .A(n122), .B(n17667), .Z(n17775) );
  XOR U17586 ( .A(n17774), .B(n17665), .Z(n17667) );
  XOR U17587 ( .A(n17776), .B(n17777), .Z(n17730) );
  AND U17588 ( .A(n17778), .B(n17779), .Z(n17777) );
  XNOR U17589 ( .A(n17776), .B(n17675), .Z(n17779) );
  XOR U17590 ( .A(n17780), .B(n17744), .Z(n17675) );
  XNOR U17591 ( .A(n17781), .B(n17751), .Z(n17744) );
  XOR U17592 ( .A(n17740), .B(n17739), .Z(n17751) );
  XNOR U17593 ( .A(n17782), .B(n17736), .Z(n17739) );
  XOR U17594 ( .A(n17783), .B(n17784), .Z(n17736) );
  AND U17595 ( .A(n17785), .B(n17786), .Z(n17784) );
  XNOR U17596 ( .A(n17787), .B(n17788), .Z(n17785) );
  IV U17597 ( .A(n17783), .Z(n17787) );
  XNOR U17598 ( .A(n17789), .B(n17790), .Z(n17782) );
  NOR U17599 ( .A(n17791), .B(n17792), .Z(n17790) );
  XNOR U17600 ( .A(n17789), .B(n17793), .Z(n17791) );
  XOR U17601 ( .A(n17794), .B(n17795), .Z(n17740) );
  NOR U17602 ( .A(n17796), .B(n17797), .Z(n17795) );
  XNOR U17603 ( .A(n17794), .B(n17798), .Z(n17796) );
  XNOR U17604 ( .A(n17750), .B(n17741), .Z(n17781) );
  XOR U17605 ( .A(n17799), .B(n17800), .Z(n17741) );
  AND U17606 ( .A(n17801), .B(n17802), .Z(n17800) );
  XOR U17607 ( .A(n17799), .B(n17803), .Z(n17801) );
  XOR U17608 ( .A(n17804), .B(n17756), .Z(n17750) );
  XOR U17609 ( .A(n17805), .B(n17806), .Z(n17756) );
  NOR U17610 ( .A(n17807), .B(n17808), .Z(n17806) );
  XOR U17611 ( .A(n17805), .B(n17809), .Z(n17807) );
  XNOR U17612 ( .A(n17755), .B(n17747), .Z(n17804) );
  XOR U17613 ( .A(n17810), .B(n17811), .Z(n17747) );
  AND U17614 ( .A(n17812), .B(n17813), .Z(n17811) );
  XOR U17615 ( .A(n17810), .B(n17814), .Z(n17812) );
  XNOR U17616 ( .A(n17815), .B(n17752), .Z(n17755) );
  XOR U17617 ( .A(n17816), .B(n17817), .Z(n17752) );
  AND U17618 ( .A(n17818), .B(n17819), .Z(n17817) );
  XNOR U17619 ( .A(n17820), .B(n17821), .Z(n17818) );
  IV U17620 ( .A(n17816), .Z(n17820) );
  XNOR U17621 ( .A(n17822), .B(n17823), .Z(n17815) );
  NOR U17622 ( .A(n17824), .B(n17825), .Z(n17823) );
  XNOR U17623 ( .A(n17822), .B(n17826), .Z(n17824) );
  XOR U17624 ( .A(n17745), .B(n17757), .Z(n17780) );
  NOR U17625 ( .A(n17683), .B(n17827), .Z(n17757) );
  XNOR U17626 ( .A(n17763), .B(n17762), .Z(n17745) );
  XNOR U17627 ( .A(n17828), .B(n17768), .Z(n17762) );
  XNOR U17628 ( .A(n17829), .B(n17830), .Z(n17768) );
  NOR U17629 ( .A(n17831), .B(n17832), .Z(n17830) );
  XOR U17630 ( .A(n17829), .B(n17833), .Z(n17831) );
  XNOR U17631 ( .A(n17767), .B(n17759), .Z(n17828) );
  XOR U17632 ( .A(n17834), .B(n17835), .Z(n17759) );
  AND U17633 ( .A(n17836), .B(n17837), .Z(n17835) );
  XOR U17634 ( .A(n17834), .B(n17838), .Z(n17836) );
  XNOR U17635 ( .A(n17839), .B(n17764), .Z(n17767) );
  XOR U17636 ( .A(n17840), .B(n17841), .Z(n17764) );
  AND U17637 ( .A(n17842), .B(n17843), .Z(n17841) );
  XNOR U17638 ( .A(n17844), .B(n17845), .Z(n17842) );
  IV U17639 ( .A(n17840), .Z(n17844) );
  XNOR U17640 ( .A(n17846), .B(n17847), .Z(n17839) );
  NOR U17641 ( .A(n17848), .B(n17849), .Z(n17847) );
  XNOR U17642 ( .A(n17846), .B(n17850), .Z(n17848) );
  XOR U17643 ( .A(n17773), .B(n17772), .Z(n17763) );
  XNOR U17644 ( .A(n17851), .B(n17769), .Z(n17772) );
  XOR U17645 ( .A(n17852), .B(n17853), .Z(n17769) );
  AND U17646 ( .A(n17854), .B(n17855), .Z(n17853) );
  XNOR U17647 ( .A(n17856), .B(n17857), .Z(n17854) );
  IV U17648 ( .A(n17852), .Z(n17856) );
  XNOR U17649 ( .A(n17858), .B(n17859), .Z(n17851) );
  NOR U17650 ( .A(n17860), .B(n17861), .Z(n17859) );
  XNOR U17651 ( .A(n17858), .B(n17862), .Z(n17860) );
  XOR U17652 ( .A(n17863), .B(n17864), .Z(n17773) );
  NOR U17653 ( .A(n17865), .B(n17866), .Z(n17864) );
  XNOR U17654 ( .A(n17863), .B(n17867), .Z(n17865) );
  XNOR U17655 ( .A(n17672), .B(n17776), .Z(n17778) );
  XNOR U17656 ( .A(n17868), .B(n17869), .Z(n17672) );
  AND U17657 ( .A(n122), .B(n17679), .Z(n17869) );
  XOR U17658 ( .A(n17868), .B(n17677), .Z(n17679) );
  AND U17659 ( .A(n17680), .B(n17683), .Z(n17776) );
  XOR U17660 ( .A(n17870), .B(n17827), .Z(n17683) );
  XNOR U17661 ( .A(p_input[160]), .B(p_input[2048]), .Z(n17827) );
  XNOR U17662 ( .A(n17803), .B(n17802), .Z(n17870) );
  XNOR U17663 ( .A(n17871), .B(n17814), .Z(n17802) );
  XOR U17664 ( .A(n17788), .B(n17786), .Z(n17814) );
  XNOR U17665 ( .A(n17872), .B(n17793), .Z(n17786) );
  XOR U17666 ( .A(p_input[184]), .B(p_input[2072]), .Z(n17793) );
  XOR U17667 ( .A(n17783), .B(n17792), .Z(n17872) );
  XOR U17668 ( .A(n17873), .B(n17789), .Z(n17792) );
  XOR U17669 ( .A(p_input[182]), .B(p_input[2070]), .Z(n17789) );
  XOR U17670 ( .A(p_input[183]), .B(n17295), .Z(n17873) );
  XOR U17671 ( .A(p_input[178]), .B(p_input[2066]), .Z(n17783) );
  XNOR U17672 ( .A(n17798), .B(n17797), .Z(n17788) );
  XOR U17673 ( .A(n17874), .B(n17794), .Z(n17797) );
  XOR U17674 ( .A(p_input[179]), .B(p_input[2067]), .Z(n17794) );
  XOR U17675 ( .A(p_input[180]), .B(n17297), .Z(n17874) );
  XOR U17676 ( .A(p_input[181]), .B(p_input[2069]), .Z(n17798) );
  XOR U17677 ( .A(n17813), .B(n17875), .Z(n17871) );
  IV U17678 ( .A(n17799), .Z(n17875) );
  XOR U17679 ( .A(p_input[161]), .B(p_input[2049]), .Z(n17799) );
  XNOR U17680 ( .A(n17876), .B(n17821), .Z(n17813) );
  XNOR U17681 ( .A(n17809), .B(n17808), .Z(n17821) );
  XNOR U17682 ( .A(n17877), .B(n17805), .Z(n17808) );
  XNOR U17683 ( .A(p_input[186]), .B(p_input[2074]), .Z(n17805) );
  XOR U17684 ( .A(p_input[187]), .B(n17300), .Z(n17877) );
  XOR U17685 ( .A(p_input[188]), .B(p_input[2076]), .Z(n17809) );
  XOR U17686 ( .A(n17819), .B(n17878), .Z(n17876) );
  IV U17687 ( .A(n17810), .Z(n17878) );
  XOR U17688 ( .A(p_input[177]), .B(p_input[2065]), .Z(n17810) );
  XNOR U17689 ( .A(n17879), .B(n17826), .Z(n17819) );
  XNOR U17690 ( .A(p_input[191]), .B(n17303), .Z(n17826) );
  XOR U17691 ( .A(n17816), .B(n17825), .Z(n17879) );
  XOR U17692 ( .A(n17880), .B(n17822), .Z(n17825) );
  XOR U17693 ( .A(p_input[189]), .B(p_input[2077]), .Z(n17822) );
  XOR U17694 ( .A(p_input[190]), .B(n17305), .Z(n17880) );
  XOR U17695 ( .A(p_input[185]), .B(p_input[2073]), .Z(n17816) );
  XOR U17696 ( .A(n17838), .B(n17837), .Z(n17803) );
  XNOR U17697 ( .A(n17881), .B(n17845), .Z(n17837) );
  XNOR U17698 ( .A(n17833), .B(n17832), .Z(n17845) );
  XNOR U17699 ( .A(n17882), .B(n17829), .Z(n17832) );
  XNOR U17700 ( .A(p_input[171]), .B(p_input[2059]), .Z(n17829) );
  XOR U17701 ( .A(p_input[172]), .B(n16451), .Z(n17882) );
  XOR U17702 ( .A(p_input[173]), .B(p_input[2061]), .Z(n17833) );
  XOR U17703 ( .A(n17843), .B(n17883), .Z(n17881) );
  IV U17704 ( .A(n17834), .Z(n17883) );
  XOR U17705 ( .A(p_input[162]), .B(p_input[2050]), .Z(n17834) );
  XNOR U17706 ( .A(n17884), .B(n17850), .Z(n17843) );
  XNOR U17707 ( .A(p_input[176]), .B(n16454), .Z(n17850) );
  XOR U17708 ( .A(n17840), .B(n17849), .Z(n17884) );
  XOR U17709 ( .A(n17885), .B(n17846), .Z(n17849) );
  XOR U17710 ( .A(p_input[174]), .B(p_input[2062]), .Z(n17846) );
  XOR U17711 ( .A(p_input[175]), .B(n16456), .Z(n17885) );
  XOR U17712 ( .A(p_input[170]), .B(p_input[2058]), .Z(n17840) );
  XOR U17713 ( .A(n17857), .B(n17855), .Z(n17838) );
  XNOR U17714 ( .A(n17886), .B(n17862), .Z(n17855) );
  XOR U17715 ( .A(p_input[169]), .B(p_input[2057]), .Z(n17862) );
  XOR U17716 ( .A(n17852), .B(n17861), .Z(n17886) );
  XOR U17717 ( .A(n17887), .B(n17858), .Z(n17861) );
  XOR U17718 ( .A(p_input[167]), .B(p_input[2055]), .Z(n17858) );
  XOR U17719 ( .A(p_input[168]), .B(n17312), .Z(n17887) );
  XOR U17720 ( .A(p_input[163]), .B(p_input[2051]), .Z(n17852) );
  XNOR U17721 ( .A(n17867), .B(n17866), .Z(n17857) );
  XOR U17722 ( .A(n17888), .B(n17863), .Z(n17866) );
  XOR U17723 ( .A(p_input[164]), .B(p_input[2052]), .Z(n17863) );
  XOR U17724 ( .A(p_input[165]), .B(n17314), .Z(n17888) );
  XOR U17725 ( .A(p_input[166]), .B(p_input[2054]), .Z(n17867) );
  XNOR U17726 ( .A(n17889), .B(n17890), .Z(n17680) );
  AND U17727 ( .A(n122), .B(n17891), .Z(n17890) );
  XNOR U17728 ( .A(n17892), .B(n17893), .Z(n122) );
  AND U17729 ( .A(n17894), .B(n17895), .Z(n17893) );
  XOR U17730 ( .A(n17892), .B(n17690), .Z(n17895) );
  XNOR U17731 ( .A(n17892), .B(n17632), .Z(n17894) );
  XOR U17732 ( .A(n17896), .B(n17897), .Z(n17892) );
  AND U17733 ( .A(n17898), .B(n17899), .Z(n17897) );
  XNOR U17734 ( .A(n17703), .B(n17896), .Z(n17899) );
  XOR U17735 ( .A(n17896), .B(n17644), .Z(n17898) );
  XOR U17736 ( .A(n17900), .B(n17901), .Z(n17896) );
  AND U17737 ( .A(n17902), .B(n17903), .Z(n17901) );
  XNOR U17738 ( .A(n17728), .B(n17900), .Z(n17903) );
  XOR U17739 ( .A(n17900), .B(n17655), .Z(n17902) );
  XOR U17740 ( .A(n17904), .B(n17905), .Z(n17900) );
  AND U17741 ( .A(n17906), .B(n17907), .Z(n17905) );
  XOR U17742 ( .A(n17904), .B(n17665), .Z(n17906) );
  XOR U17743 ( .A(n17908), .B(n17909), .Z(n17621) );
  AND U17744 ( .A(n126), .B(n17891), .Z(n17909) );
  XNOR U17745 ( .A(n17889), .B(n17908), .Z(n17891) );
  XNOR U17746 ( .A(n17910), .B(n17911), .Z(n126) );
  AND U17747 ( .A(n17912), .B(n17913), .Z(n17911) );
  XNOR U17748 ( .A(n17914), .B(n17910), .Z(n17913) );
  IV U17749 ( .A(n17690), .Z(n17914) );
  XNOR U17750 ( .A(n17915), .B(n17916), .Z(n17690) );
  AND U17751 ( .A(n129), .B(n17917), .Z(n17916) );
  XNOR U17752 ( .A(n17915), .B(n17918), .Z(n17917) );
  XNOR U17753 ( .A(n17632), .B(n17910), .Z(n17912) );
  XOR U17754 ( .A(n17919), .B(n17920), .Z(n17632) );
  AND U17755 ( .A(n137), .B(n17921), .Z(n17920) );
  XOR U17756 ( .A(n17922), .B(n17923), .Z(n17910) );
  AND U17757 ( .A(n17924), .B(n17925), .Z(n17923) );
  XNOR U17758 ( .A(n17922), .B(n17703), .Z(n17925) );
  XNOR U17759 ( .A(n17926), .B(n17927), .Z(n17703) );
  AND U17760 ( .A(n129), .B(n17928), .Z(n17927) );
  XOR U17761 ( .A(n17929), .B(n17926), .Z(n17928) );
  XNOR U17762 ( .A(n17930), .B(n17922), .Z(n17924) );
  IV U17763 ( .A(n17644), .Z(n17930) );
  XOR U17764 ( .A(n17931), .B(n17932), .Z(n17644) );
  AND U17765 ( .A(n137), .B(n17933), .Z(n17932) );
  XOR U17766 ( .A(n17934), .B(n17935), .Z(n17922) );
  AND U17767 ( .A(n17936), .B(n17937), .Z(n17935) );
  XNOR U17768 ( .A(n17934), .B(n17728), .Z(n17937) );
  XNOR U17769 ( .A(n17938), .B(n17939), .Z(n17728) );
  AND U17770 ( .A(n129), .B(n17940), .Z(n17939) );
  XNOR U17771 ( .A(n17941), .B(n17938), .Z(n17940) );
  XOR U17772 ( .A(n17655), .B(n17934), .Z(n17936) );
  XOR U17773 ( .A(n17942), .B(n17943), .Z(n17655) );
  AND U17774 ( .A(n137), .B(n17944), .Z(n17943) );
  XOR U17775 ( .A(n17904), .B(n17945), .Z(n17934) );
  AND U17776 ( .A(n17946), .B(n17907), .Z(n17945) );
  XNOR U17777 ( .A(n17774), .B(n17904), .Z(n17907) );
  XNOR U17778 ( .A(n17947), .B(n17948), .Z(n17774) );
  AND U17779 ( .A(n129), .B(n17949), .Z(n17948) );
  XOR U17780 ( .A(n17950), .B(n17947), .Z(n17949) );
  XNOR U17781 ( .A(n17951), .B(n17904), .Z(n17946) );
  IV U17782 ( .A(n17665), .Z(n17951) );
  XOR U17783 ( .A(n17952), .B(n17953), .Z(n17665) );
  AND U17784 ( .A(n137), .B(n17954), .Z(n17953) );
  XOR U17785 ( .A(n17955), .B(n17956), .Z(n17904) );
  AND U17786 ( .A(n17957), .B(n17958), .Z(n17956) );
  XNOR U17787 ( .A(n17955), .B(n17868), .Z(n17958) );
  XNOR U17788 ( .A(n17959), .B(n17960), .Z(n17868) );
  AND U17789 ( .A(n129), .B(n17961), .Z(n17960) );
  XNOR U17790 ( .A(n17962), .B(n17959), .Z(n17961) );
  XNOR U17791 ( .A(n17963), .B(n17955), .Z(n17957) );
  IV U17792 ( .A(n17677), .Z(n17963) );
  XOR U17793 ( .A(n17964), .B(n17965), .Z(n17677) );
  AND U17794 ( .A(n137), .B(n17966), .Z(n17965) );
  AND U17795 ( .A(n17908), .B(n17889), .Z(n17955) );
  XNOR U17796 ( .A(n17967), .B(n17968), .Z(n17889) );
  AND U17797 ( .A(n129), .B(n17969), .Z(n17968) );
  XNOR U17798 ( .A(n17970), .B(n17967), .Z(n17969) );
  XNOR U17799 ( .A(n17971), .B(n17972), .Z(n129) );
  AND U17800 ( .A(n17973), .B(n17974), .Z(n17972) );
  XOR U17801 ( .A(n17918), .B(n17971), .Z(n17974) );
  AND U17802 ( .A(n17975), .B(n17976), .Z(n17918) );
  XOR U17803 ( .A(n17971), .B(n17915), .Z(n17973) );
  XNOR U17804 ( .A(n17977), .B(n17978), .Z(n17915) );
  AND U17805 ( .A(n133), .B(n17921), .Z(n17978) );
  XOR U17806 ( .A(n17919), .B(n17977), .Z(n17921) );
  XOR U17807 ( .A(n17979), .B(n17980), .Z(n17971) );
  AND U17808 ( .A(n17981), .B(n17982), .Z(n17980) );
  XNOR U17809 ( .A(n17979), .B(n17975), .Z(n17982) );
  IV U17810 ( .A(n17929), .Z(n17975) );
  XOR U17811 ( .A(n17983), .B(n17984), .Z(n17929) );
  XOR U17812 ( .A(n17985), .B(n17976), .Z(n17984) );
  AND U17813 ( .A(n17941), .B(n17986), .Z(n17976) );
  AND U17814 ( .A(n17987), .B(n17988), .Z(n17985) );
  XOR U17815 ( .A(n17989), .B(n17983), .Z(n17987) );
  XNOR U17816 ( .A(n17926), .B(n17979), .Z(n17981) );
  XNOR U17817 ( .A(n17990), .B(n17991), .Z(n17926) );
  AND U17818 ( .A(n133), .B(n17933), .Z(n17991) );
  XOR U17819 ( .A(n17990), .B(n17931), .Z(n17933) );
  XOR U17820 ( .A(n17992), .B(n17993), .Z(n17979) );
  AND U17821 ( .A(n17994), .B(n17995), .Z(n17993) );
  XNOR U17822 ( .A(n17992), .B(n17941), .Z(n17995) );
  XOR U17823 ( .A(n17996), .B(n17988), .Z(n17941) );
  XNOR U17824 ( .A(n17997), .B(n17983), .Z(n17988) );
  XOR U17825 ( .A(n17998), .B(n17999), .Z(n17983) );
  AND U17826 ( .A(n18000), .B(n18001), .Z(n17999) );
  XOR U17827 ( .A(n18002), .B(n17998), .Z(n18000) );
  XNOR U17828 ( .A(n18003), .B(n18004), .Z(n17997) );
  AND U17829 ( .A(n18005), .B(n18006), .Z(n18004) );
  XOR U17830 ( .A(n18003), .B(n18007), .Z(n18005) );
  XNOR U17831 ( .A(n17989), .B(n17986), .Z(n17996) );
  AND U17832 ( .A(n18008), .B(n18009), .Z(n17986) );
  XOR U17833 ( .A(n18010), .B(n18011), .Z(n17989) );
  AND U17834 ( .A(n18012), .B(n18013), .Z(n18011) );
  XOR U17835 ( .A(n18010), .B(n18014), .Z(n18012) );
  XNOR U17836 ( .A(n17938), .B(n17992), .Z(n17994) );
  XNOR U17837 ( .A(n18015), .B(n18016), .Z(n17938) );
  AND U17838 ( .A(n133), .B(n17944), .Z(n18016) );
  XOR U17839 ( .A(n18015), .B(n17942), .Z(n17944) );
  XOR U17840 ( .A(n18017), .B(n18018), .Z(n17992) );
  AND U17841 ( .A(n18019), .B(n18020), .Z(n18018) );
  XNOR U17842 ( .A(n18017), .B(n18008), .Z(n18020) );
  IV U17843 ( .A(n17950), .Z(n18008) );
  XNOR U17844 ( .A(n18021), .B(n18001), .Z(n17950) );
  XNOR U17845 ( .A(n18022), .B(n18007), .Z(n18001) );
  XOR U17846 ( .A(n18023), .B(n18024), .Z(n18007) );
  AND U17847 ( .A(n18025), .B(n18026), .Z(n18024) );
  XOR U17848 ( .A(n18023), .B(n18027), .Z(n18025) );
  XNOR U17849 ( .A(n18006), .B(n17998), .Z(n18022) );
  XOR U17850 ( .A(n18028), .B(n18029), .Z(n17998) );
  AND U17851 ( .A(n18030), .B(n18031), .Z(n18029) );
  XNOR U17852 ( .A(n18032), .B(n18028), .Z(n18030) );
  XNOR U17853 ( .A(n18033), .B(n18003), .Z(n18006) );
  XOR U17854 ( .A(n18034), .B(n18035), .Z(n18003) );
  AND U17855 ( .A(n18036), .B(n18037), .Z(n18035) );
  XOR U17856 ( .A(n18034), .B(n18038), .Z(n18036) );
  XNOR U17857 ( .A(n18039), .B(n18040), .Z(n18033) );
  AND U17858 ( .A(n18041), .B(n18042), .Z(n18040) );
  XNOR U17859 ( .A(n18039), .B(n18043), .Z(n18041) );
  XNOR U17860 ( .A(n18002), .B(n18009), .Z(n18021) );
  AND U17861 ( .A(n17962), .B(n18044), .Z(n18009) );
  XOR U17862 ( .A(n18014), .B(n18013), .Z(n18002) );
  XNOR U17863 ( .A(n18045), .B(n18010), .Z(n18013) );
  XOR U17864 ( .A(n18046), .B(n18047), .Z(n18010) );
  AND U17865 ( .A(n18048), .B(n18049), .Z(n18047) );
  XOR U17866 ( .A(n18046), .B(n18050), .Z(n18048) );
  XNOR U17867 ( .A(n18051), .B(n18052), .Z(n18045) );
  AND U17868 ( .A(n18053), .B(n18054), .Z(n18052) );
  XOR U17869 ( .A(n18051), .B(n18055), .Z(n18053) );
  XOR U17870 ( .A(n18056), .B(n18057), .Z(n18014) );
  AND U17871 ( .A(n18058), .B(n18059), .Z(n18057) );
  XOR U17872 ( .A(n18056), .B(n18060), .Z(n18058) );
  XNOR U17873 ( .A(n17947), .B(n18017), .Z(n18019) );
  XNOR U17874 ( .A(n18061), .B(n18062), .Z(n17947) );
  AND U17875 ( .A(n133), .B(n17954), .Z(n18062) );
  XOR U17876 ( .A(n18061), .B(n17952), .Z(n17954) );
  XOR U17877 ( .A(n18063), .B(n18064), .Z(n18017) );
  AND U17878 ( .A(n18065), .B(n18066), .Z(n18064) );
  XNOR U17879 ( .A(n18063), .B(n17962), .Z(n18066) );
  XOR U17880 ( .A(n18067), .B(n18031), .Z(n17962) );
  XNOR U17881 ( .A(n18068), .B(n18038), .Z(n18031) );
  XOR U17882 ( .A(n18027), .B(n18026), .Z(n18038) );
  XNOR U17883 ( .A(n18069), .B(n18023), .Z(n18026) );
  XOR U17884 ( .A(n18070), .B(n18071), .Z(n18023) );
  AND U17885 ( .A(n18072), .B(n18073), .Z(n18071) );
  XOR U17886 ( .A(n18070), .B(n18074), .Z(n18072) );
  XNOR U17887 ( .A(n18075), .B(n18076), .Z(n18069) );
  NOR U17888 ( .A(n18077), .B(n18078), .Z(n18076) );
  XNOR U17889 ( .A(n18075), .B(n18079), .Z(n18077) );
  XOR U17890 ( .A(n18080), .B(n18081), .Z(n18027) );
  NOR U17891 ( .A(n18082), .B(n18083), .Z(n18081) );
  XNOR U17892 ( .A(n18080), .B(n18084), .Z(n18082) );
  XNOR U17893 ( .A(n18037), .B(n18028), .Z(n18068) );
  XOR U17894 ( .A(n18085), .B(n18086), .Z(n18028) );
  NOR U17895 ( .A(n18087), .B(n18088), .Z(n18086) );
  XOR U17896 ( .A(n18089), .B(n18090), .Z(n18087) );
  XOR U17897 ( .A(n18091), .B(n18043), .Z(n18037) );
  XNOR U17898 ( .A(n18092), .B(n18093), .Z(n18043) );
  NOR U17899 ( .A(n18094), .B(n18095), .Z(n18093) );
  XNOR U17900 ( .A(n18092), .B(n18096), .Z(n18094) );
  XNOR U17901 ( .A(n18042), .B(n18034), .Z(n18091) );
  XOR U17902 ( .A(n18097), .B(n18098), .Z(n18034) );
  AND U17903 ( .A(n18099), .B(n18100), .Z(n18098) );
  XOR U17904 ( .A(n18097), .B(n18101), .Z(n18099) );
  XNOR U17905 ( .A(n18102), .B(n18039), .Z(n18042) );
  XOR U17906 ( .A(n18103), .B(n18104), .Z(n18039) );
  AND U17907 ( .A(n18105), .B(n18106), .Z(n18104) );
  XOR U17908 ( .A(n18103), .B(n18107), .Z(n18105) );
  XNOR U17909 ( .A(n18108), .B(n18109), .Z(n18102) );
  NOR U17910 ( .A(n18110), .B(n18111), .Z(n18109) );
  XOR U17911 ( .A(n18108), .B(n18112), .Z(n18110) );
  XOR U17912 ( .A(n18032), .B(n18044), .Z(n18067) );
  NOR U17913 ( .A(n17970), .B(n18113), .Z(n18044) );
  XNOR U17914 ( .A(n18050), .B(n18049), .Z(n18032) );
  XNOR U17915 ( .A(n18114), .B(n18055), .Z(n18049) );
  XNOR U17916 ( .A(n18115), .B(n18116), .Z(n18055) );
  NOR U17917 ( .A(n18117), .B(n18118), .Z(n18116) );
  XOR U17918 ( .A(n18115), .B(n18119), .Z(n18117) );
  XNOR U17919 ( .A(n18054), .B(n18046), .Z(n18114) );
  XOR U17920 ( .A(n18120), .B(n18121), .Z(n18046) );
  AND U17921 ( .A(n18122), .B(n18123), .Z(n18121) );
  XOR U17922 ( .A(n18120), .B(n18124), .Z(n18122) );
  XNOR U17923 ( .A(n18125), .B(n18051), .Z(n18054) );
  XOR U17924 ( .A(n18126), .B(n18127), .Z(n18051) );
  AND U17925 ( .A(n18128), .B(n18129), .Z(n18127) );
  XNOR U17926 ( .A(n18130), .B(n18131), .Z(n18128) );
  IV U17927 ( .A(n18126), .Z(n18130) );
  XNOR U17928 ( .A(n18132), .B(n18133), .Z(n18125) );
  NOR U17929 ( .A(n18134), .B(n18135), .Z(n18133) );
  XOR U17930 ( .A(n18132), .B(n18136), .Z(n18134) );
  XOR U17931 ( .A(n18060), .B(n18059), .Z(n18050) );
  XNOR U17932 ( .A(n18137), .B(n18056), .Z(n18059) );
  XOR U17933 ( .A(n18138), .B(n18139), .Z(n18056) );
  AND U17934 ( .A(n18140), .B(n18141), .Z(n18139) );
  XNOR U17935 ( .A(n18142), .B(n18143), .Z(n18140) );
  IV U17936 ( .A(n18138), .Z(n18142) );
  XNOR U17937 ( .A(n18144), .B(n18145), .Z(n18137) );
  NOR U17938 ( .A(n18146), .B(n18147), .Z(n18145) );
  XNOR U17939 ( .A(n18144), .B(n18148), .Z(n18146) );
  XOR U17940 ( .A(n18149), .B(n18150), .Z(n18060) );
  NOR U17941 ( .A(n18151), .B(n18152), .Z(n18150) );
  XNOR U17942 ( .A(n18149), .B(n18153), .Z(n18151) );
  XNOR U17943 ( .A(n17959), .B(n18063), .Z(n18065) );
  XNOR U17944 ( .A(n18154), .B(n18155), .Z(n17959) );
  AND U17945 ( .A(n133), .B(n17966), .Z(n18155) );
  XOR U17946 ( .A(n18154), .B(n17964), .Z(n17966) );
  AND U17947 ( .A(n17967), .B(n17970), .Z(n18063) );
  XOR U17948 ( .A(n18156), .B(n18113), .Z(n17970) );
  XNOR U17949 ( .A(p_input[192]), .B(p_input[2048]), .Z(n18113) );
  XOR U17950 ( .A(n18090), .B(n18088), .Z(n18156) );
  XOR U17951 ( .A(n18157), .B(n18101), .Z(n18088) );
  XOR U17952 ( .A(n18074), .B(n18073), .Z(n18101) );
  XNOR U17953 ( .A(n18158), .B(n18079), .Z(n18073) );
  XOR U17954 ( .A(p_input[2072]), .B(p_input[216]), .Z(n18079) );
  XOR U17955 ( .A(n18070), .B(n18078), .Z(n18158) );
  XOR U17956 ( .A(n18159), .B(n18075), .Z(n18078) );
  XOR U17957 ( .A(p_input[2070]), .B(p_input[214]), .Z(n18075) );
  XNOR U17958 ( .A(p_input[2071]), .B(p_input[215]), .Z(n18159) );
  XNOR U17959 ( .A(n16727), .B(p_input[210]), .Z(n18070) );
  XNOR U17960 ( .A(n18084), .B(n18083), .Z(n18074) );
  XOR U17961 ( .A(n18160), .B(n18080), .Z(n18083) );
  XOR U17962 ( .A(p_input[2067]), .B(p_input[211]), .Z(n18080) );
  XNOR U17963 ( .A(p_input[2068]), .B(p_input[212]), .Z(n18160) );
  XOR U17964 ( .A(p_input[2069]), .B(p_input[213]), .Z(n18084) );
  XOR U17965 ( .A(n18100), .B(n18089), .Z(n18157) );
  IV U17966 ( .A(n18085), .Z(n18089) );
  XOR U17967 ( .A(p_input[193]), .B(p_input[2049]), .Z(n18085) );
  XNOR U17968 ( .A(n18161), .B(n18107), .Z(n18100) );
  XNOR U17969 ( .A(n18096), .B(n18095), .Z(n18107) );
  XOR U17970 ( .A(n18162), .B(n18092), .Z(n18095) );
  XNOR U17971 ( .A(n16444), .B(p_input[218]), .Z(n18092) );
  XNOR U17972 ( .A(p_input[2075]), .B(p_input[219]), .Z(n18162) );
  XOR U17973 ( .A(p_input[2076]), .B(p_input[220]), .Z(n18096) );
  XNOR U17974 ( .A(n18106), .B(n18097), .Z(n18161) );
  XNOR U17975 ( .A(n16732), .B(p_input[209]), .Z(n18097) );
  XOR U17976 ( .A(n18163), .B(n18112), .Z(n18106) );
  XNOR U17977 ( .A(p_input[2079]), .B(p_input[223]), .Z(n18112) );
  XOR U17978 ( .A(n18103), .B(n18111), .Z(n18163) );
  XOR U17979 ( .A(n18164), .B(n18108), .Z(n18111) );
  XOR U17980 ( .A(p_input[2077]), .B(p_input[221]), .Z(n18108) );
  XNOR U17981 ( .A(p_input[2078]), .B(p_input[222]), .Z(n18164) );
  XNOR U17982 ( .A(n16448), .B(p_input[217]), .Z(n18103) );
  XOR U17983 ( .A(n18124), .B(n18123), .Z(n18090) );
  XNOR U17984 ( .A(n18165), .B(n18131), .Z(n18123) );
  XNOR U17985 ( .A(n18119), .B(n18118), .Z(n18131) );
  XNOR U17986 ( .A(n18166), .B(n18115), .Z(n18118) );
  XNOR U17987 ( .A(p_input[203]), .B(p_input[2059]), .Z(n18115) );
  XOR U17988 ( .A(p_input[204]), .B(n16451), .Z(n18166) );
  XOR U17989 ( .A(p_input[205]), .B(p_input[2061]), .Z(n18119) );
  XOR U17990 ( .A(n18129), .B(n18167), .Z(n18165) );
  IV U17991 ( .A(n18120), .Z(n18167) );
  XOR U17992 ( .A(p_input[194]), .B(p_input[2050]), .Z(n18120) );
  XOR U17993 ( .A(n18168), .B(n18136), .Z(n18129) );
  XNOR U17994 ( .A(p_input[2064]), .B(p_input[208]), .Z(n18136) );
  XOR U17995 ( .A(n18126), .B(n18135), .Z(n18168) );
  XOR U17996 ( .A(n18169), .B(n18132), .Z(n18135) );
  XOR U17997 ( .A(p_input[2062]), .B(p_input[206]), .Z(n18132) );
  XNOR U17998 ( .A(p_input[2063]), .B(p_input[207]), .Z(n18169) );
  XOR U17999 ( .A(p_input[202]), .B(p_input[2058]), .Z(n18126) );
  XOR U18000 ( .A(n18143), .B(n18141), .Z(n18124) );
  XNOR U18001 ( .A(n18170), .B(n18148), .Z(n18141) );
  XOR U18002 ( .A(p_input[201]), .B(p_input[2057]), .Z(n18148) );
  XOR U18003 ( .A(n18138), .B(n18147), .Z(n18170) );
  XOR U18004 ( .A(n18171), .B(n18144), .Z(n18147) );
  XOR U18005 ( .A(p_input[199]), .B(p_input[2055]), .Z(n18144) );
  XOR U18006 ( .A(p_input[200]), .B(n17312), .Z(n18171) );
  XOR U18007 ( .A(p_input[195]), .B(p_input[2051]), .Z(n18138) );
  XNOR U18008 ( .A(n18153), .B(n18152), .Z(n18143) );
  XOR U18009 ( .A(n18172), .B(n18149), .Z(n18152) );
  XOR U18010 ( .A(p_input[196]), .B(p_input[2052]), .Z(n18149) );
  XOR U18011 ( .A(p_input[197]), .B(n17314), .Z(n18172) );
  XOR U18012 ( .A(p_input[198]), .B(p_input[2054]), .Z(n18153) );
  XNOR U18013 ( .A(n18173), .B(n18174), .Z(n17967) );
  AND U18014 ( .A(n133), .B(n18175), .Z(n18174) );
  XNOR U18015 ( .A(n18176), .B(n18177), .Z(n133) );
  AND U18016 ( .A(n18178), .B(n18179), .Z(n18177) );
  XOR U18017 ( .A(n18176), .B(n17977), .Z(n18179) );
  XNOR U18018 ( .A(n18176), .B(n17919), .Z(n18178) );
  XOR U18019 ( .A(n18180), .B(n18181), .Z(n18176) );
  AND U18020 ( .A(n18182), .B(n18183), .Z(n18181) );
  XNOR U18021 ( .A(n17990), .B(n18180), .Z(n18183) );
  XOR U18022 ( .A(n18180), .B(n17931), .Z(n18182) );
  XOR U18023 ( .A(n18184), .B(n18185), .Z(n18180) );
  AND U18024 ( .A(n18186), .B(n18187), .Z(n18185) );
  XNOR U18025 ( .A(n18015), .B(n18184), .Z(n18187) );
  XOR U18026 ( .A(n18184), .B(n17942), .Z(n18186) );
  XOR U18027 ( .A(n18188), .B(n18189), .Z(n18184) );
  AND U18028 ( .A(n18190), .B(n18191), .Z(n18189) );
  XOR U18029 ( .A(n18188), .B(n17952), .Z(n18190) );
  XOR U18030 ( .A(n18192), .B(n18193), .Z(n17908) );
  AND U18031 ( .A(n137), .B(n18175), .Z(n18193) );
  XNOR U18032 ( .A(n18173), .B(n18192), .Z(n18175) );
  XNOR U18033 ( .A(n18194), .B(n18195), .Z(n137) );
  AND U18034 ( .A(n18196), .B(n18197), .Z(n18195) );
  XNOR U18035 ( .A(n18198), .B(n18194), .Z(n18197) );
  IV U18036 ( .A(n17977), .Z(n18198) );
  XNOR U18037 ( .A(n18199), .B(n18200), .Z(n17977) );
  AND U18038 ( .A(n140), .B(n18201), .Z(n18200) );
  XNOR U18039 ( .A(n18199), .B(n18202), .Z(n18201) );
  XNOR U18040 ( .A(n17919), .B(n18194), .Z(n18196) );
  XOR U18041 ( .A(n18203), .B(n18204), .Z(n17919) );
  AND U18042 ( .A(n148), .B(n18205), .Z(n18204) );
  XOR U18043 ( .A(n18206), .B(n18207), .Z(n18194) );
  AND U18044 ( .A(n18208), .B(n18209), .Z(n18207) );
  XNOR U18045 ( .A(n18206), .B(n17990), .Z(n18209) );
  XNOR U18046 ( .A(n18210), .B(n18211), .Z(n17990) );
  AND U18047 ( .A(n140), .B(n18212), .Z(n18211) );
  XOR U18048 ( .A(n18213), .B(n18210), .Z(n18212) );
  XNOR U18049 ( .A(n18214), .B(n18206), .Z(n18208) );
  IV U18050 ( .A(n17931), .Z(n18214) );
  XOR U18051 ( .A(n18215), .B(n18216), .Z(n17931) );
  AND U18052 ( .A(n148), .B(n18217), .Z(n18216) );
  XOR U18053 ( .A(n18218), .B(n18219), .Z(n18206) );
  AND U18054 ( .A(n18220), .B(n18221), .Z(n18219) );
  XNOR U18055 ( .A(n18218), .B(n18015), .Z(n18221) );
  XNOR U18056 ( .A(n18222), .B(n18223), .Z(n18015) );
  AND U18057 ( .A(n140), .B(n18224), .Z(n18223) );
  XNOR U18058 ( .A(n18225), .B(n18222), .Z(n18224) );
  XOR U18059 ( .A(n17942), .B(n18218), .Z(n18220) );
  XOR U18060 ( .A(n18226), .B(n18227), .Z(n17942) );
  AND U18061 ( .A(n148), .B(n18228), .Z(n18227) );
  XOR U18062 ( .A(n18188), .B(n18229), .Z(n18218) );
  AND U18063 ( .A(n18230), .B(n18191), .Z(n18229) );
  XNOR U18064 ( .A(n18061), .B(n18188), .Z(n18191) );
  XNOR U18065 ( .A(n18231), .B(n18232), .Z(n18061) );
  AND U18066 ( .A(n140), .B(n18233), .Z(n18232) );
  XOR U18067 ( .A(n18234), .B(n18231), .Z(n18233) );
  XNOR U18068 ( .A(n18235), .B(n18188), .Z(n18230) );
  IV U18069 ( .A(n17952), .Z(n18235) );
  XOR U18070 ( .A(n18236), .B(n18237), .Z(n17952) );
  AND U18071 ( .A(n148), .B(n18238), .Z(n18237) );
  XOR U18072 ( .A(n18239), .B(n18240), .Z(n18188) );
  AND U18073 ( .A(n18241), .B(n18242), .Z(n18240) );
  XNOR U18074 ( .A(n18239), .B(n18154), .Z(n18242) );
  XNOR U18075 ( .A(n18243), .B(n18244), .Z(n18154) );
  AND U18076 ( .A(n140), .B(n18245), .Z(n18244) );
  XNOR U18077 ( .A(n18246), .B(n18243), .Z(n18245) );
  XNOR U18078 ( .A(n18247), .B(n18239), .Z(n18241) );
  IV U18079 ( .A(n17964), .Z(n18247) );
  XOR U18080 ( .A(n18248), .B(n18249), .Z(n17964) );
  AND U18081 ( .A(n148), .B(n18250), .Z(n18249) );
  AND U18082 ( .A(n18192), .B(n18173), .Z(n18239) );
  XNOR U18083 ( .A(n18251), .B(n18252), .Z(n18173) );
  AND U18084 ( .A(n140), .B(n18253), .Z(n18252) );
  XNOR U18085 ( .A(n18254), .B(n18251), .Z(n18253) );
  XNOR U18086 ( .A(n18255), .B(n18256), .Z(n140) );
  AND U18087 ( .A(n18257), .B(n18258), .Z(n18256) );
  XOR U18088 ( .A(n18202), .B(n18255), .Z(n18258) );
  AND U18089 ( .A(n18259), .B(n18260), .Z(n18202) );
  XOR U18090 ( .A(n18255), .B(n18199), .Z(n18257) );
  XNOR U18091 ( .A(n18261), .B(n18262), .Z(n18199) );
  AND U18092 ( .A(n144), .B(n18205), .Z(n18262) );
  XOR U18093 ( .A(n18203), .B(n18261), .Z(n18205) );
  XOR U18094 ( .A(n18263), .B(n18264), .Z(n18255) );
  AND U18095 ( .A(n18265), .B(n18266), .Z(n18264) );
  XNOR U18096 ( .A(n18263), .B(n18259), .Z(n18266) );
  IV U18097 ( .A(n18213), .Z(n18259) );
  XOR U18098 ( .A(n18267), .B(n18268), .Z(n18213) );
  XOR U18099 ( .A(n18269), .B(n18260), .Z(n18268) );
  AND U18100 ( .A(n18225), .B(n18270), .Z(n18260) );
  AND U18101 ( .A(n18271), .B(n18272), .Z(n18269) );
  XOR U18102 ( .A(n18273), .B(n18267), .Z(n18271) );
  XNOR U18103 ( .A(n18210), .B(n18263), .Z(n18265) );
  XNOR U18104 ( .A(n18274), .B(n18275), .Z(n18210) );
  AND U18105 ( .A(n144), .B(n18217), .Z(n18275) );
  XOR U18106 ( .A(n18274), .B(n18215), .Z(n18217) );
  XOR U18107 ( .A(n18276), .B(n18277), .Z(n18263) );
  AND U18108 ( .A(n18278), .B(n18279), .Z(n18277) );
  XNOR U18109 ( .A(n18276), .B(n18225), .Z(n18279) );
  XOR U18110 ( .A(n18280), .B(n18272), .Z(n18225) );
  XNOR U18111 ( .A(n18281), .B(n18267), .Z(n18272) );
  XOR U18112 ( .A(n18282), .B(n18283), .Z(n18267) );
  AND U18113 ( .A(n18284), .B(n18285), .Z(n18283) );
  XOR U18114 ( .A(n18286), .B(n18282), .Z(n18284) );
  XNOR U18115 ( .A(n18287), .B(n18288), .Z(n18281) );
  AND U18116 ( .A(n18289), .B(n18290), .Z(n18288) );
  XOR U18117 ( .A(n18287), .B(n18291), .Z(n18289) );
  XNOR U18118 ( .A(n18273), .B(n18270), .Z(n18280) );
  AND U18119 ( .A(n18292), .B(n18293), .Z(n18270) );
  XOR U18120 ( .A(n18294), .B(n18295), .Z(n18273) );
  AND U18121 ( .A(n18296), .B(n18297), .Z(n18295) );
  XOR U18122 ( .A(n18294), .B(n18298), .Z(n18296) );
  XNOR U18123 ( .A(n18222), .B(n18276), .Z(n18278) );
  XNOR U18124 ( .A(n18299), .B(n18300), .Z(n18222) );
  AND U18125 ( .A(n144), .B(n18228), .Z(n18300) );
  XOR U18126 ( .A(n18299), .B(n18226), .Z(n18228) );
  XOR U18127 ( .A(n18301), .B(n18302), .Z(n18276) );
  AND U18128 ( .A(n18303), .B(n18304), .Z(n18302) );
  XNOR U18129 ( .A(n18301), .B(n18292), .Z(n18304) );
  IV U18130 ( .A(n18234), .Z(n18292) );
  XNOR U18131 ( .A(n18305), .B(n18285), .Z(n18234) );
  XNOR U18132 ( .A(n18306), .B(n18291), .Z(n18285) );
  XOR U18133 ( .A(n18307), .B(n18308), .Z(n18291) );
  AND U18134 ( .A(n18309), .B(n18310), .Z(n18308) );
  XOR U18135 ( .A(n18307), .B(n18311), .Z(n18309) );
  XNOR U18136 ( .A(n18290), .B(n18282), .Z(n18306) );
  XOR U18137 ( .A(n18312), .B(n18313), .Z(n18282) );
  AND U18138 ( .A(n18314), .B(n18315), .Z(n18313) );
  XNOR U18139 ( .A(n18316), .B(n18312), .Z(n18314) );
  XNOR U18140 ( .A(n18317), .B(n18287), .Z(n18290) );
  XOR U18141 ( .A(n18318), .B(n18319), .Z(n18287) );
  AND U18142 ( .A(n18320), .B(n18321), .Z(n18319) );
  XOR U18143 ( .A(n18318), .B(n18322), .Z(n18320) );
  XNOR U18144 ( .A(n18323), .B(n18324), .Z(n18317) );
  AND U18145 ( .A(n18325), .B(n18326), .Z(n18324) );
  XNOR U18146 ( .A(n18323), .B(n18327), .Z(n18325) );
  XNOR U18147 ( .A(n18286), .B(n18293), .Z(n18305) );
  AND U18148 ( .A(n18246), .B(n18328), .Z(n18293) );
  XOR U18149 ( .A(n18298), .B(n18297), .Z(n18286) );
  XNOR U18150 ( .A(n18329), .B(n18294), .Z(n18297) );
  XOR U18151 ( .A(n18330), .B(n18331), .Z(n18294) );
  AND U18152 ( .A(n18332), .B(n18333), .Z(n18331) );
  XOR U18153 ( .A(n18330), .B(n18334), .Z(n18332) );
  XNOR U18154 ( .A(n18335), .B(n18336), .Z(n18329) );
  AND U18155 ( .A(n18337), .B(n18338), .Z(n18336) );
  XOR U18156 ( .A(n18335), .B(n18339), .Z(n18337) );
  XOR U18157 ( .A(n18340), .B(n18341), .Z(n18298) );
  AND U18158 ( .A(n18342), .B(n18343), .Z(n18341) );
  XOR U18159 ( .A(n18340), .B(n18344), .Z(n18342) );
  XNOR U18160 ( .A(n18231), .B(n18301), .Z(n18303) );
  XNOR U18161 ( .A(n18345), .B(n18346), .Z(n18231) );
  AND U18162 ( .A(n144), .B(n18238), .Z(n18346) );
  XOR U18163 ( .A(n18345), .B(n18236), .Z(n18238) );
  XOR U18164 ( .A(n18347), .B(n18348), .Z(n18301) );
  AND U18165 ( .A(n18349), .B(n18350), .Z(n18348) );
  XNOR U18166 ( .A(n18347), .B(n18246), .Z(n18350) );
  XOR U18167 ( .A(n18351), .B(n18315), .Z(n18246) );
  XNOR U18168 ( .A(n18352), .B(n18322), .Z(n18315) );
  XOR U18169 ( .A(n18311), .B(n18310), .Z(n18322) );
  XNOR U18170 ( .A(n18353), .B(n18307), .Z(n18310) );
  XOR U18171 ( .A(n18354), .B(n18355), .Z(n18307) );
  AND U18172 ( .A(n18356), .B(n18357), .Z(n18355) );
  XOR U18173 ( .A(n18354), .B(n18358), .Z(n18356) );
  XNOR U18174 ( .A(n18359), .B(n18360), .Z(n18353) );
  NOR U18175 ( .A(n18361), .B(n18362), .Z(n18360) );
  XNOR U18176 ( .A(n18359), .B(n18363), .Z(n18361) );
  XOR U18177 ( .A(n18364), .B(n18365), .Z(n18311) );
  NOR U18178 ( .A(n18366), .B(n18367), .Z(n18365) );
  XNOR U18179 ( .A(n18364), .B(n18368), .Z(n18366) );
  XNOR U18180 ( .A(n18321), .B(n18312), .Z(n18352) );
  XOR U18181 ( .A(n18369), .B(n18370), .Z(n18312) );
  NOR U18182 ( .A(n18371), .B(n18372), .Z(n18370) );
  XNOR U18183 ( .A(n18369), .B(n18373), .Z(n18371) );
  XOR U18184 ( .A(n18374), .B(n18327), .Z(n18321) );
  XNOR U18185 ( .A(n18375), .B(n18376), .Z(n18327) );
  NOR U18186 ( .A(n18377), .B(n18378), .Z(n18376) );
  XNOR U18187 ( .A(n18375), .B(n18379), .Z(n18377) );
  XNOR U18188 ( .A(n18326), .B(n18318), .Z(n18374) );
  XOR U18189 ( .A(n18380), .B(n18381), .Z(n18318) );
  AND U18190 ( .A(n18382), .B(n18383), .Z(n18381) );
  XOR U18191 ( .A(n18380), .B(n18384), .Z(n18382) );
  XNOR U18192 ( .A(n18385), .B(n18323), .Z(n18326) );
  XOR U18193 ( .A(n18386), .B(n18387), .Z(n18323) );
  AND U18194 ( .A(n18388), .B(n18389), .Z(n18387) );
  XOR U18195 ( .A(n18386), .B(n18390), .Z(n18388) );
  XNOR U18196 ( .A(n18391), .B(n18392), .Z(n18385) );
  NOR U18197 ( .A(n18393), .B(n18394), .Z(n18392) );
  XOR U18198 ( .A(n18391), .B(n18395), .Z(n18393) );
  XOR U18199 ( .A(n18316), .B(n18328), .Z(n18351) );
  NOR U18200 ( .A(n18254), .B(n18396), .Z(n18328) );
  XNOR U18201 ( .A(n18334), .B(n18333), .Z(n18316) );
  XNOR U18202 ( .A(n18397), .B(n18339), .Z(n18333) );
  XOR U18203 ( .A(n18398), .B(n18399), .Z(n18339) );
  NOR U18204 ( .A(n18400), .B(n18401), .Z(n18399) );
  XNOR U18205 ( .A(n18398), .B(n18402), .Z(n18400) );
  XNOR U18206 ( .A(n18338), .B(n18330), .Z(n18397) );
  XOR U18207 ( .A(n18403), .B(n18404), .Z(n18330) );
  AND U18208 ( .A(n18405), .B(n18406), .Z(n18404) );
  XNOR U18209 ( .A(n18403), .B(n18407), .Z(n18405) );
  XNOR U18210 ( .A(n18408), .B(n18335), .Z(n18338) );
  XOR U18211 ( .A(n18409), .B(n18410), .Z(n18335) );
  AND U18212 ( .A(n18411), .B(n18412), .Z(n18410) );
  XOR U18213 ( .A(n18409), .B(n18413), .Z(n18411) );
  XNOR U18214 ( .A(n18414), .B(n18415), .Z(n18408) );
  NOR U18215 ( .A(n18416), .B(n18417), .Z(n18415) );
  XOR U18216 ( .A(n18414), .B(n18418), .Z(n18416) );
  XOR U18217 ( .A(n18344), .B(n18343), .Z(n18334) );
  XNOR U18218 ( .A(n18419), .B(n18340), .Z(n18343) );
  XOR U18219 ( .A(n18420), .B(n18421), .Z(n18340) );
  AND U18220 ( .A(n18422), .B(n18423), .Z(n18421) );
  XOR U18221 ( .A(n18420), .B(n18424), .Z(n18422) );
  XNOR U18222 ( .A(n18425), .B(n18426), .Z(n18419) );
  NOR U18223 ( .A(n18427), .B(n18428), .Z(n18426) );
  XNOR U18224 ( .A(n18425), .B(n18429), .Z(n18427) );
  XOR U18225 ( .A(n18430), .B(n18431), .Z(n18344) );
  NOR U18226 ( .A(n18432), .B(n18433), .Z(n18431) );
  XNOR U18227 ( .A(n18430), .B(n18434), .Z(n18432) );
  XNOR U18228 ( .A(n18243), .B(n18347), .Z(n18349) );
  XNOR U18229 ( .A(n18435), .B(n18436), .Z(n18243) );
  AND U18230 ( .A(n144), .B(n18250), .Z(n18436) );
  XOR U18231 ( .A(n18435), .B(n18248), .Z(n18250) );
  AND U18232 ( .A(n18251), .B(n18254), .Z(n18347) );
  XOR U18233 ( .A(n18437), .B(n18396), .Z(n18254) );
  XNOR U18234 ( .A(p_input[2048]), .B(p_input[224]), .Z(n18396) );
  XOR U18235 ( .A(n18373), .B(n18372), .Z(n18437) );
  XOR U18236 ( .A(n18438), .B(n18384), .Z(n18372) );
  XOR U18237 ( .A(n18358), .B(n18357), .Z(n18384) );
  XNOR U18238 ( .A(n18439), .B(n18363), .Z(n18357) );
  XOR U18239 ( .A(p_input[2072]), .B(p_input[248]), .Z(n18363) );
  XOR U18240 ( .A(n18354), .B(n18362), .Z(n18439) );
  XOR U18241 ( .A(n18440), .B(n18359), .Z(n18362) );
  XOR U18242 ( .A(p_input[2070]), .B(p_input[246]), .Z(n18359) );
  XNOR U18243 ( .A(p_input[2071]), .B(p_input[247]), .Z(n18440) );
  XNOR U18244 ( .A(n16727), .B(p_input[242]), .Z(n18354) );
  XNOR U18245 ( .A(n18368), .B(n18367), .Z(n18358) );
  XOR U18246 ( .A(n18441), .B(n18364), .Z(n18367) );
  XOR U18247 ( .A(p_input[2067]), .B(p_input[243]), .Z(n18364) );
  XNOR U18248 ( .A(p_input[2068]), .B(p_input[244]), .Z(n18441) );
  XOR U18249 ( .A(p_input[2069]), .B(p_input[245]), .Z(n18368) );
  XNOR U18250 ( .A(n18383), .B(n18369), .Z(n18438) );
  XNOR U18251 ( .A(n16729), .B(p_input[225]), .Z(n18369) );
  XNOR U18252 ( .A(n18442), .B(n18390), .Z(n18383) );
  XNOR U18253 ( .A(n18379), .B(n18378), .Z(n18390) );
  XOR U18254 ( .A(n18443), .B(n18375), .Z(n18378) );
  XNOR U18255 ( .A(n16444), .B(p_input[250]), .Z(n18375) );
  XNOR U18256 ( .A(p_input[2075]), .B(p_input[251]), .Z(n18443) );
  XOR U18257 ( .A(p_input[2076]), .B(p_input[252]), .Z(n18379) );
  XNOR U18258 ( .A(n18389), .B(n18380), .Z(n18442) );
  XNOR U18259 ( .A(n16732), .B(p_input[241]), .Z(n18380) );
  XOR U18260 ( .A(n18444), .B(n18395), .Z(n18389) );
  XNOR U18261 ( .A(p_input[2079]), .B(p_input[255]), .Z(n18395) );
  XOR U18262 ( .A(n18386), .B(n18394), .Z(n18444) );
  XOR U18263 ( .A(n18445), .B(n18391), .Z(n18394) );
  XOR U18264 ( .A(p_input[2077]), .B(p_input[253]), .Z(n18391) );
  XNOR U18265 ( .A(p_input[2078]), .B(p_input[254]), .Z(n18445) );
  XNOR U18266 ( .A(n16448), .B(p_input[249]), .Z(n18386) );
  XNOR U18267 ( .A(n18407), .B(n18406), .Z(n18373) );
  XNOR U18268 ( .A(n18446), .B(n18413), .Z(n18406) );
  XNOR U18269 ( .A(n18402), .B(n18401), .Z(n18413) );
  XOR U18270 ( .A(n18447), .B(n18398), .Z(n18401) );
  XNOR U18271 ( .A(n16737), .B(p_input[235]), .Z(n18398) );
  XNOR U18272 ( .A(p_input[2060]), .B(p_input[236]), .Z(n18447) );
  XOR U18273 ( .A(p_input[2061]), .B(p_input[237]), .Z(n18402) );
  XNOR U18274 ( .A(n18412), .B(n18403), .Z(n18446) );
  XNOR U18275 ( .A(n16452), .B(p_input[226]), .Z(n18403) );
  XOR U18276 ( .A(n18448), .B(n18418), .Z(n18412) );
  XNOR U18277 ( .A(p_input[2064]), .B(p_input[240]), .Z(n18418) );
  XOR U18278 ( .A(n18409), .B(n18417), .Z(n18448) );
  XOR U18279 ( .A(n18449), .B(n18414), .Z(n18417) );
  XOR U18280 ( .A(p_input[2062]), .B(p_input[238]), .Z(n18414) );
  XNOR U18281 ( .A(p_input[2063]), .B(p_input[239]), .Z(n18449) );
  XNOR U18282 ( .A(n16740), .B(p_input[234]), .Z(n18409) );
  XNOR U18283 ( .A(n18424), .B(n18423), .Z(n18407) );
  XNOR U18284 ( .A(n18450), .B(n18429), .Z(n18423) );
  XOR U18285 ( .A(p_input[2057]), .B(p_input[233]), .Z(n18429) );
  XOR U18286 ( .A(n18420), .B(n18428), .Z(n18450) );
  XOR U18287 ( .A(n18451), .B(n18425), .Z(n18428) );
  XOR U18288 ( .A(p_input[2055]), .B(p_input[231]), .Z(n18425) );
  XNOR U18289 ( .A(p_input[2056]), .B(p_input[232]), .Z(n18451) );
  XNOR U18290 ( .A(n16459), .B(p_input[227]), .Z(n18420) );
  XNOR U18291 ( .A(n18434), .B(n18433), .Z(n18424) );
  XOR U18292 ( .A(n18452), .B(n18430), .Z(n18433) );
  XOR U18293 ( .A(p_input[2052]), .B(p_input[228]), .Z(n18430) );
  XNOR U18294 ( .A(p_input[2053]), .B(p_input[229]), .Z(n18452) );
  XOR U18295 ( .A(p_input[2054]), .B(p_input[230]), .Z(n18434) );
  XNOR U18296 ( .A(n18453), .B(n18454), .Z(n18251) );
  AND U18297 ( .A(n144), .B(n18455), .Z(n18454) );
  XNOR U18298 ( .A(n18456), .B(n18457), .Z(n144) );
  AND U18299 ( .A(n18458), .B(n18459), .Z(n18457) );
  XOR U18300 ( .A(n18456), .B(n18261), .Z(n18459) );
  XNOR U18301 ( .A(n18456), .B(n18203), .Z(n18458) );
  XOR U18302 ( .A(n18460), .B(n18461), .Z(n18456) );
  AND U18303 ( .A(n18462), .B(n18463), .Z(n18461) );
  XNOR U18304 ( .A(n18274), .B(n18460), .Z(n18463) );
  XOR U18305 ( .A(n18460), .B(n18215), .Z(n18462) );
  XOR U18306 ( .A(n18464), .B(n18465), .Z(n18460) );
  AND U18307 ( .A(n18466), .B(n18467), .Z(n18465) );
  XNOR U18308 ( .A(n18299), .B(n18464), .Z(n18467) );
  XOR U18309 ( .A(n18464), .B(n18226), .Z(n18466) );
  XOR U18310 ( .A(n18468), .B(n18469), .Z(n18464) );
  AND U18311 ( .A(n18470), .B(n18471), .Z(n18469) );
  XOR U18312 ( .A(n18468), .B(n18236), .Z(n18470) );
  XOR U18313 ( .A(n18472), .B(n18473), .Z(n18192) );
  AND U18314 ( .A(n148), .B(n18455), .Z(n18473) );
  XNOR U18315 ( .A(n18453), .B(n18472), .Z(n18455) );
  XNOR U18316 ( .A(n18474), .B(n18475), .Z(n148) );
  AND U18317 ( .A(n18476), .B(n18477), .Z(n18475) );
  XNOR U18318 ( .A(n18478), .B(n18474), .Z(n18477) );
  IV U18319 ( .A(n18261), .Z(n18478) );
  XNOR U18320 ( .A(n18479), .B(n18480), .Z(n18261) );
  AND U18321 ( .A(n151), .B(n18481), .Z(n18480) );
  XNOR U18322 ( .A(n18479), .B(n18482), .Z(n18481) );
  XNOR U18323 ( .A(n18203), .B(n18474), .Z(n18476) );
  XOR U18324 ( .A(n18483), .B(n18484), .Z(n18203) );
  AND U18325 ( .A(n159), .B(n18485), .Z(n18484) );
  XOR U18326 ( .A(n18486), .B(n18487), .Z(n18474) );
  AND U18327 ( .A(n18488), .B(n18489), .Z(n18487) );
  XNOR U18328 ( .A(n18486), .B(n18274), .Z(n18489) );
  XNOR U18329 ( .A(n18490), .B(n18491), .Z(n18274) );
  AND U18330 ( .A(n151), .B(n18492), .Z(n18491) );
  XOR U18331 ( .A(n18493), .B(n18490), .Z(n18492) );
  XNOR U18332 ( .A(n18494), .B(n18486), .Z(n18488) );
  IV U18333 ( .A(n18215), .Z(n18494) );
  XOR U18334 ( .A(n18495), .B(n18496), .Z(n18215) );
  AND U18335 ( .A(n159), .B(n18497), .Z(n18496) );
  XOR U18336 ( .A(n18498), .B(n18499), .Z(n18486) );
  AND U18337 ( .A(n18500), .B(n18501), .Z(n18499) );
  XNOR U18338 ( .A(n18498), .B(n18299), .Z(n18501) );
  XNOR U18339 ( .A(n18502), .B(n18503), .Z(n18299) );
  AND U18340 ( .A(n151), .B(n18504), .Z(n18503) );
  XNOR U18341 ( .A(n18505), .B(n18502), .Z(n18504) );
  XOR U18342 ( .A(n18226), .B(n18498), .Z(n18500) );
  XOR U18343 ( .A(n18506), .B(n18507), .Z(n18226) );
  AND U18344 ( .A(n159), .B(n18508), .Z(n18507) );
  XOR U18345 ( .A(n18468), .B(n18509), .Z(n18498) );
  AND U18346 ( .A(n18510), .B(n18471), .Z(n18509) );
  XNOR U18347 ( .A(n18345), .B(n18468), .Z(n18471) );
  XNOR U18348 ( .A(n18511), .B(n18512), .Z(n18345) );
  AND U18349 ( .A(n151), .B(n18513), .Z(n18512) );
  XOR U18350 ( .A(n18514), .B(n18511), .Z(n18513) );
  XNOR U18351 ( .A(n18515), .B(n18468), .Z(n18510) );
  IV U18352 ( .A(n18236), .Z(n18515) );
  XOR U18353 ( .A(n18516), .B(n18517), .Z(n18236) );
  AND U18354 ( .A(n159), .B(n18518), .Z(n18517) );
  XOR U18355 ( .A(n18519), .B(n18520), .Z(n18468) );
  AND U18356 ( .A(n18521), .B(n18522), .Z(n18520) );
  XNOR U18357 ( .A(n18519), .B(n18435), .Z(n18522) );
  XNOR U18358 ( .A(n18523), .B(n18524), .Z(n18435) );
  AND U18359 ( .A(n151), .B(n18525), .Z(n18524) );
  XNOR U18360 ( .A(n18526), .B(n18523), .Z(n18525) );
  XNOR U18361 ( .A(n18527), .B(n18519), .Z(n18521) );
  IV U18362 ( .A(n18248), .Z(n18527) );
  XOR U18363 ( .A(n18528), .B(n18529), .Z(n18248) );
  AND U18364 ( .A(n159), .B(n18530), .Z(n18529) );
  AND U18365 ( .A(n18472), .B(n18453), .Z(n18519) );
  XNOR U18366 ( .A(n18531), .B(n18532), .Z(n18453) );
  AND U18367 ( .A(n151), .B(n18533), .Z(n18532) );
  XNOR U18368 ( .A(n18534), .B(n18531), .Z(n18533) );
  XNOR U18369 ( .A(n18535), .B(n18536), .Z(n151) );
  AND U18370 ( .A(n18537), .B(n18538), .Z(n18536) );
  XOR U18371 ( .A(n18482), .B(n18535), .Z(n18538) );
  AND U18372 ( .A(n18539), .B(n18540), .Z(n18482) );
  XOR U18373 ( .A(n18535), .B(n18479), .Z(n18537) );
  XNOR U18374 ( .A(n18541), .B(n18542), .Z(n18479) );
  AND U18375 ( .A(n155), .B(n18485), .Z(n18542) );
  XOR U18376 ( .A(n18483), .B(n18541), .Z(n18485) );
  XOR U18377 ( .A(n18543), .B(n18544), .Z(n18535) );
  AND U18378 ( .A(n18545), .B(n18546), .Z(n18544) );
  XNOR U18379 ( .A(n18543), .B(n18539), .Z(n18546) );
  IV U18380 ( .A(n18493), .Z(n18539) );
  XOR U18381 ( .A(n18547), .B(n18548), .Z(n18493) );
  XOR U18382 ( .A(n18549), .B(n18540), .Z(n18548) );
  AND U18383 ( .A(n18505), .B(n18550), .Z(n18540) );
  AND U18384 ( .A(n18551), .B(n18552), .Z(n18549) );
  XOR U18385 ( .A(n18553), .B(n18547), .Z(n18551) );
  XNOR U18386 ( .A(n18490), .B(n18543), .Z(n18545) );
  XNOR U18387 ( .A(n18554), .B(n18555), .Z(n18490) );
  AND U18388 ( .A(n155), .B(n18497), .Z(n18555) );
  XOR U18389 ( .A(n18554), .B(n18495), .Z(n18497) );
  XOR U18390 ( .A(n18556), .B(n18557), .Z(n18543) );
  AND U18391 ( .A(n18558), .B(n18559), .Z(n18557) );
  XNOR U18392 ( .A(n18556), .B(n18505), .Z(n18559) );
  XOR U18393 ( .A(n18560), .B(n18552), .Z(n18505) );
  XNOR U18394 ( .A(n18561), .B(n18547), .Z(n18552) );
  XOR U18395 ( .A(n18562), .B(n18563), .Z(n18547) );
  AND U18396 ( .A(n18564), .B(n18565), .Z(n18563) );
  XOR U18397 ( .A(n18566), .B(n18562), .Z(n18564) );
  XNOR U18398 ( .A(n18567), .B(n18568), .Z(n18561) );
  AND U18399 ( .A(n18569), .B(n18570), .Z(n18568) );
  XOR U18400 ( .A(n18567), .B(n18571), .Z(n18569) );
  XNOR U18401 ( .A(n18553), .B(n18550), .Z(n18560) );
  AND U18402 ( .A(n18572), .B(n18573), .Z(n18550) );
  XOR U18403 ( .A(n18574), .B(n18575), .Z(n18553) );
  AND U18404 ( .A(n18576), .B(n18577), .Z(n18575) );
  XOR U18405 ( .A(n18574), .B(n18578), .Z(n18576) );
  XNOR U18406 ( .A(n18502), .B(n18556), .Z(n18558) );
  XNOR U18407 ( .A(n18579), .B(n18580), .Z(n18502) );
  AND U18408 ( .A(n155), .B(n18508), .Z(n18580) );
  XOR U18409 ( .A(n18579), .B(n18506), .Z(n18508) );
  XOR U18410 ( .A(n18581), .B(n18582), .Z(n18556) );
  AND U18411 ( .A(n18583), .B(n18584), .Z(n18582) );
  XNOR U18412 ( .A(n18581), .B(n18572), .Z(n18584) );
  IV U18413 ( .A(n18514), .Z(n18572) );
  XNOR U18414 ( .A(n18585), .B(n18565), .Z(n18514) );
  XNOR U18415 ( .A(n18586), .B(n18571), .Z(n18565) );
  XOR U18416 ( .A(n18587), .B(n18588), .Z(n18571) );
  AND U18417 ( .A(n18589), .B(n18590), .Z(n18588) );
  XOR U18418 ( .A(n18587), .B(n18591), .Z(n18589) );
  XNOR U18419 ( .A(n18570), .B(n18562), .Z(n18586) );
  XOR U18420 ( .A(n18592), .B(n18593), .Z(n18562) );
  AND U18421 ( .A(n18594), .B(n18595), .Z(n18593) );
  XNOR U18422 ( .A(n18596), .B(n18592), .Z(n18594) );
  XNOR U18423 ( .A(n18597), .B(n18567), .Z(n18570) );
  XOR U18424 ( .A(n18598), .B(n18599), .Z(n18567) );
  AND U18425 ( .A(n18600), .B(n18601), .Z(n18599) );
  XOR U18426 ( .A(n18598), .B(n18602), .Z(n18600) );
  XNOR U18427 ( .A(n18603), .B(n18604), .Z(n18597) );
  AND U18428 ( .A(n18605), .B(n18606), .Z(n18604) );
  XNOR U18429 ( .A(n18603), .B(n18607), .Z(n18605) );
  XNOR U18430 ( .A(n18566), .B(n18573), .Z(n18585) );
  AND U18431 ( .A(n18526), .B(n18608), .Z(n18573) );
  XOR U18432 ( .A(n18578), .B(n18577), .Z(n18566) );
  XNOR U18433 ( .A(n18609), .B(n18574), .Z(n18577) );
  XOR U18434 ( .A(n18610), .B(n18611), .Z(n18574) );
  AND U18435 ( .A(n18612), .B(n18613), .Z(n18611) );
  XOR U18436 ( .A(n18610), .B(n18614), .Z(n18612) );
  XNOR U18437 ( .A(n18615), .B(n18616), .Z(n18609) );
  AND U18438 ( .A(n18617), .B(n18618), .Z(n18616) );
  XOR U18439 ( .A(n18615), .B(n18619), .Z(n18617) );
  XOR U18440 ( .A(n18620), .B(n18621), .Z(n18578) );
  AND U18441 ( .A(n18622), .B(n18623), .Z(n18621) );
  XOR U18442 ( .A(n18620), .B(n18624), .Z(n18622) );
  XNOR U18443 ( .A(n18511), .B(n18581), .Z(n18583) );
  XNOR U18444 ( .A(n18625), .B(n18626), .Z(n18511) );
  AND U18445 ( .A(n155), .B(n18518), .Z(n18626) );
  XOR U18446 ( .A(n18625), .B(n18516), .Z(n18518) );
  XOR U18447 ( .A(n18627), .B(n18628), .Z(n18581) );
  AND U18448 ( .A(n18629), .B(n18630), .Z(n18628) );
  XNOR U18449 ( .A(n18627), .B(n18526), .Z(n18630) );
  XOR U18450 ( .A(n18631), .B(n18595), .Z(n18526) );
  XNOR U18451 ( .A(n18632), .B(n18602), .Z(n18595) );
  XOR U18452 ( .A(n18591), .B(n18590), .Z(n18602) );
  XNOR U18453 ( .A(n18633), .B(n18587), .Z(n18590) );
  XOR U18454 ( .A(n18634), .B(n18635), .Z(n18587) );
  AND U18455 ( .A(n18636), .B(n18637), .Z(n18635) );
  XOR U18456 ( .A(n18634), .B(n18638), .Z(n18636) );
  XNOR U18457 ( .A(n18639), .B(n18640), .Z(n18633) );
  NOR U18458 ( .A(n18641), .B(n18642), .Z(n18640) );
  XNOR U18459 ( .A(n18639), .B(n18643), .Z(n18641) );
  XOR U18460 ( .A(n18644), .B(n18645), .Z(n18591) );
  NOR U18461 ( .A(n18646), .B(n18647), .Z(n18645) );
  XNOR U18462 ( .A(n18644), .B(n18648), .Z(n18646) );
  XNOR U18463 ( .A(n18601), .B(n18592), .Z(n18632) );
  XOR U18464 ( .A(n18649), .B(n18650), .Z(n18592) );
  NOR U18465 ( .A(n18651), .B(n18652), .Z(n18650) );
  XNOR U18466 ( .A(n18649), .B(n18653), .Z(n18651) );
  XOR U18467 ( .A(n18654), .B(n18607), .Z(n18601) );
  XNOR U18468 ( .A(n18655), .B(n18656), .Z(n18607) );
  NOR U18469 ( .A(n18657), .B(n18658), .Z(n18656) );
  XNOR U18470 ( .A(n18655), .B(n18659), .Z(n18657) );
  XNOR U18471 ( .A(n18606), .B(n18598), .Z(n18654) );
  XOR U18472 ( .A(n18660), .B(n18661), .Z(n18598) );
  AND U18473 ( .A(n18662), .B(n18663), .Z(n18661) );
  XOR U18474 ( .A(n18660), .B(n18664), .Z(n18662) );
  XNOR U18475 ( .A(n18665), .B(n18603), .Z(n18606) );
  XOR U18476 ( .A(n18666), .B(n18667), .Z(n18603) );
  AND U18477 ( .A(n18668), .B(n18669), .Z(n18667) );
  XOR U18478 ( .A(n18666), .B(n18670), .Z(n18668) );
  XNOR U18479 ( .A(n18671), .B(n18672), .Z(n18665) );
  NOR U18480 ( .A(n18673), .B(n18674), .Z(n18672) );
  XOR U18481 ( .A(n18671), .B(n18675), .Z(n18673) );
  XOR U18482 ( .A(n18596), .B(n18608), .Z(n18631) );
  NOR U18483 ( .A(n18534), .B(n18676), .Z(n18608) );
  XNOR U18484 ( .A(n18614), .B(n18613), .Z(n18596) );
  XNOR U18485 ( .A(n18677), .B(n18619), .Z(n18613) );
  XOR U18486 ( .A(n18678), .B(n18679), .Z(n18619) );
  NOR U18487 ( .A(n18680), .B(n18681), .Z(n18679) );
  XNOR U18488 ( .A(n18678), .B(n18682), .Z(n18680) );
  XNOR U18489 ( .A(n18618), .B(n18610), .Z(n18677) );
  XOR U18490 ( .A(n18683), .B(n18684), .Z(n18610) );
  AND U18491 ( .A(n18685), .B(n18686), .Z(n18684) );
  XNOR U18492 ( .A(n18683), .B(n18687), .Z(n18685) );
  XNOR U18493 ( .A(n18688), .B(n18615), .Z(n18618) );
  XOR U18494 ( .A(n18689), .B(n18690), .Z(n18615) );
  AND U18495 ( .A(n18691), .B(n18692), .Z(n18690) );
  XOR U18496 ( .A(n18689), .B(n18693), .Z(n18691) );
  XNOR U18497 ( .A(n18694), .B(n18695), .Z(n18688) );
  NOR U18498 ( .A(n18696), .B(n18697), .Z(n18695) );
  XOR U18499 ( .A(n18694), .B(n18698), .Z(n18696) );
  XOR U18500 ( .A(n18624), .B(n18623), .Z(n18614) );
  XNOR U18501 ( .A(n18699), .B(n18620), .Z(n18623) );
  XOR U18502 ( .A(n18700), .B(n18701), .Z(n18620) );
  AND U18503 ( .A(n18702), .B(n18703), .Z(n18701) );
  XOR U18504 ( .A(n18700), .B(n18704), .Z(n18702) );
  XNOR U18505 ( .A(n18705), .B(n18706), .Z(n18699) );
  NOR U18506 ( .A(n18707), .B(n18708), .Z(n18706) );
  XNOR U18507 ( .A(n18705), .B(n18709), .Z(n18707) );
  XOR U18508 ( .A(n18710), .B(n18711), .Z(n18624) );
  NOR U18509 ( .A(n18712), .B(n18713), .Z(n18711) );
  XNOR U18510 ( .A(n18710), .B(n18714), .Z(n18712) );
  XNOR U18511 ( .A(n18523), .B(n18627), .Z(n18629) );
  XNOR U18512 ( .A(n18715), .B(n18716), .Z(n18523) );
  AND U18513 ( .A(n155), .B(n18530), .Z(n18716) );
  XOR U18514 ( .A(n18715), .B(n18528), .Z(n18530) );
  AND U18515 ( .A(n18531), .B(n18534), .Z(n18627) );
  XOR U18516 ( .A(n18717), .B(n18676), .Z(n18534) );
  XNOR U18517 ( .A(p_input[2048]), .B(p_input[256]), .Z(n18676) );
  XOR U18518 ( .A(n18653), .B(n18652), .Z(n18717) );
  XOR U18519 ( .A(n18718), .B(n18664), .Z(n18652) );
  XOR U18520 ( .A(n18638), .B(n18637), .Z(n18664) );
  XNOR U18521 ( .A(n18719), .B(n18643), .Z(n18637) );
  XOR U18522 ( .A(p_input[2072]), .B(p_input[280]), .Z(n18643) );
  XOR U18523 ( .A(n18634), .B(n18642), .Z(n18719) );
  XOR U18524 ( .A(n18720), .B(n18639), .Z(n18642) );
  XOR U18525 ( .A(p_input[2070]), .B(p_input[278]), .Z(n18639) );
  XNOR U18526 ( .A(p_input[2071]), .B(p_input[279]), .Z(n18720) );
  XNOR U18527 ( .A(n16727), .B(p_input[274]), .Z(n18634) );
  XNOR U18528 ( .A(n18648), .B(n18647), .Z(n18638) );
  XOR U18529 ( .A(n18721), .B(n18644), .Z(n18647) );
  XOR U18530 ( .A(p_input[2067]), .B(p_input[275]), .Z(n18644) );
  XNOR U18531 ( .A(p_input[2068]), .B(p_input[276]), .Z(n18721) );
  XOR U18532 ( .A(p_input[2069]), .B(p_input[277]), .Z(n18648) );
  XNOR U18533 ( .A(n18663), .B(n18649), .Z(n18718) );
  XNOR U18534 ( .A(n16729), .B(p_input[257]), .Z(n18649) );
  XNOR U18535 ( .A(n18722), .B(n18670), .Z(n18663) );
  XNOR U18536 ( .A(n18659), .B(n18658), .Z(n18670) );
  XOR U18537 ( .A(n18723), .B(n18655), .Z(n18658) );
  XNOR U18538 ( .A(n16444), .B(p_input[282]), .Z(n18655) );
  XNOR U18539 ( .A(p_input[2075]), .B(p_input[283]), .Z(n18723) );
  XOR U18540 ( .A(p_input[2076]), .B(p_input[284]), .Z(n18659) );
  XNOR U18541 ( .A(n18669), .B(n18660), .Z(n18722) );
  XNOR U18542 ( .A(n16732), .B(p_input[273]), .Z(n18660) );
  XOR U18543 ( .A(n18724), .B(n18675), .Z(n18669) );
  XNOR U18544 ( .A(p_input[2079]), .B(p_input[287]), .Z(n18675) );
  XOR U18545 ( .A(n18666), .B(n18674), .Z(n18724) );
  XOR U18546 ( .A(n18725), .B(n18671), .Z(n18674) );
  XOR U18547 ( .A(p_input[2077]), .B(p_input[285]), .Z(n18671) );
  XNOR U18548 ( .A(p_input[2078]), .B(p_input[286]), .Z(n18725) );
  XNOR U18549 ( .A(n16448), .B(p_input[281]), .Z(n18666) );
  XNOR U18550 ( .A(n18687), .B(n18686), .Z(n18653) );
  XNOR U18551 ( .A(n18726), .B(n18693), .Z(n18686) );
  XNOR U18552 ( .A(n18682), .B(n18681), .Z(n18693) );
  XOR U18553 ( .A(n18727), .B(n18678), .Z(n18681) );
  XNOR U18554 ( .A(n16737), .B(p_input[267]), .Z(n18678) );
  XNOR U18555 ( .A(p_input[2060]), .B(p_input[268]), .Z(n18727) );
  XOR U18556 ( .A(p_input[2061]), .B(p_input[269]), .Z(n18682) );
  XNOR U18557 ( .A(n18692), .B(n18683), .Z(n18726) );
  XNOR U18558 ( .A(n16452), .B(p_input[258]), .Z(n18683) );
  XOR U18559 ( .A(n18728), .B(n18698), .Z(n18692) );
  XNOR U18560 ( .A(p_input[2064]), .B(p_input[272]), .Z(n18698) );
  XOR U18561 ( .A(n18689), .B(n18697), .Z(n18728) );
  XOR U18562 ( .A(n18729), .B(n18694), .Z(n18697) );
  XOR U18563 ( .A(p_input[2062]), .B(p_input[270]), .Z(n18694) );
  XNOR U18564 ( .A(p_input[2063]), .B(p_input[271]), .Z(n18729) );
  XNOR U18565 ( .A(n16740), .B(p_input[266]), .Z(n18689) );
  XNOR U18566 ( .A(n18704), .B(n18703), .Z(n18687) );
  XNOR U18567 ( .A(n18730), .B(n18709), .Z(n18703) );
  XOR U18568 ( .A(p_input[2057]), .B(p_input[265]), .Z(n18709) );
  XOR U18569 ( .A(n18700), .B(n18708), .Z(n18730) );
  XOR U18570 ( .A(n18731), .B(n18705), .Z(n18708) );
  XOR U18571 ( .A(p_input[2055]), .B(p_input[263]), .Z(n18705) );
  XNOR U18572 ( .A(p_input[2056]), .B(p_input[264]), .Z(n18731) );
  XNOR U18573 ( .A(n16459), .B(p_input[259]), .Z(n18700) );
  XNOR U18574 ( .A(n18714), .B(n18713), .Z(n18704) );
  XOR U18575 ( .A(n18732), .B(n18710), .Z(n18713) );
  XOR U18576 ( .A(p_input[2052]), .B(p_input[260]), .Z(n18710) );
  XNOR U18577 ( .A(p_input[2053]), .B(p_input[261]), .Z(n18732) );
  XOR U18578 ( .A(p_input[2054]), .B(p_input[262]), .Z(n18714) );
  XNOR U18579 ( .A(n18733), .B(n18734), .Z(n18531) );
  AND U18580 ( .A(n155), .B(n18735), .Z(n18734) );
  XNOR U18581 ( .A(n18736), .B(n18737), .Z(n155) );
  AND U18582 ( .A(n18738), .B(n18739), .Z(n18737) );
  XOR U18583 ( .A(n18736), .B(n18541), .Z(n18739) );
  XNOR U18584 ( .A(n18736), .B(n18483), .Z(n18738) );
  XOR U18585 ( .A(n18740), .B(n18741), .Z(n18736) );
  AND U18586 ( .A(n18742), .B(n18743), .Z(n18741) );
  XNOR U18587 ( .A(n18554), .B(n18740), .Z(n18743) );
  XOR U18588 ( .A(n18740), .B(n18495), .Z(n18742) );
  XOR U18589 ( .A(n18744), .B(n18745), .Z(n18740) );
  AND U18590 ( .A(n18746), .B(n18747), .Z(n18745) );
  XNOR U18591 ( .A(n18579), .B(n18744), .Z(n18747) );
  XOR U18592 ( .A(n18744), .B(n18506), .Z(n18746) );
  XOR U18593 ( .A(n18748), .B(n18749), .Z(n18744) );
  AND U18594 ( .A(n18750), .B(n18751), .Z(n18749) );
  XOR U18595 ( .A(n18748), .B(n18516), .Z(n18750) );
  XOR U18596 ( .A(n18752), .B(n18753), .Z(n18472) );
  AND U18597 ( .A(n159), .B(n18735), .Z(n18753) );
  XNOR U18598 ( .A(n18733), .B(n18752), .Z(n18735) );
  XNOR U18599 ( .A(n18754), .B(n18755), .Z(n159) );
  AND U18600 ( .A(n18756), .B(n18757), .Z(n18755) );
  XNOR U18601 ( .A(n18758), .B(n18754), .Z(n18757) );
  IV U18602 ( .A(n18541), .Z(n18758) );
  XNOR U18603 ( .A(n18759), .B(n18760), .Z(n18541) );
  AND U18604 ( .A(n162), .B(n18761), .Z(n18760) );
  XNOR U18605 ( .A(n18759), .B(n18762), .Z(n18761) );
  XNOR U18606 ( .A(n18483), .B(n18754), .Z(n18756) );
  XOR U18607 ( .A(n18763), .B(n18764), .Z(n18483) );
  AND U18608 ( .A(n170), .B(n18765), .Z(n18764) );
  XOR U18609 ( .A(n18766), .B(n18767), .Z(n18754) );
  AND U18610 ( .A(n18768), .B(n18769), .Z(n18767) );
  XNOR U18611 ( .A(n18766), .B(n18554), .Z(n18769) );
  XNOR U18612 ( .A(n18770), .B(n18771), .Z(n18554) );
  AND U18613 ( .A(n162), .B(n18772), .Z(n18771) );
  XOR U18614 ( .A(n18773), .B(n18770), .Z(n18772) );
  XNOR U18615 ( .A(n18774), .B(n18766), .Z(n18768) );
  IV U18616 ( .A(n18495), .Z(n18774) );
  XOR U18617 ( .A(n18775), .B(n18776), .Z(n18495) );
  AND U18618 ( .A(n170), .B(n18777), .Z(n18776) );
  XOR U18619 ( .A(n18778), .B(n18779), .Z(n18766) );
  AND U18620 ( .A(n18780), .B(n18781), .Z(n18779) );
  XNOR U18621 ( .A(n18778), .B(n18579), .Z(n18781) );
  XNOR U18622 ( .A(n18782), .B(n18783), .Z(n18579) );
  AND U18623 ( .A(n162), .B(n18784), .Z(n18783) );
  XNOR U18624 ( .A(n18785), .B(n18782), .Z(n18784) );
  XOR U18625 ( .A(n18506), .B(n18778), .Z(n18780) );
  XOR U18626 ( .A(n18786), .B(n18787), .Z(n18506) );
  AND U18627 ( .A(n170), .B(n18788), .Z(n18787) );
  XOR U18628 ( .A(n18748), .B(n18789), .Z(n18778) );
  AND U18629 ( .A(n18790), .B(n18751), .Z(n18789) );
  XNOR U18630 ( .A(n18625), .B(n18748), .Z(n18751) );
  XNOR U18631 ( .A(n18791), .B(n18792), .Z(n18625) );
  AND U18632 ( .A(n162), .B(n18793), .Z(n18792) );
  XOR U18633 ( .A(n18794), .B(n18791), .Z(n18793) );
  XNOR U18634 ( .A(n18795), .B(n18748), .Z(n18790) );
  IV U18635 ( .A(n18516), .Z(n18795) );
  XOR U18636 ( .A(n18796), .B(n18797), .Z(n18516) );
  AND U18637 ( .A(n170), .B(n18798), .Z(n18797) );
  XOR U18638 ( .A(n18799), .B(n18800), .Z(n18748) );
  AND U18639 ( .A(n18801), .B(n18802), .Z(n18800) );
  XNOR U18640 ( .A(n18799), .B(n18715), .Z(n18802) );
  XNOR U18641 ( .A(n18803), .B(n18804), .Z(n18715) );
  AND U18642 ( .A(n162), .B(n18805), .Z(n18804) );
  XNOR U18643 ( .A(n18806), .B(n18803), .Z(n18805) );
  XNOR U18644 ( .A(n18807), .B(n18799), .Z(n18801) );
  IV U18645 ( .A(n18528), .Z(n18807) );
  XOR U18646 ( .A(n18808), .B(n18809), .Z(n18528) );
  AND U18647 ( .A(n170), .B(n18810), .Z(n18809) );
  AND U18648 ( .A(n18752), .B(n18733), .Z(n18799) );
  XNOR U18649 ( .A(n18811), .B(n18812), .Z(n18733) );
  AND U18650 ( .A(n162), .B(n18813), .Z(n18812) );
  XNOR U18651 ( .A(n18814), .B(n18811), .Z(n18813) );
  XNOR U18652 ( .A(n18815), .B(n18816), .Z(n162) );
  AND U18653 ( .A(n18817), .B(n18818), .Z(n18816) );
  XOR U18654 ( .A(n18762), .B(n18815), .Z(n18818) );
  AND U18655 ( .A(n18819), .B(n18820), .Z(n18762) );
  XOR U18656 ( .A(n18815), .B(n18759), .Z(n18817) );
  XNOR U18657 ( .A(n18821), .B(n18822), .Z(n18759) );
  AND U18658 ( .A(n166), .B(n18765), .Z(n18822) );
  XOR U18659 ( .A(n18763), .B(n18821), .Z(n18765) );
  XOR U18660 ( .A(n18823), .B(n18824), .Z(n18815) );
  AND U18661 ( .A(n18825), .B(n18826), .Z(n18824) );
  XNOR U18662 ( .A(n18823), .B(n18819), .Z(n18826) );
  IV U18663 ( .A(n18773), .Z(n18819) );
  XOR U18664 ( .A(n18827), .B(n18828), .Z(n18773) );
  XOR U18665 ( .A(n18829), .B(n18820), .Z(n18828) );
  AND U18666 ( .A(n18785), .B(n18830), .Z(n18820) );
  AND U18667 ( .A(n18831), .B(n18832), .Z(n18829) );
  XOR U18668 ( .A(n18833), .B(n18827), .Z(n18831) );
  XNOR U18669 ( .A(n18770), .B(n18823), .Z(n18825) );
  XNOR U18670 ( .A(n18834), .B(n18835), .Z(n18770) );
  AND U18671 ( .A(n166), .B(n18777), .Z(n18835) );
  XOR U18672 ( .A(n18834), .B(n18775), .Z(n18777) );
  XOR U18673 ( .A(n18836), .B(n18837), .Z(n18823) );
  AND U18674 ( .A(n18838), .B(n18839), .Z(n18837) );
  XNOR U18675 ( .A(n18836), .B(n18785), .Z(n18839) );
  XOR U18676 ( .A(n18840), .B(n18832), .Z(n18785) );
  XNOR U18677 ( .A(n18841), .B(n18827), .Z(n18832) );
  XOR U18678 ( .A(n18842), .B(n18843), .Z(n18827) );
  AND U18679 ( .A(n18844), .B(n18845), .Z(n18843) );
  XOR U18680 ( .A(n18846), .B(n18842), .Z(n18844) );
  XNOR U18681 ( .A(n18847), .B(n18848), .Z(n18841) );
  AND U18682 ( .A(n18849), .B(n18850), .Z(n18848) );
  XOR U18683 ( .A(n18847), .B(n18851), .Z(n18849) );
  XNOR U18684 ( .A(n18833), .B(n18830), .Z(n18840) );
  AND U18685 ( .A(n18852), .B(n18853), .Z(n18830) );
  XOR U18686 ( .A(n18854), .B(n18855), .Z(n18833) );
  AND U18687 ( .A(n18856), .B(n18857), .Z(n18855) );
  XOR U18688 ( .A(n18854), .B(n18858), .Z(n18856) );
  XNOR U18689 ( .A(n18782), .B(n18836), .Z(n18838) );
  XNOR U18690 ( .A(n18859), .B(n18860), .Z(n18782) );
  AND U18691 ( .A(n166), .B(n18788), .Z(n18860) );
  XOR U18692 ( .A(n18859), .B(n18786), .Z(n18788) );
  XOR U18693 ( .A(n18861), .B(n18862), .Z(n18836) );
  AND U18694 ( .A(n18863), .B(n18864), .Z(n18862) );
  XNOR U18695 ( .A(n18861), .B(n18852), .Z(n18864) );
  IV U18696 ( .A(n18794), .Z(n18852) );
  XNOR U18697 ( .A(n18865), .B(n18845), .Z(n18794) );
  XNOR U18698 ( .A(n18866), .B(n18851), .Z(n18845) );
  XOR U18699 ( .A(n18867), .B(n18868), .Z(n18851) );
  AND U18700 ( .A(n18869), .B(n18870), .Z(n18868) );
  XOR U18701 ( .A(n18867), .B(n18871), .Z(n18869) );
  XNOR U18702 ( .A(n18850), .B(n18842), .Z(n18866) );
  XOR U18703 ( .A(n18872), .B(n18873), .Z(n18842) );
  AND U18704 ( .A(n18874), .B(n18875), .Z(n18873) );
  XNOR U18705 ( .A(n18876), .B(n18872), .Z(n18874) );
  XNOR U18706 ( .A(n18877), .B(n18847), .Z(n18850) );
  XOR U18707 ( .A(n18878), .B(n18879), .Z(n18847) );
  AND U18708 ( .A(n18880), .B(n18881), .Z(n18879) );
  XOR U18709 ( .A(n18878), .B(n18882), .Z(n18880) );
  XNOR U18710 ( .A(n18883), .B(n18884), .Z(n18877) );
  AND U18711 ( .A(n18885), .B(n18886), .Z(n18884) );
  XNOR U18712 ( .A(n18883), .B(n18887), .Z(n18885) );
  XNOR U18713 ( .A(n18846), .B(n18853), .Z(n18865) );
  AND U18714 ( .A(n18806), .B(n18888), .Z(n18853) );
  XOR U18715 ( .A(n18858), .B(n18857), .Z(n18846) );
  XNOR U18716 ( .A(n18889), .B(n18854), .Z(n18857) );
  XOR U18717 ( .A(n18890), .B(n18891), .Z(n18854) );
  AND U18718 ( .A(n18892), .B(n18893), .Z(n18891) );
  XOR U18719 ( .A(n18890), .B(n18894), .Z(n18892) );
  XNOR U18720 ( .A(n18895), .B(n18896), .Z(n18889) );
  AND U18721 ( .A(n18897), .B(n18898), .Z(n18896) );
  XOR U18722 ( .A(n18895), .B(n18899), .Z(n18897) );
  XOR U18723 ( .A(n18900), .B(n18901), .Z(n18858) );
  AND U18724 ( .A(n18902), .B(n18903), .Z(n18901) );
  XOR U18725 ( .A(n18900), .B(n18904), .Z(n18902) );
  XNOR U18726 ( .A(n18791), .B(n18861), .Z(n18863) );
  XNOR U18727 ( .A(n18905), .B(n18906), .Z(n18791) );
  AND U18728 ( .A(n166), .B(n18798), .Z(n18906) );
  XOR U18729 ( .A(n18905), .B(n18796), .Z(n18798) );
  XOR U18730 ( .A(n18907), .B(n18908), .Z(n18861) );
  AND U18731 ( .A(n18909), .B(n18910), .Z(n18908) );
  XNOR U18732 ( .A(n18907), .B(n18806), .Z(n18910) );
  XOR U18733 ( .A(n18911), .B(n18875), .Z(n18806) );
  XNOR U18734 ( .A(n18912), .B(n18882), .Z(n18875) );
  XOR U18735 ( .A(n18871), .B(n18870), .Z(n18882) );
  XNOR U18736 ( .A(n18913), .B(n18867), .Z(n18870) );
  XOR U18737 ( .A(n18914), .B(n18915), .Z(n18867) );
  AND U18738 ( .A(n18916), .B(n18917), .Z(n18915) );
  XOR U18739 ( .A(n18914), .B(n18918), .Z(n18916) );
  XNOR U18740 ( .A(n18919), .B(n18920), .Z(n18913) );
  NOR U18741 ( .A(n18921), .B(n18922), .Z(n18920) );
  XNOR U18742 ( .A(n18919), .B(n18923), .Z(n18921) );
  XOR U18743 ( .A(n18924), .B(n18925), .Z(n18871) );
  NOR U18744 ( .A(n18926), .B(n18927), .Z(n18925) );
  XNOR U18745 ( .A(n18924), .B(n18928), .Z(n18926) );
  XNOR U18746 ( .A(n18881), .B(n18872), .Z(n18912) );
  XOR U18747 ( .A(n18929), .B(n18930), .Z(n18872) );
  NOR U18748 ( .A(n18931), .B(n18932), .Z(n18930) );
  XNOR U18749 ( .A(n18929), .B(n18933), .Z(n18931) );
  XOR U18750 ( .A(n18934), .B(n18887), .Z(n18881) );
  XNOR U18751 ( .A(n18935), .B(n18936), .Z(n18887) );
  NOR U18752 ( .A(n18937), .B(n18938), .Z(n18936) );
  XNOR U18753 ( .A(n18935), .B(n18939), .Z(n18937) );
  XNOR U18754 ( .A(n18886), .B(n18878), .Z(n18934) );
  XOR U18755 ( .A(n18940), .B(n18941), .Z(n18878) );
  AND U18756 ( .A(n18942), .B(n18943), .Z(n18941) );
  XOR U18757 ( .A(n18940), .B(n18944), .Z(n18942) );
  XNOR U18758 ( .A(n18945), .B(n18883), .Z(n18886) );
  XOR U18759 ( .A(n18946), .B(n18947), .Z(n18883) );
  AND U18760 ( .A(n18948), .B(n18949), .Z(n18947) );
  XOR U18761 ( .A(n18946), .B(n18950), .Z(n18948) );
  XNOR U18762 ( .A(n18951), .B(n18952), .Z(n18945) );
  NOR U18763 ( .A(n18953), .B(n18954), .Z(n18952) );
  XOR U18764 ( .A(n18951), .B(n18955), .Z(n18953) );
  XOR U18765 ( .A(n18876), .B(n18888), .Z(n18911) );
  NOR U18766 ( .A(n18814), .B(n18956), .Z(n18888) );
  XNOR U18767 ( .A(n18894), .B(n18893), .Z(n18876) );
  XNOR U18768 ( .A(n18957), .B(n18899), .Z(n18893) );
  XOR U18769 ( .A(n18958), .B(n18959), .Z(n18899) );
  NOR U18770 ( .A(n18960), .B(n18961), .Z(n18959) );
  XNOR U18771 ( .A(n18958), .B(n18962), .Z(n18960) );
  XNOR U18772 ( .A(n18898), .B(n18890), .Z(n18957) );
  XOR U18773 ( .A(n18963), .B(n18964), .Z(n18890) );
  AND U18774 ( .A(n18965), .B(n18966), .Z(n18964) );
  XNOR U18775 ( .A(n18963), .B(n18967), .Z(n18965) );
  XNOR U18776 ( .A(n18968), .B(n18895), .Z(n18898) );
  XOR U18777 ( .A(n18969), .B(n18970), .Z(n18895) );
  AND U18778 ( .A(n18971), .B(n18972), .Z(n18970) );
  XOR U18779 ( .A(n18969), .B(n18973), .Z(n18971) );
  XNOR U18780 ( .A(n18974), .B(n18975), .Z(n18968) );
  NOR U18781 ( .A(n18976), .B(n18977), .Z(n18975) );
  XOR U18782 ( .A(n18974), .B(n18978), .Z(n18976) );
  XOR U18783 ( .A(n18904), .B(n18903), .Z(n18894) );
  XNOR U18784 ( .A(n18979), .B(n18900), .Z(n18903) );
  XOR U18785 ( .A(n18980), .B(n18981), .Z(n18900) );
  AND U18786 ( .A(n18982), .B(n18983), .Z(n18981) );
  XOR U18787 ( .A(n18980), .B(n18984), .Z(n18982) );
  XNOR U18788 ( .A(n18985), .B(n18986), .Z(n18979) );
  NOR U18789 ( .A(n18987), .B(n18988), .Z(n18986) );
  XNOR U18790 ( .A(n18985), .B(n18989), .Z(n18987) );
  XOR U18791 ( .A(n18990), .B(n18991), .Z(n18904) );
  NOR U18792 ( .A(n18992), .B(n18993), .Z(n18991) );
  XNOR U18793 ( .A(n18990), .B(n18994), .Z(n18992) );
  XNOR U18794 ( .A(n18803), .B(n18907), .Z(n18909) );
  XNOR U18795 ( .A(n18995), .B(n18996), .Z(n18803) );
  AND U18796 ( .A(n166), .B(n18810), .Z(n18996) );
  XOR U18797 ( .A(n18995), .B(n18808), .Z(n18810) );
  AND U18798 ( .A(n18811), .B(n18814), .Z(n18907) );
  XOR U18799 ( .A(n18997), .B(n18956), .Z(n18814) );
  XNOR U18800 ( .A(p_input[2048]), .B(p_input[288]), .Z(n18956) );
  XOR U18801 ( .A(n18933), .B(n18932), .Z(n18997) );
  XOR U18802 ( .A(n18998), .B(n18944), .Z(n18932) );
  XOR U18803 ( .A(n18918), .B(n18917), .Z(n18944) );
  XNOR U18804 ( .A(n18999), .B(n18923), .Z(n18917) );
  XOR U18805 ( .A(p_input[2072]), .B(p_input[312]), .Z(n18923) );
  XOR U18806 ( .A(n18914), .B(n18922), .Z(n18999) );
  XOR U18807 ( .A(n19000), .B(n18919), .Z(n18922) );
  XOR U18808 ( .A(p_input[2070]), .B(p_input[310]), .Z(n18919) );
  XNOR U18809 ( .A(p_input[2071]), .B(p_input[311]), .Z(n19000) );
  XNOR U18810 ( .A(n16727), .B(p_input[306]), .Z(n18914) );
  XNOR U18811 ( .A(n18928), .B(n18927), .Z(n18918) );
  XOR U18812 ( .A(n19001), .B(n18924), .Z(n18927) );
  XOR U18813 ( .A(p_input[2067]), .B(p_input[307]), .Z(n18924) );
  XNOR U18814 ( .A(p_input[2068]), .B(p_input[308]), .Z(n19001) );
  XOR U18815 ( .A(p_input[2069]), .B(p_input[309]), .Z(n18928) );
  XNOR U18816 ( .A(n18943), .B(n18929), .Z(n18998) );
  XNOR U18817 ( .A(n16729), .B(p_input[289]), .Z(n18929) );
  XNOR U18818 ( .A(n19002), .B(n18950), .Z(n18943) );
  XNOR U18819 ( .A(n18939), .B(n18938), .Z(n18950) );
  XOR U18820 ( .A(n19003), .B(n18935), .Z(n18938) );
  XNOR U18821 ( .A(n16444), .B(p_input[314]), .Z(n18935) );
  XNOR U18822 ( .A(p_input[2075]), .B(p_input[315]), .Z(n19003) );
  XOR U18823 ( .A(p_input[2076]), .B(p_input[316]), .Z(n18939) );
  XNOR U18824 ( .A(n18949), .B(n18940), .Z(n19002) );
  XNOR U18825 ( .A(n16732), .B(p_input[305]), .Z(n18940) );
  XOR U18826 ( .A(n19004), .B(n18955), .Z(n18949) );
  XNOR U18827 ( .A(p_input[2079]), .B(p_input[319]), .Z(n18955) );
  XOR U18828 ( .A(n18946), .B(n18954), .Z(n19004) );
  XOR U18829 ( .A(n19005), .B(n18951), .Z(n18954) );
  XOR U18830 ( .A(p_input[2077]), .B(p_input[317]), .Z(n18951) );
  XNOR U18831 ( .A(p_input[2078]), .B(p_input[318]), .Z(n19005) );
  XNOR U18832 ( .A(n16448), .B(p_input[313]), .Z(n18946) );
  XNOR U18833 ( .A(n18967), .B(n18966), .Z(n18933) );
  XNOR U18834 ( .A(n19006), .B(n18973), .Z(n18966) );
  XNOR U18835 ( .A(n18962), .B(n18961), .Z(n18973) );
  XOR U18836 ( .A(n19007), .B(n18958), .Z(n18961) );
  XNOR U18837 ( .A(n16737), .B(p_input[299]), .Z(n18958) );
  XNOR U18838 ( .A(p_input[2060]), .B(p_input[300]), .Z(n19007) );
  XOR U18839 ( .A(p_input[2061]), .B(p_input[301]), .Z(n18962) );
  XNOR U18840 ( .A(n18972), .B(n18963), .Z(n19006) );
  XNOR U18841 ( .A(n16452), .B(p_input[290]), .Z(n18963) );
  XOR U18842 ( .A(n19008), .B(n18978), .Z(n18972) );
  XNOR U18843 ( .A(p_input[2064]), .B(p_input[304]), .Z(n18978) );
  XOR U18844 ( .A(n18969), .B(n18977), .Z(n19008) );
  XOR U18845 ( .A(n19009), .B(n18974), .Z(n18977) );
  XOR U18846 ( .A(p_input[2062]), .B(p_input[302]), .Z(n18974) );
  XNOR U18847 ( .A(p_input[2063]), .B(p_input[303]), .Z(n19009) );
  XNOR U18848 ( .A(n16740), .B(p_input[298]), .Z(n18969) );
  XNOR U18849 ( .A(n18984), .B(n18983), .Z(n18967) );
  XNOR U18850 ( .A(n19010), .B(n18989), .Z(n18983) );
  XOR U18851 ( .A(p_input[2057]), .B(p_input[297]), .Z(n18989) );
  XOR U18852 ( .A(n18980), .B(n18988), .Z(n19010) );
  XOR U18853 ( .A(n19011), .B(n18985), .Z(n18988) );
  XOR U18854 ( .A(p_input[2055]), .B(p_input[295]), .Z(n18985) );
  XNOR U18855 ( .A(p_input[2056]), .B(p_input[296]), .Z(n19011) );
  XNOR U18856 ( .A(n16459), .B(p_input[291]), .Z(n18980) );
  XNOR U18857 ( .A(n18994), .B(n18993), .Z(n18984) );
  XOR U18858 ( .A(n19012), .B(n18990), .Z(n18993) );
  XOR U18859 ( .A(p_input[2052]), .B(p_input[292]), .Z(n18990) );
  XNOR U18860 ( .A(p_input[2053]), .B(p_input[293]), .Z(n19012) );
  XOR U18861 ( .A(p_input[2054]), .B(p_input[294]), .Z(n18994) );
  XNOR U18862 ( .A(n19013), .B(n19014), .Z(n18811) );
  AND U18863 ( .A(n166), .B(n19015), .Z(n19014) );
  XNOR U18864 ( .A(n19016), .B(n19017), .Z(n166) );
  AND U18865 ( .A(n19018), .B(n19019), .Z(n19017) );
  XOR U18866 ( .A(n19016), .B(n18821), .Z(n19019) );
  XNOR U18867 ( .A(n19016), .B(n18763), .Z(n19018) );
  XOR U18868 ( .A(n19020), .B(n19021), .Z(n19016) );
  AND U18869 ( .A(n19022), .B(n19023), .Z(n19021) );
  XNOR U18870 ( .A(n18834), .B(n19020), .Z(n19023) );
  XOR U18871 ( .A(n19020), .B(n18775), .Z(n19022) );
  XOR U18872 ( .A(n19024), .B(n19025), .Z(n19020) );
  AND U18873 ( .A(n19026), .B(n19027), .Z(n19025) );
  XNOR U18874 ( .A(n18859), .B(n19024), .Z(n19027) );
  XOR U18875 ( .A(n19024), .B(n18786), .Z(n19026) );
  XOR U18876 ( .A(n19028), .B(n19029), .Z(n19024) );
  AND U18877 ( .A(n19030), .B(n19031), .Z(n19029) );
  XOR U18878 ( .A(n19028), .B(n18796), .Z(n19030) );
  XOR U18879 ( .A(n19032), .B(n19033), .Z(n18752) );
  AND U18880 ( .A(n170), .B(n19015), .Z(n19033) );
  XNOR U18881 ( .A(n19013), .B(n19032), .Z(n19015) );
  XNOR U18882 ( .A(n19034), .B(n19035), .Z(n170) );
  AND U18883 ( .A(n19036), .B(n19037), .Z(n19035) );
  XNOR U18884 ( .A(n19038), .B(n19034), .Z(n19037) );
  IV U18885 ( .A(n18821), .Z(n19038) );
  XNOR U18886 ( .A(n19039), .B(n19040), .Z(n18821) );
  AND U18887 ( .A(n173), .B(n19041), .Z(n19040) );
  XNOR U18888 ( .A(n19039), .B(n19042), .Z(n19041) );
  XNOR U18889 ( .A(n18763), .B(n19034), .Z(n19036) );
  XOR U18890 ( .A(n19043), .B(n19044), .Z(n18763) );
  AND U18891 ( .A(n181), .B(n19045), .Z(n19044) );
  XOR U18892 ( .A(n19046), .B(n19047), .Z(n19034) );
  AND U18893 ( .A(n19048), .B(n19049), .Z(n19047) );
  XNOR U18894 ( .A(n19046), .B(n18834), .Z(n19049) );
  XNOR U18895 ( .A(n19050), .B(n19051), .Z(n18834) );
  AND U18896 ( .A(n173), .B(n19052), .Z(n19051) );
  XOR U18897 ( .A(n19053), .B(n19050), .Z(n19052) );
  XNOR U18898 ( .A(n19054), .B(n19046), .Z(n19048) );
  IV U18899 ( .A(n18775), .Z(n19054) );
  XOR U18900 ( .A(n19055), .B(n19056), .Z(n18775) );
  AND U18901 ( .A(n181), .B(n19057), .Z(n19056) );
  XOR U18902 ( .A(n19058), .B(n19059), .Z(n19046) );
  AND U18903 ( .A(n19060), .B(n19061), .Z(n19059) );
  XNOR U18904 ( .A(n19058), .B(n18859), .Z(n19061) );
  XNOR U18905 ( .A(n19062), .B(n19063), .Z(n18859) );
  AND U18906 ( .A(n173), .B(n19064), .Z(n19063) );
  XNOR U18907 ( .A(n19065), .B(n19062), .Z(n19064) );
  XOR U18908 ( .A(n18786), .B(n19058), .Z(n19060) );
  XOR U18909 ( .A(n19066), .B(n19067), .Z(n18786) );
  AND U18910 ( .A(n181), .B(n19068), .Z(n19067) );
  XOR U18911 ( .A(n19028), .B(n19069), .Z(n19058) );
  AND U18912 ( .A(n19070), .B(n19031), .Z(n19069) );
  XNOR U18913 ( .A(n18905), .B(n19028), .Z(n19031) );
  XNOR U18914 ( .A(n19071), .B(n19072), .Z(n18905) );
  AND U18915 ( .A(n173), .B(n19073), .Z(n19072) );
  XOR U18916 ( .A(n19074), .B(n19071), .Z(n19073) );
  XNOR U18917 ( .A(n19075), .B(n19028), .Z(n19070) );
  IV U18918 ( .A(n18796), .Z(n19075) );
  XOR U18919 ( .A(n19076), .B(n19077), .Z(n18796) );
  AND U18920 ( .A(n181), .B(n19078), .Z(n19077) );
  XOR U18921 ( .A(n19079), .B(n19080), .Z(n19028) );
  AND U18922 ( .A(n19081), .B(n19082), .Z(n19080) );
  XNOR U18923 ( .A(n19079), .B(n18995), .Z(n19082) );
  XNOR U18924 ( .A(n19083), .B(n19084), .Z(n18995) );
  AND U18925 ( .A(n173), .B(n19085), .Z(n19084) );
  XNOR U18926 ( .A(n19086), .B(n19083), .Z(n19085) );
  XNOR U18927 ( .A(n19087), .B(n19079), .Z(n19081) );
  IV U18928 ( .A(n18808), .Z(n19087) );
  XOR U18929 ( .A(n19088), .B(n19089), .Z(n18808) );
  AND U18930 ( .A(n181), .B(n19090), .Z(n19089) );
  AND U18931 ( .A(n19032), .B(n19013), .Z(n19079) );
  XNOR U18932 ( .A(n19091), .B(n19092), .Z(n19013) );
  AND U18933 ( .A(n173), .B(n19093), .Z(n19092) );
  XNOR U18934 ( .A(n19094), .B(n19091), .Z(n19093) );
  XNOR U18935 ( .A(n19095), .B(n19096), .Z(n173) );
  AND U18936 ( .A(n19097), .B(n19098), .Z(n19096) );
  XOR U18937 ( .A(n19042), .B(n19095), .Z(n19098) );
  AND U18938 ( .A(n19099), .B(n19100), .Z(n19042) );
  XOR U18939 ( .A(n19095), .B(n19039), .Z(n19097) );
  XNOR U18940 ( .A(n19101), .B(n19102), .Z(n19039) );
  AND U18941 ( .A(n177), .B(n19045), .Z(n19102) );
  XOR U18942 ( .A(n19043), .B(n19101), .Z(n19045) );
  XOR U18943 ( .A(n19103), .B(n19104), .Z(n19095) );
  AND U18944 ( .A(n19105), .B(n19106), .Z(n19104) );
  XNOR U18945 ( .A(n19103), .B(n19099), .Z(n19106) );
  IV U18946 ( .A(n19053), .Z(n19099) );
  XOR U18947 ( .A(n19107), .B(n19108), .Z(n19053) );
  XOR U18948 ( .A(n19109), .B(n19100), .Z(n19108) );
  AND U18949 ( .A(n19065), .B(n19110), .Z(n19100) );
  AND U18950 ( .A(n19111), .B(n19112), .Z(n19109) );
  XOR U18951 ( .A(n19113), .B(n19107), .Z(n19111) );
  XNOR U18952 ( .A(n19050), .B(n19103), .Z(n19105) );
  XNOR U18953 ( .A(n19114), .B(n19115), .Z(n19050) );
  AND U18954 ( .A(n177), .B(n19057), .Z(n19115) );
  XOR U18955 ( .A(n19114), .B(n19055), .Z(n19057) );
  XOR U18956 ( .A(n19116), .B(n19117), .Z(n19103) );
  AND U18957 ( .A(n19118), .B(n19119), .Z(n19117) );
  XNOR U18958 ( .A(n19116), .B(n19065), .Z(n19119) );
  XOR U18959 ( .A(n19120), .B(n19112), .Z(n19065) );
  XNOR U18960 ( .A(n19121), .B(n19107), .Z(n19112) );
  XOR U18961 ( .A(n19122), .B(n19123), .Z(n19107) );
  AND U18962 ( .A(n19124), .B(n19125), .Z(n19123) );
  XOR U18963 ( .A(n19126), .B(n19122), .Z(n19124) );
  XNOR U18964 ( .A(n19127), .B(n19128), .Z(n19121) );
  AND U18965 ( .A(n19129), .B(n19130), .Z(n19128) );
  XOR U18966 ( .A(n19127), .B(n19131), .Z(n19129) );
  XNOR U18967 ( .A(n19113), .B(n19110), .Z(n19120) );
  AND U18968 ( .A(n19132), .B(n19133), .Z(n19110) );
  XOR U18969 ( .A(n19134), .B(n19135), .Z(n19113) );
  AND U18970 ( .A(n19136), .B(n19137), .Z(n19135) );
  XOR U18971 ( .A(n19134), .B(n19138), .Z(n19136) );
  XNOR U18972 ( .A(n19062), .B(n19116), .Z(n19118) );
  XNOR U18973 ( .A(n19139), .B(n19140), .Z(n19062) );
  AND U18974 ( .A(n177), .B(n19068), .Z(n19140) );
  XOR U18975 ( .A(n19139), .B(n19066), .Z(n19068) );
  XOR U18976 ( .A(n19141), .B(n19142), .Z(n19116) );
  AND U18977 ( .A(n19143), .B(n19144), .Z(n19142) );
  XNOR U18978 ( .A(n19141), .B(n19132), .Z(n19144) );
  IV U18979 ( .A(n19074), .Z(n19132) );
  XNOR U18980 ( .A(n19145), .B(n19125), .Z(n19074) );
  XNOR U18981 ( .A(n19146), .B(n19131), .Z(n19125) );
  XOR U18982 ( .A(n19147), .B(n19148), .Z(n19131) );
  AND U18983 ( .A(n19149), .B(n19150), .Z(n19148) );
  XOR U18984 ( .A(n19147), .B(n19151), .Z(n19149) );
  XNOR U18985 ( .A(n19130), .B(n19122), .Z(n19146) );
  XOR U18986 ( .A(n19152), .B(n19153), .Z(n19122) );
  AND U18987 ( .A(n19154), .B(n19155), .Z(n19153) );
  XNOR U18988 ( .A(n19156), .B(n19152), .Z(n19154) );
  XNOR U18989 ( .A(n19157), .B(n19127), .Z(n19130) );
  XOR U18990 ( .A(n19158), .B(n19159), .Z(n19127) );
  AND U18991 ( .A(n19160), .B(n19161), .Z(n19159) );
  XOR U18992 ( .A(n19158), .B(n19162), .Z(n19160) );
  XNOR U18993 ( .A(n19163), .B(n19164), .Z(n19157) );
  AND U18994 ( .A(n19165), .B(n19166), .Z(n19164) );
  XNOR U18995 ( .A(n19163), .B(n19167), .Z(n19165) );
  XNOR U18996 ( .A(n19126), .B(n19133), .Z(n19145) );
  AND U18997 ( .A(n19086), .B(n19168), .Z(n19133) );
  XOR U18998 ( .A(n19138), .B(n19137), .Z(n19126) );
  XNOR U18999 ( .A(n19169), .B(n19134), .Z(n19137) );
  XOR U19000 ( .A(n19170), .B(n19171), .Z(n19134) );
  AND U19001 ( .A(n19172), .B(n19173), .Z(n19171) );
  XOR U19002 ( .A(n19170), .B(n19174), .Z(n19172) );
  XNOR U19003 ( .A(n19175), .B(n19176), .Z(n19169) );
  AND U19004 ( .A(n19177), .B(n19178), .Z(n19176) );
  XOR U19005 ( .A(n19175), .B(n19179), .Z(n19177) );
  XOR U19006 ( .A(n19180), .B(n19181), .Z(n19138) );
  AND U19007 ( .A(n19182), .B(n19183), .Z(n19181) );
  XOR U19008 ( .A(n19180), .B(n19184), .Z(n19182) );
  XNOR U19009 ( .A(n19071), .B(n19141), .Z(n19143) );
  XNOR U19010 ( .A(n19185), .B(n19186), .Z(n19071) );
  AND U19011 ( .A(n177), .B(n19078), .Z(n19186) );
  XOR U19012 ( .A(n19185), .B(n19076), .Z(n19078) );
  XOR U19013 ( .A(n19187), .B(n19188), .Z(n19141) );
  AND U19014 ( .A(n19189), .B(n19190), .Z(n19188) );
  XNOR U19015 ( .A(n19187), .B(n19086), .Z(n19190) );
  XOR U19016 ( .A(n19191), .B(n19155), .Z(n19086) );
  XNOR U19017 ( .A(n19192), .B(n19162), .Z(n19155) );
  XOR U19018 ( .A(n19151), .B(n19150), .Z(n19162) );
  XNOR U19019 ( .A(n19193), .B(n19147), .Z(n19150) );
  XOR U19020 ( .A(n19194), .B(n19195), .Z(n19147) );
  AND U19021 ( .A(n19196), .B(n19197), .Z(n19195) );
  XOR U19022 ( .A(n19194), .B(n19198), .Z(n19196) );
  XNOR U19023 ( .A(n19199), .B(n19200), .Z(n19193) );
  NOR U19024 ( .A(n19201), .B(n19202), .Z(n19200) );
  XNOR U19025 ( .A(n19199), .B(n19203), .Z(n19201) );
  XOR U19026 ( .A(n19204), .B(n19205), .Z(n19151) );
  NOR U19027 ( .A(n19206), .B(n19207), .Z(n19205) );
  XNOR U19028 ( .A(n19204), .B(n19208), .Z(n19206) );
  XNOR U19029 ( .A(n19161), .B(n19152), .Z(n19192) );
  XOR U19030 ( .A(n19209), .B(n19210), .Z(n19152) );
  NOR U19031 ( .A(n19211), .B(n19212), .Z(n19210) );
  XNOR U19032 ( .A(n19209), .B(n19213), .Z(n19211) );
  XOR U19033 ( .A(n19214), .B(n19167), .Z(n19161) );
  XNOR U19034 ( .A(n19215), .B(n19216), .Z(n19167) );
  NOR U19035 ( .A(n19217), .B(n19218), .Z(n19216) );
  XNOR U19036 ( .A(n19215), .B(n19219), .Z(n19217) );
  XNOR U19037 ( .A(n19166), .B(n19158), .Z(n19214) );
  XOR U19038 ( .A(n19220), .B(n19221), .Z(n19158) );
  AND U19039 ( .A(n19222), .B(n19223), .Z(n19221) );
  XOR U19040 ( .A(n19220), .B(n19224), .Z(n19222) );
  XNOR U19041 ( .A(n19225), .B(n19163), .Z(n19166) );
  XOR U19042 ( .A(n19226), .B(n19227), .Z(n19163) );
  AND U19043 ( .A(n19228), .B(n19229), .Z(n19227) );
  XOR U19044 ( .A(n19226), .B(n19230), .Z(n19228) );
  XNOR U19045 ( .A(n19231), .B(n19232), .Z(n19225) );
  NOR U19046 ( .A(n19233), .B(n19234), .Z(n19232) );
  XOR U19047 ( .A(n19231), .B(n19235), .Z(n19233) );
  XOR U19048 ( .A(n19156), .B(n19168), .Z(n19191) );
  NOR U19049 ( .A(n19094), .B(n19236), .Z(n19168) );
  XNOR U19050 ( .A(n19174), .B(n19173), .Z(n19156) );
  XNOR U19051 ( .A(n19237), .B(n19179), .Z(n19173) );
  XOR U19052 ( .A(n19238), .B(n19239), .Z(n19179) );
  NOR U19053 ( .A(n19240), .B(n19241), .Z(n19239) );
  XNOR U19054 ( .A(n19238), .B(n19242), .Z(n19240) );
  XNOR U19055 ( .A(n19178), .B(n19170), .Z(n19237) );
  XOR U19056 ( .A(n19243), .B(n19244), .Z(n19170) );
  AND U19057 ( .A(n19245), .B(n19246), .Z(n19244) );
  XNOR U19058 ( .A(n19243), .B(n19247), .Z(n19245) );
  XNOR U19059 ( .A(n19248), .B(n19175), .Z(n19178) );
  XOR U19060 ( .A(n19249), .B(n19250), .Z(n19175) );
  AND U19061 ( .A(n19251), .B(n19252), .Z(n19250) );
  XOR U19062 ( .A(n19249), .B(n19253), .Z(n19251) );
  XNOR U19063 ( .A(n19254), .B(n19255), .Z(n19248) );
  NOR U19064 ( .A(n19256), .B(n19257), .Z(n19255) );
  XOR U19065 ( .A(n19254), .B(n19258), .Z(n19256) );
  XOR U19066 ( .A(n19184), .B(n19183), .Z(n19174) );
  XNOR U19067 ( .A(n19259), .B(n19180), .Z(n19183) );
  XOR U19068 ( .A(n19260), .B(n19261), .Z(n19180) );
  AND U19069 ( .A(n19262), .B(n19263), .Z(n19261) );
  XOR U19070 ( .A(n19260), .B(n19264), .Z(n19262) );
  XNOR U19071 ( .A(n19265), .B(n19266), .Z(n19259) );
  NOR U19072 ( .A(n19267), .B(n19268), .Z(n19266) );
  XNOR U19073 ( .A(n19265), .B(n19269), .Z(n19267) );
  XOR U19074 ( .A(n19270), .B(n19271), .Z(n19184) );
  NOR U19075 ( .A(n19272), .B(n19273), .Z(n19271) );
  XNOR U19076 ( .A(n19270), .B(n19274), .Z(n19272) );
  XNOR U19077 ( .A(n19083), .B(n19187), .Z(n19189) );
  XNOR U19078 ( .A(n19275), .B(n19276), .Z(n19083) );
  AND U19079 ( .A(n177), .B(n19090), .Z(n19276) );
  XOR U19080 ( .A(n19275), .B(n19088), .Z(n19090) );
  AND U19081 ( .A(n19091), .B(n19094), .Z(n19187) );
  XOR U19082 ( .A(n19277), .B(n19236), .Z(n19094) );
  XNOR U19083 ( .A(p_input[2048]), .B(p_input[320]), .Z(n19236) );
  XOR U19084 ( .A(n19213), .B(n19212), .Z(n19277) );
  XOR U19085 ( .A(n19278), .B(n19224), .Z(n19212) );
  XOR U19086 ( .A(n19198), .B(n19197), .Z(n19224) );
  XNOR U19087 ( .A(n19279), .B(n19203), .Z(n19197) );
  XOR U19088 ( .A(p_input[2072]), .B(p_input[344]), .Z(n19203) );
  XOR U19089 ( .A(n19194), .B(n19202), .Z(n19279) );
  XOR U19090 ( .A(n19280), .B(n19199), .Z(n19202) );
  XOR U19091 ( .A(p_input[2070]), .B(p_input[342]), .Z(n19199) );
  XNOR U19092 ( .A(p_input[2071]), .B(p_input[343]), .Z(n19280) );
  XNOR U19093 ( .A(n16727), .B(p_input[338]), .Z(n19194) );
  XNOR U19094 ( .A(n19208), .B(n19207), .Z(n19198) );
  XOR U19095 ( .A(n19281), .B(n19204), .Z(n19207) );
  XOR U19096 ( .A(p_input[2067]), .B(p_input[339]), .Z(n19204) );
  XNOR U19097 ( .A(p_input[2068]), .B(p_input[340]), .Z(n19281) );
  XOR U19098 ( .A(p_input[2069]), .B(p_input[341]), .Z(n19208) );
  XNOR U19099 ( .A(n19223), .B(n19209), .Z(n19278) );
  XNOR U19100 ( .A(n16729), .B(p_input[321]), .Z(n19209) );
  XNOR U19101 ( .A(n19282), .B(n19230), .Z(n19223) );
  XNOR U19102 ( .A(n19219), .B(n19218), .Z(n19230) );
  XOR U19103 ( .A(n19283), .B(n19215), .Z(n19218) );
  XNOR U19104 ( .A(n16444), .B(p_input[346]), .Z(n19215) );
  XNOR U19105 ( .A(p_input[2075]), .B(p_input[347]), .Z(n19283) );
  XOR U19106 ( .A(p_input[2076]), .B(p_input[348]), .Z(n19219) );
  XNOR U19107 ( .A(n19229), .B(n19220), .Z(n19282) );
  XNOR U19108 ( .A(n16732), .B(p_input[337]), .Z(n19220) );
  XOR U19109 ( .A(n19284), .B(n19235), .Z(n19229) );
  XNOR U19110 ( .A(p_input[2079]), .B(p_input[351]), .Z(n19235) );
  XOR U19111 ( .A(n19226), .B(n19234), .Z(n19284) );
  XOR U19112 ( .A(n19285), .B(n19231), .Z(n19234) );
  XOR U19113 ( .A(p_input[2077]), .B(p_input[349]), .Z(n19231) );
  XNOR U19114 ( .A(p_input[2078]), .B(p_input[350]), .Z(n19285) );
  XNOR U19115 ( .A(n16448), .B(p_input[345]), .Z(n19226) );
  XNOR U19116 ( .A(n19247), .B(n19246), .Z(n19213) );
  XNOR U19117 ( .A(n19286), .B(n19253), .Z(n19246) );
  XNOR U19118 ( .A(n19242), .B(n19241), .Z(n19253) );
  XOR U19119 ( .A(n19287), .B(n19238), .Z(n19241) );
  XNOR U19120 ( .A(n16737), .B(p_input[331]), .Z(n19238) );
  XNOR U19121 ( .A(p_input[2060]), .B(p_input[332]), .Z(n19287) );
  XOR U19122 ( .A(p_input[2061]), .B(p_input[333]), .Z(n19242) );
  XNOR U19123 ( .A(n19252), .B(n19243), .Z(n19286) );
  XNOR U19124 ( .A(n16452), .B(p_input[322]), .Z(n19243) );
  XOR U19125 ( .A(n19288), .B(n19258), .Z(n19252) );
  XNOR U19126 ( .A(p_input[2064]), .B(p_input[336]), .Z(n19258) );
  XOR U19127 ( .A(n19249), .B(n19257), .Z(n19288) );
  XOR U19128 ( .A(n19289), .B(n19254), .Z(n19257) );
  XOR U19129 ( .A(p_input[2062]), .B(p_input[334]), .Z(n19254) );
  XNOR U19130 ( .A(p_input[2063]), .B(p_input[335]), .Z(n19289) );
  XNOR U19131 ( .A(n16740), .B(p_input[330]), .Z(n19249) );
  XNOR U19132 ( .A(n19264), .B(n19263), .Z(n19247) );
  XNOR U19133 ( .A(n19290), .B(n19269), .Z(n19263) );
  XOR U19134 ( .A(p_input[2057]), .B(p_input[329]), .Z(n19269) );
  XOR U19135 ( .A(n19260), .B(n19268), .Z(n19290) );
  XOR U19136 ( .A(n19291), .B(n19265), .Z(n19268) );
  XOR U19137 ( .A(p_input[2055]), .B(p_input[327]), .Z(n19265) );
  XNOR U19138 ( .A(p_input[2056]), .B(p_input[328]), .Z(n19291) );
  XNOR U19139 ( .A(n16459), .B(p_input[323]), .Z(n19260) );
  XNOR U19140 ( .A(n19274), .B(n19273), .Z(n19264) );
  XOR U19141 ( .A(n19292), .B(n19270), .Z(n19273) );
  XOR U19142 ( .A(p_input[2052]), .B(p_input[324]), .Z(n19270) );
  XNOR U19143 ( .A(p_input[2053]), .B(p_input[325]), .Z(n19292) );
  XOR U19144 ( .A(p_input[2054]), .B(p_input[326]), .Z(n19274) );
  XNOR U19145 ( .A(n19293), .B(n19294), .Z(n19091) );
  AND U19146 ( .A(n177), .B(n19295), .Z(n19294) );
  XNOR U19147 ( .A(n19296), .B(n19297), .Z(n177) );
  AND U19148 ( .A(n19298), .B(n19299), .Z(n19297) );
  XOR U19149 ( .A(n19296), .B(n19101), .Z(n19299) );
  XNOR U19150 ( .A(n19296), .B(n19043), .Z(n19298) );
  XOR U19151 ( .A(n19300), .B(n19301), .Z(n19296) );
  AND U19152 ( .A(n19302), .B(n19303), .Z(n19301) );
  XNOR U19153 ( .A(n19114), .B(n19300), .Z(n19303) );
  XOR U19154 ( .A(n19300), .B(n19055), .Z(n19302) );
  XOR U19155 ( .A(n19304), .B(n19305), .Z(n19300) );
  AND U19156 ( .A(n19306), .B(n19307), .Z(n19305) );
  XNOR U19157 ( .A(n19139), .B(n19304), .Z(n19307) );
  XOR U19158 ( .A(n19304), .B(n19066), .Z(n19306) );
  XOR U19159 ( .A(n19308), .B(n19309), .Z(n19304) );
  AND U19160 ( .A(n19310), .B(n19311), .Z(n19309) );
  XOR U19161 ( .A(n19308), .B(n19076), .Z(n19310) );
  XOR U19162 ( .A(n19312), .B(n19313), .Z(n19032) );
  AND U19163 ( .A(n181), .B(n19295), .Z(n19313) );
  XNOR U19164 ( .A(n19293), .B(n19312), .Z(n19295) );
  XNOR U19165 ( .A(n19314), .B(n19315), .Z(n181) );
  AND U19166 ( .A(n19316), .B(n19317), .Z(n19315) );
  XNOR U19167 ( .A(n19318), .B(n19314), .Z(n19317) );
  IV U19168 ( .A(n19101), .Z(n19318) );
  XNOR U19169 ( .A(n19319), .B(n19320), .Z(n19101) );
  AND U19170 ( .A(n184), .B(n19321), .Z(n19320) );
  XNOR U19171 ( .A(n19319), .B(n19322), .Z(n19321) );
  XNOR U19172 ( .A(n19043), .B(n19314), .Z(n19316) );
  XOR U19173 ( .A(n19323), .B(n19324), .Z(n19043) );
  AND U19174 ( .A(n192), .B(n19325), .Z(n19324) );
  XOR U19175 ( .A(n19326), .B(n19327), .Z(n19314) );
  AND U19176 ( .A(n19328), .B(n19329), .Z(n19327) );
  XNOR U19177 ( .A(n19326), .B(n19114), .Z(n19329) );
  XNOR U19178 ( .A(n19330), .B(n19331), .Z(n19114) );
  AND U19179 ( .A(n184), .B(n19332), .Z(n19331) );
  XOR U19180 ( .A(n19333), .B(n19330), .Z(n19332) );
  XNOR U19181 ( .A(n19334), .B(n19326), .Z(n19328) );
  IV U19182 ( .A(n19055), .Z(n19334) );
  XOR U19183 ( .A(n19335), .B(n19336), .Z(n19055) );
  AND U19184 ( .A(n192), .B(n19337), .Z(n19336) );
  XOR U19185 ( .A(n19338), .B(n19339), .Z(n19326) );
  AND U19186 ( .A(n19340), .B(n19341), .Z(n19339) );
  XNOR U19187 ( .A(n19338), .B(n19139), .Z(n19341) );
  XNOR U19188 ( .A(n19342), .B(n19343), .Z(n19139) );
  AND U19189 ( .A(n184), .B(n19344), .Z(n19343) );
  XNOR U19190 ( .A(n19345), .B(n19342), .Z(n19344) );
  XOR U19191 ( .A(n19066), .B(n19338), .Z(n19340) );
  XOR U19192 ( .A(n19346), .B(n19347), .Z(n19066) );
  AND U19193 ( .A(n192), .B(n19348), .Z(n19347) );
  XOR U19194 ( .A(n19308), .B(n19349), .Z(n19338) );
  AND U19195 ( .A(n19350), .B(n19311), .Z(n19349) );
  XNOR U19196 ( .A(n19185), .B(n19308), .Z(n19311) );
  XNOR U19197 ( .A(n19351), .B(n19352), .Z(n19185) );
  AND U19198 ( .A(n184), .B(n19353), .Z(n19352) );
  XOR U19199 ( .A(n19354), .B(n19351), .Z(n19353) );
  XNOR U19200 ( .A(n19355), .B(n19308), .Z(n19350) );
  IV U19201 ( .A(n19076), .Z(n19355) );
  XOR U19202 ( .A(n19356), .B(n19357), .Z(n19076) );
  AND U19203 ( .A(n192), .B(n19358), .Z(n19357) );
  XOR U19204 ( .A(n19359), .B(n19360), .Z(n19308) );
  AND U19205 ( .A(n19361), .B(n19362), .Z(n19360) );
  XNOR U19206 ( .A(n19359), .B(n19275), .Z(n19362) );
  XNOR U19207 ( .A(n19363), .B(n19364), .Z(n19275) );
  AND U19208 ( .A(n184), .B(n19365), .Z(n19364) );
  XNOR U19209 ( .A(n19366), .B(n19363), .Z(n19365) );
  XNOR U19210 ( .A(n19367), .B(n19359), .Z(n19361) );
  IV U19211 ( .A(n19088), .Z(n19367) );
  XOR U19212 ( .A(n19368), .B(n19369), .Z(n19088) );
  AND U19213 ( .A(n192), .B(n19370), .Z(n19369) );
  AND U19214 ( .A(n19312), .B(n19293), .Z(n19359) );
  XNOR U19215 ( .A(n19371), .B(n19372), .Z(n19293) );
  AND U19216 ( .A(n184), .B(n19373), .Z(n19372) );
  XNOR U19217 ( .A(n19374), .B(n19371), .Z(n19373) );
  XNOR U19218 ( .A(n19375), .B(n19376), .Z(n184) );
  AND U19219 ( .A(n19377), .B(n19378), .Z(n19376) );
  XOR U19220 ( .A(n19322), .B(n19375), .Z(n19378) );
  AND U19221 ( .A(n19379), .B(n19380), .Z(n19322) );
  XOR U19222 ( .A(n19375), .B(n19319), .Z(n19377) );
  XNOR U19223 ( .A(n19381), .B(n19382), .Z(n19319) );
  AND U19224 ( .A(n188), .B(n19325), .Z(n19382) );
  XOR U19225 ( .A(n19323), .B(n19381), .Z(n19325) );
  XOR U19226 ( .A(n19383), .B(n19384), .Z(n19375) );
  AND U19227 ( .A(n19385), .B(n19386), .Z(n19384) );
  XNOR U19228 ( .A(n19383), .B(n19379), .Z(n19386) );
  IV U19229 ( .A(n19333), .Z(n19379) );
  XOR U19230 ( .A(n19387), .B(n19388), .Z(n19333) );
  XOR U19231 ( .A(n19389), .B(n19380), .Z(n19388) );
  AND U19232 ( .A(n19345), .B(n19390), .Z(n19380) );
  AND U19233 ( .A(n19391), .B(n19392), .Z(n19389) );
  XOR U19234 ( .A(n19393), .B(n19387), .Z(n19391) );
  XNOR U19235 ( .A(n19330), .B(n19383), .Z(n19385) );
  XNOR U19236 ( .A(n19394), .B(n19395), .Z(n19330) );
  AND U19237 ( .A(n188), .B(n19337), .Z(n19395) );
  XOR U19238 ( .A(n19394), .B(n19335), .Z(n19337) );
  XOR U19239 ( .A(n19396), .B(n19397), .Z(n19383) );
  AND U19240 ( .A(n19398), .B(n19399), .Z(n19397) );
  XNOR U19241 ( .A(n19396), .B(n19345), .Z(n19399) );
  XOR U19242 ( .A(n19400), .B(n19392), .Z(n19345) );
  XNOR U19243 ( .A(n19401), .B(n19387), .Z(n19392) );
  XOR U19244 ( .A(n19402), .B(n19403), .Z(n19387) );
  AND U19245 ( .A(n19404), .B(n19405), .Z(n19403) );
  XOR U19246 ( .A(n19406), .B(n19402), .Z(n19404) );
  XNOR U19247 ( .A(n19407), .B(n19408), .Z(n19401) );
  AND U19248 ( .A(n19409), .B(n19410), .Z(n19408) );
  XOR U19249 ( .A(n19407), .B(n19411), .Z(n19409) );
  XNOR U19250 ( .A(n19393), .B(n19390), .Z(n19400) );
  AND U19251 ( .A(n19412), .B(n19413), .Z(n19390) );
  XOR U19252 ( .A(n19414), .B(n19415), .Z(n19393) );
  AND U19253 ( .A(n19416), .B(n19417), .Z(n19415) );
  XOR U19254 ( .A(n19414), .B(n19418), .Z(n19416) );
  XNOR U19255 ( .A(n19342), .B(n19396), .Z(n19398) );
  XNOR U19256 ( .A(n19419), .B(n19420), .Z(n19342) );
  AND U19257 ( .A(n188), .B(n19348), .Z(n19420) );
  XOR U19258 ( .A(n19419), .B(n19346), .Z(n19348) );
  XOR U19259 ( .A(n19421), .B(n19422), .Z(n19396) );
  AND U19260 ( .A(n19423), .B(n19424), .Z(n19422) );
  XNOR U19261 ( .A(n19421), .B(n19412), .Z(n19424) );
  IV U19262 ( .A(n19354), .Z(n19412) );
  XNOR U19263 ( .A(n19425), .B(n19405), .Z(n19354) );
  XNOR U19264 ( .A(n19426), .B(n19411), .Z(n19405) );
  XOR U19265 ( .A(n19427), .B(n19428), .Z(n19411) );
  AND U19266 ( .A(n19429), .B(n19430), .Z(n19428) );
  XOR U19267 ( .A(n19427), .B(n19431), .Z(n19429) );
  XNOR U19268 ( .A(n19410), .B(n19402), .Z(n19426) );
  XOR U19269 ( .A(n19432), .B(n19433), .Z(n19402) );
  AND U19270 ( .A(n19434), .B(n19435), .Z(n19433) );
  XNOR U19271 ( .A(n19436), .B(n19432), .Z(n19434) );
  XNOR U19272 ( .A(n19437), .B(n19407), .Z(n19410) );
  XOR U19273 ( .A(n19438), .B(n19439), .Z(n19407) );
  AND U19274 ( .A(n19440), .B(n19441), .Z(n19439) );
  XOR U19275 ( .A(n19438), .B(n19442), .Z(n19440) );
  XNOR U19276 ( .A(n19443), .B(n19444), .Z(n19437) );
  AND U19277 ( .A(n19445), .B(n19446), .Z(n19444) );
  XNOR U19278 ( .A(n19443), .B(n19447), .Z(n19445) );
  XNOR U19279 ( .A(n19406), .B(n19413), .Z(n19425) );
  AND U19280 ( .A(n19366), .B(n19448), .Z(n19413) );
  XOR U19281 ( .A(n19418), .B(n19417), .Z(n19406) );
  XNOR U19282 ( .A(n19449), .B(n19414), .Z(n19417) );
  XOR U19283 ( .A(n19450), .B(n19451), .Z(n19414) );
  AND U19284 ( .A(n19452), .B(n19453), .Z(n19451) );
  XOR U19285 ( .A(n19450), .B(n19454), .Z(n19452) );
  XNOR U19286 ( .A(n19455), .B(n19456), .Z(n19449) );
  AND U19287 ( .A(n19457), .B(n19458), .Z(n19456) );
  XOR U19288 ( .A(n19455), .B(n19459), .Z(n19457) );
  XOR U19289 ( .A(n19460), .B(n19461), .Z(n19418) );
  AND U19290 ( .A(n19462), .B(n19463), .Z(n19461) );
  XOR U19291 ( .A(n19460), .B(n19464), .Z(n19462) );
  XNOR U19292 ( .A(n19351), .B(n19421), .Z(n19423) );
  XNOR U19293 ( .A(n19465), .B(n19466), .Z(n19351) );
  AND U19294 ( .A(n188), .B(n19358), .Z(n19466) );
  XOR U19295 ( .A(n19465), .B(n19356), .Z(n19358) );
  XOR U19296 ( .A(n19467), .B(n19468), .Z(n19421) );
  AND U19297 ( .A(n19469), .B(n19470), .Z(n19468) );
  XNOR U19298 ( .A(n19467), .B(n19366), .Z(n19470) );
  XOR U19299 ( .A(n19471), .B(n19435), .Z(n19366) );
  XNOR U19300 ( .A(n19472), .B(n19442), .Z(n19435) );
  XOR U19301 ( .A(n19431), .B(n19430), .Z(n19442) );
  XNOR U19302 ( .A(n19473), .B(n19427), .Z(n19430) );
  XOR U19303 ( .A(n19474), .B(n19475), .Z(n19427) );
  AND U19304 ( .A(n19476), .B(n19477), .Z(n19475) );
  XOR U19305 ( .A(n19474), .B(n19478), .Z(n19476) );
  XNOR U19306 ( .A(n19479), .B(n19480), .Z(n19473) );
  NOR U19307 ( .A(n19481), .B(n19482), .Z(n19480) );
  XNOR U19308 ( .A(n19479), .B(n19483), .Z(n19481) );
  XOR U19309 ( .A(n19484), .B(n19485), .Z(n19431) );
  NOR U19310 ( .A(n19486), .B(n19487), .Z(n19485) );
  XNOR U19311 ( .A(n19484), .B(n19488), .Z(n19486) );
  XNOR U19312 ( .A(n19441), .B(n19432), .Z(n19472) );
  XOR U19313 ( .A(n19489), .B(n19490), .Z(n19432) );
  NOR U19314 ( .A(n19491), .B(n19492), .Z(n19490) );
  XNOR U19315 ( .A(n19489), .B(n19493), .Z(n19491) );
  XOR U19316 ( .A(n19494), .B(n19447), .Z(n19441) );
  XNOR U19317 ( .A(n19495), .B(n19496), .Z(n19447) );
  NOR U19318 ( .A(n19497), .B(n19498), .Z(n19496) );
  XNOR U19319 ( .A(n19495), .B(n19499), .Z(n19497) );
  XNOR U19320 ( .A(n19446), .B(n19438), .Z(n19494) );
  XOR U19321 ( .A(n19500), .B(n19501), .Z(n19438) );
  AND U19322 ( .A(n19502), .B(n19503), .Z(n19501) );
  XOR U19323 ( .A(n19500), .B(n19504), .Z(n19502) );
  XNOR U19324 ( .A(n19505), .B(n19443), .Z(n19446) );
  XOR U19325 ( .A(n19506), .B(n19507), .Z(n19443) );
  AND U19326 ( .A(n19508), .B(n19509), .Z(n19507) );
  XOR U19327 ( .A(n19506), .B(n19510), .Z(n19508) );
  XNOR U19328 ( .A(n19511), .B(n19512), .Z(n19505) );
  NOR U19329 ( .A(n19513), .B(n19514), .Z(n19512) );
  XOR U19330 ( .A(n19511), .B(n19515), .Z(n19513) );
  XOR U19331 ( .A(n19436), .B(n19448), .Z(n19471) );
  NOR U19332 ( .A(n19374), .B(n19516), .Z(n19448) );
  XNOR U19333 ( .A(n19454), .B(n19453), .Z(n19436) );
  XNOR U19334 ( .A(n19517), .B(n19459), .Z(n19453) );
  XOR U19335 ( .A(n19518), .B(n19519), .Z(n19459) );
  NOR U19336 ( .A(n19520), .B(n19521), .Z(n19519) );
  XNOR U19337 ( .A(n19518), .B(n19522), .Z(n19520) );
  XNOR U19338 ( .A(n19458), .B(n19450), .Z(n19517) );
  XOR U19339 ( .A(n19523), .B(n19524), .Z(n19450) );
  AND U19340 ( .A(n19525), .B(n19526), .Z(n19524) );
  XNOR U19341 ( .A(n19523), .B(n19527), .Z(n19525) );
  XNOR U19342 ( .A(n19528), .B(n19455), .Z(n19458) );
  XOR U19343 ( .A(n19529), .B(n19530), .Z(n19455) );
  AND U19344 ( .A(n19531), .B(n19532), .Z(n19530) );
  XOR U19345 ( .A(n19529), .B(n19533), .Z(n19531) );
  XNOR U19346 ( .A(n19534), .B(n19535), .Z(n19528) );
  NOR U19347 ( .A(n19536), .B(n19537), .Z(n19535) );
  XOR U19348 ( .A(n19534), .B(n19538), .Z(n19536) );
  XOR U19349 ( .A(n19464), .B(n19463), .Z(n19454) );
  XNOR U19350 ( .A(n19539), .B(n19460), .Z(n19463) );
  XOR U19351 ( .A(n19540), .B(n19541), .Z(n19460) );
  AND U19352 ( .A(n19542), .B(n19543), .Z(n19541) );
  XOR U19353 ( .A(n19540), .B(n19544), .Z(n19542) );
  XNOR U19354 ( .A(n19545), .B(n19546), .Z(n19539) );
  NOR U19355 ( .A(n19547), .B(n19548), .Z(n19546) );
  XNOR U19356 ( .A(n19545), .B(n19549), .Z(n19547) );
  XOR U19357 ( .A(n19550), .B(n19551), .Z(n19464) );
  NOR U19358 ( .A(n19552), .B(n19553), .Z(n19551) );
  XNOR U19359 ( .A(n19550), .B(n19554), .Z(n19552) );
  XNOR U19360 ( .A(n19363), .B(n19467), .Z(n19469) );
  XNOR U19361 ( .A(n19555), .B(n19556), .Z(n19363) );
  AND U19362 ( .A(n188), .B(n19370), .Z(n19556) );
  XOR U19363 ( .A(n19555), .B(n19368), .Z(n19370) );
  AND U19364 ( .A(n19371), .B(n19374), .Z(n19467) );
  XOR U19365 ( .A(n19557), .B(n19516), .Z(n19374) );
  XNOR U19366 ( .A(p_input[2048]), .B(p_input[352]), .Z(n19516) );
  XOR U19367 ( .A(n19493), .B(n19492), .Z(n19557) );
  XOR U19368 ( .A(n19558), .B(n19504), .Z(n19492) );
  XOR U19369 ( .A(n19478), .B(n19477), .Z(n19504) );
  XNOR U19370 ( .A(n19559), .B(n19483), .Z(n19477) );
  XOR U19371 ( .A(p_input[2072]), .B(p_input[376]), .Z(n19483) );
  XOR U19372 ( .A(n19474), .B(n19482), .Z(n19559) );
  XOR U19373 ( .A(n19560), .B(n19479), .Z(n19482) );
  XOR U19374 ( .A(p_input[2070]), .B(p_input[374]), .Z(n19479) );
  XNOR U19375 ( .A(p_input[2071]), .B(p_input[375]), .Z(n19560) );
  XNOR U19376 ( .A(n16727), .B(p_input[370]), .Z(n19474) );
  XNOR U19377 ( .A(n19488), .B(n19487), .Z(n19478) );
  XOR U19378 ( .A(n19561), .B(n19484), .Z(n19487) );
  XOR U19379 ( .A(p_input[2067]), .B(p_input[371]), .Z(n19484) );
  XNOR U19380 ( .A(p_input[2068]), .B(p_input[372]), .Z(n19561) );
  XOR U19381 ( .A(p_input[2069]), .B(p_input[373]), .Z(n19488) );
  XNOR U19382 ( .A(n19503), .B(n19489), .Z(n19558) );
  XNOR U19383 ( .A(n16729), .B(p_input[353]), .Z(n19489) );
  XNOR U19384 ( .A(n19562), .B(n19510), .Z(n19503) );
  XNOR U19385 ( .A(n19499), .B(n19498), .Z(n19510) );
  XOR U19386 ( .A(n19563), .B(n19495), .Z(n19498) );
  XNOR U19387 ( .A(n16444), .B(p_input[378]), .Z(n19495) );
  XNOR U19388 ( .A(p_input[2075]), .B(p_input[379]), .Z(n19563) );
  XOR U19389 ( .A(p_input[2076]), .B(p_input[380]), .Z(n19499) );
  XNOR U19390 ( .A(n19509), .B(n19500), .Z(n19562) );
  XNOR U19391 ( .A(n16732), .B(p_input[369]), .Z(n19500) );
  XOR U19392 ( .A(n19564), .B(n19515), .Z(n19509) );
  XNOR U19393 ( .A(p_input[2079]), .B(p_input[383]), .Z(n19515) );
  XOR U19394 ( .A(n19506), .B(n19514), .Z(n19564) );
  XOR U19395 ( .A(n19565), .B(n19511), .Z(n19514) );
  XOR U19396 ( .A(p_input[2077]), .B(p_input[381]), .Z(n19511) );
  XNOR U19397 ( .A(p_input[2078]), .B(p_input[382]), .Z(n19565) );
  XNOR U19398 ( .A(n16448), .B(p_input[377]), .Z(n19506) );
  XNOR U19399 ( .A(n19527), .B(n19526), .Z(n19493) );
  XNOR U19400 ( .A(n19566), .B(n19533), .Z(n19526) );
  XNOR U19401 ( .A(n19522), .B(n19521), .Z(n19533) );
  XOR U19402 ( .A(n19567), .B(n19518), .Z(n19521) );
  XNOR U19403 ( .A(n16737), .B(p_input[363]), .Z(n19518) );
  XNOR U19404 ( .A(p_input[2060]), .B(p_input[364]), .Z(n19567) );
  XOR U19405 ( .A(p_input[2061]), .B(p_input[365]), .Z(n19522) );
  XNOR U19406 ( .A(n19532), .B(n19523), .Z(n19566) );
  XNOR U19407 ( .A(n16452), .B(p_input[354]), .Z(n19523) );
  XOR U19408 ( .A(n19568), .B(n19538), .Z(n19532) );
  XNOR U19409 ( .A(p_input[2064]), .B(p_input[368]), .Z(n19538) );
  XOR U19410 ( .A(n19529), .B(n19537), .Z(n19568) );
  XOR U19411 ( .A(n19569), .B(n19534), .Z(n19537) );
  XOR U19412 ( .A(p_input[2062]), .B(p_input[366]), .Z(n19534) );
  XNOR U19413 ( .A(p_input[2063]), .B(p_input[367]), .Z(n19569) );
  XNOR U19414 ( .A(n16740), .B(p_input[362]), .Z(n19529) );
  XNOR U19415 ( .A(n19544), .B(n19543), .Z(n19527) );
  XNOR U19416 ( .A(n19570), .B(n19549), .Z(n19543) );
  XOR U19417 ( .A(p_input[2057]), .B(p_input[361]), .Z(n19549) );
  XOR U19418 ( .A(n19540), .B(n19548), .Z(n19570) );
  XOR U19419 ( .A(n19571), .B(n19545), .Z(n19548) );
  XOR U19420 ( .A(p_input[2055]), .B(p_input[359]), .Z(n19545) );
  XNOR U19421 ( .A(p_input[2056]), .B(p_input[360]), .Z(n19571) );
  XNOR U19422 ( .A(n16459), .B(p_input[355]), .Z(n19540) );
  XNOR U19423 ( .A(n19554), .B(n19553), .Z(n19544) );
  XOR U19424 ( .A(n19572), .B(n19550), .Z(n19553) );
  XOR U19425 ( .A(p_input[2052]), .B(p_input[356]), .Z(n19550) );
  XNOR U19426 ( .A(p_input[2053]), .B(p_input[357]), .Z(n19572) );
  XOR U19427 ( .A(p_input[2054]), .B(p_input[358]), .Z(n19554) );
  XNOR U19428 ( .A(n19573), .B(n19574), .Z(n19371) );
  AND U19429 ( .A(n188), .B(n19575), .Z(n19574) );
  XNOR U19430 ( .A(n19576), .B(n19577), .Z(n188) );
  AND U19431 ( .A(n19578), .B(n19579), .Z(n19577) );
  XOR U19432 ( .A(n19576), .B(n19381), .Z(n19579) );
  XNOR U19433 ( .A(n19576), .B(n19323), .Z(n19578) );
  XOR U19434 ( .A(n19580), .B(n19581), .Z(n19576) );
  AND U19435 ( .A(n19582), .B(n19583), .Z(n19581) );
  XNOR U19436 ( .A(n19394), .B(n19580), .Z(n19583) );
  XOR U19437 ( .A(n19580), .B(n19335), .Z(n19582) );
  XOR U19438 ( .A(n19584), .B(n19585), .Z(n19580) );
  AND U19439 ( .A(n19586), .B(n19587), .Z(n19585) );
  XNOR U19440 ( .A(n19419), .B(n19584), .Z(n19587) );
  XOR U19441 ( .A(n19584), .B(n19346), .Z(n19586) );
  XOR U19442 ( .A(n19588), .B(n19589), .Z(n19584) );
  AND U19443 ( .A(n19590), .B(n19591), .Z(n19589) );
  XOR U19444 ( .A(n19588), .B(n19356), .Z(n19590) );
  XOR U19445 ( .A(n19592), .B(n19593), .Z(n19312) );
  AND U19446 ( .A(n192), .B(n19575), .Z(n19593) );
  XNOR U19447 ( .A(n19573), .B(n19592), .Z(n19575) );
  XNOR U19448 ( .A(n19594), .B(n19595), .Z(n192) );
  AND U19449 ( .A(n19596), .B(n19597), .Z(n19595) );
  XNOR U19450 ( .A(n19598), .B(n19594), .Z(n19597) );
  IV U19451 ( .A(n19381), .Z(n19598) );
  XNOR U19452 ( .A(n19599), .B(n19600), .Z(n19381) );
  AND U19453 ( .A(n195), .B(n19601), .Z(n19600) );
  XNOR U19454 ( .A(n19599), .B(n19602), .Z(n19601) );
  XNOR U19455 ( .A(n19323), .B(n19594), .Z(n19596) );
  XOR U19456 ( .A(n19603), .B(n19604), .Z(n19323) );
  AND U19457 ( .A(n203), .B(n19605), .Z(n19604) );
  XOR U19458 ( .A(n19606), .B(n19607), .Z(n19594) );
  AND U19459 ( .A(n19608), .B(n19609), .Z(n19607) );
  XNOR U19460 ( .A(n19606), .B(n19394), .Z(n19609) );
  XNOR U19461 ( .A(n19610), .B(n19611), .Z(n19394) );
  AND U19462 ( .A(n195), .B(n19612), .Z(n19611) );
  XOR U19463 ( .A(n19613), .B(n19610), .Z(n19612) );
  XNOR U19464 ( .A(n19614), .B(n19606), .Z(n19608) );
  IV U19465 ( .A(n19335), .Z(n19614) );
  XOR U19466 ( .A(n19615), .B(n19616), .Z(n19335) );
  AND U19467 ( .A(n203), .B(n19617), .Z(n19616) );
  XOR U19468 ( .A(n19618), .B(n19619), .Z(n19606) );
  AND U19469 ( .A(n19620), .B(n19621), .Z(n19619) );
  XNOR U19470 ( .A(n19618), .B(n19419), .Z(n19621) );
  XNOR U19471 ( .A(n19622), .B(n19623), .Z(n19419) );
  AND U19472 ( .A(n195), .B(n19624), .Z(n19623) );
  XNOR U19473 ( .A(n19625), .B(n19622), .Z(n19624) );
  XOR U19474 ( .A(n19346), .B(n19618), .Z(n19620) );
  XOR U19475 ( .A(n19626), .B(n19627), .Z(n19346) );
  AND U19476 ( .A(n203), .B(n19628), .Z(n19627) );
  XOR U19477 ( .A(n19588), .B(n19629), .Z(n19618) );
  AND U19478 ( .A(n19630), .B(n19591), .Z(n19629) );
  XNOR U19479 ( .A(n19465), .B(n19588), .Z(n19591) );
  XNOR U19480 ( .A(n19631), .B(n19632), .Z(n19465) );
  AND U19481 ( .A(n195), .B(n19633), .Z(n19632) );
  XOR U19482 ( .A(n19634), .B(n19631), .Z(n19633) );
  XNOR U19483 ( .A(n19635), .B(n19588), .Z(n19630) );
  IV U19484 ( .A(n19356), .Z(n19635) );
  XOR U19485 ( .A(n19636), .B(n19637), .Z(n19356) );
  AND U19486 ( .A(n203), .B(n19638), .Z(n19637) );
  XOR U19487 ( .A(n19639), .B(n19640), .Z(n19588) );
  AND U19488 ( .A(n19641), .B(n19642), .Z(n19640) );
  XNOR U19489 ( .A(n19639), .B(n19555), .Z(n19642) );
  XNOR U19490 ( .A(n19643), .B(n19644), .Z(n19555) );
  AND U19491 ( .A(n195), .B(n19645), .Z(n19644) );
  XNOR U19492 ( .A(n19646), .B(n19643), .Z(n19645) );
  XNOR U19493 ( .A(n19647), .B(n19639), .Z(n19641) );
  IV U19494 ( .A(n19368), .Z(n19647) );
  XOR U19495 ( .A(n19648), .B(n19649), .Z(n19368) );
  AND U19496 ( .A(n203), .B(n19650), .Z(n19649) );
  AND U19497 ( .A(n19592), .B(n19573), .Z(n19639) );
  XNOR U19498 ( .A(n19651), .B(n19652), .Z(n19573) );
  AND U19499 ( .A(n195), .B(n19653), .Z(n19652) );
  XNOR U19500 ( .A(n19654), .B(n19651), .Z(n19653) );
  XNOR U19501 ( .A(n19655), .B(n19656), .Z(n195) );
  AND U19502 ( .A(n19657), .B(n19658), .Z(n19656) );
  XOR U19503 ( .A(n19602), .B(n19655), .Z(n19658) );
  AND U19504 ( .A(n19659), .B(n19660), .Z(n19602) );
  XOR U19505 ( .A(n19655), .B(n19599), .Z(n19657) );
  XNOR U19506 ( .A(n19661), .B(n19662), .Z(n19599) );
  AND U19507 ( .A(n199), .B(n19605), .Z(n19662) );
  XOR U19508 ( .A(n19603), .B(n19661), .Z(n19605) );
  XOR U19509 ( .A(n19663), .B(n19664), .Z(n19655) );
  AND U19510 ( .A(n19665), .B(n19666), .Z(n19664) );
  XNOR U19511 ( .A(n19663), .B(n19659), .Z(n19666) );
  IV U19512 ( .A(n19613), .Z(n19659) );
  XOR U19513 ( .A(n19667), .B(n19668), .Z(n19613) );
  XOR U19514 ( .A(n19669), .B(n19660), .Z(n19668) );
  AND U19515 ( .A(n19625), .B(n19670), .Z(n19660) );
  AND U19516 ( .A(n19671), .B(n19672), .Z(n19669) );
  XOR U19517 ( .A(n19673), .B(n19667), .Z(n19671) );
  XNOR U19518 ( .A(n19610), .B(n19663), .Z(n19665) );
  XNOR U19519 ( .A(n19674), .B(n19675), .Z(n19610) );
  AND U19520 ( .A(n199), .B(n19617), .Z(n19675) );
  XOR U19521 ( .A(n19674), .B(n19615), .Z(n19617) );
  XOR U19522 ( .A(n19676), .B(n19677), .Z(n19663) );
  AND U19523 ( .A(n19678), .B(n19679), .Z(n19677) );
  XNOR U19524 ( .A(n19676), .B(n19625), .Z(n19679) );
  XOR U19525 ( .A(n19680), .B(n19672), .Z(n19625) );
  XNOR U19526 ( .A(n19681), .B(n19667), .Z(n19672) );
  XOR U19527 ( .A(n19682), .B(n19683), .Z(n19667) );
  AND U19528 ( .A(n19684), .B(n19685), .Z(n19683) );
  XOR U19529 ( .A(n19686), .B(n19682), .Z(n19684) );
  XNOR U19530 ( .A(n19687), .B(n19688), .Z(n19681) );
  AND U19531 ( .A(n19689), .B(n19690), .Z(n19688) );
  XOR U19532 ( .A(n19687), .B(n19691), .Z(n19689) );
  XNOR U19533 ( .A(n19673), .B(n19670), .Z(n19680) );
  AND U19534 ( .A(n19692), .B(n19693), .Z(n19670) );
  XOR U19535 ( .A(n19694), .B(n19695), .Z(n19673) );
  AND U19536 ( .A(n19696), .B(n19697), .Z(n19695) );
  XOR U19537 ( .A(n19694), .B(n19698), .Z(n19696) );
  XNOR U19538 ( .A(n19622), .B(n19676), .Z(n19678) );
  XNOR U19539 ( .A(n19699), .B(n19700), .Z(n19622) );
  AND U19540 ( .A(n199), .B(n19628), .Z(n19700) );
  XOR U19541 ( .A(n19699), .B(n19626), .Z(n19628) );
  XOR U19542 ( .A(n19701), .B(n19702), .Z(n19676) );
  AND U19543 ( .A(n19703), .B(n19704), .Z(n19702) );
  XNOR U19544 ( .A(n19701), .B(n19692), .Z(n19704) );
  IV U19545 ( .A(n19634), .Z(n19692) );
  XNOR U19546 ( .A(n19705), .B(n19685), .Z(n19634) );
  XNOR U19547 ( .A(n19706), .B(n19691), .Z(n19685) );
  XOR U19548 ( .A(n19707), .B(n19708), .Z(n19691) );
  AND U19549 ( .A(n19709), .B(n19710), .Z(n19708) );
  XOR U19550 ( .A(n19707), .B(n19711), .Z(n19709) );
  XNOR U19551 ( .A(n19690), .B(n19682), .Z(n19706) );
  XOR U19552 ( .A(n19712), .B(n19713), .Z(n19682) );
  AND U19553 ( .A(n19714), .B(n19715), .Z(n19713) );
  XNOR U19554 ( .A(n19716), .B(n19712), .Z(n19714) );
  XNOR U19555 ( .A(n19717), .B(n19687), .Z(n19690) );
  XOR U19556 ( .A(n19718), .B(n19719), .Z(n19687) );
  AND U19557 ( .A(n19720), .B(n19721), .Z(n19719) );
  XOR U19558 ( .A(n19718), .B(n19722), .Z(n19720) );
  XNOR U19559 ( .A(n19723), .B(n19724), .Z(n19717) );
  AND U19560 ( .A(n19725), .B(n19726), .Z(n19724) );
  XNOR U19561 ( .A(n19723), .B(n19727), .Z(n19725) );
  XNOR U19562 ( .A(n19686), .B(n19693), .Z(n19705) );
  AND U19563 ( .A(n19646), .B(n19728), .Z(n19693) );
  XOR U19564 ( .A(n19698), .B(n19697), .Z(n19686) );
  XNOR U19565 ( .A(n19729), .B(n19694), .Z(n19697) );
  XOR U19566 ( .A(n19730), .B(n19731), .Z(n19694) );
  AND U19567 ( .A(n19732), .B(n19733), .Z(n19731) );
  XOR U19568 ( .A(n19730), .B(n19734), .Z(n19732) );
  XNOR U19569 ( .A(n19735), .B(n19736), .Z(n19729) );
  AND U19570 ( .A(n19737), .B(n19738), .Z(n19736) );
  XOR U19571 ( .A(n19735), .B(n19739), .Z(n19737) );
  XOR U19572 ( .A(n19740), .B(n19741), .Z(n19698) );
  AND U19573 ( .A(n19742), .B(n19743), .Z(n19741) );
  XOR U19574 ( .A(n19740), .B(n19744), .Z(n19742) );
  XNOR U19575 ( .A(n19631), .B(n19701), .Z(n19703) );
  XNOR U19576 ( .A(n19745), .B(n19746), .Z(n19631) );
  AND U19577 ( .A(n199), .B(n19638), .Z(n19746) );
  XOR U19578 ( .A(n19745), .B(n19636), .Z(n19638) );
  XOR U19579 ( .A(n19747), .B(n19748), .Z(n19701) );
  AND U19580 ( .A(n19749), .B(n19750), .Z(n19748) );
  XNOR U19581 ( .A(n19747), .B(n19646), .Z(n19750) );
  XOR U19582 ( .A(n19751), .B(n19715), .Z(n19646) );
  XNOR U19583 ( .A(n19752), .B(n19722), .Z(n19715) );
  XOR U19584 ( .A(n19711), .B(n19710), .Z(n19722) );
  XNOR U19585 ( .A(n19753), .B(n19707), .Z(n19710) );
  XOR U19586 ( .A(n19754), .B(n19755), .Z(n19707) );
  AND U19587 ( .A(n19756), .B(n19757), .Z(n19755) );
  XOR U19588 ( .A(n19754), .B(n19758), .Z(n19756) );
  XNOR U19589 ( .A(n19759), .B(n19760), .Z(n19753) );
  NOR U19590 ( .A(n19761), .B(n19762), .Z(n19760) );
  XNOR U19591 ( .A(n19759), .B(n19763), .Z(n19761) );
  XOR U19592 ( .A(n19764), .B(n19765), .Z(n19711) );
  NOR U19593 ( .A(n19766), .B(n19767), .Z(n19765) );
  XNOR U19594 ( .A(n19764), .B(n19768), .Z(n19766) );
  XNOR U19595 ( .A(n19721), .B(n19712), .Z(n19752) );
  XOR U19596 ( .A(n19769), .B(n19770), .Z(n19712) );
  NOR U19597 ( .A(n19771), .B(n19772), .Z(n19770) );
  XNOR U19598 ( .A(n19769), .B(n19773), .Z(n19771) );
  XOR U19599 ( .A(n19774), .B(n19727), .Z(n19721) );
  XNOR U19600 ( .A(n19775), .B(n19776), .Z(n19727) );
  NOR U19601 ( .A(n19777), .B(n19778), .Z(n19776) );
  XNOR U19602 ( .A(n19775), .B(n19779), .Z(n19777) );
  XNOR U19603 ( .A(n19726), .B(n19718), .Z(n19774) );
  XOR U19604 ( .A(n19780), .B(n19781), .Z(n19718) );
  AND U19605 ( .A(n19782), .B(n19783), .Z(n19781) );
  XOR U19606 ( .A(n19780), .B(n19784), .Z(n19782) );
  XNOR U19607 ( .A(n19785), .B(n19723), .Z(n19726) );
  XOR U19608 ( .A(n19786), .B(n19787), .Z(n19723) );
  AND U19609 ( .A(n19788), .B(n19789), .Z(n19787) );
  XOR U19610 ( .A(n19786), .B(n19790), .Z(n19788) );
  XNOR U19611 ( .A(n19791), .B(n19792), .Z(n19785) );
  NOR U19612 ( .A(n19793), .B(n19794), .Z(n19792) );
  XOR U19613 ( .A(n19791), .B(n19795), .Z(n19793) );
  XOR U19614 ( .A(n19716), .B(n19728), .Z(n19751) );
  NOR U19615 ( .A(n19654), .B(n19796), .Z(n19728) );
  XNOR U19616 ( .A(n19734), .B(n19733), .Z(n19716) );
  XNOR U19617 ( .A(n19797), .B(n19739), .Z(n19733) );
  XOR U19618 ( .A(n19798), .B(n19799), .Z(n19739) );
  NOR U19619 ( .A(n19800), .B(n19801), .Z(n19799) );
  XNOR U19620 ( .A(n19798), .B(n19802), .Z(n19800) );
  XNOR U19621 ( .A(n19738), .B(n19730), .Z(n19797) );
  XOR U19622 ( .A(n19803), .B(n19804), .Z(n19730) );
  AND U19623 ( .A(n19805), .B(n19806), .Z(n19804) );
  XNOR U19624 ( .A(n19803), .B(n19807), .Z(n19805) );
  XNOR U19625 ( .A(n19808), .B(n19735), .Z(n19738) );
  XOR U19626 ( .A(n19809), .B(n19810), .Z(n19735) );
  AND U19627 ( .A(n19811), .B(n19812), .Z(n19810) );
  XOR U19628 ( .A(n19809), .B(n19813), .Z(n19811) );
  XNOR U19629 ( .A(n19814), .B(n19815), .Z(n19808) );
  NOR U19630 ( .A(n19816), .B(n19817), .Z(n19815) );
  XOR U19631 ( .A(n19814), .B(n19818), .Z(n19816) );
  XOR U19632 ( .A(n19744), .B(n19743), .Z(n19734) );
  XNOR U19633 ( .A(n19819), .B(n19740), .Z(n19743) );
  XOR U19634 ( .A(n19820), .B(n19821), .Z(n19740) );
  AND U19635 ( .A(n19822), .B(n19823), .Z(n19821) );
  XOR U19636 ( .A(n19820), .B(n19824), .Z(n19822) );
  XNOR U19637 ( .A(n19825), .B(n19826), .Z(n19819) );
  NOR U19638 ( .A(n19827), .B(n19828), .Z(n19826) );
  XNOR U19639 ( .A(n19825), .B(n19829), .Z(n19827) );
  XOR U19640 ( .A(n19830), .B(n19831), .Z(n19744) );
  NOR U19641 ( .A(n19832), .B(n19833), .Z(n19831) );
  XNOR U19642 ( .A(n19830), .B(n19834), .Z(n19832) );
  XNOR U19643 ( .A(n19643), .B(n19747), .Z(n19749) );
  XNOR U19644 ( .A(n19835), .B(n19836), .Z(n19643) );
  AND U19645 ( .A(n199), .B(n19650), .Z(n19836) );
  XOR U19646 ( .A(n19835), .B(n19648), .Z(n19650) );
  AND U19647 ( .A(n19651), .B(n19654), .Z(n19747) );
  XOR U19648 ( .A(n19837), .B(n19796), .Z(n19654) );
  XNOR U19649 ( .A(p_input[2048]), .B(p_input[384]), .Z(n19796) );
  XOR U19650 ( .A(n19773), .B(n19772), .Z(n19837) );
  XOR U19651 ( .A(n19838), .B(n19784), .Z(n19772) );
  XOR U19652 ( .A(n19758), .B(n19757), .Z(n19784) );
  XNOR U19653 ( .A(n19839), .B(n19763), .Z(n19757) );
  XOR U19654 ( .A(p_input[2072]), .B(p_input[408]), .Z(n19763) );
  XOR U19655 ( .A(n19754), .B(n19762), .Z(n19839) );
  XOR U19656 ( .A(n19840), .B(n19759), .Z(n19762) );
  XOR U19657 ( .A(p_input[2070]), .B(p_input[406]), .Z(n19759) );
  XNOR U19658 ( .A(p_input[2071]), .B(p_input[407]), .Z(n19840) );
  XNOR U19659 ( .A(n16727), .B(p_input[402]), .Z(n19754) );
  XNOR U19660 ( .A(n19768), .B(n19767), .Z(n19758) );
  XOR U19661 ( .A(n19841), .B(n19764), .Z(n19767) );
  XOR U19662 ( .A(p_input[2067]), .B(p_input[403]), .Z(n19764) );
  XNOR U19663 ( .A(p_input[2068]), .B(p_input[404]), .Z(n19841) );
  XOR U19664 ( .A(p_input[2069]), .B(p_input[405]), .Z(n19768) );
  XNOR U19665 ( .A(n19783), .B(n19769), .Z(n19838) );
  XNOR U19666 ( .A(n16729), .B(p_input[385]), .Z(n19769) );
  XNOR U19667 ( .A(n19842), .B(n19790), .Z(n19783) );
  XNOR U19668 ( .A(n19779), .B(n19778), .Z(n19790) );
  XOR U19669 ( .A(n19843), .B(n19775), .Z(n19778) );
  XNOR U19670 ( .A(n16444), .B(p_input[410]), .Z(n19775) );
  XNOR U19671 ( .A(p_input[2075]), .B(p_input[411]), .Z(n19843) );
  XOR U19672 ( .A(p_input[2076]), .B(p_input[412]), .Z(n19779) );
  XNOR U19673 ( .A(n19789), .B(n19780), .Z(n19842) );
  XNOR U19674 ( .A(n16732), .B(p_input[401]), .Z(n19780) );
  XOR U19675 ( .A(n19844), .B(n19795), .Z(n19789) );
  XNOR U19676 ( .A(p_input[2079]), .B(p_input[415]), .Z(n19795) );
  XOR U19677 ( .A(n19786), .B(n19794), .Z(n19844) );
  XOR U19678 ( .A(n19845), .B(n19791), .Z(n19794) );
  XOR U19679 ( .A(p_input[2077]), .B(p_input[413]), .Z(n19791) );
  XNOR U19680 ( .A(p_input[2078]), .B(p_input[414]), .Z(n19845) );
  XNOR U19681 ( .A(n16448), .B(p_input[409]), .Z(n19786) );
  XNOR U19682 ( .A(n19807), .B(n19806), .Z(n19773) );
  XNOR U19683 ( .A(n19846), .B(n19813), .Z(n19806) );
  XNOR U19684 ( .A(n19802), .B(n19801), .Z(n19813) );
  XOR U19685 ( .A(n19847), .B(n19798), .Z(n19801) );
  XNOR U19686 ( .A(n16737), .B(p_input[395]), .Z(n19798) );
  XNOR U19687 ( .A(p_input[2060]), .B(p_input[396]), .Z(n19847) );
  XOR U19688 ( .A(p_input[2061]), .B(p_input[397]), .Z(n19802) );
  XNOR U19689 ( .A(n19812), .B(n19803), .Z(n19846) );
  XNOR U19690 ( .A(n16452), .B(p_input[386]), .Z(n19803) );
  XOR U19691 ( .A(n19848), .B(n19818), .Z(n19812) );
  XNOR U19692 ( .A(p_input[2064]), .B(p_input[400]), .Z(n19818) );
  XOR U19693 ( .A(n19809), .B(n19817), .Z(n19848) );
  XOR U19694 ( .A(n19849), .B(n19814), .Z(n19817) );
  XOR U19695 ( .A(p_input[2062]), .B(p_input[398]), .Z(n19814) );
  XNOR U19696 ( .A(p_input[2063]), .B(p_input[399]), .Z(n19849) );
  XNOR U19697 ( .A(n16740), .B(p_input[394]), .Z(n19809) );
  XNOR U19698 ( .A(n19824), .B(n19823), .Z(n19807) );
  XNOR U19699 ( .A(n19850), .B(n19829), .Z(n19823) );
  XOR U19700 ( .A(p_input[2057]), .B(p_input[393]), .Z(n19829) );
  XOR U19701 ( .A(n19820), .B(n19828), .Z(n19850) );
  XOR U19702 ( .A(n19851), .B(n19825), .Z(n19828) );
  XOR U19703 ( .A(p_input[2055]), .B(p_input[391]), .Z(n19825) );
  XNOR U19704 ( .A(p_input[2056]), .B(p_input[392]), .Z(n19851) );
  XNOR U19705 ( .A(n16459), .B(p_input[387]), .Z(n19820) );
  XNOR U19706 ( .A(n19834), .B(n19833), .Z(n19824) );
  XOR U19707 ( .A(n19852), .B(n19830), .Z(n19833) );
  XOR U19708 ( .A(p_input[2052]), .B(p_input[388]), .Z(n19830) );
  XNOR U19709 ( .A(p_input[2053]), .B(p_input[389]), .Z(n19852) );
  XOR U19710 ( .A(p_input[2054]), .B(p_input[390]), .Z(n19834) );
  XNOR U19711 ( .A(n19853), .B(n19854), .Z(n19651) );
  AND U19712 ( .A(n199), .B(n19855), .Z(n19854) );
  XNOR U19713 ( .A(n19856), .B(n19857), .Z(n199) );
  AND U19714 ( .A(n19858), .B(n19859), .Z(n19857) );
  XOR U19715 ( .A(n19856), .B(n19661), .Z(n19859) );
  XNOR U19716 ( .A(n19856), .B(n19603), .Z(n19858) );
  XOR U19717 ( .A(n19860), .B(n19861), .Z(n19856) );
  AND U19718 ( .A(n19862), .B(n19863), .Z(n19861) );
  XNOR U19719 ( .A(n19674), .B(n19860), .Z(n19863) );
  XOR U19720 ( .A(n19860), .B(n19615), .Z(n19862) );
  XOR U19721 ( .A(n19864), .B(n19865), .Z(n19860) );
  AND U19722 ( .A(n19866), .B(n19867), .Z(n19865) );
  XNOR U19723 ( .A(n19699), .B(n19864), .Z(n19867) );
  XOR U19724 ( .A(n19864), .B(n19626), .Z(n19866) );
  XOR U19725 ( .A(n19868), .B(n19869), .Z(n19864) );
  AND U19726 ( .A(n19870), .B(n19871), .Z(n19869) );
  XOR U19727 ( .A(n19868), .B(n19636), .Z(n19870) );
  XOR U19728 ( .A(n19872), .B(n19873), .Z(n19592) );
  AND U19729 ( .A(n203), .B(n19855), .Z(n19873) );
  XNOR U19730 ( .A(n19853), .B(n19872), .Z(n19855) );
  XNOR U19731 ( .A(n19874), .B(n19875), .Z(n203) );
  AND U19732 ( .A(n19876), .B(n19877), .Z(n19875) );
  XNOR U19733 ( .A(n19878), .B(n19874), .Z(n19877) );
  IV U19734 ( .A(n19661), .Z(n19878) );
  XNOR U19735 ( .A(n19879), .B(n19880), .Z(n19661) );
  AND U19736 ( .A(n206), .B(n19881), .Z(n19880) );
  XNOR U19737 ( .A(n19879), .B(n19882), .Z(n19881) );
  XNOR U19738 ( .A(n19603), .B(n19874), .Z(n19876) );
  XOR U19739 ( .A(n19883), .B(n19884), .Z(n19603) );
  AND U19740 ( .A(n214), .B(n19885), .Z(n19884) );
  XOR U19741 ( .A(n19886), .B(n19887), .Z(n19874) );
  AND U19742 ( .A(n19888), .B(n19889), .Z(n19887) );
  XNOR U19743 ( .A(n19886), .B(n19674), .Z(n19889) );
  XNOR U19744 ( .A(n19890), .B(n19891), .Z(n19674) );
  AND U19745 ( .A(n206), .B(n19892), .Z(n19891) );
  XOR U19746 ( .A(n19893), .B(n19890), .Z(n19892) );
  XNOR U19747 ( .A(n19894), .B(n19886), .Z(n19888) );
  IV U19748 ( .A(n19615), .Z(n19894) );
  XOR U19749 ( .A(n19895), .B(n19896), .Z(n19615) );
  AND U19750 ( .A(n214), .B(n19897), .Z(n19896) );
  XOR U19751 ( .A(n19898), .B(n19899), .Z(n19886) );
  AND U19752 ( .A(n19900), .B(n19901), .Z(n19899) );
  XNOR U19753 ( .A(n19898), .B(n19699), .Z(n19901) );
  XNOR U19754 ( .A(n19902), .B(n19903), .Z(n19699) );
  AND U19755 ( .A(n206), .B(n19904), .Z(n19903) );
  XNOR U19756 ( .A(n19905), .B(n19902), .Z(n19904) );
  XOR U19757 ( .A(n19626), .B(n19898), .Z(n19900) );
  XOR U19758 ( .A(n19906), .B(n19907), .Z(n19626) );
  AND U19759 ( .A(n214), .B(n19908), .Z(n19907) );
  XOR U19760 ( .A(n19868), .B(n19909), .Z(n19898) );
  AND U19761 ( .A(n19910), .B(n19871), .Z(n19909) );
  XNOR U19762 ( .A(n19745), .B(n19868), .Z(n19871) );
  XNOR U19763 ( .A(n19911), .B(n19912), .Z(n19745) );
  AND U19764 ( .A(n206), .B(n19913), .Z(n19912) );
  XOR U19765 ( .A(n19914), .B(n19911), .Z(n19913) );
  XNOR U19766 ( .A(n19915), .B(n19868), .Z(n19910) );
  IV U19767 ( .A(n19636), .Z(n19915) );
  XOR U19768 ( .A(n19916), .B(n19917), .Z(n19636) );
  AND U19769 ( .A(n214), .B(n19918), .Z(n19917) );
  XOR U19770 ( .A(n19919), .B(n19920), .Z(n19868) );
  AND U19771 ( .A(n19921), .B(n19922), .Z(n19920) );
  XNOR U19772 ( .A(n19919), .B(n19835), .Z(n19922) );
  XNOR U19773 ( .A(n19923), .B(n19924), .Z(n19835) );
  AND U19774 ( .A(n206), .B(n19925), .Z(n19924) );
  XNOR U19775 ( .A(n19926), .B(n19923), .Z(n19925) );
  XNOR U19776 ( .A(n19927), .B(n19919), .Z(n19921) );
  IV U19777 ( .A(n19648), .Z(n19927) );
  XOR U19778 ( .A(n19928), .B(n19929), .Z(n19648) );
  AND U19779 ( .A(n214), .B(n19930), .Z(n19929) );
  AND U19780 ( .A(n19872), .B(n19853), .Z(n19919) );
  XNOR U19781 ( .A(n19931), .B(n19932), .Z(n19853) );
  AND U19782 ( .A(n206), .B(n19933), .Z(n19932) );
  XNOR U19783 ( .A(n19934), .B(n19931), .Z(n19933) );
  XNOR U19784 ( .A(n19935), .B(n19936), .Z(n206) );
  AND U19785 ( .A(n19937), .B(n19938), .Z(n19936) );
  XOR U19786 ( .A(n19882), .B(n19935), .Z(n19938) );
  AND U19787 ( .A(n19939), .B(n19940), .Z(n19882) );
  XOR U19788 ( .A(n19935), .B(n19879), .Z(n19937) );
  XNOR U19789 ( .A(n19941), .B(n19942), .Z(n19879) );
  AND U19790 ( .A(n210), .B(n19885), .Z(n19942) );
  XOR U19791 ( .A(n19883), .B(n19941), .Z(n19885) );
  XOR U19792 ( .A(n19943), .B(n19944), .Z(n19935) );
  AND U19793 ( .A(n19945), .B(n19946), .Z(n19944) );
  XNOR U19794 ( .A(n19943), .B(n19939), .Z(n19946) );
  IV U19795 ( .A(n19893), .Z(n19939) );
  XOR U19796 ( .A(n19947), .B(n19948), .Z(n19893) );
  XOR U19797 ( .A(n19949), .B(n19940), .Z(n19948) );
  AND U19798 ( .A(n19905), .B(n19950), .Z(n19940) );
  AND U19799 ( .A(n19951), .B(n19952), .Z(n19949) );
  XOR U19800 ( .A(n19953), .B(n19947), .Z(n19951) );
  XNOR U19801 ( .A(n19890), .B(n19943), .Z(n19945) );
  XNOR U19802 ( .A(n19954), .B(n19955), .Z(n19890) );
  AND U19803 ( .A(n210), .B(n19897), .Z(n19955) );
  XOR U19804 ( .A(n19954), .B(n19895), .Z(n19897) );
  XOR U19805 ( .A(n19956), .B(n19957), .Z(n19943) );
  AND U19806 ( .A(n19958), .B(n19959), .Z(n19957) );
  XNOR U19807 ( .A(n19956), .B(n19905), .Z(n19959) );
  XOR U19808 ( .A(n19960), .B(n19952), .Z(n19905) );
  XNOR U19809 ( .A(n19961), .B(n19947), .Z(n19952) );
  XOR U19810 ( .A(n19962), .B(n19963), .Z(n19947) );
  AND U19811 ( .A(n19964), .B(n19965), .Z(n19963) );
  XOR U19812 ( .A(n19966), .B(n19962), .Z(n19964) );
  XNOR U19813 ( .A(n19967), .B(n19968), .Z(n19961) );
  AND U19814 ( .A(n19969), .B(n19970), .Z(n19968) );
  XOR U19815 ( .A(n19967), .B(n19971), .Z(n19969) );
  XNOR U19816 ( .A(n19953), .B(n19950), .Z(n19960) );
  AND U19817 ( .A(n19972), .B(n19973), .Z(n19950) );
  XOR U19818 ( .A(n19974), .B(n19975), .Z(n19953) );
  AND U19819 ( .A(n19976), .B(n19977), .Z(n19975) );
  XOR U19820 ( .A(n19974), .B(n19978), .Z(n19976) );
  XNOR U19821 ( .A(n19902), .B(n19956), .Z(n19958) );
  XNOR U19822 ( .A(n19979), .B(n19980), .Z(n19902) );
  AND U19823 ( .A(n210), .B(n19908), .Z(n19980) );
  XOR U19824 ( .A(n19979), .B(n19906), .Z(n19908) );
  XOR U19825 ( .A(n19981), .B(n19982), .Z(n19956) );
  AND U19826 ( .A(n19983), .B(n19984), .Z(n19982) );
  XNOR U19827 ( .A(n19981), .B(n19972), .Z(n19984) );
  IV U19828 ( .A(n19914), .Z(n19972) );
  XNOR U19829 ( .A(n19985), .B(n19965), .Z(n19914) );
  XNOR U19830 ( .A(n19986), .B(n19971), .Z(n19965) );
  XOR U19831 ( .A(n19987), .B(n19988), .Z(n19971) );
  AND U19832 ( .A(n19989), .B(n19990), .Z(n19988) );
  XOR U19833 ( .A(n19987), .B(n19991), .Z(n19989) );
  XNOR U19834 ( .A(n19970), .B(n19962), .Z(n19986) );
  XOR U19835 ( .A(n19992), .B(n19993), .Z(n19962) );
  AND U19836 ( .A(n19994), .B(n19995), .Z(n19993) );
  XNOR U19837 ( .A(n19996), .B(n19992), .Z(n19994) );
  XNOR U19838 ( .A(n19997), .B(n19967), .Z(n19970) );
  XOR U19839 ( .A(n19998), .B(n19999), .Z(n19967) );
  AND U19840 ( .A(n20000), .B(n20001), .Z(n19999) );
  XOR U19841 ( .A(n19998), .B(n20002), .Z(n20000) );
  XNOR U19842 ( .A(n20003), .B(n20004), .Z(n19997) );
  AND U19843 ( .A(n20005), .B(n20006), .Z(n20004) );
  XNOR U19844 ( .A(n20003), .B(n20007), .Z(n20005) );
  XNOR U19845 ( .A(n19966), .B(n19973), .Z(n19985) );
  AND U19846 ( .A(n19926), .B(n20008), .Z(n19973) );
  XOR U19847 ( .A(n19978), .B(n19977), .Z(n19966) );
  XNOR U19848 ( .A(n20009), .B(n19974), .Z(n19977) );
  XOR U19849 ( .A(n20010), .B(n20011), .Z(n19974) );
  AND U19850 ( .A(n20012), .B(n20013), .Z(n20011) );
  XOR U19851 ( .A(n20010), .B(n20014), .Z(n20012) );
  XNOR U19852 ( .A(n20015), .B(n20016), .Z(n20009) );
  AND U19853 ( .A(n20017), .B(n20018), .Z(n20016) );
  XOR U19854 ( .A(n20015), .B(n20019), .Z(n20017) );
  XOR U19855 ( .A(n20020), .B(n20021), .Z(n19978) );
  AND U19856 ( .A(n20022), .B(n20023), .Z(n20021) );
  XOR U19857 ( .A(n20020), .B(n20024), .Z(n20022) );
  XNOR U19858 ( .A(n19911), .B(n19981), .Z(n19983) );
  XNOR U19859 ( .A(n20025), .B(n20026), .Z(n19911) );
  AND U19860 ( .A(n210), .B(n19918), .Z(n20026) );
  XOR U19861 ( .A(n20025), .B(n19916), .Z(n19918) );
  XOR U19862 ( .A(n20027), .B(n20028), .Z(n19981) );
  AND U19863 ( .A(n20029), .B(n20030), .Z(n20028) );
  XNOR U19864 ( .A(n20027), .B(n19926), .Z(n20030) );
  XOR U19865 ( .A(n20031), .B(n19995), .Z(n19926) );
  XNOR U19866 ( .A(n20032), .B(n20002), .Z(n19995) );
  XOR U19867 ( .A(n19991), .B(n19990), .Z(n20002) );
  XNOR U19868 ( .A(n20033), .B(n19987), .Z(n19990) );
  XOR U19869 ( .A(n20034), .B(n20035), .Z(n19987) );
  AND U19870 ( .A(n20036), .B(n20037), .Z(n20035) );
  XOR U19871 ( .A(n20034), .B(n20038), .Z(n20036) );
  XNOR U19872 ( .A(n20039), .B(n20040), .Z(n20033) );
  NOR U19873 ( .A(n20041), .B(n20042), .Z(n20040) );
  XNOR U19874 ( .A(n20039), .B(n20043), .Z(n20041) );
  XOR U19875 ( .A(n20044), .B(n20045), .Z(n19991) );
  NOR U19876 ( .A(n20046), .B(n20047), .Z(n20045) );
  XNOR U19877 ( .A(n20044), .B(n20048), .Z(n20046) );
  XNOR U19878 ( .A(n20001), .B(n19992), .Z(n20032) );
  XOR U19879 ( .A(n20049), .B(n20050), .Z(n19992) );
  NOR U19880 ( .A(n20051), .B(n20052), .Z(n20050) );
  XNOR U19881 ( .A(n20049), .B(n20053), .Z(n20051) );
  XOR U19882 ( .A(n20054), .B(n20007), .Z(n20001) );
  XNOR U19883 ( .A(n20055), .B(n20056), .Z(n20007) );
  NOR U19884 ( .A(n20057), .B(n20058), .Z(n20056) );
  XNOR U19885 ( .A(n20055), .B(n20059), .Z(n20057) );
  XNOR U19886 ( .A(n20006), .B(n19998), .Z(n20054) );
  XOR U19887 ( .A(n20060), .B(n20061), .Z(n19998) );
  AND U19888 ( .A(n20062), .B(n20063), .Z(n20061) );
  XOR U19889 ( .A(n20060), .B(n20064), .Z(n20062) );
  XNOR U19890 ( .A(n20065), .B(n20003), .Z(n20006) );
  XOR U19891 ( .A(n20066), .B(n20067), .Z(n20003) );
  AND U19892 ( .A(n20068), .B(n20069), .Z(n20067) );
  XOR U19893 ( .A(n20066), .B(n20070), .Z(n20068) );
  XNOR U19894 ( .A(n20071), .B(n20072), .Z(n20065) );
  NOR U19895 ( .A(n20073), .B(n20074), .Z(n20072) );
  XOR U19896 ( .A(n20071), .B(n20075), .Z(n20073) );
  XOR U19897 ( .A(n19996), .B(n20008), .Z(n20031) );
  NOR U19898 ( .A(n19934), .B(n20076), .Z(n20008) );
  XNOR U19899 ( .A(n20014), .B(n20013), .Z(n19996) );
  XNOR U19900 ( .A(n20077), .B(n20019), .Z(n20013) );
  XOR U19901 ( .A(n20078), .B(n20079), .Z(n20019) );
  NOR U19902 ( .A(n20080), .B(n20081), .Z(n20079) );
  XNOR U19903 ( .A(n20078), .B(n20082), .Z(n20080) );
  XNOR U19904 ( .A(n20018), .B(n20010), .Z(n20077) );
  XOR U19905 ( .A(n20083), .B(n20084), .Z(n20010) );
  AND U19906 ( .A(n20085), .B(n20086), .Z(n20084) );
  XNOR U19907 ( .A(n20083), .B(n20087), .Z(n20085) );
  XNOR U19908 ( .A(n20088), .B(n20015), .Z(n20018) );
  XOR U19909 ( .A(n20089), .B(n20090), .Z(n20015) );
  AND U19910 ( .A(n20091), .B(n20092), .Z(n20090) );
  XOR U19911 ( .A(n20089), .B(n20093), .Z(n20091) );
  XNOR U19912 ( .A(n20094), .B(n20095), .Z(n20088) );
  NOR U19913 ( .A(n20096), .B(n20097), .Z(n20095) );
  XOR U19914 ( .A(n20094), .B(n20098), .Z(n20096) );
  XOR U19915 ( .A(n20024), .B(n20023), .Z(n20014) );
  XNOR U19916 ( .A(n20099), .B(n20020), .Z(n20023) );
  XOR U19917 ( .A(n20100), .B(n20101), .Z(n20020) );
  AND U19918 ( .A(n20102), .B(n20103), .Z(n20101) );
  XOR U19919 ( .A(n20100), .B(n20104), .Z(n20102) );
  XNOR U19920 ( .A(n20105), .B(n20106), .Z(n20099) );
  NOR U19921 ( .A(n20107), .B(n20108), .Z(n20106) );
  XNOR U19922 ( .A(n20105), .B(n20109), .Z(n20107) );
  XOR U19923 ( .A(n20110), .B(n20111), .Z(n20024) );
  NOR U19924 ( .A(n20112), .B(n20113), .Z(n20111) );
  XNOR U19925 ( .A(n20110), .B(n20114), .Z(n20112) );
  XNOR U19926 ( .A(n19923), .B(n20027), .Z(n20029) );
  XNOR U19927 ( .A(n20115), .B(n20116), .Z(n19923) );
  AND U19928 ( .A(n210), .B(n19930), .Z(n20116) );
  XOR U19929 ( .A(n20115), .B(n19928), .Z(n19930) );
  AND U19930 ( .A(n19931), .B(n19934), .Z(n20027) );
  XOR U19931 ( .A(n20117), .B(n20076), .Z(n19934) );
  XNOR U19932 ( .A(p_input[2048]), .B(p_input[416]), .Z(n20076) );
  XOR U19933 ( .A(n20053), .B(n20052), .Z(n20117) );
  XOR U19934 ( .A(n20118), .B(n20064), .Z(n20052) );
  XOR U19935 ( .A(n20038), .B(n20037), .Z(n20064) );
  XNOR U19936 ( .A(n20119), .B(n20043), .Z(n20037) );
  XOR U19937 ( .A(p_input[2072]), .B(p_input[440]), .Z(n20043) );
  XOR U19938 ( .A(n20034), .B(n20042), .Z(n20119) );
  XOR U19939 ( .A(n20120), .B(n20039), .Z(n20042) );
  XOR U19940 ( .A(p_input[2070]), .B(p_input[438]), .Z(n20039) );
  XNOR U19941 ( .A(p_input[2071]), .B(p_input[439]), .Z(n20120) );
  XNOR U19942 ( .A(n16727), .B(p_input[434]), .Z(n20034) );
  XNOR U19943 ( .A(n20048), .B(n20047), .Z(n20038) );
  XOR U19944 ( .A(n20121), .B(n20044), .Z(n20047) );
  XOR U19945 ( .A(p_input[2067]), .B(p_input[435]), .Z(n20044) );
  XNOR U19946 ( .A(p_input[2068]), .B(p_input[436]), .Z(n20121) );
  XOR U19947 ( .A(p_input[2069]), .B(p_input[437]), .Z(n20048) );
  XNOR U19948 ( .A(n20063), .B(n20049), .Z(n20118) );
  XNOR U19949 ( .A(n16729), .B(p_input[417]), .Z(n20049) );
  XNOR U19950 ( .A(n20122), .B(n20070), .Z(n20063) );
  XNOR U19951 ( .A(n20059), .B(n20058), .Z(n20070) );
  XOR U19952 ( .A(n20123), .B(n20055), .Z(n20058) );
  XNOR U19953 ( .A(n16444), .B(p_input[442]), .Z(n20055) );
  XNOR U19954 ( .A(p_input[2075]), .B(p_input[443]), .Z(n20123) );
  XOR U19955 ( .A(p_input[2076]), .B(p_input[444]), .Z(n20059) );
  XNOR U19956 ( .A(n20069), .B(n20060), .Z(n20122) );
  XNOR U19957 ( .A(n16732), .B(p_input[433]), .Z(n20060) );
  XOR U19958 ( .A(n20124), .B(n20075), .Z(n20069) );
  XNOR U19959 ( .A(p_input[2079]), .B(p_input[447]), .Z(n20075) );
  XOR U19960 ( .A(n20066), .B(n20074), .Z(n20124) );
  XOR U19961 ( .A(n20125), .B(n20071), .Z(n20074) );
  XOR U19962 ( .A(p_input[2077]), .B(p_input[445]), .Z(n20071) );
  XNOR U19963 ( .A(p_input[2078]), .B(p_input[446]), .Z(n20125) );
  XNOR U19964 ( .A(n16448), .B(p_input[441]), .Z(n20066) );
  XNOR U19965 ( .A(n20087), .B(n20086), .Z(n20053) );
  XNOR U19966 ( .A(n20126), .B(n20093), .Z(n20086) );
  XNOR U19967 ( .A(n20082), .B(n20081), .Z(n20093) );
  XOR U19968 ( .A(n20127), .B(n20078), .Z(n20081) );
  XNOR U19969 ( .A(n16737), .B(p_input[427]), .Z(n20078) );
  XNOR U19970 ( .A(p_input[2060]), .B(p_input[428]), .Z(n20127) );
  XOR U19971 ( .A(p_input[2061]), .B(p_input[429]), .Z(n20082) );
  XNOR U19972 ( .A(n20092), .B(n20083), .Z(n20126) );
  XNOR U19973 ( .A(n16452), .B(p_input[418]), .Z(n20083) );
  XOR U19974 ( .A(n20128), .B(n20098), .Z(n20092) );
  XNOR U19975 ( .A(p_input[2064]), .B(p_input[432]), .Z(n20098) );
  XOR U19976 ( .A(n20089), .B(n20097), .Z(n20128) );
  XOR U19977 ( .A(n20129), .B(n20094), .Z(n20097) );
  XOR U19978 ( .A(p_input[2062]), .B(p_input[430]), .Z(n20094) );
  XNOR U19979 ( .A(p_input[2063]), .B(p_input[431]), .Z(n20129) );
  XNOR U19980 ( .A(n16740), .B(p_input[426]), .Z(n20089) );
  XNOR U19981 ( .A(n20104), .B(n20103), .Z(n20087) );
  XNOR U19982 ( .A(n20130), .B(n20109), .Z(n20103) );
  XOR U19983 ( .A(p_input[2057]), .B(p_input[425]), .Z(n20109) );
  XOR U19984 ( .A(n20100), .B(n20108), .Z(n20130) );
  XOR U19985 ( .A(n20131), .B(n20105), .Z(n20108) );
  XOR U19986 ( .A(p_input[2055]), .B(p_input[423]), .Z(n20105) );
  XNOR U19987 ( .A(p_input[2056]), .B(p_input[424]), .Z(n20131) );
  XNOR U19988 ( .A(n16459), .B(p_input[419]), .Z(n20100) );
  XNOR U19989 ( .A(n20114), .B(n20113), .Z(n20104) );
  XOR U19990 ( .A(n20132), .B(n20110), .Z(n20113) );
  XOR U19991 ( .A(p_input[2052]), .B(p_input[420]), .Z(n20110) );
  XNOR U19992 ( .A(p_input[2053]), .B(p_input[421]), .Z(n20132) );
  XOR U19993 ( .A(p_input[2054]), .B(p_input[422]), .Z(n20114) );
  XNOR U19994 ( .A(n20133), .B(n20134), .Z(n19931) );
  AND U19995 ( .A(n210), .B(n20135), .Z(n20134) );
  XNOR U19996 ( .A(n20136), .B(n20137), .Z(n210) );
  AND U19997 ( .A(n20138), .B(n20139), .Z(n20137) );
  XOR U19998 ( .A(n20136), .B(n19941), .Z(n20139) );
  XNOR U19999 ( .A(n20136), .B(n19883), .Z(n20138) );
  XOR U20000 ( .A(n20140), .B(n20141), .Z(n20136) );
  AND U20001 ( .A(n20142), .B(n20143), .Z(n20141) );
  XNOR U20002 ( .A(n19954), .B(n20140), .Z(n20143) );
  XOR U20003 ( .A(n20140), .B(n19895), .Z(n20142) );
  XOR U20004 ( .A(n20144), .B(n20145), .Z(n20140) );
  AND U20005 ( .A(n20146), .B(n20147), .Z(n20145) );
  XNOR U20006 ( .A(n19979), .B(n20144), .Z(n20147) );
  XOR U20007 ( .A(n20144), .B(n19906), .Z(n20146) );
  XOR U20008 ( .A(n20148), .B(n20149), .Z(n20144) );
  AND U20009 ( .A(n20150), .B(n20151), .Z(n20149) );
  XOR U20010 ( .A(n20148), .B(n19916), .Z(n20150) );
  XOR U20011 ( .A(n20152), .B(n20153), .Z(n19872) );
  AND U20012 ( .A(n214), .B(n20135), .Z(n20153) );
  XNOR U20013 ( .A(n20133), .B(n20152), .Z(n20135) );
  XNOR U20014 ( .A(n20154), .B(n20155), .Z(n214) );
  AND U20015 ( .A(n20156), .B(n20157), .Z(n20155) );
  XNOR U20016 ( .A(n20158), .B(n20154), .Z(n20157) );
  IV U20017 ( .A(n19941), .Z(n20158) );
  XNOR U20018 ( .A(n20159), .B(n20160), .Z(n19941) );
  AND U20019 ( .A(n217), .B(n20161), .Z(n20160) );
  XNOR U20020 ( .A(n20159), .B(n20162), .Z(n20161) );
  XNOR U20021 ( .A(n19883), .B(n20154), .Z(n20156) );
  XOR U20022 ( .A(n20163), .B(n20164), .Z(n19883) );
  AND U20023 ( .A(n225), .B(n20165), .Z(n20164) );
  XOR U20024 ( .A(n20166), .B(n20167), .Z(n20154) );
  AND U20025 ( .A(n20168), .B(n20169), .Z(n20167) );
  XNOR U20026 ( .A(n20166), .B(n19954), .Z(n20169) );
  XNOR U20027 ( .A(n20170), .B(n20171), .Z(n19954) );
  AND U20028 ( .A(n217), .B(n20172), .Z(n20171) );
  XOR U20029 ( .A(n20173), .B(n20170), .Z(n20172) );
  XNOR U20030 ( .A(n20174), .B(n20166), .Z(n20168) );
  IV U20031 ( .A(n19895), .Z(n20174) );
  XOR U20032 ( .A(n20175), .B(n20176), .Z(n19895) );
  AND U20033 ( .A(n225), .B(n20177), .Z(n20176) );
  XOR U20034 ( .A(n20178), .B(n20179), .Z(n20166) );
  AND U20035 ( .A(n20180), .B(n20181), .Z(n20179) );
  XNOR U20036 ( .A(n20178), .B(n19979), .Z(n20181) );
  XNOR U20037 ( .A(n20182), .B(n20183), .Z(n19979) );
  AND U20038 ( .A(n217), .B(n20184), .Z(n20183) );
  XNOR U20039 ( .A(n20185), .B(n20182), .Z(n20184) );
  XOR U20040 ( .A(n19906), .B(n20178), .Z(n20180) );
  XOR U20041 ( .A(n20186), .B(n20187), .Z(n19906) );
  AND U20042 ( .A(n225), .B(n20188), .Z(n20187) );
  XOR U20043 ( .A(n20148), .B(n20189), .Z(n20178) );
  AND U20044 ( .A(n20190), .B(n20151), .Z(n20189) );
  XNOR U20045 ( .A(n20025), .B(n20148), .Z(n20151) );
  XNOR U20046 ( .A(n20191), .B(n20192), .Z(n20025) );
  AND U20047 ( .A(n217), .B(n20193), .Z(n20192) );
  XOR U20048 ( .A(n20194), .B(n20191), .Z(n20193) );
  XNOR U20049 ( .A(n20195), .B(n20148), .Z(n20190) );
  IV U20050 ( .A(n19916), .Z(n20195) );
  XOR U20051 ( .A(n20196), .B(n20197), .Z(n19916) );
  AND U20052 ( .A(n225), .B(n20198), .Z(n20197) );
  XOR U20053 ( .A(n20199), .B(n20200), .Z(n20148) );
  AND U20054 ( .A(n20201), .B(n20202), .Z(n20200) );
  XNOR U20055 ( .A(n20199), .B(n20115), .Z(n20202) );
  XNOR U20056 ( .A(n20203), .B(n20204), .Z(n20115) );
  AND U20057 ( .A(n217), .B(n20205), .Z(n20204) );
  XNOR U20058 ( .A(n20206), .B(n20203), .Z(n20205) );
  XNOR U20059 ( .A(n20207), .B(n20199), .Z(n20201) );
  IV U20060 ( .A(n19928), .Z(n20207) );
  XOR U20061 ( .A(n20208), .B(n20209), .Z(n19928) );
  AND U20062 ( .A(n225), .B(n20210), .Z(n20209) );
  AND U20063 ( .A(n20152), .B(n20133), .Z(n20199) );
  XNOR U20064 ( .A(n20211), .B(n20212), .Z(n20133) );
  AND U20065 ( .A(n217), .B(n20213), .Z(n20212) );
  XNOR U20066 ( .A(n20214), .B(n20211), .Z(n20213) );
  XNOR U20067 ( .A(n20215), .B(n20216), .Z(n217) );
  AND U20068 ( .A(n20217), .B(n20218), .Z(n20216) );
  XOR U20069 ( .A(n20162), .B(n20215), .Z(n20218) );
  AND U20070 ( .A(n20219), .B(n20220), .Z(n20162) );
  XOR U20071 ( .A(n20215), .B(n20159), .Z(n20217) );
  XNOR U20072 ( .A(n20221), .B(n20222), .Z(n20159) );
  AND U20073 ( .A(n221), .B(n20165), .Z(n20222) );
  XOR U20074 ( .A(n20163), .B(n20221), .Z(n20165) );
  XOR U20075 ( .A(n20223), .B(n20224), .Z(n20215) );
  AND U20076 ( .A(n20225), .B(n20226), .Z(n20224) );
  XNOR U20077 ( .A(n20223), .B(n20219), .Z(n20226) );
  IV U20078 ( .A(n20173), .Z(n20219) );
  XOR U20079 ( .A(n20227), .B(n20228), .Z(n20173) );
  XOR U20080 ( .A(n20229), .B(n20220), .Z(n20228) );
  AND U20081 ( .A(n20185), .B(n20230), .Z(n20220) );
  AND U20082 ( .A(n20231), .B(n20232), .Z(n20229) );
  XOR U20083 ( .A(n20233), .B(n20227), .Z(n20231) );
  XNOR U20084 ( .A(n20170), .B(n20223), .Z(n20225) );
  XNOR U20085 ( .A(n20234), .B(n20235), .Z(n20170) );
  AND U20086 ( .A(n221), .B(n20177), .Z(n20235) );
  XOR U20087 ( .A(n20234), .B(n20175), .Z(n20177) );
  XOR U20088 ( .A(n20236), .B(n20237), .Z(n20223) );
  AND U20089 ( .A(n20238), .B(n20239), .Z(n20237) );
  XNOR U20090 ( .A(n20236), .B(n20185), .Z(n20239) );
  XOR U20091 ( .A(n20240), .B(n20232), .Z(n20185) );
  XNOR U20092 ( .A(n20241), .B(n20227), .Z(n20232) );
  XOR U20093 ( .A(n20242), .B(n20243), .Z(n20227) );
  AND U20094 ( .A(n20244), .B(n20245), .Z(n20243) );
  XOR U20095 ( .A(n20246), .B(n20242), .Z(n20244) );
  XNOR U20096 ( .A(n20247), .B(n20248), .Z(n20241) );
  AND U20097 ( .A(n20249), .B(n20250), .Z(n20248) );
  XOR U20098 ( .A(n20247), .B(n20251), .Z(n20249) );
  XNOR U20099 ( .A(n20233), .B(n20230), .Z(n20240) );
  AND U20100 ( .A(n20252), .B(n20253), .Z(n20230) );
  XOR U20101 ( .A(n20254), .B(n20255), .Z(n20233) );
  AND U20102 ( .A(n20256), .B(n20257), .Z(n20255) );
  XOR U20103 ( .A(n20254), .B(n20258), .Z(n20256) );
  XNOR U20104 ( .A(n20182), .B(n20236), .Z(n20238) );
  XNOR U20105 ( .A(n20259), .B(n20260), .Z(n20182) );
  AND U20106 ( .A(n221), .B(n20188), .Z(n20260) );
  XOR U20107 ( .A(n20259), .B(n20186), .Z(n20188) );
  XOR U20108 ( .A(n20261), .B(n20262), .Z(n20236) );
  AND U20109 ( .A(n20263), .B(n20264), .Z(n20262) );
  XNOR U20110 ( .A(n20261), .B(n20252), .Z(n20264) );
  IV U20111 ( .A(n20194), .Z(n20252) );
  XNOR U20112 ( .A(n20265), .B(n20245), .Z(n20194) );
  XNOR U20113 ( .A(n20266), .B(n20251), .Z(n20245) );
  XOR U20114 ( .A(n20267), .B(n20268), .Z(n20251) );
  AND U20115 ( .A(n20269), .B(n20270), .Z(n20268) );
  XOR U20116 ( .A(n20267), .B(n20271), .Z(n20269) );
  XNOR U20117 ( .A(n20250), .B(n20242), .Z(n20266) );
  XOR U20118 ( .A(n20272), .B(n20273), .Z(n20242) );
  AND U20119 ( .A(n20274), .B(n20275), .Z(n20273) );
  XNOR U20120 ( .A(n20276), .B(n20272), .Z(n20274) );
  XNOR U20121 ( .A(n20277), .B(n20247), .Z(n20250) );
  XOR U20122 ( .A(n20278), .B(n20279), .Z(n20247) );
  AND U20123 ( .A(n20280), .B(n20281), .Z(n20279) );
  XOR U20124 ( .A(n20278), .B(n20282), .Z(n20280) );
  XNOR U20125 ( .A(n20283), .B(n20284), .Z(n20277) );
  AND U20126 ( .A(n20285), .B(n20286), .Z(n20284) );
  XNOR U20127 ( .A(n20283), .B(n20287), .Z(n20285) );
  XNOR U20128 ( .A(n20246), .B(n20253), .Z(n20265) );
  AND U20129 ( .A(n20206), .B(n20288), .Z(n20253) );
  XOR U20130 ( .A(n20258), .B(n20257), .Z(n20246) );
  XNOR U20131 ( .A(n20289), .B(n20254), .Z(n20257) );
  XOR U20132 ( .A(n20290), .B(n20291), .Z(n20254) );
  AND U20133 ( .A(n20292), .B(n20293), .Z(n20291) );
  XOR U20134 ( .A(n20290), .B(n20294), .Z(n20292) );
  XNOR U20135 ( .A(n20295), .B(n20296), .Z(n20289) );
  AND U20136 ( .A(n20297), .B(n20298), .Z(n20296) );
  XOR U20137 ( .A(n20295), .B(n20299), .Z(n20297) );
  XOR U20138 ( .A(n20300), .B(n20301), .Z(n20258) );
  AND U20139 ( .A(n20302), .B(n20303), .Z(n20301) );
  XOR U20140 ( .A(n20300), .B(n20304), .Z(n20302) );
  XNOR U20141 ( .A(n20191), .B(n20261), .Z(n20263) );
  XNOR U20142 ( .A(n20305), .B(n20306), .Z(n20191) );
  AND U20143 ( .A(n221), .B(n20198), .Z(n20306) );
  XOR U20144 ( .A(n20305), .B(n20196), .Z(n20198) );
  XOR U20145 ( .A(n20307), .B(n20308), .Z(n20261) );
  AND U20146 ( .A(n20309), .B(n20310), .Z(n20308) );
  XNOR U20147 ( .A(n20307), .B(n20206), .Z(n20310) );
  XOR U20148 ( .A(n20311), .B(n20275), .Z(n20206) );
  XNOR U20149 ( .A(n20312), .B(n20282), .Z(n20275) );
  XOR U20150 ( .A(n20271), .B(n20270), .Z(n20282) );
  XNOR U20151 ( .A(n20313), .B(n20267), .Z(n20270) );
  XOR U20152 ( .A(n20314), .B(n20315), .Z(n20267) );
  AND U20153 ( .A(n20316), .B(n20317), .Z(n20315) );
  XOR U20154 ( .A(n20314), .B(n20318), .Z(n20316) );
  XNOR U20155 ( .A(n20319), .B(n20320), .Z(n20313) );
  NOR U20156 ( .A(n20321), .B(n20322), .Z(n20320) );
  XNOR U20157 ( .A(n20319), .B(n20323), .Z(n20321) );
  XOR U20158 ( .A(n20324), .B(n20325), .Z(n20271) );
  NOR U20159 ( .A(n20326), .B(n20327), .Z(n20325) );
  XNOR U20160 ( .A(n20324), .B(n20328), .Z(n20326) );
  XNOR U20161 ( .A(n20281), .B(n20272), .Z(n20312) );
  XOR U20162 ( .A(n20329), .B(n20330), .Z(n20272) );
  NOR U20163 ( .A(n20331), .B(n20332), .Z(n20330) );
  XNOR U20164 ( .A(n20329), .B(n20333), .Z(n20331) );
  XOR U20165 ( .A(n20334), .B(n20287), .Z(n20281) );
  XNOR U20166 ( .A(n20335), .B(n20336), .Z(n20287) );
  NOR U20167 ( .A(n20337), .B(n20338), .Z(n20336) );
  XNOR U20168 ( .A(n20335), .B(n20339), .Z(n20337) );
  XNOR U20169 ( .A(n20286), .B(n20278), .Z(n20334) );
  XOR U20170 ( .A(n20340), .B(n20341), .Z(n20278) );
  AND U20171 ( .A(n20342), .B(n20343), .Z(n20341) );
  XOR U20172 ( .A(n20340), .B(n20344), .Z(n20342) );
  XNOR U20173 ( .A(n20345), .B(n20283), .Z(n20286) );
  XOR U20174 ( .A(n20346), .B(n20347), .Z(n20283) );
  AND U20175 ( .A(n20348), .B(n20349), .Z(n20347) );
  XOR U20176 ( .A(n20346), .B(n20350), .Z(n20348) );
  XNOR U20177 ( .A(n20351), .B(n20352), .Z(n20345) );
  NOR U20178 ( .A(n20353), .B(n20354), .Z(n20352) );
  XOR U20179 ( .A(n20351), .B(n20355), .Z(n20353) );
  XOR U20180 ( .A(n20276), .B(n20288), .Z(n20311) );
  NOR U20181 ( .A(n20214), .B(n20356), .Z(n20288) );
  XNOR U20182 ( .A(n20294), .B(n20293), .Z(n20276) );
  XNOR U20183 ( .A(n20357), .B(n20299), .Z(n20293) );
  XOR U20184 ( .A(n20358), .B(n20359), .Z(n20299) );
  NOR U20185 ( .A(n20360), .B(n20361), .Z(n20359) );
  XNOR U20186 ( .A(n20358), .B(n20362), .Z(n20360) );
  XNOR U20187 ( .A(n20298), .B(n20290), .Z(n20357) );
  XOR U20188 ( .A(n20363), .B(n20364), .Z(n20290) );
  AND U20189 ( .A(n20365), .B(n20366), .Z(n20364) );
  XNOR U20190 ( .A(n20363), .B(n20367), .Z(n20365) );
  XNOR U20191 ( .A(n20368), .B(n20295), .Z(n20298) );
  XOR U20192 ( .A(n20369), .B(n20370), .Z(n20295) );
  AND U20193 ( .A(n20371), .B(n20372), .Z(n20370) );
  XOR U20194 ( .A(n20369), .B(n20373), .Z(n20371) );
  XNOR U20195 ( .A(n20374), .B(n20375), .Z(n20368) );
  NOR U20196 ( .A(n20376), .B(n20377), .Z(n20375) );
  XOR U20197 ( .A(n20374), .B(n20378), .Z(n20376) );
  XOR U20198 ( .A(n20304), .B(n20303), .Z(n20294) );
  XNOR U20199 ( .A(n20379), .B(n20300), .Z(n20303) );
  XOR U20200 ( .A(n20380), .B(n20381), .Z(n20300) );
  AND U20201 ( .A(n20382), .B(n20383), .Z(n20381) );
  XOR U20202 ( .A(n20380), .B(n20384), .Z(n20382) );
  XNOR U20203 ( .A(n20385), .B(n20386), .Z(n20379) );
  NOR U20204 ( .A(n20387), .B(n20388), .Z(n20386) );
  XNOR U20205 ( .A(n20385), .B(n20389), .Z(n20387) );
  XOR U20206 ( .A(n20390), .B(n20391), .Z(n20304) );
  NOR U20207 ( .A(n20392), .B(n20393), .Z(n20391) );
  XNOR U20208 ( .A(n20390), .B(n20394), .Z(n20392) );
  XNOR U20209 ( .A(n20203), .B(n20307), .Z(n20309) );
  XNOR U20210 ( .A(n20395), .B(n20396), .Z(n20203) );
  AND U20211 ( .A(n221), .B(n20210), .Z(n20396) );
  XOR U20212 ( .A(n20395), .B(n20208), .Z(n20210) );
  AND U20213 ( .A(n20211), .B(n20214), .Z(n20307) );
  XOR U20214 ( .A(n20397), .B(n20356), .Z(n20214) );
  XNOR U20215 ( .A(p_input[2048]), .B(p_input[448]), .Z(n20356) );
  XOR U20216 ( .A(n20333), .B(n20332), .Z(n20397) );
  XOR U20217 ( .A(n20398), .B(n20344), .Z(n20332) );
  XOR U20218 ( .A(n20318), .B(n20317), .Z(n20344) );
  XNOR U20219 ( .A(n20399), .B(n20323), .Z(n20317) );
  XOR U20220 ( .A(p_input[2072]), .B(p_input[472]), .Z(n20323) );
  XOR U20221 ( .A(n20314), .B(n20322), .Z(n20399) );
  XOR U20222 ( .A(n20400), .B(n20319), .Z(n20322) );
  XOR U20223 ( .A(p_input[2070]), .B(p_input[470]), .Z(n20319) );
  XNOR U20224 ( .A(p_input[2071]), .B(p_input[471]), .Z(n20400) );
  XNOR U20225 ( .A(n16727), .B(p_input[466]), .Z(n20314) );
  XNOR U20226 ( .A(n20328), .B(n20327), .Z(n20318) );
  XOR U20227 ( .A(n20401), .B(n20324), .Z(n20327) );
  XOR U20228 ( .A(p_input[2067]), .B(p_input[467]), .Z(n20324) );
  XNOR U20229 ( .A(p_input[2068]), .B(p_input[468]), .Z(n20401) );
  XOR U20230 ( .A(p_input[2069]), .B(p_input[469]), .Z(n20328) );
  XNOR U20231 ( .A(n20343), .B(n20329), .Z(n20398) );
  XNOR U20232 ( .A(n16729), .B(p_input[449]), .Z(n20329) );
  XNOR U20233 ( .A(n20402), .B(n20350), .Z(n20343) );
  XNOR U20234 ( .A(n20339), .B(n20338), .Z(n20350) );
  XOR U20235 ( .A(n20403), .B(n20335), .Z(n20338) );
  XNOR U20236 ( .A(n16444), .B(p_input[474]), .Z(n20335) );
  XNOR U20237 ( .A(p_input[2075]), .B(p_input[475]), .Z(n20403) );
  XOR U20238 ( .A(p_input[2076]), .B(p_input[476]), .Z(n20339) );
  XNOR U20239 ( .A(n20349), .B(n20340), .Z(n20402) );
  XNOR U20240 ( .A(n16732), .B(p_input[465]), .Z(n20340) );
  XOR U20241 ( .A(n20404), .B(n20355), .Z(n20349) );
  XNOR U20242 ( .A(p_input[2079]), .B(p_input[479]), .Z(n20355) );
  XOR U20243 ( .A(n20346), .B(n20354), .Z(n20404) );
  XOR U20244 ( .A(n20405), .B(n20351), .Z(n20354) );
  XOR U20245 ( .A(p_input[2077]), .B(p_input[477]), .Z(n20351) );
  XNOR U20246 ( .A(p_input[2078]), .B(p_input[478]), .Z(n20405) );
  XNOR U20247 ( .A(n16448), .B(p_input[473]), .Z(n20346) );
  XNOR U20248 ( .A(n20367), .B(n20366), .Z(n20333) );
  XNOR U20249 ( .A(n20406), .B(n20373), .Z(n20366) );
  XNOR U20250 ( .A(n20362), .B(n20361), .Z(n20373) );
  XOR U20251 ( .A(n20407), .B(n20358), .Z(n20361) );
  XNOR U20252 ( .A(n16737), .B(p_input[459]), .Z(n20358) );
  XNOR U20253 ( .A(p_input[2060]), .B(p_input[460]), .Z(n20407) );
  XOR U20254 ( .A(p_input[2061]), .B(p_input[461]), .Z(n20362) );
  XNOR U20255 ( .A(n20372), .B(n20363), .Z(n20406) );
  XNOR U20256 ( .A(n16452), .B(p_input[450]), .Z(n20363) );
  XOR U20257 ( .A(n20408), .B(n20378), .Z(n20372) );
  XNOR U20258 ( .A(p_input[2064]), .B(p_input[464]), .Z(n20378) );
  XOR U20259 ( .A(n20369), .B(n20377), .Z(n20408) );
  XOR U20260 ( .A(n20409), .B(n20374), .Z(n20377) );
  XOR U20261 ( .A(p_input[2062]), .B(p_input[462]), .Z(n20374) );
  XNOR U20262 ( .A(p_input[2063]), .B(p_input[463]), .Z(n20409) );
  XNOR U20263 ( .A(n16740), .B(p_input[458]), .Z(n20369) );
  XNOR U20264 ( .A(n20384), .B(n20383), .Z(n20367) );
  XNOR U20265 ( .A(n20410), .B(n20389), .Z(n20383) );
  XOR U20266 ( .A(p_input[2057]), .B(p_input[457]), .Z(n20389) );
  XOR U20267 ( .A(n20380), .B(n20388), .Z(n20410) );
  XOR U20268 ( .A(n20411), .B(n20385), .Z(n20388) );
  XOR U20269 ( .A(p_input[2055]), .B(p_input[455]), .Z(n20385) );
  XNOR U20270 ( .A(p_input[2056]), .B(p_input[456]), .Z(n20411) );
  XNOR U20271 ( .A(n16459), .B(p_input[451]), .Z(n20380) );
  XNOR U20272 ( .A(n20394), .B(n20393), .Z(n20384) );
  XOR U20273 ( .A(n20412), .B(n20390), .Z(n20393) );
  XOR U20274 ( .A(p_input[2052]), .B(p_input[452]), .Z(n20390) );
  XNOR U20275 ( .A(p_input[2053]), .B(p_input[453]), .Z(n20412) );
  XOR U20276 ( .A(p_input[2054]), .B(p_input[454]), .Z(n20394) );
  XNOR U20277 ( .A(n20413), .B(n20414), .Z(n20211) );
  AND U20278 ( .A(n221), .B(n20415), .Z(n20414) );
  XNOR U20279 ( .A(n20416), .B(n20417), .Z(n221) );
  AND U20280 ( .A(n20418), .B(n20419), .Z(n20417) );
  XOR U20281 ( .A(n20416), .B(n20221), .Z(n20419) );
  XNOR U20282 ( .A(n20416), .B(n20163), .Z(n20418) );
  XOR U20283 ( .A(n20420), .B(n20421), .Z(n20416) );
  AND U20284 ( .A(n20422), .B(n20423), .Z(n20421) );
  XNOR U20285 ( .A(n20234), .B(n20420), .Z(n20423) );
  XOR U20286 ( .A(n20420), .B(n20175), .Z(n20422) );
  XOR U20287 ( .A(n20424), .B(n20425), .Z(n20420) );
  AND U20288 ( .A(n20426), .B(n20427), .Z(n20425) );
  XNOR U20289 ( .A(n20259), .B(n20424), .Z(n20427) );
  XOR U20290 ( .A(n20424), .B(n20186), .Z(n20426) );
  XOR U20291 ( .A(n20428), .B(n20429), .Z(n20424) );
  AND U20292 ( .A(n20430), .B(n20431), .Z(n20429) );
  XOR U20293 ( .A(n20428), .B(n20196), .Z(n20430) );
  XOR U20294 ( .A(n20432), .B(n20433), .Z(n20152) );
  AND U20295 ( .A(n225), .B(n20415), .Z(n20433) );
  XNOR U20296 ( .A(n20413), .B(n20432), .Z(n20415) );
  XNOR U20297 ( .A(n20434), .B(n20435), .Z(n225) );
  AND U20298 ( .A(n20436), .B(n20437), .Z(n20435) );
  XNOR U20299 ( .A(n20438), .B(n20434), .Z(n20437) );
  IV U20300 ( .A(n20221), .Z(n20438) );
  XNOR U20301 ( .A(n20439), .B(n20440), .Z(n20221) );
  AND U20302 ( .A(n228), .B(n20441), .Z(n20440) );
  XNOR U20303 ( .A(n20439), .B(n20442), .Z(n20441) );
  XNOR U20304 ( .A(n20163), .B(n20434), .Z(n20436) );
  XOR U20305 ( .A(n20443), .B(n20444), .Z(n20163) );
  AND U20306 ( .A(n236), .B(n20445), .Z(n20444) );
  XOR U20307 ( .A(n20446), .B(n20447), .Z(n20434) );
  AND U20308 ( .A(n20448), .B(n20449), .Z(n20447) );
  XNOR U20309 ( .A(n20446), .B(n20234), .Z(n20449) );
  XNOR U20310 ( .A(n20450), .B(n20451), .Z(n20234) );
  AND U20311 ( .A(n228), .B(n20452), .Z(n20451) );
  XOR U20312 ( .A(n20453), .B(n20450), .Z(n20452) );
  XNOR U20313 ( .A(n20454), .B(n20446), .Z(n20448) );
  IV U20314 ( .A(n20175), .Z(n20454) );
  XOR U20315 ( .A(n20455), .B(n20456), .Z(n20175) );
  AND U20316 ( .A(n236), .B(n20457), .Z(n20456) );
  XOR U20317 ( .A(n20458), .B(n20459), .Z(n20446) );
  AND U20318 ( .A(n20460), .B(n20461), .Z(n20459) );
  XNOR U20319 ( .A(n20458), .B(n20259), .Z(n20461) );
  XNOR U20320 ( .A(n20462), .B(n20463), .Z(n20259) );
  AND U20321 ( .A(n228), .B(n20464), .Z(n20463) );
  XNOR U20322 ( .A(n20465), .B(n20462), .Z(n20464) );
  XOR U20323 ( .A(n20186), .B(n20458), .Z(n20460) );
  XOR U20324 ( .A(n20466), .B(n20467), .Z(n20186) );
  AND U20325 ( .A(n236), .B(n20468), .Z(n20467) );
  XOR U20326 ( .A(n20428), .B(n20469), .Z(n20458) );
  AND U20327 ( .A(n20470), .B(n20431), .Z(n20469) );
  XNOR U20328 ( .A(n20305), .B(n20428), .Z(n20431) );
  XNOR U20329 ( .A(n20471), .B(n20472), .Z(n20305) );
  AND U20330 ( .A(n228), .B(n20473), .Z(n20472) );
  XOR U20331 ( .A(n20474), .B(n20471), .Z(n20473) );
  XNOR U20332 ( .A(n20475), .B(n20428), .Z(n20470) );
  IV U20333 ( .A(n20196), .Z(n20475) );
  XOR U20334 ( .A(n20476), .B(n20477), .Z(n20196) );
  AND U20335 ( .A(n236), .B(n20478), .Z(n20477) );
  XOR U20336 ( .A(n20479), .B(n20480), .Z(n20428) );
  AND U20337 ( .A(n20481), .B(n20482), .Z(n20480) );
  XNOR U20338 ( .A(n20479), .B(n20395), .Z(n20482) );
  XNOR U20339 ( .A(n20483), .B(n20484), .Z(n20395) );
  AND U20340 ( .A(n228), .B(n20485), .Z(n20484) );
  XNOR U20341 ( .A(n20486), .B(n20483), .Z(n20485) );
  XNOR U20342 ( .A(n20487), .B(n20479), .Z(n20481) );
  IV U20343 ( .A(n20208), .Z(n20487) );
  XOR U20344 ( .A(n20488), .B(n20489), .Z(n20208) );
  AND U20345 ( .A(n236), .B(n20490), .Z(n20489) );
  AND U20346 ( .A(n20432), .B(n20413), .Z(n20479) );
  XNOR U20347 ( .A(n20491), .B(n20492), .Z(n20413) );
  AND U20348 ( .A(n228), .B(n20493), .Z(n20492) );
  XNOR U20349 ( .A(n20494), .B(n20491), .Z(n20493) );
  XNOR U20350 ( .A(n20495), .B(n20496), .Z(n228) );
  AND U20351 ( .A(n20497), .B(n20498), .Z(n20496) );
  XOR U20352 ( .A(n20442), .B(n20495), .Z(n20498) );
  AND U20353 ( .A(n20499), .B(n20500), .Z(n20442) );
  XOR U20354 ( .A(n20495), .B(n20439), .Z(n20497) );
  XNOR U20355 ( .A(n20501), .B(n20502), .Z(n20439) );
  AND U20356 ( .A(n232), .B(n20445), .Z(n20502) );
  XOR U20357 ( .A(n20443), .B(n20501), .Z(n20445) );
  XOR U20358 ( .A(n20503), .B(n20504), .Z(n20495) );
  AND U20359 ( .A(n20505), .B(n20506), .Z(n20504) );
  XNOR U20360 ( .A(n20503), .B(n20499), .Z(n20506) );
  IV U20361 ( .A(n20453), .Z(n20499) );
  XOR U20362 ( .A(n20507), .B(n20508), .Z(n20453) );
  XOR U20363 ( .A(n20509), .B(n20500), .Z(n20508) );
  AND U20364 ( .A(n20465), .B(n20510), .Z(n20500) );
  AND U20365 ( .A(n20511), .B(n20512), .Z(n20509) );
  XOR U20366 ( .A(n20513), .B(n20507), .Z(n20511) );
  XNOR U20367 ( .A(n20450), .B(n20503), .Z(n20505) );
  XNOR U20368 ( .A(n20514), .B(n20515), .Z(n20450) );
  AND U20369 ( .A(n232), .B(n20457), .Z(n20515) );
  XOR U20370 ( .A(n20514), .B(n20455), .Z(n20457) );
  XOR U20371 ( .A(n20516), .B(n20517), .Z(n20503) );
  AND U20372 ( .A(n20518), .B(n20519), .Z(n20517) );
  XNOR U20373 ( .A(n20516), .B(n20465), .Z(n20519) );
  XOR U20374 ( .A(n20520), .B(n20512), .Z(n20465) );
  XNOR U20375 ( .A(n20521), .B(n20507), .Z(n20512) );
  XOR U20376 ( .A(n20522), .B(n20523), .Z(n20507) );
  AND U20377 ( .A(n20524), .B(n20525), .Z(n20523) );
  XOR U20378 ( .A(n20526), .B(n20522), .Z(n20524) );
  XNOR U20379 ( .A(n20527), .B(n20528), .Z(n20521) );
  AND U20380 ( .A(n20529), .B(n20530), .Z(n20528) );
  XOR U20381 ( .A(n20527), .B(n20531), .Z(n20529) );
  XNOR U20382 ( .A(n20513), .B(n20510), .Z(n20520) );
  AND U20383 ( .A(n20532), .B(n20533), .Z(n20510) );
  XOR U20384 ( .A(n20534), .B(n20535), .Z(n20513) );
  AND U20385 ( .A(n20536), .B(n20537), .Z(n20535) );
  XOR U20386 ( .A(n20534), .B(n20538), .Z(n20536) );
  XNOR U20387 ( .A(n20462), .B(n20516), .Z(n20518) );
  XNOR U20388 ( .A(n20539), .B(n20540), .Z(n20462) );
  AND U20389 ( .A(n232), .B(n20468), .Z(n20540) );
  XOR U20390 ( .A(n20539), .B(n20466), .Z(n20468) );
  XOR U20391 ( .A(n20541), .B(n20542), .Z(n20516) );
  AND U20392 ( .A(n20543), .B(n20544), .Z(n20542) );
  XNOR U20393 ( .A(n20541), .B(n20532), .Z(n20544) );
  IV U20394 ( .A(n20474), .Z(n20532) );
  XNOR U20395 ( .A(n20545), .B(n20525), .Z(n20474) );
  XNOR U20396 ( .A(n20546), .B(n20531), .Z(n20525) );
  XOR U20397 ( .A(n20547), .B(n20548), .Z(n20531) );
  AND U20398 ( .A(n20549), .B(n20550), .Z(n20548) );
  XOR U20399 ( .A(n20547), .B(n20551), .Z(n20549) );
  XNOR U20400 ( .A(n20530), .B(n20522), .Z(n20546) );
  XOR U20401 ( .A(n20552), .B(n20553), .Z(n20522) );
  AND U20402 ( .A(n20554), .B(n20555), .Z(n20553) );
  XNOR U20403 ( .A(n20556), .B(n20552), .Z(n20554) );
  XNOR U20404 ( .A(n20557), .B(n20527), .Z(n20530) );
  XOR U20405 ( .A(n20558), .B(n20559), .Z(n20527) );
  AND U20406 ( .A(n20560), .B(n20561), .Z(n20559) );
  XOR U20407 ( .A(n20558), .B(n20562), .Z(n20560) );
  XNOR U20408 ( .A(n20563), .B(n20564), .Z(n20557) );
  AND U20409 ( .A(n20565), .B(n20566), .Z(n20564) );
  XNOR U20410 ( .A(n20563), .B(n20567), .Z(n20565) );
  XNOR U20411 ( .A(n20526), .B(n20533), .Z(n20545) );
  AND U20412 ( .A(n20486), .B(n20568), .Z(n20533) );
  XOR U20413 ( .A(n20538), .B(n20537), .Z(n20526) );
  XNOR U20414 ( .A(n20569), .B(n20534), .Z(n20537) );
  XOR U20415 ( .A(n20570), .B(n20571), .Z(n20534) );
  AND U20416 ( .A(n20572), .B(n20573), .Z(n20571) );
  XOR U20417 ( .A(n20570), .B(n20574), .Z(n20572) );
  XNOR U20418 ( .A(n20575), .B(n20576), .Z(n20569) );
  AND U20419 ( .A(n20577), .B(n20578), .Z(n20576) );
  XOR U20420 ( .A(n20575), .B(n20579), .Z(n20577) );
  XOR U20421 ( .A(n20580), .B(n20581), .Z(n20538) );
  AND U20422 ( .A(n20582), .B(n20583), .Z(n20581) );
  XOR U20423 ( .A(n20580), .B(n20584), .Z(n20582) );
  XNOR U20424 ( .A(n20471), .B(n20541), .Z(n20543) );
  XNOR U20425 ( .A(n20585), .B(n20586), .Z(n20471) );
  AND U20426 ( .A(n232), .B(n20478), .Z(n20586) );
  XOR U20427 ( .A(n20585), .B(n20476), .Z(n20478) );
  XOR U20428 ( .A(n20587), .B(n20588), .Z(n20541) );
  AND U20429 ( .A(n20589), .B(n20590), .Z(n20588) );
  XNOR U20430 ( .A(n20587), .B(n20486), .Z(n20590) );
  XOR U20431 ( .A(n20591), .B(n20555), .Z(n20486) );
  XNOR U20432 ( .A(n20592), .B(n20562), .Z(n20555) );
  XOR U20433 ( .A(n20551), .B(n20550), .Z(n20562) );
  XNOR U20434 ( .A(n20593), .B(n20547), .Z(n20550) );
  XOR U20435 ( .A(n20594), .B(n20595), .Z(n20547) );
  AND U20436 ( .A(n20596), .B(n20597), .Z(n20595) );
  XOR U20437 ( .A(n20594), .B(n20598), .Z(n20596) );
  XNOR U20438 ( .A(n20599), .B(n20600), .Z(n20593) );
  NOR U20439 ( .A(n20601), .B(n20602), .Z(n20600) );
  XNOR U20440 ( .A(n20599), .B(n20603), .Z(n20601) );
  XOR U20441 ( .A(n20604), .B(n20605), .Z(n20551) );
  NOR U20442 ( .A(n20606), .B(n20607), .Z(n20605) );
  XNOR U20443 ( .A(n20604), .B(n20608), .Z(n20606) );
  XNOR U20444 ( .A(n20561), .B(n20552), .Z(n20592) );
  XOR U20445 ( .A(n20609), .B(n20610), .Z(n20552) );
  NOR U20446 ( .A(n20611), .B(n20612), .Z(n20610) );
  XNOR U20447 ( .A(n20609), .B(n20613), .Z(n20611) );
  XOR U20448 ( .A(n20614), .B(n20567), .Z(n20561) );
  XNOR U20449 ( .A(n20615), .B(n20616), .Z(n20567) );
  NOR U20450 ( .A(n20617), .B(n20618), .Z(n20616) );
  XNOR U20451 ( .A(n20615), .B(n20619), .Z(n20617) );
  XNOR U20452 ( .A(n20566), .B(n20558), .Z(n20614) );
  XOR U20453 ( .A(n20620), .B(n20621), .Z(n20558) );
  AND U20454 ( .A(n20622), .B(n20623), .Z(n20621) );
  XOR U20455 ( .A(n20620), .B(n20624), .Z(n20622) );
  XNOR U20456 ( .A(n20625), .B(n20563), .Z(n20566) );
  XOR U20457 ( .A(n20626), .B(n20627), .Z(n20563) );
  AND U20458 ( .A(n20628), .B(n20629), .Z(n20627) );
  XOR U20459 ( .A(n20626), .B(n20630), .Z(n20628) );
  XNOR U20460 ( .A(n20631), .B(n20632), .Z(n20625) );
  NOR U20461 ( .A(n20633), .B(n20634), .Z(n20632) );
  XOR U20462 ( .A(n20631), .B(n20635), .Z(n20633) );
  XOR U20463 ( .A(n20556), .B(n20568), .Z(n20591) );
  NOR U20464 ( .A(n20494), .B(n20636), .Z(n20568) );
  XNOR U20465 ( .A(n20574), .B(n20573), .Z(n20556) );
  XNOR U20466 ( .A(n20637), .B(n20579), .Z(n20573) );
  XOR U20467 ( .A(n20638), .B(n20639), .Z(n20579) );
  NOR U20468 ( .A(n20640), .B(n20641), .Z(n20639) );
  XNOR U20469 ( .A(n20638), .B(n20642), .Z(n20640) );
  XNOR U20470 ( .A(n20578), .B(n20570), .Z(n20637) );
  XOR U20471 ( .A(n20643), .B(n20644), .Z(n20570) );
  AND U20472 ( .A(n20645), .B(n20646), .Z(n20644) );
  XNOR U20473 ( .A(n20643), .B(n20647), .Z(n20645) );
  XNOR U20474 ( .A(n20648), .B(n20575), .Z(n20578) );
  XOR U20475 ( .A(n20649), .B(n20650), .Z(n20575) );
  AND U20476 ( .A(n20651), .B(n20652), .Z(n20650) );
  XOR U20477 ( .A(n20649), .B(n20653), .Z(n20651) );
  XNOR U20478 ( .A(n20654), .B(n20655), .Z(n20648) );
  NOR U20479 ( .A(n20656), .B(n20657), .Z(n20655) );
  XOR U20480 ( .A(n20654), .B(n20658), .Z(n20656) );
  XOR U20481 ( .A(n20584), .B(n20583), .Z(n20574) );
  XNOR U20482 ( .A(n20659), .B(n20580), .Z(n20583) );
  XOR U20483 ( .A(n20660), .B(n20661), .Z(n20580) );
  AND U20484 ( .A(n20662), .B(n20663), .Z(n20661) );
  XOR U20485 ( .A(n20660), .B(n20664), .Z(n20662) );
  XNOR U20486 ( .A(n20665), .B(n20666), .Z(n20659) );
  NOR U20487 ( .A(n20667), .B(n20668), .Z(n20666) );
  XNOR U20488 ( .A(n20665), .B(n20669), .Z(n20667) );
  XOR U20489 ( .A(n20670), .B(n20671), .Z(n20584) );
  NOR U20490 ( .A(n20672), .B(n20673), .Z(n20671) );
  XNOR U20491 ( .A(n20670), .B(n20674), .Z(n20672) );
  XNOR U20492 ( .A(n20483), .B(n20587), .Z(n20589) );
  XNOR U20493 ( .A(n20675), .B(n20676), .Z(n20483) );
  AND U20494 ( .A(n232), .B(n20490), .Z(n20676) );
  XOR U20495 ( .A(n20675), .B(n20488), .Z(n20490) );
  AND U20496 ( .A(n20491), .B(n20494), .Z(n20587) );
  XOR U20497 ( .A(n20677), .B(n20636), .Z(n20494) );
  XNOR U20498 ( .A(p_input[2048]), .B(p_input[480]), .Z(n20636) );
  XOR U20499 ( .A(n20613), .B(n20612), .Z(n20677) );
  XOR U20500 ( .A(n20678), .B(n20624), .Z(n20612) );
  XOR U20501 ( .A(n20598), .B(n20597), .Z(n20624) );
  XNOR U20502 ( .A(n20679), .B(n20603), .Z(n20597) );
  XOR U20503 ( .A(p_input[2072]), .B(p_input[504]), .Z(n20603) );
  XOR U20504 ( .A(n20594), .B(n20602), .Z(n20679) );
  XOR U20505 ( .A(n20680), .B(n20599), .Z(n20602) );
  XOR U20506 ( .A(p_input[2070]), .B(p_input[502]), .Z(n20599) );
  XNOR U20507 ( .A(p_input[2071]), .B(p_input[503]), .Z(n20680) );
  XNOR U20508 ( .A(n16727), .B(p_input[498]), .Z(n20594) );
  XNOR U20509 ( .A(n20608), .B(n20607), .Z(n20598) );
  XOR U20510 ( .A(n20681), .B(n20604), .Z(n20607) );
  XOR U20511 ( .A(p_input[2067]), .B(p_input[499]), .Z(n20604) );
  XNOR U20512 ( .A(p_input[2068]), .B(p_input[500]), .Z(n20681) );
  XOR U20513 ( .A(p_input[2069]), .B(p_input[501]), .Z(n20608) );
  XNOR U20514 ( .A(n20623), .B(n20609), .Z(n20678) );
  XNOR U20515 ( .A(n16729), .B(p_input[481]), .Z(n20609) );
  XNOR U20516 ( .A(n20682), .B(n20630), .Z(n20623) );
  XNOR U20517 ( .A(n20619), .B(n20618), .Z(n20630) );
  XOR U20518 ( .A(n20683), .B(n20615), .Z(n20618) );
  XNOR U20519 ( .A(n16444), .B(p_input[506]), .Z(n20615) );
  XNOR U20520 ( .A(p_input[2075]), .B(p_input[507]), .Z(n20683) );
  XOR U20521 ( .A(p_input[2076]), .B(p_input[508]), .Z(n20619) );
  XNOR U20522 ( .A(n20629), .B(n20620), .Z(n20682) );
  XNOR U20523 ( .A(n16732), .B(p_input[497]), .Z(n20620) );
  XOR U20524 ( .A(n20684), .B(n20635), .Z(n20629) );
  XNOR U20525 ( .A(p_input[2079]), .B(p_input[511]), .Z(n20635) );
  XOR U20526 ( .A(n20626), .B(n20634), .Z(n20684) );
  XOR U20527 ( .A(n20685), .B(n20631), .Z(n20634) );
  XOR U20528 ( .A(p_input[2077]), .B(p_input[509]), .Z(n20631) );
  XNOR U20529 ( .A(p_input[2078]), .B(p_input[510]), .Z(n20685) );
  XNOR U20530 ( .A(n16448), .B(p_input[505]), .Z(n20626) );
  XNOR U20531 ( .A(n20647), .B(n20646), .Z(n20613) );
  XNOR U20532 ( .A(n20686), .B(n20653), .Z(n20646) );
  XNOR U20533 ( .A(n20642), .B(n20641), .Z(n20653) );
  XOR U20534 ( .A(n20687), .B(n20638), .Z(n20641) );
  XNOR U20535 ( .A(n16737), .B(p_input[491]), .Z(n20638) );
  XNOR U20536 ( .A(p_input[2060]), .B(p_input[492]), .Z(n20687) );
  XOR U20537 ( .A(p_input[2061]), .B(p_input[493]), .Z(n20642) );
  XNOR U20538 ( .A(n20652), .B(n20643), .Z(n20686) );
  XNOR U20539 ( .A(n16452), .B(p_input[482]), .Z(n20643) );
  XOR U20540 ( .A(n20688), .B(n20658), .Z(n20652) );
  XNOR U20541 ( .A(p_input[2064]), .B(p_input[496]), .Z(n20658) );
  XOR U20542 ( .A(n20649), .B(n20657), .Z(n20688) );
  XOR U20543 ( .A(n20689), .B(n20654), .Z(n20657) );
  XOR U20544 ( .A(p_input[2062]), .B(p_input[494]), .Z(n20654) );
  XNOR U20545 ( .A(p_input[2063]), .B(p_input[495]), .Z(n20689) );
  XNOR U20546 ( .A(n16740), .B(p_input[490]), .Z(n20649) );
  XNOR U20547 ( .A(n20664), .B(n20663), .Z(n20647) );
  XNOR U20548 ( .A(n20690), .B(n20669), .Z(n20663) );
  XOR U20549 ( .A(p_input[2057]), .B(p_input[489]), .Z(n20669) );
  XOR U20550 ( .A(n20660), .B(n20668), .Z(n20690) );
  XOR U20551 ( .A(n20691), .B(n20665), .Z(n20668) );
  XOR U20552 ( .A(p_input[2055]), .B(p_input[487]), .Z(n20665) );
  XNOR U20553 ( .A(p_input[2056]), .B(p_input[488]), .Z(n20691) );
  XNOR U20554 ( .A(n16459), .B(p_input[483]), .Z(n20660) );
  XNOR U20555 ( .A(n20674), .B(n20673), .Z(n20664) );
  XOR U20556 ( .A(n20692), .B(n20670), .Z(n20673) );
  XOR U20557 ( .A(p_input[2052]), .B(p_input[484]), .Z(n20670) );
  XNOR U20558 ( .A(p_input[2053]), .B(p_input[485]), .Z(n20692) );
  XOR U20559 ( .A(p_input[2054]), .B(p_input[486]), .Z(n20674) );
  XNOR U20560 ( .A(n20693), .B(n20694), .Z(n20491) );
  AND U20561 ( .A(n232), .B(n20695), .Z(n20694) );
  XNOR U20562 ( .A(n20696), .B(n20697), .Z(n232) );
  AND U20563 ( .A(n20698), .B(n20699), .Z(n20697) );
  XOR U20564 ( .A(n20696), .B(n20501), .Z(n20699) );
  XNOR U20565 ( .A(n20696), .B(n20443), .Z(n20698) );
  XOR U20566 ( .A(n20700), .B(n20701), .Z(n20696) );
  AND U20567 ( .A(n20702), .B(n20703), .Z(n20701) );
  XNOR U20568 ( .A(n20514), .B(n20700), .Z(n20703) );
  XOR U20569 ( .A(n20700), .B(n20455), .Z(n20702) );
  XOR U20570 ( .A(n20704), .B(n20705), .Z(n20700) );
  AND U20571 ( .A(n20706), .B(n20707), .Z(n20705) );
  XNOR U20572 ( .A(n20539), .B(n20704), .Z(n20707) );
  XOR U20573 ( .A(n20704), .B(n20466), .Z(n20706) );
  XOR U20574 ( .A(n20708), .B(n20709), .Z(n20704) );
  AND U20575 ( .A(n20710), .B(n20711), .Z(n20709) );
  XOR U20576 ( .A(n20708), .B(n20476), .Z(n20710) );
  XOR U20577 ( .A(n20712), .B(n20713), .Z(n20432) );
  AND U20578 ( .A(n236), .B(n20695), .Z(n20713) );
  XNOR U20579 ( .A(n20693), .B(n20712), .Z(n20695) );
  XNOR U20580 ( .A(n20714), .B(n20715), .Z(n236) );
  AND U20581 ( .A(n20716), .B(n20717), .Z(n20715) );
  XNOR U20582 ( .A(n20718), .B(n20714), .Z(n20717) );
  IV U20583 ( .A(n20501), .Z(n20718) );
  XNOR U20584 ( .A(n20719), .B(n20720), .Z(n20501) );
  AND U20585 ( .A(n239), .B(n20721), .Z(n20720) );
  XNOR U20586 ( .A(n20719), .B(n20722), .Z(n20721) );
  XNOR U20587 ( .A(n20443), .B(n20714), .Z(n20716) );
  XOR U20588 ( .A(n20723), .B(n20724), .Z(n20443) );
  AND U20589 ( .A(n247), .B(n20725), .Z(n20724) );
  XOR U20590 ( .A(n20726), .B(n20727), .Z(n20714) );
  AND U20591 ( .A(n20728), .B(n20729), .Z(n20727) );
  XNOR U20592 ( .A(n20726), .B(n20514), .Z(n20729) );
  XNOR U20593 ( .A(n20730), .B(n20731), .Z(n20514) );
  AND U20594 ( .A(n239), .B(n20732), .Z(n20731) );
  XOR U20595 ( .A(n20733), .B(n20730), .Z(n20732) );
  XNOR U20596 ( .A(n20734), .B(n20726), .Z(n20728) );
  IV U20597 ( .A(n20455), .Z(n20734) );
  XOR U20598 ( .A(n20735), .B(n20736), .Z(n20455) );
  AND U20599 ( .A(n247), .B(n20737), .Z(n20736) );
  XOR U20600 ( .A(n20738), .B(n20739), .Z(n20726) );
  AND U20601 ( .A(n20740), .B(n20741), .Z(n20739) );
  XNOR U20602 ( .A(n20738), .B(n20539), .Z(n20741) );
  XNOR U20603 ( .A(n20742), .B(n20743), .Z(n20539) );
  AND U20604 ( .A(n239), .B(n20744), .Z(n20743) );
  XNOR U20605 ( .A(n20745), .B(n20742), .Z(n20744) );
  XOR U20606 ( .A(n20466), .B(n20738), .Z(n20740) );
  XOR U20607 ( .A(n20746), .B(n20747), .Z(n20466) );
  AND U20608 ( .A(n247), .B(n20748), .Z(n20747) );
  XOR U20609 ( .A(n20708), .B(n20749), .Z(n20738) );
  AND U20610 ( .A(n20750), .B(n20711), .Z(n20749) );
  XNOR U20611 ( .A(n20585), .B(n20708), .Z(n20711) );
  XNOR U20612 ( .A(n20751), .B(n20752), .Z(n20585) );
  AND U20613 ( .A(n239), .B(n20753), .Z(n20752) );
  XOR U20614 ( .A(n20754), .B(n20751), .Z(n20753) );
  XNOR U20615 ( .A(n20755), .B(n20708), .Z(n20750) );
  IV U20616 ( .A(n20476), .Z(n20755) );
  XOR U20617 ( .A(n20756), .B(n20757), .Z(n20476) );
  AND U20618 ( .A(n247), .B(n20758), .Z(n20757) );
  XOR U20619 ( .A(n20759), .B(n20760), .Z(n20708) );
  AND U20620 ( .A(n20761), .B(n20762), .Z(n20760) );
  XNOR U20621 ( .A(n20759), .B(n20675), .Z(n20762) );
  XNOR U20622 ( .A(n20763), .B(n20764), .Z(n20675) );
  AND U20623 ( .A(n239), .B(n20765), .Z(n20764) );
  XNOR U20624 ( .A(n20766), .B(n20763), .Z(n20765) );
  XNOR U20625 ( .A(n20767), .B(n20759), .Z(n20761) );
  IV U20626 ( .A(n20488), .Z(n20767) );
  XOR U20627 ( .A(n20768), .B(n20769), .Z(n20488) );
  AND U20628 ( .A(n247), .B(n20770), .Z(n20769) );
  AND U20629 ( .A(n20712), .B(n20693), .Z(n20759) );
  XNOR U20630 ( .A(n20771), .B(n20772), .Z(n20693) );
  AND U20631 ( .A(n239), .B(n20773), .Z(n20772) );
  XNOR U20632 ( .A(n20774), .B(n20771), .Z(n20773) );
  XNOR U20633 ( .A(n20775), .B(n20776), .Z(n239) );
  AND U20634 ( .A(n20777), .B(n20778), .Z(n20776) );
  XOR U20635 ( .A(n20722), .B(n20775), .Z(n20778) );
  AND U20636 ( .A(n20779), .B(n20780), .Z(n20722) );
  XOR U20637 ( .A(n20775), .B(n20719), .Z(n20777) );
  XNOR U20638 ( .A(n20781), .B(n20782), .Z(n20719) );
  AND U20639 ( .A(n243), .B(n20725), .Z(n20782) );
  XOR U20640 ( .A(n20723), .B(n20781), .Z(n20725) );
  XOR U20641 ( .A(n20783), .B(n20784), .Z(n20775) );
  AND U20642 ( .A(n20785), .B(n20786), .Z(n20784) );
  XNOR U20643 ( .A(n20783), .B(n20779), .Z(n20786) );
  IV U20644 ( .A(n20733), .Z(n20779) );
  XOR U20645 ( .A(n20787), .B(n20788), .Z(n20733) );
  XOR U20646 ( .A(n20789), .B(n20780), .Z(n20788) );
  AND U20647 ( .A(n20745), .B(n20790), .Z(n20780) );
  AND U20648 ( .A(n20791), .B(n20792), .Z(n20789) );
  XOR U20649 ( .A(n20793), .B(n20787), .Z(n20791) );
  XNOR U20650 ( .A(n20730), .B(n20783), .Z(n20785) );
  XNOR U20651 ( .A(n20794), .B(n20795), .Z(n20730) );
  AND U20652 ( .A(n243), .B(n20737), .Z(n20795) );
  XOR U20653 ( .A(n20794), .B(n20735), .Z(n20737) );
  XOR U20654 ( .A(n20796), .B(n20797), .Z(n20783) );
  AND U20655 ( .A(n20798), .B(n20799), .Z(n20797) );
  XNOR U20656 ( .A(n20796), .B(n20745), .Z(n20799) );
  XOR U20657 ( .A(n20800), .B(n20792), .Z(n20745) );
  XNOR U20658 ( .A(n20801), .B(n20787), .Z(n20792) );
  XOR U20659 ( .A(n20802), .B(n20803), .Z(n20787) );
  AND U20660 ( .A(n20804), .B(n20805), .Z(n20803) );
  XOR U20661 ( .A(n20806), .B(n20802), .Z(n20804) );
  XNOR U20662 ( .A(n20807), .B(n20808), .Z(n20801) );
  AND U20663 ( .A(n20809), .B(n20810), .Z(n20808) );
  XOR U20664 ( .A(n20807), .B(n20811), .Z(n20809) );
  XNOR U20665 ( .A(n20793), .B(n20790), .Z(n20800) );
  AND U20666 ( .A(n20812), .B(n20813), .Z(n20790) );
  XOR U20667 ( .A(n20814), .B(n20815), .Z(n20793) );
  AND U20668 ( .A(n20816), .B(n20817), .Z(n20815) );
  XOR U20669 ( .A(n20814), .B(n20818), .Z(n20816) );
  XNOR U20670 ( .A(n20742), .B(n20796), .Z(n20798) );
  XNOR U20671 ( .A(n20819), .B(n20820), .Z(n20742) );
  AND U20672 ( .A(n243), .B(n20748), .Z(n20820) );
  XOR U20673 ( .A(n20819), .B(n20746), .Z(n20748) );
  XOR U20674 ( .A(n20821), .B(n20822), .Z(n20796) );
  AND U20675 ( .A(n20823), .B(n20824), .Z(n20822) );
  XNOR U20676 ( .A(n20821), .B(n20812), .Z(n20824) );
  IV U20677 ( .A(n20754), .Z(n20812) );
  XNOR U20678 ( .A(n20825), .B(n20805), .Z(n20754) );
  XNOR U20679 ( .A(n20826), .B(n20811), .Z(n20805) );
  XOR U20680 ( .A(n20827), .B(n20828), .Z(n20811) );
  AND U20681 ( .A(n20829), .B(n20830), .Z(n20828) );
  XOR U20682 ( .A(n20827), .B(n20831), .Z(n20829) );
  XNOR U20683 ( .A(n20810), .B(n20802), .Z(n20826) );
  XOR U20684 ( .A(n20832), .B(n20833), .Z(n20802) );
  AND U20685 ( .A(n20834), .B(n20835), .Z(n20833) );
  XNOR U20686 ( .A(n20836), .B(n20832), .Z(n20834) );
  XNOR U20687 ( .A(n20837), .B(n20807), .Z(n20810) );
  XOR U20688 ( .A(n20838), .B(n20839), .Z(n20807) );
  AND U20689 ( .A(n20840), .B(n20841), .Z(n20839) );
  XOR U20690 ( .A(n20838), .B(n20842), .Z(n20840) );
  XNOR U20691 ( .A(n20843), .B(n20844), .Z(n20837) );
  AND U20692 ( .A(n20845), .B(n20846), .Z(n20844) );
  XNOR U20693 ( .A(n20843), .B(n20847), .Z(n20845) );
  XNOR U20694 ( .A(n20806), .B(n20813), .Z(n20825) );
  AND U20695 ( .A(n20766), .B(n20848), .Z(n20813) );
  XOR U20696 ( .A(n20818), .B(n20817), .Z(n20806) );
  XNOR U20697 ( .A(n20849), .B(n20814), .Z(n20817) );
  XOR U20698 ( .A(n20850), .B(n20851), .Z(n20814) );
  AND U20699 ( .A(n20852), .B(n20853), .Z(n20851) );
  XOR U20700 ( .A(n20850), .B(n20854), .Z(n20852) );
  XNOR U20701 ( .A(n20855), .B(n20856), .Z(n20849) );
  AND U20702 ( .A(n20857), .B(n20858), .Z(n20856) );
  XOR U20703 ( .A(n20855), .B(n20859), .Z(n20857) );
  XOR U20704 ( .A(n20860), .B(n20861), .Z(n20818) );
  AND U20705 ( .A(n20862), .B(n20863), .Z(n20861) );
  XOR U20706 ( .A(n20860), .B(n20864), .Z(n20862) );
  XNOR U20707 ( .A(n20751), .B(n20821), .Z(n20823) );
  XNOR U20708 ( .A(n20865), .B(n20866), .Z(n20751) );
  AND U20709 ( .A(n243), .B(n20758), .Z(n20866) );
  XOR U20710 ( .A(n20865), .B(n20756), .Z(n20758) );
  XOR U20711 ( .A(n20867), .B(n20868), .Z(n20821) );
  AND U20712 ( .A(n20869), .B(n20870), .Z(n20868) );
  XNOR U20713 ( .A(n20867), .B(n20766), .Z(n20870) );
  XOR U20714 ( .A(n20871), .B(n20835), .Z(n20766) );
  XNOR U20715 ( .A(n20872), .B(n20842), .Z(n20835) );
  XOR U20716 ( .A(n20831), .B(n20830), .Z(n20842) );
  XNOR U20717 ( .A(n20873), .B(n20827), .Z(n20830) );
  XOR U20718 ( .A(n20874), .B(n20875), .Z(n20827) );
  AND U20719 ( .A(n20876), .B(n20877), .Z(n20875) );
  XOR U20720 ( .A(n20874), .B(n20878), .Z(n20876) );
  XNOR U20721 ( .A(n20879), .B(n20880), .Z(n20873) );
  NOR U20722 ( .A(n20881), .B(n20882), .Z(n20880) );
  XNOR U20723 ( .A(n20879), .B(n20883), .Z(n20881) );
  XOR U20724 ( .A(n20884), .B(n20885), .Z(n20831) );
  NOR U20725 ( .A(n20886), .B(n20887), .Z(n20885) );
  XNOR U20726 ( .A(n20884), .B(n20888), .Z(n20886) );
  XNOR U20727 ( .A(n20841), .B(n20832), .Z(n20872) );
  XOR U20728 ( .A(n20889), .B(n20890), .Z(n20832) );
  NOR U20729 ( .A(n20891), .B(n20892), .Z(n20890) );
  XNOR U20730 ( .A(n20889), .B(n20893), .Z(n20891) );
  XOR U20731 ( .A(n20894), .B(n20847), .Z(n20841) );
  XNOR U20732 ( .A(n20895), .B(n20896), .Z(n20847) );
  NOR U20733 ( .A(n20897), .B(n20898), .Z(n20896) );
  XNOR U20734 ( .A(n20895), .B(n20899), .Z(n20897) );
  XNOR U20735 ( .A(n20846), .B(n20838), .Z(n20894) );
  XOR U20736 ( .A(n20900), .B(n20901), .Z(n20838) );
  AND U20737 ( .A(n20902), .B(n20903), .Z(n20901) );
  XOR U20738 ( .A(n20900), .B(n20904), .Z(n20902) );
  XNOR U20739 ( .A(n20905), .B(n20843), .Z(n20846) );
  XOR U20740 ( .A(n20906), .B(n20907), .Z(n20843) );
  AND U20741 ( .A(n20908), .B(n20909), .Z(n20907) );
  XOR U20742 ( .A(n20906), .B(n20910), .Z(n20908) );
  XNOR U20743 ( .A(n20911), .B(n20912), .Z(n20905) );
  NOR U20744 ( .A(n20913), .B(n20914), .Z(n20912) );
  XOR U20745 ( .A(n20911), .B(n20915), .Z(n20913) );
  XOR U20746 ( .A(n20836), .B(n20848), .Z(n20871) );
  NOR U20747 ( .A(n20774), .B(n20916), .Z(n20848) );
  XNOR U20748 ( .A(n20854), .B(n20853), .Z(n20836) );
  XNOR U20749 ( .A(n20917), .B(n20859), .Z(n20853) );
  XOR U20750 ( .A(n20918), .B(n20919), .Z(n20859) );
  NOR U20751 ( .A(n20920), .B(n20921), .Z(n20919) );
  XNOR U20752 ( .A(n20918), .B(n20922), .Z(n20920) );
  XNOR U20753 ( .A(n20858), .B(n20850), .Z(n20917) );
  XOR U20754 ( .A(n20923), .B(n20924), .Z(n20850) );
  AND U20755 ( .A(n20925), .B(n20926), .Z(n20924) );
  XNOR U20756 ( .A(n20923), .B(n20927), .Z(n20925) );
  XNOR U20757 ( .A(n20928), .B(n20855), .Z(n20858) );
  XOR U20758 ( .A(n20929), .B(n20930), .Z(n20855) );
  AND U20759 ( .A(n20931), .B(n20932), .Z(n20930) );
  XOR U20760 ( .A(n20929), .B(n20933), .Z(n20931) );
  XNOR U20761 ( .A(n20934), .B(n20935), .Z(n20928) );
  NOR U20762 ( .A(n20936), .B(n20937), .Z(n20935) );
  XOR U20763 ( .A(n20934), .B(n20938), .Z(n20936) );
  XOR U20764 ( .A(n20864), .B(n20863), .Z(n20854) );
  XNOR U20765 ( .A(n20939), .B(n20860), .Z(n20863) );
  XOR U20766 ( .A(n20940), .B(n20941), .Z(n20860) );
  AND U20767 ( .A(n20942), .B(n20943), .Z(n20941) );
  XOR U20768 ( .A(n20940), .B(n20944), .Z(n20942) );
  XNOR U20769 ( .A(n20945), .B(n20946), .Z(n20939) );
  NOR U20770 ( .A(n20947), .B(n20948), .Z(n20946) );
  XNOR U20771 ( .A(n20945), .B(n20949), .Z(n20947) );
  XOR U20772 ( .A(n20950), .B(n20951), .Z(n20864) );
  NOR U20773 ( .A(n20952), .B(n20953), .Z(n20951) );
  XNOR U20774 ( .A(n20950), .B(n20954), .Z(n20952) );
  XNOR U20775 ( .A(n20763), .B(n20867), .Z(n20869) );
  XNOR U20776 ( .A(n20955), .B(n20956), .Z(n20763) );
  AND U20777 ( .A(n243), .B(n20770), .Z(n20956) );
  XOR U20778 ( .A(n20955), .B(n20768), .Z(n20770) );
  AND U20779 ( .A(n20771), .B(n20774), .Z(n20867) );
  XOR U20780 ( .A(n20957), .B(n20916), .Z(n20774) );
  XNOR U20781 ( .A(p_input[2048]), .B(p_input[512]), .Z(n20916) );
  XOR U20782 ( .A(n20893), .B(n20892), .Z(n20957) );
  XOR U20783 ( .A(n20958), .B(n20904), .Z(n20892) );
  XOR U20784 ( .A(n20878), .B(n20877), .Z(n20904) );
  XNOR U20785 ( .A(n20959), .B(n20883), .Z(n20877) );
  XOR U20786 ( .A(p_input[2072]), .B(p_input[536]), .Z(n20883) );
  XOR U20787 ( .A(n20874), .B(n20882), .Z(n20959) );
  XOR U20788 ( .A(n20960), .B(n20879), .Z(n20882) );
  XOR U20789 ( .A(p_input[2070]), .B(p_input[534]), .Z(n20879) );
  XNOR U20790 ( .A(p_input[2071]), .B(p_input[535]), .Z(n20960) );
  XNOR U20791 ( .A(n16727), .B(p_input[530]), .Z(n20874) );
  XNOR U20792 ( .A(n20888), .B(n20887), .Z(n20878) );
  XOR U20793 ( .A(n20961), .B(n20884), .Z(n20887) );
  XOR U20794 ( .A(p_input[2067]), .B(p_input[531]), .Z(n20884) );
  XNOR U20795 ( .A(p_input[2068]), .B(p_input[532]), .Z(n20961) );
  XOR U20796 ( .A(p_input[2069]), .B(p_input[533]), .Z(n20888) );
  XNOR U20797 ( .A(n20903), .B(n20889), .Z(n20958) );
  XNOR U20798 ( .A(n16729), .B(p_input[513]), .Z(n20889) );
  XNOR U20799 ( .A(n20962), .B(n20910), .Z(n20903) );
  XNOR U20800 ( .A(n20899), .B(n20898), .Z(n20910) );
  XOR U20801 ( .A(n20963), .B(n20895), .Z(n20898) );
  XNOR U20802 ( .A(n16444), .B(p_input[538]), .Z(n20895) );
  XNOR U20803 ( .A(p_input[2075]), .B(p_input[539]), .Z(n20963) );
  XOR U20804 ( .A(p_input[2076]), .B(p_input[540]), .Z(n20899) );
  XNOR U20805 ( .A(n20909), .B(n20900), .Z(n20962) );
  XNOR U20806 ( .A(n16732), .B(p_input[529]), .Z(n20900) );
  XOR U20807 ( .A(n20964), .B(n20915), .Z(n20909) );
  XNOR U20808 ( .A(p_input[2079]), .B(p_input[543]), .Z(n20915) );
  XOR U20809 ( .A(n20906), .B(n20914), .Z(n20964) );
  XOR U20810 ( .A(n20965), .B(n20911), .Z(n20914) );
  XOR U20811 ( .A(p_input[2077]), .B(p_input[541]), .Z(n20911) );
  XNOR U20812 ( .A(p_input[2078]), .B(p_input[542]), .Z(n20965) );
  XNOR U20813 ( .A(n16448), .B(p_input[537]), .Z(n20906) );
  XNOR U20814 ( .A(n20927), .B(n20926), .Z(n20893) );
  XNOR U20815 ( .A(n20966), .B(n20933), .Z(n20926) );
  XNOR U20816 ( .A(n20922), .B(n20921), .Z(n20933) );
  XOR U20817 ( .A(n20967), .B(n20918), .Z(n20921) );
  XNOR U20818 ( .A(n16737), .B(p_input[523]), .Z(n20918) );
  XNOR U20819 ( .A(p_input[2060]), .B(p_input[524]), .Z(n20967) );
  XOR U20820 ( .A(p_input[2061]), .B(p_input[525]), .Z(n20922) );
  XNOR U20821 ( .A(n20932), .B(n20923), .Z(n20966) );
  XNOR U20822 ( .A(n16452), .B(p_input[514]), .Z(n20923) );
  XOR U20823 ( .A(n20968), .B(n20938), .Z(n20932) );
  XNOR U20824 ( .A(p_input[2064]), .B(p_input[528]), .Z(n20938) );
  XOR U20825 ( .A(n20929), .B(n20937), .Z(n20968) );
  XOR U20826 ( .A(n20969), .B(n20934), .Z(n20937) );
  XOR U20827 ( .A(p_input[2062]), .B(p_input[526]), .Z(n20934) );
  XNOR U20828 ( .A(p_input[2063]), .B(p_input[527]), .Z(n20969) );
  XNOR U20829 ( .A(n16740), .B(p_input[522]), .Z(n20929) );
  XNOR U20830 ( .A(n20944), .B(n20943), .Z(n20927) );
  XNOR U20831 ( .A(n20970), .B(n20949), .Z(n20943) );
  XOR U20832 ( .A(p_input[2057]), .B(p_input[521]), .Z(n20949) );
  XOR U20833 ( .A(n20940), .B(n20948), .Z(n20970) );
  XOR U20834 ( .A(n20971), .B(n20945), .Z(n20948) );
  XOR U20835 ( .A(p_input[2055]), .B(p_input[519]), .Z(n20945) );
  XNOR U20836 ( .A(p_input[2056]), .B(p_input[520]), .Z(n20971) );
  XNOR U20837 ( .A(n16459), .B(p_input[515]), .Z(n20940) );
  XNOR U20838 ( .A(n20954), .B(n20953), .Z(n20944) );
  XOR U20839 ( .A(n20972), .B(n20950), .Z(n20953) );
  XOR U20840 ( .A(p_input[2052]), .B(p_input[516]), .Z(n20950) );
  XNOR U20841 ( .A(p_input[2053]), .B(p_input[517]), .Z(n20972) );
  XOR U20842 ( .A(p_input[2054]), .B(p_input[518]), .Z(n20954) );
  XNOR U20843 ( .A(n20973), .B(n20974), .Z(n20771) );
  AND U20844 ( .A(n243), .B(n20975), .Z(n20974) );
  XNOR U20845 ( .A(n20976), .B(n20977), .Z(n243) );
  AND U20846 ( .A(n20978), .B(n20979), .Z(n20977) );
  XOR U20847 ( .A(n20976), .B(n20781), .Z(n20979) );
  XNOR U20848 ( .A(n20976), .B(n20723), .Z(n20978) );
  XOR U20849 ( .A(n20980), .B(n20981), .Z(n20976) );
  AND U20850 ( .A(n20982), .B(n20983), .Z(n20981) );
  XNOR U20851 ( .A(n20794), .B(n20980), .Z(n20983) );
  XOR U20852 ( .A(n20980), .B(n20735), .Z(n20982) );
  XOR U20853 ( .A(n20984), .B(n20985), .Z(n20980) );
  AND U20854 ( .A(n20986), .B(n20987), .Z(n20985) );
  XNOR U20855 ( .A(n20819), .B(n20984), .Z(n20987) );
  XOR U20856 ( .A(n20984), .B(n20746), .Z(n20986) );
  XOR U20857 ( .A(n20988), .B(n20989), .Z(n20984) );
  AND U20858 ( .A(n20990), .B(n20991), .Z(n20989) );
  XOR U20859 ( .A(n20988), .B(n20756), .Z(n20990) );
  XOR U20860 ( .A(n20992), .B(n20993), .Z(n20712) );
  AND U20861 ( .A(n247), .B(n20975), .Z(n20993) );
  XNOR U20862 ( .A(n20973), .B(n20992), .Z(n20975) );
  XNOR U20863 ( .A(n20994), .B(n20995), .Z(n247) );
  AND U20864 ( .A(n20996), .B(n20997), .Z(n20995) );
  XNOR U20865 ( .A(n20998), .B(n20994), .Z(n20997) );
  IV U20866 ( .A(n20781), .Z(n20998) );
  XNOR U20867 ( .A(n20999), .B(n21000), .Z(n20781) );
  AND U20868 ( .A(n250), .B(n21001), .Z(n21000) );
  XNOR U20869 ( .A(n20999), .B(n21002), .Z(n21001) );
  XNOR U20870 ( .A(n20723), .B(n20994), .Z(n20996) );
  XOR U20871 ( .A(n21003), .B(n21004), .Z(n20723) );
  AND U20872 ( .A(n258), .B(n21005), .Z(n21004) );
  XOR U20873 ( .A(n21006), .B(n21007), .Z(n20994) );
  AND U20874 ( .A(n21008), .B(n21009), .Z(n21007) );
  XNOR U20875 ( .A(n21006), .B(n20794), .Z(n21009) );
  XNOR U20876 ( .A(n21010), .B(n21011), .Z(n20794) );
  AND U20877 ( .A(n250), .B(n21012), .Z(n21011) );
  XOR U20878 ( .A(n21013), .B(n21010), .Z(n21012) );
  XNOR U20879 ( .A(n21014), .B(n21006), .Z(n21008) );
  IV U20880 ( .A(n20735), .Z(n21014) );
  XOR U20881 ( .A(n21015), .B(n21016), .Z(n20735) );
  AND U20882 ( .A(n258), .B(n21017), .Z(n21016) );
  XOR U20883 ( .A(n21018), .B(n21019), .Z(n21006) );
  AND U20884 ( .A(n21020), .B(n21021), .Z(n21019) );
  XNOR U20885 ( .A(n21018), .B(n20819), .Z(n21021) );
  XNOR U20886 ( .A(n21022), .B(n21023), .Z(n20819) );
  AND U20887 ( .A(n250), .B(n21024), .Z(n21023) );
  XNOR U20888 ( .A(n21025), .B(n21022), .Z(n21024) );
  XOR U20889 ( .A(n20746), .B(n21018), .Z(n21020) );
  XOR U20890 ( .A(n21026), .B(n21027), .Z(n20746) );
  AND U20891 ( .A(n258), .B(n21028), .Z(n21027) );
  XOR U20892 ( .A(n20988), .B(n21029), .Z(n21018) );
  AND U20893 ( .A(n21030), .B(n20991), .Z(n21029) );
  XNOR U20894 ( .A(n20865), .B(n20988), .Z(n20991) );
  XNOR U20895 ( .A(n21031), .B(n21032), .Z(n20865) );
  AND U20896 ( .A(n250), .B(n21033), .Z(n21032) );
  XOR U20897 ( .A(n21034), .B(n21031), .Z(n21033) );
  XNOR U20898 ( .A(n21035), .B(n20988), .Z(n21030) );
  IV U20899 ( .A(n20756), .Z(n21035) );
  XOR U20900 ( .A(n21036), .B(n21037), .Z(n20756) );
  AND U20901 ( .A(n258), .B(n21038), .Z(n21037) );
  XOR U20902 ( .A(n21039), .B(n21040), .Z(n20988) );
  AND U20903 ( .A(n21041), .B(n21042), .Z(n21040) );
  XNOR U20904 ( .A(n21039), .B(n20955), .Z(n21042) );
  XNOR U20905 ( .A(n21043), .B(n21044), .Z(n20955) );
  AND U20906 ( .A(n250), .B(n21045), .Z(n21044) );
  XNOR U20907 ( .A(n21046), .B(n21043), .Z(n21045) );
  XNOR U20908 ( .A(n21047), .B(n21039), .Z(n21041) );
  IV U20909 ( .A(n20768), .Z(n21047) );
  XOR U20910 ( .A(n21048), .B(n21049), .Z(n20768) );
  AND U20911 ( .A(n258), .B(n21050), .Z(n21049) );
  AND U20912 ( .A(n20992), .B(n20973), .Z(n21039) );
  XNOR U20913 ( .A(n21051), .B(n21052), .Z(n20973) );
  AND U20914 ( .A(n250), .B(n21053), .Z(n21052) );
  XNOR U20915 ( .A(n21054), .B(n21051), .Z(n21053) );
  XNOR U20916 ( .A(n21055), .B(n21056), .Z(n250) );
  AND U20917 ( .A(n21057), .B(n21058), .Z(n21056) );
  XOR U20918 ( .A(n21002), .B(n21055), .Z(n21058) );
  AND U20919 ( .A(n21059), .B(n21060), .Z(n21002) );
  XOR U20920 ( .A(n21055), .B(n20999), .Z(n21057) );
  XNOR U20921 ( .A(n21061), .B(n21062), .Z(n20999) );
  AND U20922 ( .A(n254), .B(n21005), .Z(n21062) );
  XOR U20923 ( .A(n21003), .B(n21061), .Z(n21005) );
  XOR U20924 ( .A(n21063), .B(n21064), .Z(n21055) );
  AND U20925 ( .A(n21065), .B(n21066), .Z(n21064) );
  XNOR U20926 ( .A(n21063), .B(n21059), .Z(n21066) );
  IV U20927 ( .A(n21013), .Z(n21059) );
  XOR U20928 ( .A(n21067), .B(n21068), .Z(n21013) );
  XOR U20929 ( .A(n21069), .B(n21060), .Z(n21068) );
  AND U20930 ( .A(n21025), .B(n21070), .Z(n21060) );
  AND U20931 ( .A(n21071), .B(n21072), .Z(n21069) );
  XOR U20932 ( .A(n21073), .B(n21067), .Z(n21071) );
  XNOR U20933 ( .A(n21010), .B(n21063), .Z(n21065) );
  XNOR U20934 ( .A(n21074), .B(n21075), .Z(n21010) );
  AND U20935 ( .A(n254), .B(n21017), .Z(n21075) );
  XOR U20936 ( .A(n21074), .B(n21015), .Z(n21017) );
  XOR U20937 ( .A(n21076), .B(n21077), .Z(n21063) );
  AND U20938 ( .A(n21078), .B(n21079), .Z(n21077) );
  XNOR U20939 ( .A(n21076), .B(n21025), .Z(n21079) );
  XOR U20940 ( .A(n21080), .B(n21072), .Z(n21025) );
  XNOR U20941 ( .A(n21081), .B(n21067), .Z(n21072) );
  XOR U20942 ( .A(n21082), .B(n21083), .Z(n21067) );
  AND U20943 ( .A(n21084), .B(n21085), .Z(n21083) );
  XOR U20944 ( .A(n21086), .B(n21082), .Z(n21084) );
  XNOR U20945 ( .A(n21087), .B(n21088), .Z(n21081) );
  AND U20946 ( .A(n21089), .B(n21090), .Z(n21088) );
  XOR U20947 ( .A(n21087), .B(n21091), .Z(n21089) );
  XNOR U20948 ( .A(n21073), .B(n21070), .Z(n21080) );
  AND U20949 ( .A(n21092), .B(n21093), .Z(n21070) );
  XOR U20950 ( .A(n21094), .B(n21095), .Z(n21073) );
  AND U20951 ( .A(n21096), .B(n21097), .Z(n21095) );
  XOR U20952 ( .A(n21094), .B(n21098), .Z(n21096) );
  XNOR U20953 ( .A(n21022), .B(n21076), .Z(n21078) );
  XNOR U20954 ( .A(n21099), .B(n21100), .Z(n21022) );
  AND U20955 ( .A(n254), .B(n21028), .Z(n21100) );
  XOR U20956 ( .A(n21099), .B(n21026), .Z(n21028) );
  XOR U20957 ( .A(n21101), .B(n21102), .Z(n21076) );
  AND U20958 ( .A(n21103), .B(n21104), .Z(n21102) );
  XNOR U20959 ( .A(n21101), .B(n21092), .Z(n21104) );
  IV U20960 ( .A(n21034), .Z(n21092) );
  XNOR U20961 ( .A(n21105), .B(n21085), .Z(n21034) );
  XNOR U20962 ( .A(n21106), .B(n21091), .Z(n21085) );
  XOR U20963 ( .A(n21107), .B(n21108), .Z(n21091) );
  AND U20964 ( .A(n21109), .B(n21110), .Z(n21108) );
  XOR U20965 ( .A(n21107), .B(n21111), .Z(n21109) );
  XNOR U20966 ( .A(n21090), .B(n21082), .Z(n21106) );
  XOR U20967 ( .A(n21112), .B(n21113), .Z(n21082) );
  AND U20968 ( .A(n21114), .B(n21115), .Z(n21113) );
  XNOR U20969 ( .A(n21116), .B(n21112), .Z(n21114) );
  XNOR U20970 ( .A(n21117), .B(n21087), .Z(n21090) );
  XOR U20971 ( .A(n21118), .B(n21119), .Z(n21087) );
  AND U20972 ( .A(n21120), .B(n21121), .Z(n21119) );
  XOR U20973 ( .A(n21118), .B(n21122), .Z(n21120) );
  XNOR U20974 ( .A(n21123), .B(n21124), .Z(n21117) );
  AND U20975 ( .A(n21125), .B(n21126), .Z(n21124) );
  XNOR U20976 ( .A(n21123), .B(n21127), .Z(n21125) );
  XNOR U20977 ( .A(n21086), .B(n21093), .Z(n21105) );
  AND U20978 ( .A(n21046), .B(n21128), .Z(n21093) );
  XOR U20979 ( .A(n21098), .B(n21097), .Z(n21086) );
  XNOR U20980 ( .A(n21129), .B(n21094), .Z(n21097) );
  XOR U20981 ( .A(n21130), .B(n21131), .Z(n21094) );
  AND U20982 ( .A(n21132), .B(n21133), .Z(n21131) );
  XOR U20983 ( .A(n21130), .B(n21134), .Z(n21132) );
  XNOR U20984 ( .A(n21135), .B(n21136), .Z(n21129) );
  AND U20985 ( .A(n21137), .B(n21138), .Z(n21136) );
  XOR U20986 ( .A(n21135), .B(n21139), .Z(n21137) );
  XOR U20987 ( .A(n21140), .B(n21141), .Z(n21098) );
  AND U20988 ( .A(n21142), .B(n21143), .Z(n21141) );
  XOR U20989 ( .A(n21140), .B(n21144), .Z(n21142) );
  XNOR U20990 ( .A(n21031), .B(n21101), .Z(n21103) );
  XNOR U20991 ( .A(n21145), .B(n21146), .Z(n21031) );
  AND U20992 ( .A(n254), .B(n21038), .Z(n21146) );
  XOR U20993 ( .A(n21145), .B(n21036), .Z(n21038) );
  XOR U20994 ( .A(n21147), .B(n21148), .Z(n21101) );
  AND U20995 ( .A(n21149), .B(n21150), .Z(n21148) );
  XNOR U20996 ( .A(n21147), .B(n21046), .Z(n21150) );
  XOR U20997 ( .A(n21151), .B(n21115), .Z(n21046) );
  XNOR U20998 ( .A(n21152), .B(n21122), .Z(n21115) );
  XOR U20999 ( .A(n21111), .B(n21110), .Z(n21122) );
  XNOR U21000 ( .A(n21153), .B(n21107), .Z(n21110) );
  XOR U21001 ( .A(n21154), .B(n21155), .Z(n21107) );
  AND U21002 ( .A(n21156), .B(n21157), .Z(n21155) );
  XOR U21003 ( .A(n21154), .B(n21158), .Z(n21156) );
  XNOR U21004 ( .A(n21159), .B(n21160), .Z(n21153) );
  NOR U21005 ( .A(n21161), .B(n21162), .Z(n21160) );
  XNOR U21006 ( .A(n21159), .B(n21163), .Z(n21161) );
  XOR U21007 ( .A(n21164), .B(n21165), .Z(n21111) );
  NOR U21008 ( .A(n21166), .B(n21167), .Z(n21165) );
  XNOR U21009 ( .A(n21164), .B(n21168), .Z(n21166) );
  XNOR U21010 ( .A(n21121), .B(n21112), .Z(n21152) );
  XOR U21011 ( .A(n21169), .B(n21170), .Z(n21112) );
  NOR U21012 ( .A(n21171), .B(n21172), .Z(n21170) );
  XNOR U21013 ( .A(n21169), .B(n21173), .Z(n21171) );
  XOR U21014 ( .A(n21174), .B(n21127), .Z(n21121) );
  XNOR U21015 ( .A(n21175), .B(n21176), .Z(n21127) );
  NOR U21016 ( .A(n21177), .B(n21178), .Z(n21176) );
  XNOR U21017 ( .A(n21175), .B(n21179), .Z(n21177) );
  XNOR U21018 ( .A(n21126), .B(n21118), .Z(n21174) );
  XOR U21019 ( .A(n21180), .B(n21181), .Z(n21118) );
  AND U21020 ( .A(n21182), .B(n21183), .Z(n21181) );
  XOR U21021 ( .A(n21180), .B(n21184), .Z(n21182) );
  XNOR U21022 ( .A(n21185), .B(n21123), .Z(n21126) );
  XOR U21023 ( .A(n21186), .B(n21187), .Z(n21123) );
  AND U21024 ( .A(n21188), .B(n21189), .Z(n21187) );
  XOR U21025 ( .A(n21186), .B(n21190), .Z(n21188) );
  XNOR U21026 ( .A(n21191), .B(n21192), .Z(n21185) );
  NOR U21027 ( .A(n21193), .B(n21194), .Z(n21192) );
  XOR U21028 ( .A(n21191), .B(n21195), .Z(n21193) );
  XOR U21029 ( .A(n21116), .B(n21128), .Z(n21151) );
  NOR U21030 ( .A(n21054), .B(n21196), .Z(n21128) );
  XNOR U21031 ( .A(n21134), .B(n21133), .Z(n21116) );
  XNOR U21032 ( .A(n21197), .B(n21139), .Z(n21133) );
  XOR U21033 ( .A(n21198), .B(n21199), .Z(n21139) );
  NOR U21034 ( .A(n21200), .B(n21201), .Z(n21199) );
  XNOR U21035 ( .A(n21198), .B(n21202), .Z(n21200) );
  XNOR U21036 ( .A(n21138), .B(n21130), .Z(n21197) );
  XOR U21037 ( .A(n21203), .B(n21204), .Z(n21130) );
  AND U21038 ( .A(n21205), .B(n21206), .Z(n21204) );
  XNOR U21039 ( .A(n21203), .B(n21207), .Z(n21205) );
  XNOR U21040 ( .A(n21208), .B(n21135), .Z(n21138) );
  XOR U21041 ( .A(n21209), .B(n21210), .Z(n21135) );
  AND U21042 ( .A(n21211), .B(n21212), .Z(n21210) );
  XOR U21043 ( .A(n21209), .B(n21213), .Z(n21211) );
  XNOR U21044 ( .A(n21214), .B(n21215), .Z(n21208) );
  NOR U21045 ( .A(n21216), .B(n21217), .Z(n21215) );
  XOR U21046 ( .A(n21214), .B(n21218), .Z(n21216) );
  XOR U21047 ( .A(n21144), .B(n21143), .Z(n21134) );
  XNOR U21048 ( .A(n21219), .B(n21140), .Z(n21143) );
  XOR U21049 ( .A(n21220), .B(n21221), .Z(n21140) );
  AND U21050 ( .A(n21222), .B(n21223), .Z(n21221) );
  XOR U21051 ( .A(n21220), .B(n21224), .Z(n21222) );
  XNOR U21052 ( .A(n21225), .B(n21226), .Z(n21219) );
  NOR U21053 ( .A(n21227), .B(n21228), .Z(n21226) );
  XNOR U21054 ( .A(n21225), .B(n21229), .Z(n21227) );
  XOR U21055 ( .A(n21230), .B(n21231), .Z(n21144) );
  NOR U21056 ( .A(n21232), .B(n21233), .Z(n21231) );
  XNOR U21057 ( .A(n21230), .B(n21234), .Z(n21232) );
  XNOR U21058 ( .A(n21043), .B(n21147), .Z(n21149) );
  XNOR U21059 ( .A(n21235), .B(n21236), .Z(n21043) );
  AND U21060 ( .A(n254), .B(n21050), .Z(n21236) );
  XOR U21061 ( .A(n21235), .B(n21048), .Z(n21050) );
  AND U21062 ( .A(n21051), .B(n21054), .Z(n21147) );
  XOR U21063 ( .A(n21237), .B(n21196), .Z(n21054) );
  XNOR U21064 ( .A(p_input[2048]), .B(p_input[544]), .Z(n21196) );
  XOR U21065 ( .A(n21173), .B(n21172), .Z(n21237) );
  XOR U21066 ( .A(n21238), .B(n21184), .Z(n21172) );
  XOR U21067 ( .A(n21158), .B(n21157), .Z(n21184) );
  XNOR U21068 ( .A(n21239), .B(n21163), .Z(n21157) );
  XOR U21069 ( .A(p_input[2072]), .B(p_input[568]), .Z(n21163) );
  XOR U21070 ( .A(n21154), .B(n21162), .Z(n21239) );
  XOR U21071 ( .A(n21240), .B(n21159), .Z(n21162) );
  XOR U21072 ( .A(p_input[2070]), .B(p_input[566]), .Z(n21159) );
  XNOR U21073 ( .A(p_input[2071]), .B(p_input[567]), .Z(n21240) );
  XNOR U21074 ( .A(n16727), .B(p_input[562]), .Z(n21154) );
  XNOR U21075 ( .A(n21168), .B(n21167), .Z(n21158) );
  XOR U21076 ( .A(n21241), .B(n21164), .Z(n21167) );
  XOR U21077 ( .A(p_input[2067]), .B(p_input[563]), .Z(n21164) );
  XNOR U21078 ( .A(p_input[2068]), .B(p_input[564]), .Z(n21241) );
  XOR U21079 ( .A(p_input[2069]), .B(p_input[565]), .Z(n21168) );
  XNOR U21080 ( .A(n21183), .B(n21169), .Z(n21238) );
  XNOR U21081 ( .A(n16729), .B(p_input[545]), .Z(n21169) );
  XNOR U21082 ( .A(n21242), .B(n21190), .Z(n21183) );
  XNOR U21083 ( .A(n21179), .B(n21178), .Z(n21190) );
  XOR U21084 ( .A(n21243), .B(n21175), .Z(n21178) );
  XNOR U21085 ( .A(n16444), .B(p_input[570]), .Z(n21175) );
  XNOR U21086 ( .A(p_input[2075]), .B(p_input[571]), .Z(n21243) );
  XOR U21087 ( .A(p_input[2076]), .B(p_input[572]), .Z(n21179) );
  XNOR U21088 ( .A(n21189), .B(n21180), .Z(n21242) );
  XNOR U21089 ( .A(n16732), .B(p_input[561]), .Z(n21180) );
  XOR U21090 ( .A(n21244), .B(n21195), .Z(n21189) );
  XNOR U21091 ( .A(p_input[2079]), .B(p_input[575]), .Z(n21195) );
  XOR U21092 ( .A(n21186), .B(n21194), .Z(n21244) );
  XOR U21093 ( .A(n21245), .B(n21191), .Z(n21194) );
  XOR U21094 ( .A(p_input[2077]), .B(p_input[573]), .Z(n21191) );
  XNOR U21095 ( .A(p_input[2078]), .B(p_input[574]), .Z(n21245) );
  XNOR U21096 ( .A(n16448), .B(p_input[569]), .Z(n21186) );
  XNOR U21097 ( .A(n21207), .B(n21206), .Z(n21173) );
  XNOR U21098 ( .A(n21246), .B(n21213), .Z(n21206) );
  XNOR U21099 ( .A(n21202), .B(n21201), .Z(n21213) );
  XOR U21100 ( .A(n21247), .B(n21198), .Z(n21201) );
  XNOR U21101 ( .A(n16737), .B(p_input[555]), .Z(n21198) );
  XNOR U21102 ( .A(p_input[2060]), .B(p_input[556]), .Z(n21247) );
  XOR U21103 ( .A(p_input[2061]), .B(p_input[557]), .Z(n21202) );
  XNOR U21104 ( .A(n21212), .B(n21203), .Z(n21246) );
  XNOR U21105 ( .A(n16452), .B(p_input[546]), .Z(n21203) );
  XOR U21106 ( .A(n21248), .B(n21218), .Z(n21212) );
  XNOR U21107 ( .A(p_input[2064]), .B(p_input[560]), .Z(n21218) );
  XOR U21108 ( .A(n21209), .B(n21217), .Z(n21248) );
  XOR U21109 ( .A(n21249), .B(n21214), .Z(n21217) );
  XOR U21110 ( .A(p_input[2062]), .B(p_input[558]), .Z(n21214) );
  XNOR U21111 ( .A(p_input[2063]), .B(p_input[559]), .Z(n21249) );
  XNOR U21112 ( .A(n16740), .B(p_input[554]), .Z(n21209) );
  XNOR U21113 ( .A(n21224), .B(n21223), .Z(n21207) );
  XNOR U21114 ( .A(n21250), .B(n21229), .Z(n21223) );
  XOR U21115 ( .A(p_input[2057]), .B(p_input[553]), .Z(n21229) );
  XOR U21116 ( .A(n21220), .B(n21228), .Z(n21250) );
  XOR U21117 ( .A(n21251), .B(n21225), .Z(n21228) );
  XOR U21118 ( .A(p_input[2055]), .B(p_input[551]), .Z(n21225) );
  XNOR U21119 ( .A(p_input[2056]), .B(p_input[552]), .Z(n21251) );
  XNOR U21120 ( .A(n16459), .B(p_input[547]), .Z(n21220) );
  XNOR U21121 ( .A(n21234), .B(n21233), .Z(n21224) );
  XOR U21122 ( .A(n21252), .B(n21230), .Z(n21233) );
  XOR U21123 ( .A(p_input[2052]), .B(p_input[548]), .Z(n21230) );
  XNOR U21124 ( .A(p_input[2053]), .B(p_input[549]), .Z(n21252) );
  XOR U21125 ( .A(p_input[2054]), .B(p_input[550]), .Z(n21234) );
  XNOR U21126 ( .A(n21253), .B(n21254), .Z(n21051) );
  AND U21127 ( .A(n254), .B(n21255), .Z(n21254) );
  XNOR U21128 ( .A(n21256), .B(n21257), .Z(n254) );
  AND U21129 ( .A(n21258), .B(n21259), .Z(n21257) );
  XOR U21130 ( .A(n21256), .B(n21061), .Z(n21259) );
  XNOR U21131 ( .A(n21256), .B(n21003), .Z(n21258) );
  XOR U21132 ( .A(n21260), .B(n21261), .Z(n21256) );
  AND U21133 ( .A(n21262), .B(n21263), .Z(n21261) );
  XNOR U21134 ( .A(n21074), .B(n21260), .Z(n21263) );
  XOR U21135 ( .A(n21260), .B(n21015), .Z(n21262) );
  XOR U21136 ( .A(n21264), .B(n21265), .Z(n21260) );
  AND U21137 ( .A(n21266), .B(n21267), .Z(n21265) );
  XNOR U21138 ( .A(n21099), .B(n21264), .Z(n21267) );
  XOR U21139 ( .A(n21264), .B(n21026), .Z(n21266) );
  XOR U21140 ( .A(n21268), .B(n21269), .Z(n21264) );
  AND U21141 ( .A(n21270), .B(n21271), .Z(n21269) );
  XOR U21142 ( .A(n21268), .B(n21036), .Z(n21270) );
  XOR U21143 ( .A(n21272), .B(n21273), .Z(n20992) );
  AND U21144 ( .A(n258), .B(n21255), .Z(n21273) );
  XNOR U21145 ( .A(n21253), .B(n21272), .Z(n21255) );
  XNOR U21146 ( .A(n21274), .B(n21275), .Z(n258) );
  AND U21147 ( .A(n21276), .B(n21277), .Z(n21275) );
  XNOR U21148 ( .A(n21278), .B(n21274), .Z(n21277) );
  IV U21149 ( .A(n21061), .Z(n21278) );
  XNOR U21150 ( .A(n21279), .B(n21280), .Z(n21061) );
  AND U21151 ( .A(n261), .B(n21281), .Z(n21280) );
  XNOR U21152 ( .A(n21279), .B(n21282), .Z(n21281) );
  XNOR U21153 ( .A(n21003), .B(n21274), .Z(n21276) );
  XOR U21154 ( .A(n21283), .B(n21284), .Z(n21003) );
  AND U21155 ( .A(n269), .B(n21285), .Z(n21284) );
  XOR U21156 ( .A(n21286), .B(n21287), .Z(n21274) );
  AND U21157 ( .A(n21288), .B(n21289), .Z(n21287) );
  XNOR U21158 ( .A(n21286), .B(n21074), .Z(n21289) );
  XNOR U21159 ( .A(n21290), .B(n21291), .Z(n21074) );
  AND U21160 ( .A(n261), .B(n21292), .Z(n21291) );
  XOR U21161 ( .A(n21293), .B(n21290), .Z(n21292) );
  XNOR U21162 ( .A(n21294), .B(n21286), .Z(n21288) );
  IV U21163 ( .A(n21015), .Z(n21294) );
  XOR U21164 ( .A(n21295), .B(n21296), .Z(n21015) );
  AND U21165 ( .A(n269), .B(n21297), .Z(n21296) );
  XOR U21166 ( .A(n21298), .B(n21299), .Z(n21286) );
  AND U21167 ( .A(n21300), .B(n21301), .Z(n21299) );
  XNOR U21168 ( .A(n21298), .B(n21099), .Z(n21301) );
  XNOR U21169 ( .A(n21302), .B(n21303), .Z(n21099) );
  AND U21170 ( .A(n261), .B(n21304), .Z(n21303) );
  XNOR U21171 ( .A(n21305), .B(n21302), .Z(n21304) );
  XOR U21172 ( .A(n21026), .B(n21298), .Z(n21300) );
  XOR U21173 ( .A(n21306), .B(n21307), .Z(n21026) );
  AND U21174 ( .A(n269), .B(n21308), .Z(n21307) );
  XOR U21175 ( .A(n21268), .B(n21309), .Z(n21298) );
  AND U21176 ( .A(n21310), .B(n21271), .Z(n21309) );
  XNOR U21177 ( .A(n21145), .B(n21268), .Z(n21271) );
  XNOR U21178 ( .A(n21311), .B(n21312), .Z(n21145) );
  AND U21179 ( .A(n261), .B(n21313), .Z(n21312) );
  XOR U21180 ( .A(n21314), .B(n21311), .Z(n21313) );
  XNOR U21181 ( .A(n21315), .B(n21268), .Z(n21310) );
  IV U21182 ( .A(n21036), .Z(n21315) );
  XOR U21183 ( .A(n21316), .B(n21317), .Z(n21036) );
  AND U21184 ( .A(n269), .B(n21318), .Z(n21317) );
  XOR U21185 ( .A(n21319), .B(n21320), .Z(n21268) );
  AND U21186 ( .A(n21321), .B(n21322), .Z(n21320) );
  XNOR U21187 ( .A(n21319), .B(n21235), .Z(n21322) );
  XNOR U21188 ( .A(n21323), .B(n21324), .Z(n21235) );
  AND U21189 ( .A(n261), .B(n21325), .Z(n21324) );
  XNOR U21190 ( .A(n21326), .B(n21323), .Z(n21325) );
  XNOR U21191 ( .A(n21327), .B(n21319), .Z(n21321) );
  IV U21192 ( .A(n21048), .Z(n21327) );
  XOR U21193 ( .A(n21328), .B(n21329), .Z(n21048) );
  AND U21194 ( .A(n269), .B(n21330), .Z(n21329) );
  AND U21195 ( .A(n21272), .B(n21253), .Z(n21319) );
  XNOR U21196 ( .A(n21331), .B(n21332), .Z(n21253) );
  AND U21197 ( .A(n261), .B(n21333), .Z(n21332) );
  XNOR U21198 ( .A(n21334), .B(n21331), .Z(n21333) );
  XNOR U21199 ( .A(n21335), .B(n21336), .Z(n261) );
  AND U21200 ( .A(n21337), .B(n21338), .Z(n21336) );
  XOR U21201 ( .A(n21282), .B(n21335), .Z(n21338) );
  AND U21202 ( .A(n21339), .B(n21340), .Z(n21282) );
  XOR U21203 ( .A(n21335), .B(n21279), .Z(n21337) );
  XNOR U21204 ( .A(n21341), .B(n21342), .Z(n21279) );
  AND U21205 ( .A(n265), .B(n21285), .Z(n21342) );
  XOR U21206 ( .A(n21283), .B(n21341), .Z(n21285) );
  XOR U21207 ( .A(n21343), .B(n21344), .Z(n21335) );
  AND U21208 ( .A(n21345), .B(n21346), .Z(n21344) );
  XNOR U21209 ( .A(n21343), .B(n21339), .Z(n21346) );
  IV U21210 ( .A(n21293), .Z(n21339) );
  XOR U21211 ( .A(n21347), .B(n21348), .Z(n21293) );
  XOR U21212 ( .A(n21349), .B(n21340), .Z(n21348) );
  AND U21213 ( .A(n21305), .B(n21350), .Z(n21340) );
  AND U21214 ( .A(n21351), .B(n21352), .Z(n21349) );
  XOR U21215 ( .A(n21353), .B(n21347), .Z(n21351) );
  XNOR U21216 ( .A(n21290), .B(n21343), .Z(n21345) );
  XNOR U21217 ( .A(n21354), .B(n21355), .Z(n21290) );
  AND U21218 ( .A(n265), .B(n21297), .Z(n21355) );
  XOR U21219 ( .A(n21354), .B(n21295), .Z(n21297) );
  XOR U21220 ( .A(n21356), .B(n21357), .Z(n21343) );
  AND U21221 ( .A(n21358), .B(n21359), .Z(n21357) );
  XNOR U21222 ( .A(n21356), .B(n21305), .Z(n21359) );
  XOR U21223 ( .A(n21360), .B(n21352), .Z(n21305) );
  XNOR U21224 ( .A(n21361), .B(n21347), .Z(n21352) );
  XOR U21225 ( .A(n21362), .B(n21363), .Z(n21347) );
  AND U21226 ( .A(n21364), .B(n21365), .Z(n21363) );
  XOR U21227 ( .A(n21366), .B(n21362), .Z(n21364) );
  XNOR U21228 ( .A(n21367), .B(n21368), .Z(n21361) );
  AND U21229 ( .A(n21369), .B(n21370), .Z(n21368) );
  XOR U21230 ( .A(n21367), .B(n21371), .Z(n21369) );
  XNOR U21231 ( .A(n21353), .B(n21350), .Z(n21360) );
  AND U21232 ( .A(n21372), .B(n21373), .Z(n21350) );
  XOR U21233 ( .A(n21374), .B(n21375), .Z(n21353) );
  AND U21234 ( .A(n21376), .B(n21377), .Z(n21375) );
  XOR U21235 ( .A(n21374), .B(n21378), .Z(n21376) );
  XNOR U21236 ( .A(n21302), .B(n21356), .Z(n21358) );
  XNOR U21237 ( .A(n21379), .B(n21380), .Z(n21302) );
  AND U21238 ( .A(n265), .B(n21308), .Z(n21380) );
  XOR U21239 ( .A(n21379), .B(n21306), .Z(n21308) );
  XOR U21240 ( .A(n21381), .B(n21382), .Z(n21356) );
  AND U21241 ( .A(n21383), .B(n21384), .Z(n21382) );
  XNOR U21242 ( .A(n21381), .B(n21372), .Z(n21384) );
  IV U21243 ( .A(n21314), .Z(n21372) );
  XNOR U21244 ( .A(n21385), .B(n21365), .Z(n21314) );
  XNOR U21245 ( .A(n21386), .B(n21371), .Z(n21365) );
  XOR U21246 ( .A(n21387), .B(n21388), .Z(n21371) );
  AND U21247 ( .A(n21389), .B(n21390), .Z(n21388) );
  XOR U21248 ( .A(n21387), .B(n21391), .Z(n21389) );
  XNOR U21249 ( .A(n21370), .B(n21362), .Z(n21386) );
  XOR U21250 ( .A(n21392), .B(n21393), .Z(n21362) );
  AND U21251 ( .A(n21394), .B(n21395), .Z(n21393) );
  XNOR U21252 ( .A(n21396), .B(n21392), .Z(n21394) );
  XNOR U21253 ( .A(n21397), .B(n21367), .Z(n21370) );
  XOR U21254 ( .A(n21398), .B(n21399), .Z(n21367) );
  AND U21255 ( .A(n21400), .B(n21401), .Z(n21399) );
  XOR U21256 ( .A(n21398), .B(n21402), .Z(n21400) );
  XNOR U21257 ( .A(n21403), .B(n21404), .Z(n21397) );
  AND U21258 ( .A(n21405), .B(n21406), .Z(n21404) );
  XNOR U21259 ( .A(n21403), .B(n21407), .Z(n21405) );
  XNOR U21260 ( .A(n21366), .B(n21373), .Z(n21385) );
  AND U21261 ( .A(n21326), .B(n21408), .Z(n21373) );
  XOR U21262 ( .A(n21378), .B(n21377), .Z(n21366) );
  XNOR U21263 ( .A(n21409), .B(n21374), .Z(n21377) );
  XOR U21264 ( .A(n21410), .B(n21411), .Z(n21374) );
  AND U21265 ( .A(n21412), .B(n21413), .Z(n21411) );
  XOR U21266 ( .A(n21410), .B(n21414), .Z(n21412) );
  XNOR U21267 ( .A(n21415), .B(n21416), .Z(n21409) );
  AND U21268 ( .A(n21417), .B(n21418), .Z(n21416) );
  XOR U21269 ( .A(n21415), .B(n21419), .Z(n21417) );
  XOR U21270 ( .A(n21420), .B(n21421), .Z(n21378) );
  AND U21271 ( .A(n21422), .B(n21423), .Z(n21421) );
  XOR U21272 ( .A(n21420), .B(n21424), .Z(n21422) );
  XNOR U21273 ( .A(n21311), .B(n21381), .Z(n21383) );
  XNOR U21274 ( .A(n21425), .B(n21426), .Z(n21311) );
  AND U21275 ( .A(n265), .B(n21318), .Z(n21426) );
  XOR U21276 ( .A(n21425), .B(n21316), .Z(n21318) );
  XOR U21277 ( .A(n21427), .B(n21428), .Z(n21381) );
  AND U21278 ( .A(n21429), .B(n21430), .Z(n21428) );
  XNOR U21279 ( .A(n21427), .B(n21326), .Z(n21430) );
  XOR U21280 ( .A(n21431), .B(n21395), .Z(n21326) );
  XNOR U21281 ( .A(n21432), .B(n21402), .Z(n21395) );
  XOR U21282 ( .A(n21391), .B(n21390), .Z(n21402) );
  XNOR U21283 ( .A(n21433), .B(n21387), .Z(n21390) );
  XOR U21284 ( .A(n21434), .B(n21435), .Z(n21387) );
  AND U21285 ( .A(n21436), .B(n21437), .Z(n21435) );
  XOR U21286 ( .A(n21434), .B(n21438), .Z(n21436) );
  XNOR U21287 ( .A(n21439), .B(n21440), .Z(n21433) );
  NOR U21288 ( .A(n21441), .B(n21442), .Z(n21440) );
  XNOR U21289 ( .A(n21439), .B(n21443), .Z(n21441) );
  XOR U21290 ( .A(n21444), .B(n21445), .Z(n21391) );
  NOR U21291 ( .A(n21446), .B(n21447), .Z(n21445) );
  XNOR U21292 ( .A(n21444), .B(n21448), .Z(n21446) );
  XNOR U21293 ( .A(n21401), .B(n21392), .Z(n21432) );
  XOR U21294 ( .A(n21449), .B(n21450), .Z(n21392) );
  NOR U21295 ( .A(n21451), .B(n21452), .Z(n21450) );
  XNOR U21296 ( .A(n21449), .B(n21453), .Z(n21451) );
  XOR U21297 ( .A(n21454), .B(n21407), .Z(n21401) );
  XNOR U21298 ( .A(n21455), .B(n21456), .Z(n21407) );
  NOR U21299 ( .A(n21457), .B(n21458), .Z(n21456) );
  XNOR U21300 ( .A(n21455), .B(n21459), .Z(n21457) );
  XNOR U21301 ( .A(n21406), .B(n21398), .Z(n21454) );
  XOR U21302 ( .A(n21460), .B(n21461), .Z(n21398) );
  AND U21303 ( .A(n21462), .B(n21463), .Z(n21461) );
  XOR U21304 ( .A(n21460), .B(n21464), .Z(n21462) );
  XNOR U21305 ( .A(n21465), .B(n21403), .Z(n21406) );
  XOR U21306 ( .A(n21466), .B(n21467), .Z(n21403) );
  AND U21307 ( .A(n21468), .B(n21469), .Z(n21467) );
  XOR U21308 ( .A(n21466), .B(n21470), .Z(n21468) );
  XNOR U21309 ( .A(n21471), .B(n21472), .Z(n21465) );
  NOR U21310 ( .A(n21473), .B(n21474), .Z(n21472) );
  XOR U21311 ( .A(n21471), .B(n21475), .Z(n21473) );
  XOR U21312 ( .A(n21396), .B(n21408), .Z(n21431) );
  NOR U21313 ( .A(n21334), .B(n21476), .Z(n21408) );
  XNOR U21314 ( .A(n21414), .B(n21413), .Z(n21396) );
  XNOR U21315 ( .A(n21477), .B(n21419), .Z(n21413) );
  XOR U21316 ( .A(n21478), .B(n21479), .Z(n21419) );
  NOR U21317 ( .A(n21480), .B(n21481), .Z(n21479) );
  XNOR U21318 ( .A(n21478), .B(n21482), .Z(n21480) );
  XNOR U21319 ( .A(n21418), .B(n21410), .Z(n21477) );
  XOR U21320 ( .A(n21483), .B(n21484), .Z(n21410) );
  AND U21321 ( .A(n21485), .B(n21486), .Z(n21484) );
  XNOR U21322 ( .A(n21483), .B(n21487), .Z(n21485) );
  XNOR U21323 ( .A(n21488), .B(n21415), .Z(n21418) );
  XOR U21324 ( .A(n21489), .B(n21490), .Z(n21415) );
  AND U21325 ( .A(n21491), .B(n21492), .Z(n21490) );
  XOR U21326 ( .A(n21489), .B(n21493), .Z(n21491) );
  XNOR U21327 ( .A(n21494), .B(n21495), .Z(n21488) );
  NOR U21328 ( .A(n21496), .B(n21497), .Z(n21495) );
  XOR U21329 ( .A(n21494), .B(n21498), .Z(n21496) );
  XOR U21330 ( .A(n21424), .B(n21423), .Z(n21414) );
  XNOR U21331 ( .A(n21499), .B(n21420), .Z(n21423) );
  XOR U21332 ( .A(n21500), .B(n21501), .Z(n21420) );
  AND U21333 ( .A(n21502), .B(n21503), .Z(n21501) );
  XOR U21334 ( .A(n21500), .B(n21504), .Z(n21502) );
  XNOR U21335 ( .A(n21505), .B(n21506), .Z(n21499) );
  NOR U21336 ( .A(n21507), .B(n21508), .Z(n21506) );
  XNOR U21337 ( .A(n21505), .B(n21509), .Z(n21507) );
  XOR U21338 ( .A(n21510), .B(n21511), .Z(n21424) );
  NOR U21339 ( .A(n21512), .B(n21513), .Z(n21511) );
  XNOR U21340 ( .A(n21510), .B(n21514), .Z(n21512) );
  XNOR U21341 ( .A(n21323), .B(n21427), .Z(n21429) );
  XNOR U21342 ( .A(n21515), .B(n21516), .Z(n21323) );
  AND U21343 ( .A(n265), .B(n21330), .Z(n21516) );
  XOR U21344 ( .A(n21515), .B(n21328), .Z(n21330) );
  AND U21345 ( .A(n21331), .B(n21334), .Z(n21427) );
  XOR U21346 ( .A(n21517), .B(n21476), .Z(n21334) );
  XNOR U21347 ( .A(p_input[2048]), .B(p_input[576]), .Z(n21476) );
  XOR U21348 ( .A(n21453), .B(n21452), .Z(n21517) );
  XOR U21349 ( .A(n21518), .B(n21464), .Z(n21452) );
  XOR U21350 ( .A(n21438), .B(n21437), .Z(n21464) );
  XNOR U21351 ( .A(n21519), .B(n21443), .Z(n21437) );
  XOR U21352 ( .A(p_input[2072]), .B(p_input[600]), .Z(n21443) );
  XOR U21353 ( .A(n21434), .B(n21442), .Z(n21519) );
  XOR U21354 ( .A(n21520), .B(n21439), .Z(n21442) );
  XOR U21355 ( .A(p_input[2070]), .B(p_input[598]), .Z(n21439) );
  XNOR U21356 ( .A(p_input[2071]), .B(p_input[599]), .Z(n21520) );
  XNOR U21357 ( .A(n16727), .B(p_input[594]), .Z(n21434) );
  XNOR U21358 ( .A(n21448), .B(n21447), .Z(n21438) );
  XOR U21359 ( .A(n21521), .B(n21444), .Z(n21447) );
  XOR U21360 ( .A(p_input[2067]), .B(p_input[595]), .Z(n21444) );
  XNOR U21361 ( .A(p_input[2068]), .B(p_input[596]), .Z(n21521) );
  XOR U21362 ( .A(p_input[2069]), .B(p_input[597]), .Z(n21448) );
  XNOR U21363 ( .A(n21463), .B(n21449), .Z(n21518) );
  XNOR U21364 ( .A(n16729), .B(p_input[577]), .Z(n21449) );
  XNOR U21365 ( .A(n21522), .B(n21470), .Z(n21463) );
  XNOR U21366 ( .A(n21459), .B(n21458), .Z(n21470) );
  XOR U21367 ( .A(n21523), .B(n21455), .Z(n21458) );
  XNOR U21368 ( .A(n16444), .B(p_input[602]), .Z(n21455) );
  XNOR U21369 ( .A(p_input[2075]), .B(p_input[603]), .Z(n21523) );
  XOR U21370 ( .A(p_input[2076]), .B(p_input[604]), .Z(n21459) );
  XNOR U21371 ( .A(n21469), .B(n21460), .Z(n21522) );
  XNOR U21372 ( .A(n16732), .B(p_input[593]), .Z(n21460) );
  XOR U21373 ( .A(n21524), .B(n21475), .Z(n21469) );
  XNOR U21374 ( .A(p_input[2079]), .B(p_input[607]), .Z(n21475) );
  XOR U21375 ( .A(n21466), .B(n21474), .Z(n21524) );
  XOR U21376 ( .A(n21525), .B(n21471), .Z(n21474) );
  XOR U21377 ( .A(p_input[2077]), .B(p_input[605]), .Z(n21471) );
  XNOR U21378 ( .A(p_input[2078]), .B(p_input[606]), .Z(n21525) );
  XNOR U21379 ( .A(n16448), .B(p_input[601]), .Z(n21466) );
  XNOR U21380 ( .A(n21487), .B(n21486), .Z(n21453) );
  XNOR U21381 ( .A(n21526), .B(n21493), .Z(n21486) );
  XNOR U21382 ( .A(n21482), .B(n21481), .Z(n21493) );
  XOR U21383 ( .A(n21527), .B(n21478), .Z(n21481) );
  XNOR U21384 ( .A(n16737), .B(p_input[587]), .Z(n21478) );
  XNOR U21385 ( .A(p_input[2060]), .B(p_input[588]), .Z(n21527) );
  XOR U21386 ( .A(p_input[2061]), .B(p_input[589]), .Z(n21482) );
  XNOR U21387 ( .A(n21492), .B(n21483), .Z(n21526) );
  XNOR U21388 ( .A(n16452), .B(p_input[578]), .Z(n21483) );
  XOR U21389 ( .A(n21528), .B(n21498), .Z(n21492) );
  XNOR U21390 ( .A(p_input[2064]), .B(p_input[592]), .Z(n21498) );
  XOR U21391 ( .A(n21489), .B(n21497), .Z(n21528) );
  XOR U21392 ( .A(n21529), .B(n21494), .Z(n21497) );
  XOR U21393 ( .A(p_input[2062]), .B(p_input[590]), .Z(n21494) );
  XNOR U21394 ( .A(p_input[2063]), .B(p_input[591]), .Z(n21529) );
  XNOR U21395 ( .A(n16740), .B(p_input[586]), .Z(n21489) );
  XNOR U21396 ( .A(n21504), .B(n21503), .Z(n21487) );
  XNOR U21397 ( .A(n21530), .B(n21509), .Z(n21503) );
  XOR U21398 ( .A(p_input[2057]), .B(p_input[585]), .Z(n21509) );
  XOR U21399 ( .A(n21500), .B(n21508), .Z(n21530) );
  XOR U21400 ( .A(n21531), .B(n21505), .Z(n21508) );
  XOR U21401 ( .A(p_input[2055]), .B(p_input[583]), .Z(n21505) );
  XNOR U21402 ( .A(p_input[2056]), .B(p_input[584]), .Z(n21531) );
  XNOR U21403 ( .A(n16459), .B(p_input[579]), .Z(n21500) );
  XNOR U21404 ( .A(n21514), .B(n21513), .Z(n21504) );
  XOR U21405 ( .A(n21532), .B(n21510), .Z(n21513) );
  XOR U21406 ( .A(p_input[2052]), .B(p_input[580]), .Z(n21510) );
  XNOR U21407 ( .A(p_input[2053]), .B(p_input[581]), .Z(n21532) );
  XOR U21408 ( .A(p_input[2054]), .B(p_input[582]), .Z(n21514) );
  XNOR U21409 ( .A(n21533), .B(n21534), .Z(n21331) );
  AND U21410 ( .A(n265), .B(n21535), .Z(n21534) );
  XNOR U21411 ( .A(n21536), .B(n21537), .Z(n265) );
  AND U21412 ( .A(n21538), .B(n21539), .Z(n21537) );
  XOR U21413 ( .A(n21536), .B(n21341), .Z(n21539) );
  XNOR U21414 ( .A(n21536), .B(n21283), .Z(n21538) );
  XOR U21415 ( .A(n21540), .B(n21541), .Z(n21536) );
  AND U21416 ( .A(n21542), .B(n21543), .Z(n21541) );
  XNOR U21417 ( .A(n21354), .B(n21540), .Z(n21543) );
  XOR U21418 ( .A(n21540), .B(n21295), .Z(n21542) );
  XOR U21419 ( .A(n21544), .B(n21545), .Z(n21540) );
  AND U21420 ( .A(n21546), .B(n21547), .Z(n21545) );
  XNOR U21421 ( .A(n21379), .B(n21544), .Z(n21547) );
  XOR U21422 ( .A(n21544), .B(n21306), .Z(n21546) );
  XOR U21423 ( .A(n21548), .B(n21549), .Z(n21544) );
  AND U21424 ( .A(n21550), .B(n21551), .Z(n21549) );
  XOR U21425 ( .A(n21548), .B(n21316), .Z(n21550) );
  XOR U21426 ( .A(n21552), .B(n21553), .Z(n21272) );
  AND U21427 ( .A(n269), .B(n21535), .Z(n21553) );
  XNOR U21428 ( .A(n21533), .B(n21552), .Z(n21535) );
  XNOR U21429 ( .A(n21554), .B(n21555), .Z(n269) );
  AND U21430 ( .A(n21556), .B(n21557), .Z(n21555) );
  XNOR U21431 ( .A(n21558), .B(n21554), .Z(n21557) );
  IV U21432 ( .A(n21341), .Z(n21558) );
  XNOR U21433 ( .A(n21559), .B(n21560), .Z(n21341) );
  AND U21434 ( .A(n272), .B(n21561), .Z(n21560) );
  XNOR U21435 ( .A(n21559), .B(n21562), .Z(n21561) );
  XNOR U21436 ( .A(n21283), .B(n21554), .Z(n21556) );
  XOR U21437 ( .A(n21563), .B(n21564), .Z(n21283) );
  AND U21438 ( .A(n280), .B(n21565), .Z(n21564) );
  XOR U21439 ( .A(n21566), .B(n21567), .Z(n21554) );
  AND U21440 ( .A(n21568), .B(n21569), .Z(n21567) );
  XNOR U21441 ( .A(n21566), .B(n21354), .Z(n21569) );
  XNOR U21442 ( .A(n21570), .B(n21571), .Z(n21354) );
  AND U21443 ( .A(n272), .B(n21572), .Z(n21571) );
  XOR U21444 ( .A(n21573), .B(n21570), .Z(n21572) );
  XNOR U21445 ( .A(n21574), .B(n21566), .Z(n21568) );
  IV U21446 ( .A(n21295), .Z(n21574) );
  XOR U21447 ( .A(n21575), .B(n21576), .Z(n21295) );
  AND U21448 ( .A(n280), .B(n21577), .Z(n21576) );
  XOR U21449 ( .A(n21578), .B(n21579), .Z(n21566) );
  AND U21450 ( .A(n21580), .B(n21581), .Z(n21579) );
  XNOR U21451 ( .A(n21578), .B(n21379), .Z(n21581) );
  XNOR U21452 ( .A(n21582), .B(n21583), .Z(n21379) );
  AND U21453 ( .A(n272), .B(n21584), .Z(n21583) );
  XNOR U21454 ( .A(n21585), .B(n21582), .Z(n21584) );
  XOR U21455 ( .A(n21306), .B(n21578), .Z(n21580) );
  XOR U21456 ( .A(n21586), .B(n21587), .Z(n21306) );
  AND U21457 ( .A(n280), .B(n21588), .Z(n21587) );
  XOR U21458 ( .A(n21548), .B(n21589), .Z(n21578) );
  AND U21459 ( .A(n21590), .B(n21551), .Z(n21589) );
  XNOR U21460 ( .A(n21425), .B(n21548), .Z(n21551) );
  XNOR U21461 ( .A(n21591), .B(n21592), .Z(n21425) );
  AND U21462 ( .A(n272), .B(n21593), .Z(n21592) );
  XOR U21463 ( .A(n21594), .B(n21591), .Z(n21593) );
  XNOR U21464 ( .A(n21595), .B(n21548), .Z(n21590) );
  IV U21465 ( .A(n21316), .Z(n21595) );
  XOR U21466 ( .A(n21596), .B(n21597), .Z(n21316) );
  AND U21467 ( .A(n280), .B(n21598), .Z(n21597) );
  XOR U21468 ( .A(n21599), .B(n21600), .Z(n21548) );
  AND U21469 ( .A(n21601), .B(n21602), .Z(n21600) );
  XNOR U21470 ( .A(n21599), .B(n21515), .Z(n21602) );
  XNOR U21471 ( .A(n21603), .B(n21604), .Z(n21515) );
  AND U21472 ( .A(n272), .B(n21605), .Z(n21604) );
  XNOR U21473 ( .A(n21606), .B(n21603), .Z(n21605) );
  XNOR U21474 ( .A(n21607), .B(n21599), .Z(n21601) );
  IV U21475 ( .A(n21328), .Z(n21607) );
  XOR U21476 ( .A(n21608), .B(n21609), .Z(n21328) );
  AND U21477 ( .A(n280), .B(n21610), .Z(n21609) );
  AND U21478 ( .A(n21552), .B(n21533), .Z(n21599) );
  XNOR U21479 ( .A(n21611), .B(n21612), .Z(n21533) );
  AND U21480 ( .A(n272), .B(n21613), .Z(n21612) );
  XNOR U21481 ( .A(n21614), .B(n21611), .Z(n21613) );
  XNOR U21482 ( .A(n21615), .B(n21616), .Z(n272) );
  AND U21483 ( .A(n21617), .B(n21618), .Z(n21616) );
  XOR U21484 ( .A(n21562), .B(n21615), .Z(n21618) );
  AND U21485 ( .A(n21619), .B(n21620), .Z(n21562) );
  XOR U21486 ( .A(n21615), .B(n21559), .Z(n21617) );
  XNOR U21487 ( .A(n21621), .B(n21622), .Z(n21559) );
  AND U21488 ( .A(n276), .B(n21565), .Z(n21622) );
  XOR U21489 ( .A(n21563), .B(n21621), .Z(n21565) );
  XOR U21490 ( .A(n21623), .B(n21624), .Z(n21615) );
  AND U21491 ( .A(n21625), .B(n21626), .Z(n21624) );
  XNOR U21492 ( .A(n21623), .B(n21619), .Z(n21626) );
  IV U21493 ( .A(n21573), .Z(n21619) );
  XOR U21494 ( .A(n21627), .B(n21628), .Z(n21573) );
  XOR U21495 ( .A(n21629), .B(n21620), .Z(n21628) );
  AND U21496 ( .A(n21585), .B(n21630), .Z(n21620) );
  AND U21497 ( .A(n21631), .B(n21632), .Z(n21629) );
  XOR U21498 ( .A(n21633), .B(n21627), .Z(n21631) );
  XNOR U21499 ( .A(n21570), .B(n21623), .Z(n21625) );
  XNOR U21500 ( .A(n21634), .B(n21635), .Z(n21570) );
  AND U21501 ( .A(n276), .B(n21577), .Z(n21635) );
  XOR U21502 ( .A(n21634), .B(n21575), .Z(n21577) );
  XOR U21503 ( .A(n21636), .B(n21637), .Z(n21623) );
  AND U21504 ( .A(n21638), .B(n21639), .Z(n21637) );
  XNOR U21505 ( .A(n21636), .B(n21585), .Z(n21639) );
  XOR U21506 ( .A(n21640), .B(n21632), .Z(n21585) );
  XNOR U21507 ( .A(n21641), .B(n21627), .Z(n21632) );
  XOR U21508 ( .A(n21642), .B(n21643), .Z(n21627) );
  AND U21509 ( .A(n21644), .B(n21645), .Z(n21643) );
  XOR U21510 ( .A(n21646), .B(n21642), .Z(n21644) );
  XNOR U21511 ( .A(n21647), .B(n21648), .Z(n21641) );
  AND U21512 ( .A(n21649), .B(n21650), .Z(n21648) );
  XOR U21513 ( .A(n21647), .B(n21651), .Z(n21649) );
  XNOR U21514 ( .A(n21633), .B(n21630), .Z(n21640) );
  AND U21515 ( .A(n21652), .B(n21653), .Z(n21630) );
  XOR U21516 ( .A(n21654), .B(n21655), .Z(n21633) );
  AND U21517 ( .A(n21656), .B(n21657), .Z(n21655) );
  XOR U21518 ( .A(n21654), .B(n21658), .Z(n21656) );
  XNOR U21519 ( .A(n21582), .B(n21636), .Z(n21638) );
  XNOR U21520 ( .A(n21659), .B(n21660), .Z(n21582) );
  AND U21521 ( .A(n276), .B(n21588), .Z(n21660) );
  XOR U21522 ( .A(n21659), .B(n21586), .Z(n21588) );
  XOR U21523 ( .A(n21661), .B(n21662), .Z(n21636) );
  AND U21524 ( .A(n21663), .B(n21664), .Z(n21662) );
  XNOR U21525 ( .A(n21661), .B(n21652), .Z(n21664) );
  IV U21526 ( .A(n21594), .Z(n21652) );
  XNOR U21527 ( .A(n21665), .B(n21645), .Z(n21594) );
  XNOR U21528 ( .A(n21666), .B(n21651), .Z(n21645) );
  XOR U21529 ( .A(n21667), .B(n21668), .Z(n21651) );
  AND U21530 ( .A(n21669), .B(n21670), .Z(n21668) );
  XOR U21531 ( .A(n21667), .B(n21671), .Z(n21669) );
  XNOR U21532 ( .A(n21650), .B(n21642), .Z(n21666) );
  XOR U21533 ( .A(n21672), .B(n21673), .Z(n21642) );
  AND U21534 ( .A(n21674), .B(n21675), .Z(n21673) );
  XNOR U21535 ( .A(n21676), .B(n21672), .Z(n21674) );
  XNOR U21536 ( .A(n21677), .B(n21647), .Z(n21650) );
  XOR U21537 ( .A(n21678), .B(n21679), .Z(n21647) );
  AND U21538 ( .A(n21680), .B(n21681), .Z(n21679) );
  XOR U21539 ( .A(n21678), .B(n21682), .Z(n21680) );
  XNOR U21540 ( .A(n21683), .B(n21684), .Z(n21677) );
  AND U21541 ( .A(n21685), .B(n21686), .Z(n21684) );
  XNOR U21542 ( .A(n21683), .B(n21687), .Z(n21685) );
  XNOR U21543 ( .A(n21646), .B(n21653), .Z(n21665) );
  AND U21544 ( .A(n21606), .B(n21688), .Z(n21653) );
  XOR U21545 ( .A(n21658), .B(n21657), .Z(n21646) );
  XNOR U21546 ( .A(n21689), .B(n21654), .Z(n21657) );
  XOR U21547 ( .A(n21690), .B(n21691), .Z(n21654) );
  AND U21548 ( .A(n21692), .B(n21693), .Z(n21691) );
  XOR U21549 ( .A(n21690), .B(n21694), .Z(n21692) );
  XNOR U21550 ( .A(n21695), .B(n21696), .Z(n21689) );
  AND U21551 ( .A(n21697), .B(n21698), .Z(n21696) );
  XOR U21552 ( .A(n21695), .B(n21699), .Z(n21697) );
  XOR U21553 ( .A(n21700), .B(n21701), .Z(n21658) );
  AND U21554 ( .A(n21702), .B(n21703), .Z(n21701) );
  XOR U21555 ( .A(n21700), .B(n21704), .Z(n21702) );
  XNOR U21556 ( .A(n21591), .B(n21661), .Z(n21663) );
  XNOR U21557 ( .A(n21705), .B(n21706), .Z(n21591) );
  AND U21558 ( .A(n276), .B(n21598), .Z(n21706) );
  XOR U21559 ( .A(n21705), .B(n21596), .Z(n21598) );
  XOR U21560 ( .A(n21707), .B(n21708), .Z(n21661) );
  AND U21561 ( .A(n21709), .B(n21710), .Z(n21708) );
  XNOR U21562 ( .A(n21707), .B(n21606), .Z(n21710) );
  XOR U21563 ( .A(n21711), .B(n21675), .Z(n21606) );
  XNOR U21564 ( .A(n21712), .B(n21682), .Z(n21675) );
  XOR U21565 ( .A(n21671), .B(n21670), .Z(n21682) );
  XNOR U21566 ( .A(n21713), .B(n21667), .Z(n21670) );
  XOR U21567 ( .A(n21714), .B(n21715), .Z(n21667) );
  AND U21568 ( .A(n21716), .B(n21717), .Z(n21715) );
  XOR U21569 ( .A(n21714), .B(n21718), .Z(n21716) );
  XNOR U21570 ( .A(n21719), .B(n21720), .Z(n21713) );
  NOR U21571 ( .A(n21721), .B(n21722), .Z(n21720) );
  XNOR U21572 ( .A(n21719), .B(n21723), .Z(n21721) );
  XOR U21573 ( .A(n21724), .B(n21725), .Z(n21671) );
  NOR U21574 ( .A(n21726), .B(n21727), .Z(n21725) );
  XNOR U21575 ( .A(n21724), .B(n21728), .Z(n21726) );
  XNOR U21576 ( .A(n21681), .B(n21672), .Z(n21712) );
  XOR U21577 ( .A(n21729), .B(n21730), .Z(n21672) );
  NOR U21578 ( .A(n21731), .B(n21732), .Z(n21730) );
  XNOR U21579 ( .A(n21729), .B(n21733), .Z(n21731) );
  XOR U21580 ( .A(n21734), .B(n21687), .Z(n21681) );
  XNOR U21581 ( .A(n21735), .B(n21736), .Z(n21687) );
  NOR U21582 ( .A(n21737), .B(n21738), .Z(n21736) );
  XNOR U21583 ( .A(n21735), .B(n21739), .Z(n21737) );
  XNOR U21584 ( .A(n21686), .B(n21678), .Z(n21734) );
  XOR U21585 ( .A(n21740), .B(n21741), .Z(n21678) );
  AND U21586 ( .A(n21742), .B(n21743), .Z(n21741) );
  XOR U21587 ( .A(n21740), .B(n21744), .Z(n21742) );
  XNOR U21588 ( .A(n21745), .B(n21683), .Z(n21686) );
  XOR U21589 ( .A(n21746), .B(n21747), .Z(n21683) );
  AND U21590 ( .A(n21748), .B(n21749), .Z(n21747) );
  XOR U21591 ( .A(n21746), .B(n21750), .Z(n21748) );
  XNOR U21592 ( .A(n21751), .B(n21752), .Z(n21745) );
  NOR U21593 ( .A(n21753), .B(n21754), .Z(n21752) );
  XOR U21594 ( .A(n21751), .B(n21755), .Z(n21753) );
  XOR U21595 ( .A(n21676), .B(n21688), .Z(n21711) );
  NOR U21596 ( .A(n21614), .B(n21756), .Z(n21688) );
  XNOR U21597 ( .A(n21694), .B(n21693), .Z(n21676) );
  XNOR U21598 ( .A(n21757), .B(n21699), .Z(n21693) );
  XOR U21599 ( .A(n21758), .B(n21759), .Z(n21699) );
  NOR U21600 ( .A(n21760), .B(n21761), .Z(n21759) );
  XNOR U21601 ( .A(n21758), .B(n21762), .Z(n21760) );
  XNOR U21602 ( .A(n21698), .B(n21690), .Z(n21757) );
  XOR U21603 ( .A(n21763), .B(n21764), .Z(n21690) );
  AND U21604 ( .A(n21765), .B(n21766), .Z(n21764) );
  XNOR U21605 ( .A(n21763), .B(n21767), .Z(n21765) );
  XNOR U21606 ( .A(n21768), .B(n21695), .Z(n21698) );
  XOR U21607 ( .A(n21769), .B(n21770), .Z(n21695) );
  AND U21608 ( .A(n21771), .B(n21772), .Z(n21770) );
  XOR U21609 ( .A(n21769), .B(n21773), .Z(n21771) );
  XNOR U21610 ( .A(n21774), .B(n21775), .Z(n21768) );
  NOR U21611 ( .A(n21776), .B(n21777), .Z(n21775) );
  XOR U21612 ( .A(n21774), .B(n21778), .Z(n21776) );
  XOR U21613 ( .A(n21704), .B(n21703), .Z(n21694) );
  XNOR U21614 ( .A(n21779), .B(n21700), .Z(n21703) );
  XOR U21615 ( .A(n21780), .B(n21781), .Z(n21700) );
  AND U21616 ( .A(n21782), .B(n21783), .Z(n21781) );
  XOR U21617 ( .A(n21780), .B(n21784), .Z(n21782) );
  XNOR U21618 ( .A(n21785), .B(n21786), .Z(n21779) );
  NOR U21619 ( .A(n21787), .B(n21788), .Z(n21786) );
  XNOR U21620 ( .A(n21785), .B(n21789), .Z(n21787) );
  XOR U21621 ( .A(n21790), .B(n21791), .Z(n21704) );
  NOR U21622 ( .A(n21792), .B(n21793), .Z(n21791) );
  XNOR U21623 ( .A(n21790), .B(n21794), .Z(n21792) );
  XNOR U21624 ( .A(n21603), .B(n21707), .Z(n21709) );
  XNOR U21625 ( .A(n21795), .B(n21796), .Z(n21603) );
  AND U21626 ( .A(n276), .B(n21610), .Z(n21796) );
  XOR U21627 ( .A(n21795), .B(n21608), .Z(n21610) );
  AND U21628 ( .A(n21611), .B(n21614), .Z(n21707) );
  XOR U21629 ( .A(n21797), .B(n21756), .Z(n21614) );
  XNOR U21630 ( .A(p_input[2048]), .B(p_input[608]), .Z(n21756) );
  XOR U21631 ( .A(n21733), .B(n21732), .Z(n21797) );
  XOR U21632 ( .A(n21798), .B(n21744), .Z(n21732) );
  XOR U21633 ( .A(n21718), .B(n21717), .Z(n21744) );
  XNOR U21634 ( .A(n21799), .B(n21723), .Z(n21717) );
  XOR U21635 ( .A(p_input[2072]), .B(p_input[632]), .Z(n21723) );
  XOR U21636 ( .A(n21714), .B(n21722), .Z(n21799) );
  XOR U21637 ( .A(n21800), .B(n21719), .Z(n21722) );
  XOR U21638 ( .A(p_input[2070]), .B(p_input[630]), .Z(n21719) );
  XNOR U21639 ( .A(p_input[2071]), .B(p_input[631]), .Z(n21800) );
  XNOR U21640 ( .A(n16727), .B(p_input[626]), .Z(n21714) );
  XNOR U21641 ( .A(n21728), .B(n21727), .Z(n21718) );
  XOR U21642 ( .A(n21801), .B(n21724), .Z(n21727) );
  XOR U21643 ( .A(p_input[2067]), .B(p_input[627]), .Z(n21724) );
  XNOR U21644 ( .A(p_input[2068]), .B(p_input[628]), .Z(n21801) );
  XOR U21645 ( .A(p_input[2069]), .B(p_input[629]), .Z(n21728) );
  XNOR U21646 ( .A(n21743), .B(n21729), .Z(n21798) );
  XNOR U21647 ( .A(n16729), .B(p_input[609]), .Z(n21729) );
  XNOR U21648 ( .A(n21802), .B(n21750), .Z(n21743) );
  XNOR U21649 ( .A(n21739), .B(n21738), .Z(n21750) );
  XOR U21650 ( .A(n21803), .B(n21735), .Z(n21738) );
  XNOR U21651 ( .A(n16444), .B(p_input[634]), .Z(n21735) );
  XNOR U21652 ( .A(p_input[2075]), .B(p_input[635]), .Z(n21803) );
  XOR U21653 ( .A(p_input[2076]), .B(p_input[636]), .Z(n21739) );
  XNOR U21654 ( .A(n21749), .B(n21740), .Z(n21802) );
  XNOR U21655 ( .A(n16732), .B(p_input[625]), .Z(n21740) );
  XOR U21656 ( .A(n21804), .B(n21755), .Z(n21749) );
  XNOR U21657 ( .A(p_input[2079]), .B(p_input[639]), .Z(n21755) );
  XOR U21658 ( .A(n21746), .B(n21754), .Z(n21804) );
  XOR U21659 ( .A(n21805), .B(n21751), .Z(n21754) );
  XOR U21660 ( .A(p_input[2077]), .B(p_input[637]), .Z(n21751) );
  XNOR U21661 ( .A(p_input[2078]), .B(p_input[638]), .Z(n21805) );
  XNOR U21662 ( .A(n16448), .B(p_input[633]), .Z(n21746) );
  XNOR U21663 ( .A(n21767), .B(n21766), .Z(n21733) );
  XNOR U21664 ( .A(n21806), .B(n21773), .Z(n21766) );
  XNOR U21665 ( .A(n21762), .B(n21761), .Z(n21773) );
  XOR U21666 ( .A(n21807), .B(n21758), .Z(n21761) );
  XNOR U21667 ( .A(n16737), .B(p_input[619]), .Z(n21758) );
  XNOR U21668 ( .A(p_input[2060]), .B(p_input[620]), .Z(n21807) );
  XOR U21669 ( .A(p_input[2061]), .B(p_input[621]), .Z(n21762) );
  XNOR U21670 ( .A(n21772), .B(n21763), .Z(n21806) );
  XNOR U21671 ( .A(n16452), .B(p_input[610]), .Z(n21763) );
  XOR U21672 ( .A(n21808), .B(n21778), .Z(n21772) );
  XNOR U21673 ( .A(p_input[2064]), .B(p_input[624]), .Z(n21778) );
  XOR U21674 ( .A(n21769), .B(n21777), .Z(n21808) );
  XOR U21675 ( .A(n21809), .B(n21774), .Z(n21777) );
  XOR U21676 ( .A(p_input[2062]), .B(p_input[622]), .Z(n21774) );
  XNOR U21677 ( .A(p_input[2063]), .B(p_input[623]), .Z(n21809) );
  XNOR U21678 ( .A(n16740), .B(p_input[618]), .Z(n21769) );
  XNOR U21679 ( .A(n21784), .B(n21783), .Z(n21767) );
  XNOR U21680 ( .A(n21810), .B(n21789), .Z(n21783) );
  XOR U21681 ( .A(p_input[2057]), .B(p_input[617]), .Z(n21789) );
  XOR U21682 ( .A(n21780), .B(n21788), .Z(n21810) );
  XOR U21683 ( .A(n21811), .B(n21785), .Z(n21788) );
  XOR U21684 ( .A(p_input[2055]), .B(p_input[615]), .Z(n21785) );
  XNOR U21685 ( .A(p_input[2056]), .B(p_input[616]), .Z(n21811) );
  XNOR U21686 ( .A(n16459), .B(p_input[611]), .Z(n21780) );
  XNOR U21687 ( .A(n21794), .B(n21793), .Z(n21784) );
  XOR U21688 ( .A(n21812), .B(n21790), .Z(n21793) );
  XOR U21689 ( .A(p_input[2052]), .B(p_input[612]), .Z(n21790) );
  XNOR U21690 ( .A(p_input[2053]), .B(p_input[613]), .Z(n21812) );
  XOR U21691 ( .A(p_input[2054]), .B(p_input[614]), .Z(n21794) );
  XNOR U21692 ( .A(n21813), .B(n21814), .Z(n21611) );
  AND U21693 ( .A(n276), .B(n21815), .Z(n21814) );
  XNOR U21694 ( .A(n21816), .B(n21817), .Z(n276) );
  AND U21695 ( .A(n21818), .B(n21819), .Z(n21817) );
  XOR U21696 ( .A(n21816), .B(n21621), .Z(n21819) );
  XNOR U21697 ( .A(n21816), .B(n21563), .Z(n21818) );
  XOR U21698 ( .A(n21820), .B(n21821), .Z(n21816) );
  AND U21699 ( .A(n21822), .B(n21823), .Z(n21821) );
  XNOR U21700 ( .A(n21634), .B(n21820), .Z(n21823) );
  XOR U21701 ( .A(n21820), .B(n21575), .Z(n21822) );
  XOR U21702 ( .A(n21824), .B(n21825), .Z(n21820) );
  AND U21703 ( .A(n21826), .B(n21827), .Z(n21825) );
  XNOR U21704 ( .A(n21659), .B(n21824), .Z(n21827) );
  XOR U21705 ( .A(n21824), .B(n21586), .Z(n21826) );
  XOR U21706 ( .A(n21828), .B(n21829), .Z(n21824) );
  AND U21707 ( .A(n21830), .B(n21831), .Z(n21829) );
  XOR U21708 ( .A(n21828), .B(n21596), .Z(n21830) );
  XOR U21709 ( .A(n21832), .B(n21833), .Z(n21552) );
  AND U21710 ( .A(n280), .B(n21815), .Z(n21833) );
  XNOR U21711 ( .A(n21813), .B(n21832), .Z(n21815) );
  XNOR U21712 ( .A(n21834), .B(n21835), .Z(n280) );
  AND U21713 ( .A(n21836), .B(n21837), .Z(n21835) );
  XNOR U21714 ( .A(n21838), .B(n21834), .Z(n21837) );
  IV U21715 ( .A(n21621), .Z(n21838) );
  XNOR U21716 ( .A(n21839), .B(n21840), .Z(n21621) );
  AND U21717 ( .A(n283), .B(n21841), .Z(n21840) );
  XNOR U21718 ( .A(n21839), .B(n21842), .Z(n21841) );
  XNOR U21719 ( .A(n21563), .B(n21834), .Z(n21836) );
  XOR U21720 ( .A(n21843), .B(n21844), .Z(n21563) );
  AND U21721 ( .A(n291), .B(n21845), .Z(n21844) );
  XOR U21722 ( .A(n21846), .B(n21847), .Z(n21834) );
  AND U21723 ( .A(n21848), .B(n21849), .Z(n21847) );
  XNOR U21724 ( .A(n21846), .B(n21634), .Z(n21849) );
  XNOR U21725 ( .A(n21850), .B(n21851), .Z(n21634) );
  AND U21726 ( .A(n283), .B(n21852), .Z(n21851) );
  XOR U21727 ( .A(n21853), .B(n21850), .Z(n21852) );
  XNOR U21728 ( .A(n21854), .B(n21846), .Z(n21848) );
  IV U21729 ( .A(n21575), .Z(n21854) );
  XOR U21730 ( .A(n21855), .B(n21856), .Z(n21575) );
  AND U21731 ( .A(n291), .B(n21857), .Z(n21856) );
  XOR U21732 ( .A(n21858), .B(n21859), .Z(n21846) );
  AND U21733 ( .A(n21860), .B(n21861), .Z(n21859) );
  XNOR U21734 ( .A(n21858), .B(n21659), .Z(n21861) );
  XNOR U21735 ( .A(n21862), .B(n21863), .Z(n21659) );
  AND U21736 ( .A(n283), .B(n21864), .Z(n21863) );
  XNOR U21737 ( .A(n21865), .B(n21862), .Z(n21864) );
  XOR U21738 ( .A(n21586), .B(n21858), .Z(n21860) );
  XOR U21739 ( .A(n21866), .B(n21867), .Z(n21586) );
  AND U21740 ( .A(n291), .B(n21868), .Z(n21867) );
  XOR U21741 ( .A(n21828), .B(n21869), .Z(n21858) );
  AND U21742 ( .A(n21870), .B(n21831), .Z(n21869) );
  XNOR U21743 ( .A(n21705), .B(n21828), .Z(n21831) );
  XNOR U21744 ( .A(n21871), .B(n21872), .Z(n21705) );
  AND U21745 ( .A(n283), .B(n21873), .Z(n21872) );
  XOR U21746 ( .A(n21874), .B(n21871), .Z(n21873) );
  XNOR U21747 ( .A(n21875), .B(n21828), .Z(n21870) );
  IV U21748 ( .A(n21596), .Z(n21875) );
  XOR U21749 ( .A(n21876), .B(n21877), .Z(n21596) );
  AND U21750 ( .A(n291), .B(n21878), .Z(n21877) );
  XOR U21751 ( .A(n21879), .B(n21880), .Z(n21828) );
  AND U21752 ( .A(n21881), .B(n21882), .Z(n21880) );
  XNOR U21753 ( .A(n21879), .B(n21795), .Z(n21882) );
  XNOR U21754 ( .A(n21883), .B(n21884), .Z(n21795) );
  AND U21755 ( .A(n283), .B(n21885), .Z(n21884) );
  XNOR U21756 ( .A(n21886), .B(n21883), .Z(n21885) );
  XNOR U21757 ( .A(n21887), .B(n21879), .Z(n21881) );
  IV U21758 ( .A(n21608), .Z(n21887) );
  XOR U21759 ( .A(n21888), .B(n21889), .Z(n21608) );
  AND U21760 ( .A(n291), .B(n21890), .Z(n21889) );
  AND U21761 ( .A(n21832), .B(n21813), .Z(n21879) );
  XNOR U21762 ( .A(n21891), .B(n21892), .Z(n21813) );
  AND U21763 ( .A(n283), .B(n21893), .Z(n21892) );
  XNOR U21764 ( .A(n21894), .B(n21891), .Z(n21893) );
  XNOR U21765 ( .A(n21895), .B(n21896), .Z(n283) );
  AND U21766 ( .A(n21897), .B(n21898), .Z(n21896) );
  XOR U21767 ( .A(n21842), .B(n21895), .Z(n21898) );
  AND U21768 ( .A(n21899), .B(n21900), .Z(n21842) );
  XOR U21769 ( .A(n21895), .B(n21839), .Z(n21897) );
  XNOR U21770 ( .A(n21901), .B(n21902), .Z(n21839) );
  AND U21771 ( .A(n287), .B(n21845), .Z(n21902) );
  XOR U21772 ( .A(n21843), .B(n21901), .Z(n21845) );
  XOR U21773 ( .A(n21903), .B(n21904), .Z(n21895) );
  AND U21774 ( .A(n21905), .B(n21906), .Z(n21904) );
  XNOR U21775 ( .A(n21903), .B(n21899), .Z(n21906) );
  IV U21776 ( .A(n21853), .Z(n21899) );
  XOR U21777 ( .A(n21907), .B(n21908), .Z(n21853) );
  XOR U21778 ( .A(n21909), .B(n21900), .Z(n21908) );
  AND U21779 ( .A(n21865), .B(n21910), .Z(n21900) );
  AND U21780 ( .A(n21911), .B(n21912), .Z(n21909) );
  XOR U21781 ( .A(n21913), .B(n21907), .Z(n21911) );
  XNOR U21782 ( .A(n21850), .B(n21903), .Z(n21905) );
  XNOR U21783 ( .A(n21914), .B(n21915), .Z(n21850) );
  AND U21784 ( .A(n287), .B(n21857), .Z(n21915) );
  XOR U21785 ( .A(n21914), .B(n21855), .Z(n21857) );
  XOR U21786 ( .A(n21916), .B(n21917), .Z(n21903) );
  AND U21787 ( .A(n21918), .B(n21919), .Z(n21917) );
  XNOR U21788 ( .A(n21916), .B(n21865), .Z(n21919) );
  XOR U21789 ( .A(n21920), .B(n21912), .Z(n21865) );
  XNOR U21790 ( .A(n21921), .B(n21907), .Z(n21912) );
  XOR U21791 ( .A(n21922), .B(n21923), .Z(n21907) );
  AND U21792 ( .A(n21924), .B(n21925), .Z(n21923) );
  XOR U21793 ( .A(n21926), .B(n21922), .Z(n21924) );
  XNOR U21794 ( .A(n21927), .B(n21928), .Z(n21921) );
  AND U21795 ( .A(n21929), .B(n21930), .Z(n21928) );
  XOR U21796 ( .A(n21927), .B(n21931), .Z(n21929) );
  XNOR U21797 ( .A(n21913), .B(n21910), .Z(n21920) );
  AND U21798 ( .A(n21932), .B(n21933), .Z(n21910) );
  XOR U21799 ( .A(n21934), .B(n21935), .Z(n21913) );
  AND U21800 ( .A(n21936), .B(n21937), .Z(n21935) );
  XOR U21801 ( .A(n21934), .B(n21938), .Z(n21936) );
  XNOR U21802 ( .A(n21862), .B(n21916), .Z(n21918) );
  XNOR U21803 ( .A(n21939), .B(n21940), .Z(n21862) );
  AND U21804 ( .A(n287), .B(n21868), .Z(n21940) );
  XOR U21805 ( .A(n21939), .B(n21866), .Z(n21868) );
  XOR U21806 ( .A(n21941), .B(n21942), .Z(n21916) );
  AND U21807 ( .A(n21943), .B(n21944), .Z(n21942) );
  XNOR U21808 ( .A(n21941), .B(n21932), .Z(n21944) );
  IV U21809 ( .A(n21874), .Z(n21932) );
  XNOR U21810 ( .A(n21945), .B(n21925), .Z(n21874) );
  XNOR U21811 ( .A(n21946), .B(n21931), .Z(n21925) );
  XOR U21812 ( .A(n21947), .B(n21948), .Z(n21931) );
  AND U21813 ( .A(n21949), .B(n21950), .Z(n21948) );
  XOR U21814 ( .A(n21947), .B(n21951), .Z(n21949) );
  XNOR U21815 ( .A(n21930), .B(n21922), .Z(n21946) );
  XOR U21816 ( .A(n21952), .B(n21953), .Z(n21922) );
  AND U21817 ( .A(n21954), .B(n21955), .Z(n21953) );
  XNOR U21818 ( .A(n21956), .B(n21952), .Z(n21954) );
  XNOR U21819 ( .A(n21957), .B(n21927), .Z(n21930) );
  XOR U21820 ( .A(n21958), .B(n21959), .Z(n21927) );
  AND U21821 ( .A(n21960), .B(n21961), .Z(n21959) );
  XOR U21822 ( .A(n21958), .B(n21962), .Z(n21960) );
  XNOR U21823 ( .A(n21963), .B(n21964), .Z(n21957) );
  AND U21824 ( .A(n21965), .B(n21966), .Z(n21964) );
  XNOR U21825 ( .A(n21963), .B(n21967), .Z(n21965) );
  XNOR U21826 ( .A(n21926), .B(n21933), .Z(n21945) );
  AND U21827 ( .A(n21886), .B(n21968), .Z(n21933) );
  XOR U21828 ( .A(n21938), .B(n21937), .Z(n21926) );
  XNOR U21829 ( .A(n21969), .B(n21934), .Z(n21937) );
  XOR U21830 ( .A(n21970), .B(n21971), .Z(n21934) );
  AND U21831 ( .A(n21972), .B(n21973), .Z(n21971) );
  XOR U21832 ( .A(n21970), .B(n21974), .Z(n21972) );
  XNOR U21833 ( .A(n21975), .B(n21976), .Z(n21969) );
  AND U21834 ( .A(n21977), .B(n21978), .Z(n21976) );
  XOR U21835 ( .A(n21975), .B(n21979), .Z(n21977) );
  XOR U21836 ( .A(n21980), .B(n21981), .Z(n21938) );
  AND U21837 ( .A(n21982), .B(n21983), .Z(n21981) );
  XOR U21838 ( .A(n21980), .B(n21984), .Z(n21982) );
  XNOR U21839 ( .A(n21871), .B(n21941), .Z(n21943) );
  XNOR U21840 ( .A(n21985), .B(n21986), .Z(n21871) );
  AND U21841 ( .A(n287), .B(n21878), .Z(n21986) );
  XOR U21842 ( .A(n21985), .B(n21876), .Z(n21878) );
  XOR U21843 ( .A(n21987), .B(n21988), .Z(n21941) );
  AND U21844 ( .A(n21989), .B(n21990), .Z(n21988) );
  XNOR U21845 ( .A(n21987), .B(n21886), .Z(n21990) );
  XOR U21846 ( .A(n21991), .B(n21955), .Z(n21886) );
  XNOR U21847 ( .A(n21992), .B(n21962), .Z(n21955) );
  XOR U21848 ( .A(n21951), .B(n21950), .Z(n21962) );
  XNOR U21849 ( .A(n21993), .B(n21947), .Z(n21950) );
  XOR U21850 ( .A(n21994), .B(n21995), .Z(n21947) );
  AND U21851 ( .A(n21996), .B(n21997), .Z(n21995) );
  XOR U21852 ( .A(n21994), .B(n21998), .Z(n21996) );
  XNOR U21853 ( .A(n21999), .B(n22000), .Z(n21993) );
  NOR U21854 ( .A(n22001), .B(n22002), .Z(n22000) );
  XNOR U21855 ( .A(n21999), .B(n22003), .Z(n22001) );
  XOR U21856 ( .A(n22004), .B(n22005), .Z(n21951) );
  NOR U21857 ( .A(n22006), .B(n22007), .Z(n22005) );
  XNOR U21858 ( .A(n22004), .B(n22008), .Z(n22006) );
  XNOR U21859 ( .A(n21961), .B(n21952), .Z(n21992) );
  XOR U21860 ( .A(n22009), .B(n22010), .Z(n21952) );
  NOR U21861 ( .A(n22011), .B(n22012), .Z(n22010) );
  XNOR U21862 ( .A(n22009), .B(n22013), .Z(n22011) );
  XOR U21863 ( .A(n22014), .B(n21967), .Z(n21961) );
  XNOR U21864 ( .A(n22015), .B(n22016), .Z(n21967) );
  NOR U21865 ( .A(n22017), .B(n22018), .Z(n22016) );
  XNOR U21866 ( .A(n22015), .B(n22019), .Z(n22017) );
  XNOR U21867 ( .A(n21966), .B(n21958), .Z(n22014) );
  XOR U21868 ( .A(n22020), .B(n22021), .Z(n21958) );
  AND U21869 ( .A(n22022), .B(n22023), .Z(n22021) );
  XOR U21870 ( .A(n22020), .B(n22024), .Z(n22022) );
  XNOR U21871 ( .A(n22025), .B(n21963), .Z(n21966) );
  XOR U21872 ( .A(n22026), .B(n22027), .Z(n21963) );
  AND U21873 ( .A(n22028), .B(n22029), .Z(n22027) );
  XOR U21874 ( .A(n22026), .B(n22030), .Z(n22028) );
  XNOR U21875 ( .A(n22031), .B(n22032), .Z(n22025) );
  NOR U21876 ( .A(n22033), .B(n22034), .Z(n22032) );
  XOR U21877 ( .A(n22031), .B(n22035), .Z(n22033) );
  XOR U21878 ( .A(n21956), .B(n21968), .Z(n21991) );
  NOR U21879 ( .A(n21894), .B(n22036), .Z(n21968) );
  XNOR U21880 ( .A(n21974), .B(n21973), .Z(n21956) );
  XNOR U21881 ( .A(n22037), .B(n21979), .Z(n21973) );
  XOR U21882 ( .A(n22038), .B(n22039), .Z(n21979) );
  NOR U21883 ( .A(n22040), .B(n22041), .Z(n22039) );
  XNOR U21884 ( .A(n22038), .B(n22042), .Z(n22040) );
  XNOR U21885 ( .A(n21978), .B(n21970), .Z(n22037) );
  XOR U21886 ( .A(n22043), .B(n22044), .Z(n21970) );
  AND U21887 ( .A(n22045), .B(n22046), .Z(n22044) );
  XNOR U21888 ( .A(n22043), .B(n22047), .Z(n22045) );
  XNOR U21889 ( .A(n22048), .B(n21975), .Z(n21978) );
  XOR U21890 ( .A(n22049), .B(n22050), .Z(n21975) );
  AND U21891 ( .A(n22051), .B(n22052), .Z(n22050) );
  XOR U21892 ( .A(n22049), .B(n22053), .Z(n22051) );
  XNOR U21893 ( .A(n22054), .B(n22055), .Z(n22048) );
  NOR U21894 ( .A(n22056), .B(n22057), .Z(n22055) );
  XOR U21895 ( .A(n22054), .B(n22058), .Z(n22056) );
  XOR U21896 ( .A(n21984), .B(n21983), .Z(n21974) );
  XNOR U21897 ( .A(n22059), .B(n21980), .Z(n21983) );
  XOR U21898 ( .A(n22060), .B(n22061), .Z(n21980) );
  AND U21899 ( .A(n22062), .B(n22063), .Z(n22061) );
  XOR U21900 ( .A(n22060), .B(n22064), .Z(n22062) );
  XNOR U21901 ( .A(n22065), .B(n22066), .Z(n22059) );
  NOR U21902 ( .A(n22067), .B(n22068), .Z(n22066) );
  XNOR U21903 ( .A(n22065), .B(n22069), .Z(n22067) );
  XOR U21904 ( .A(n22070), .B(n22071), .Z(n21984) );
  NOR U21905 ( .A(n22072), .B(n22073), .Z(n22071) );
  XNOR U21906 ( .A(n22070), .B(n22074), .Z(n22072) );
  XNOR U21907 ( .A(n21883), .B(n21987), .Z(n21989) );
  XNOR U21908 ( .A(n22075), .B(n22076), .Z(n21883) );
  AND U21909 ( .A(n287), .B(n21890), .Z(n22076) );
  XOR U21910 ( .A(n22075), .B(n21888), .Z(n21890) );
  AND U21911 ( .A(n21891), .B(n21894), .Z(n21987) );
  XOR U21912 ( .A(n22077), .B(n22036), .Z(n21894) );
  XNOR U21913 ( .A(p_input[2048]), .B(p_input[640]), .Z(n22036) );
  XOR U21914 ( .A(n22013), .B(n22012), .Z(n22077) );
  XOR U21915 ( .A(n22078), .B(n22024), .Z(n22012) );
  XOR U21916 ( .A(n21998), .B(n21997), .Z(n22024) );
  XNOR U21917 ( .A(n22079), .B(n22003), .Z(n21997) );
  XOR U21918 ( .A(p_input[2072]), .B(p_input[664]), .Z(n22003) );
  XOR U21919 ( .A(n21994), .B(n22002), .Z(n22079) );
  XOR U21920 ( .A(n22080), .B(n21999), .Z(n22002) );
  XOR U21921 ( .A(p_input[2070]), .B(p_input[662]), .Z(n21999) );
  XNOR U21922 ( .A(p_input[2071]), .B(p_input[663]), .Z(n22080) );
  XNOR U21923 ( .A(n16727), .B(p_input[658]), .Z(n21994) );
  XNOR U21924 ( .A(n22008), .B(n22007), .Z(n21998) );
  XOR U21925 ( .A(n22081), .B(n22004), .Z(n22007) );
  XOR U21926 ( .A(p_input[2067]), .B(p_input[659]), .Z(n22004) );
  XNOR U21927 ( .A(p_input[2068]), .B(p_input[660]), .Z(n22081) );
  XOR U21928 ( .A(p_input[2069]), .B(p_input[661]), .Z(n22008) );
  XNOR U21929 ( .A(n22023), .B(n22009), .Z(n22078) );
  XNOR U21930 ( .A(n16729), .B(p_input[641]), .Z(n22009) );
  XNOR U21931 ( .A(n22082), .B(n22030), .Z(n22023) );
  XNOR U21932 ( .A(n22019), .B(n22018), .Z(n22030) );
  XOR U21933 ( .A(n22083), .B(n22015), .Z(n22018) );
  XNOR U21934 ( .A(n16444), .B(p_input[666]), .Z(n22015) );
  XNOR U21935 ( .A(p_input[2075]), .B(p_input[667]), .Z(n22083) );
  XOR U21936 ( .A(p_input[2076]), .B(p_input[668]), .Z(n22019) );
  XNOR U21937 ( .A(n22029), .B(n22020), .Z(n22082) );
  XNOR U21938 ( .A(n16732), .B(p_input[657]), .Z(n22020) );
  XOR U21939 ( .A(n22084), .B(n22035), .Z(n22029) );
  XNOR U21940 ( .A(p_input[2079]), .B(p_input[671]), .Z(n22035) );
  XOR U21941 ( .A(n22026), .B(n22034), .Z(n22084) );
  XOR U21942 ( .A(n22085), .B(n22031), .Z(n22034) );
  XOR U21943 ( .A(p_input[2077]), .B(p_input[669]), .Z(n22031) );
  XNOR U21944 ( .A(p_input[2078]), .B(p_input[670]), .Z(n22085) );
  XNOR U21945 ( .A(n16448), .B(p_input[665]), .Z(n22026) );
  XNOR U21946 ( .A(n22047), .B(n22046), .Z(n22013) );
  XNOR U21947 ( .A(n22086), .B(n22053), .Z(n22046) );
  XNOR U21948 ( .A(n22042), .B(n22041), .Z(n22053) );
  XOR U21949 ( .A(n22087), .B(n22038), .Z(n22041) );
  XNOR U21950 ( .A(n16737), .B(p_input[651]), .Z(n22038) );
  XNOR U21951 ( .A(p_input[2060]), .B(p_input[652]), .Z(n22087) );
  XOR U21952 ( .A(p_input[2061]), .B(p_input[653]), .Z(n22042) );
  XNOR U21953 ( .A(n22052), .B(n22043), .Z(n22086) );
  XNOR U21954 ( .A(n16452), .B(p_input[642]), .Z(n22043) );
  XOR U21955 ( .A(n22088), .B(n22058), .Z(n22052) );
  XNOR U21956 ( .A(p_input[2064]), .B(p_input[656]), .Z(n22058) );
  XOR U21957 ( .A(n22049), .B(n22057), .Z(n22088) );
  XOR U21958 ( .A(n22089), .B(n22054), .Z(n22057) );
  XOR U21959 ( .A(p_input[2062]), .B(p_input[654]), .Z(n22054) );
  XNOR U21960 ( .A(p_input[2063]), .B(p_input[655]), .Z(n22089) );
  XNOR U21961 ( .A(n16740), .B(p_input[650]), .Z(n22049) );
  XNOR U21962 ( .A(n22064), .B(n22063), .Z(n22047) );
  XNOR U21963 ( .A(n22090), .B(n22069), .Z(n22063) );
  XOR U21964 ( .A(p_input[2057]), .B(p_input[649]), .Z(n22069) );
  XOR U21965 ( .A(n22060), .B(n22068), .Z(n22090) );
  XOR U21966 ( .A(n22091), .B(n22065), .Z(n22068) );
  XOR U21967 ( .A(p_input[2055]), .B(p_input[647]), .Z(n22065) );
  XNOR U21968 ( .A(p_input[2056]), .B(p_input[648]), .Z(n22091) );
  XNOR U21969 ( .A(n16459), .B(p_input[643]), .Z(n22060) );
  XNOR U21970 ( .A(n22074), .B(n22073), .Z(n22064) );
  XOR U21971 ( .A(n22092), .B(n22070), .Z(n22073) );
  XOR U21972 ( .A(p_input[2052]), .B(p_input[644]), .Z(n22070) );
  XNOR U21973 ( .A(p_input[2053]), .B(p_input[645]), .Z(n22092) );
  XOR U21974 ( .A(p_input[2054]), .B(p_input[646]), .Z(n22074) );
  XNOR U21975 ( .A(n22093), .B(n22094), .Z(n21891) );
  AND U21976 ( .A(n287), .B(n22095), .Z(n22094) );
  XNOR U21977 ( .A(n22096), .B(n22097), .Z(n287) );
  AND U21978 ( .A(n22098), .B(n22099), .Z(n22097) );
  XOR U21979 ( .A(n22096), .B(n21901), .Z(n22099) );
  XNOR U21980 ( .A(n22096), .B(n21843), .Z(n22098) );
  XOR U21981 ( .A(n22100), .B(n22101), .Z(n22096) );
  AND U21982 ( .A(n22102), .B(n22103), .Z(n22101) );
  XNOR U21983 ( .A(n21914), .B(n22100), .Z(n22103) );
  XOR U21984 ( .A(n22100), .B(n21855), .Z(n22102) );
  XOR U21985 ( .A(n22104), .B(n22105), .Z(n22100) );
  AND U21986 ( .A(n22106), .B(n22107), .Z(n22105) );
  XNOR U21987 ( .A(n21939), .B(n22104), .Z(n22107) );
  XOR U21988 ( .A(n22104), .B(n21866), .Z(n22106) );
  XOR U21989 ( .A(n22108), .B(n22109), .Z(n22104) );
  AND U21990 ( .A(n22110), .B(n22111), .Z(n22109) );
  XOR U21991 ( .A(n22108), .B(n21876), .Z(n22110) );
  XOR U21992 ( .A(n22112), .B(n22113), .Z(n21832) );
  AND U21993 ( .A(n291), .B(n22095), .Z(n22113) );
  XNOR U21994 ( .A(n22093), .B(n22112), .Z(n22095) );
  XNOR U21995 ( .A(n22114), .B(n22115), .Z(n291) );
  AND U21996 ( .A(n22116), .B(n22117), .Z(n22115) );
  XNOR U21997 ( .A(n22118), .B(n22114), .Z(n22117) );
  IV U21998 ( .A(n21901), .Z(n22118) );
  XNOR U21999 ( .A(n22119), .B(n22120), .Z(n21901) );
  AND U22000 ( .A(n294), .B(n22121), .Z(n22120) );
  XNOR U22001 ( .A(n22119), .B(n22122), .Z(n22121) );
  XNOR U22002 ( .A(n21843), .B(n22114), .Z(n22116) );
  XOR U22003 ( .A(n22123), .B(n22124), .Z(n21843) );
  AND U22004 ( .A(n302), .B(n22125), .Z(n22124) );
  XOR U22005 ( .A(n22126), .B(n22127), .Z(n22114) );
  AND U22006 ( .A(n22128), .B(n22129), .Z(n22127) );
  XNOR U22007 ( .A(n22126), .B(n21914), .Z(n22129) );
  XNOR U22008 ( .A(n22130), .B(n22131), .Z(n21914) );
  AND U22009 ( .A(n294), .B(n22132), .Z(n22131) );
  XOR U22010 ( .A(n22133), .B(n22130), .Z(n22132) );
  XNOR U22011 ( .A(n22134), .B(n22126), .Z(n22128) );
  IV U22012 ( .A(n21855), .Z(n22134) );
  XOR U22013 ( .A(n22135), .B(n22136), .Z(n21855) );
  AND U22014 ( .A(n302), .B(n22137), .Z(n22136) );
  XOR U22015 ( .A(n22138), .B(n22139), .Z(n22126) );
  AND U22016 ( .A(n22140), .B(n22141), .Z(n22139) );
  XNOR U22017 ( .A(n22138), .B(n21939), .Z(n22141) );
  XNOR U22018 ( .A(n22142), .B(n22143), .Z(n21939) );
  AND U22019 ( .A(n294), .B(n22144), .Z(n22143) );
  XNOR U22020 ( .A(n22145), .B(n22142), .Z(n22144) );
  XOR U22021 ( .A(n21866), .B(n22138), .Z(n22140) );
  XOR U22022 ( .A(n22146), .B(n22147), .Z(n21866) );
  AND U22023 ( .A(n302), .B(n22148), .Z(n22147) );
  XOR U22024 ( .A(n22108), .B(n22149), .Z(n22138) );
  AND U22025 ( .A(n22150), .B(n22111), .Z(n22149) );
  XNOR U22026 ( .A(n21985), .B(n22108), .Z(n22111) );
  XNOR U22027 ( .A(n22151), .B(n22152), .Z(n21985) );
  AND U22028 ( .A(n294), .B(n22153), .Z(n22152) );
  XOR U22029 ( .A(n22154), .B(n22151), .Z(n22153) );
  XNOR U22030 ( .A(n22155), .B(n22108), .Z(n22150) );
  IV U22031 ( .A(n21876), .Z(n22155) );
  XOR U22032 ( .A(n22156), .B(n22157), .Z(n21876) );
  AND U22033 ( .A(n302), .B(n22158), .Z(n22157) );
  XOR U22034 ( .A(n22159), .B(n22160), .Z(n22108) );
  AND U22035 ( .A(n22161), .B(n22162), .Z(n22160) );
  XNOR U22036 ( .A(n22159), .B(n22075), .Z(n22162) );
  XNOR U22037 ( .A(n22163), .B(n22164), .Z(n22075) );
  AND U22038 ( .A(n294), .B(n22165), .Z(n22164) );
  XNOR U22039 ( .A(n22166), .B(n22163), .Z(n22165) );
  XNOR U22040 ( .A(n22167), .B(n22159), .Z(n22161) );
  IV U22041 ( .A(n21888), .Z(n22167) );
  XOR U22042 ( .A(n22168), .B(n22169), .Z(n21888) );
  AND U22043 ( .A(n302), .B(n22170), .Z(n22169) );
  AND U22044 ( .A(n22112), .B(n22093), .Z(n22159) );
  XNOR U22045 ( .A(n22171), .B(n22172), .Z(n22093) );
  AND U22046 ( .A(n294), .B(n22173), .Z(n22172) );
  XNOR U22047 ( .A(n22174), .B(n22171), .Z(n22173) );
  XNOR U22048 ( .A(n22175), .B(n22176), .Z(n294) );
  AND U22049 ( .A(n22177), .B(n22178), .Z(n22176) );
  XOR U22050 ( .A(n22122), .B(n22175), .Z(n22178) );
  AND U22051 ( .A(n22179), .B(n22180), .Z(n22122) );
  XOR U22052 ( .A(n22175), .B(n22119), .Z(n22177) );
  XNOR U22053 ( .A(n22181), .B(n22182), .Z(n22119) );
  AND U22054 ( .A(n298), .B(n22125), .Z(n22182) );
  XOR U22055 ( .A(n22123), .B(n22181), .Z(n22125) );
  XOR U22056 ( .A(n22183), .B(n22184), .Z(n22175) );
  AND U22057 ( .A(n22185), .B(n22186), .Z(n22184) );
  XNOR U22058 ( .A(n22183), .B(n22179), .Z(n22186) );
  IV U22059 ( .A(n22133), .Z(n22179) );
  XOR U22060 ( .A(n22187), .B(n22188), .Z(n22133) );
  XOR U22061 ( .A(n22189), .B(n22180), .Z(n22188) );
  AND U22062 ( .A(n22145), .B(n22190), .Z(n22180) );
  AND U22063 ( .A(n22191), .B(n22192), .Z(n22189) );
  XOR U22064 ( .A(n22193), .B(n22187), .Z(n22191) );
  XNOR U22065 ( .A(n22130), .B(n22183), .Z(n22185) );
  XNOR U22066 ( .A(n22194), .B(n22195), .Z(n22130) );
  AND U22067 ( .A(n298), .B(n22137), .Z(n22195) );
  XOR U22068 ( .A(n22194), .B(n22135), .Z(n22137) );
  XOR U22069 ( .A(n22196), .B(n22197), .Z(n22183) );
  AND U22070 ( .A(n22198), .B(n22199), .Z(n22197) );
  XNOR U22071 ( .A(n22196), .B(n22145), .Z(n22199) );
  XOR U22072 ( .A(n22200), .B(n22192), .Z(n22145) );
  XNOR U22073 ( .A(n22201), .B(n22187), .Z(n22192) );
  XOR U22074 ( .A(n22202), .B(n22203), .Z(n22187) );
  AND U22075 ( .A(n22204), .B(n22205), .Z(n22203) );
  XOR U22076 ( .A(n22206), .B(n22202), .Z(n22204) );
  XNOR U22077 ( .A(n22207), .B(n22208), .Z(n22201) );
  AND U22078 ( .A(n22209), .B(n22210), .Z(n22208) );
  XOR U22079 ( .A(n22207), .B(n22211), .Z(n22209) );
  XNOR U22080 ( .A(n22193), .B(n22190), .Z(n22200) );
  AND U22081 ( .A(n22212), .B(n22213), .Z(n22190) );
  XOR U22082 ( .A(n22214), .B(n22215), .Z(n22193) );
  AND U22083 ( .A(n22216), .B(n22217), .Z(n22215) );
  XOR U22084 ( .A(n22214), .B(n22218), .Z(n22216) );
  XNOR U22085 ( .A(n22142), .B(n22196), .Z(n22198) );
  XNOR U22086 ( .A(n22219), .B(n22220), .Z(n22142) );
  AND U22087 ( .A(n298), .B(n22148), .Z(n22220) );
  XOR U22088 ( .A(n22219), .B(n22146), .Z(n22148) );
  XOR U22089 ( .A(n22221), .B(n22222), .Z(n22196) );
  AND U22090 ( .A(n22223), .B(n22224), .Z(n22222) );
  XNOR U22091 ( .A(n22221), .B(n22212), .Z(n22224) );
  IV U22092 ( .A(n22154), .Z(n22212) );
  XNOR U22093 ( .A(n22225), .B(n22205), .Z(n22154) );
  XNOR U22094 ( .A(n22226), .B(n22211), .Z(n22205) );
  XOR U22095 ( .A(n22227), .B(n22228), .Z(n22211) );
  AND U22096 ( .A(n22229), .B(n22230), .Z(n22228) );
  XOR U22097 ( .A(n22227), .B(n22231), .Z(n22229) );
  XNOR U22098 ( .A(n22210), .B(n22202), .Z(n22226) );
  XOR U22099 ( .A(n22232), .B(n22233), .Z(n22202) );
  AND U22100 ( .A(n22234), .B(n22235), .Z(n22233) );
  XNOR U22101 ( .A(n22236), .B(n22232), .Z(n22234) );
  XNOR U22102 ( .A(n22237), .B(n22207), .Z(n22210) );
  XOR U22103 ( .A(n22238), .B(n22239), .Z(n22207) );
  AND U22104 ( .A(n22240), .B(n22241), .Z(n22239) );
  XOR U22105 ( .A(n22238), .B(n22242), .Z(n22240) );
  XNOR U22106 ( .A(n22243), .B(n22244), .Z(n22237) );
  AND U22107 ( .A(n22245), .B(n22246), .Z(n22244) );
  XNOR U22108 ( .A(n22243), .B(n22247), .Z(n22245) );
  XNOR U22109 ( .A(n22206), .B(n22213), .Z(n22225) );
  AND U22110 ( .A(n22166), .B(n22248), .Z(n22213) );
  XOR U22111 ( .A(n22218), .B(n22217), .Z(n22206) );
  XNOR U22112 ( .A(n22249), .B(n22214), .Z(n22217) );
  XOR U22113 ( .A(n22250), .B(n22251), .Z(n22214) );
  AND U22114 ( .A(n22252), .B(n22253), .Z(n22251) );
  XOR U22115 ( .A(n22250), .B(n22254), .Z(n22252) );
  XNOR U22116 ( .A(n22255), .B(n22256), .Z(n22249) );
  AND U22117 ( .A(n22257), .B(n22258), .Z(n22256) );
  XOR U22118 ( .A(n22255), .B(n22259), .Z(n22257) );
  XOR U22119 ( .A(n22260), .B(n22261), .Z(n22218) );
  AND U22120 ( .A(n22262), .B(n22263), .Z(n22261) );
  XOR U22121 ( .A(n22260), .B(n22264), .Z(n22262) );
  XNOR U22122 ( .A(n22151), .B(n22221), .Z(n22223) );
  XNOR U22123 ( .A(n22265), .B(n22266), .Z(n22151) );
  AND U22124 ( .A(n298), .B(n22158), .Z(n22266) );
  XOR U22125 ( .A(n22265), .B(n22156), .Z(n22158) );
  XOR U22126 ( .A(n22267), .B(n22268), .Z(n22221) );
  AND U22127 ( .A(n22269), .B(n22270), .Z(n22268) );
  XNOR U22128 ( .A(n22267), .B(n22166), .Z(n22270) );
  XOR U22129 ( .A(n22271), .B(n22235), .Z(n22166) );
  XNOR U22130 ( .A(n22272), .B(n22242), .Z(n22235) );
  XOR U22131 ( .A(n22231), .B(n22230), .Z(n22242) );
  XNOR U22132 ( .A(n22273), .B(n22227), .Z(n22230) );
  XOR U22133 ( .A(n22274), .B(n22275), .Z(n22227) );
  AND U22134 ( .A(n22276), .B(n22277), .Z(n22275) );
  XOR U22135 ( .A(n22274), .B(n22278), .Z(n22276) );
  XNOR U22136 ( .A(n22279), .B(n22280), .Z(n22273) );
  NOR U22137 ( .A(n22281), .B(n22282), .Z(n22280) );
  XNOR U22138 ( .A(n22279), .B(n22283), .Z(n22281) );
  XOR U22139 ( .A(n22284), .B(n22285), .Z(n22231) );
  NOR U22140 ( .A(n22286), .B(n22287), .Z(n22285) );
  XNOR U22141 ( .A(n22284), .B(n22288), .Z(n22286) );
  XNOR U22142 ( .A(n22241), .B(n22232), .Z(n22272) );
  XOR U22143 ( .A(n22289), .B(n22290), .Z(n22232) );
  NOR U22144 ( .A(n22291), .B(n22292), .Z(n22290) );
  XNOR U22145 ( .A(n22289), .B(n22293), .Z(n22291) );
  XOR U22146 ( .A(n22294), .B(n22247), .Z(n22241) );
  XNOR U22147 ( .A(n22295), .B(n22296), .Z(n22247) );
  NOR U22148 ( .A(n22297), .B(n22298), .Z(n22296) );
  XNOR U22149 ( .A(n22295), .B(n22299), .Z(n22297) );
  XNOR U22150 ( .A(n22246), .B(n22238), .Z(n22294) );
  XOR U22151 ( .A(n22300), .B(n22301), .Z(n22238) );
  AND U22152 ( .A(n22302), .B(n22303), .Z(n22301) );
  XOR U22153 ( .A(n22300), .B(n22304), .Z(n22302) );
  XNOR U22154 ( .A(n22305), .B(n22243), .Z(n22246) );
  XOR U22155 ( .A(n22306), .B(n22307), .Z(n22243) );
  AND U22156 ( .A(n22308), .B(n22309), .Z(n22307) );
  XOR U22157 ( .A(n22306), .B(n22310), .Z(n22308) );
  XNOR U22158 ( .A(n22311), .B(n22312), .Z(n22305) );
  NOR U22159 ( .A(n22313), .B(n22314), .Z(n22312) );
  XOR U22160 ( .A(n22311), .B(n22315), .Z(n22313) );
  XOR U22161 ( .A(n22236), .B(n22248), .Z(n22271) );
  NOR U22162 ( .A(n22174), .B(n22316), .Z(n22248) );
  XNOR U22163 ( .A(n22254), .B(n22253), .Z(n22236) );
  XNOR U22164 ( .A(n22317), .B(n22259), .Z(n22253) );
  XOR U22165 ( .A(n22318), .B(n22319), .Z(n22259) );
  NOR U22166 ( .A(n22320), .B(n22321), .Z(n22319) );
  XNOR U22167 ( .A(n22318), .B(n22322), .Z(n22320) );
  XNOR U22168 ( .A(n22258), .B(n22250), .Z(n22317) );
  XOR U22169 ( .A(n22323), .B(n22324), .Z(n22250) );
  AND U22170 ( .A(n22325), .B(n22326), .Z(n22324) );
  XNOR U22171 ( .A(n22323), .B(n22327), .Z(n22325) );
  XNOR U22172 ( .A(n22328), .B(n22255), .Z(n22258) );
  XOR U22173 ( .A(n22329), .B(n22330), .Z(n22255) );
  AND U22174 ( .A(n22331), .B(n22332), .Z(n22330) );
  XOR U22175 ( .A(n22329), .B(n22333), .Z(n22331) );
  XNOR U22176 ( .A(n22334), .B(n22335), .Z(n22328) );
  NOR U22177 ( .A(n22336), .B(n22337), .Z(n22335) );
  XOR U22178 ( .A(n22334), .B(n22338), .Z(n22336) );
  XOR U22179 ( .A(n22264), .B(n22263), .Z(n22254) );
  XNOR U22180 ( .A(n22339), .B(n22260), .Z(n22263) );
  XOR U22181 ( .A(n22340), .B(n22341), .Z(n22260) );
  AND U22182 ( .A(n22342), .B(n22343), .Z(n22341) );
  XOR U22183 ( .A(n22340), .B(n22344), .Z(n22342) );
  XNOR U22184 ( .A(n22345), .B(n22346), .Z(n22339) );
  NOR U22185 ( .A(n22347), .B(n22348), .Z(n22346) );
  XNOR U22186 ( .A(n22345), .B(n22349), .Z(n22347) );
  XOR U22187 ( .A(n22350), .B(n22351), .Z(n22264) );
  NOR U22188 ( .A(n22352), .B(n22353), .Z(n22351) );
  XNOR U22189 ( .A(n22350), .B(n22354), .Z(n22352) );
  XNOR U22190 ( .A(n22163), .B(n22267), .Z(n22269) );
  XNOR U22191 ( .A(n22355), .B(n22356), .Z(n22163) );
  AND U22192 ( .A(n298), .B(n22170), .Z(n22356) );
  XOR U22193 ( .A(n22355), .B(n22168), .Z(n22170) );
  AND U22194 ( .A(n22171), .B(n22174), .Z(n22267) );
  XOR U22195 ( .A(n22357), .B(n22316), .Z(n22174) );
  XNOR U22196 ( .A(p_input[2048]), .B(p_input[672]), .Z(n22316) );
  XOR U22197 ( .A(n22293), .B(n22292), .Z(n22357) );
  XOR U22198 ( .A(n22358), .B(n22304), .Z(n22292) );
  XOR U22199 ( .A(n22278), .B(n22277), .Z(n22304) );
  XNOR U22200 ( .A(n22359), .B(n22283), .Z(n22277) );
  XOR U22201 ( .A(p_input[2072]), .B(p_input[696]), .Z(n22283) );
  XOR U22202 ( .A(n22274), .B(n22282), .Z(n22359) );
  XOR U22203 ( .A(n22360), .B(n22279), .Z(n22282) );
  XOR U22204 ( .A(p_input[2070]), .B(p_input[694]), .Z(n22279) );
  XNOR U22205 ( .A(p_input[2071]), .B(p_input[695]), .Z(n22360) );
  XNOR U22206 ( .A(n16727), .B(p_input[690]), .Z(n22274) );
  XNOR U22207 ( .A(n22288), .B(n22287), .Z(n22278) );
  XOR U22208 ( .A(n22361), .B(n22284), .Z(n22287) );
  XOR U22209 ( .A(p_input[2067]), .B(p_input[691]), .Z(n22284) );
  XNOR U22210 ( .A(p_input[2068]), .B(p_input[692]), .Z(n22361) );
  XOR U22211 ( .A(p_input[2069]), .B(p_input[693]), .Z(n22288) );
  XNOR U22212 ( .A(n22303), .B(n22289), .Z(n22358) );
  XNOR U22213 ( .A(n16729), .B(p_input[673]), .Z(n22289) );
  XNOR U22214 ( .A(n22362), .B(n22310), .Z(n22303) );
  XNOR U22215 ( .A(n22299), .B(n22298), .Z(n22310) );
  XOR U22216 ( .A(n22363), .B(n22295), .Z(n22298) );
  XNOR U22217 ( .A(n16444), .B(p_input[698]), .Z(n22295) );
  XNOR U22218 ( .A(p_input[2075]), .B(p_input[699]), .Z(n22363) );
  XOR U22219 ( .A(p_input[2076]), .B(p_input[700]), .Z(n22299) );
  XNOR U22220 ( .A(n22309), .B(n22300), .Z(n22362) );
  XNOR U22221 ( .A(n16732), .B(p_input[689]), .Z(n22300) );
  XOR U22222 ( .A(n22364), .B(n22315), .Z(n22309) );
  XNOR U22223 ( .A(p_input[2079]), .B(p_input[703]), .Z(n22315) );
  XOR U22224 ( .A(n22306), .B(n22314), .Z(n22364) );
  XOR U22225 ( .A(n22365), .B(n22311), .Z(n22314) );
  XOR U22226 ( .A(p_input[2077]), .B(p_input[701]), .Z(n22311) );
  XNOR U22227 ( .A(p_input[2078]), .B(p_input[702]), .Z(n22365) );
  XNOR U22228 ( .A(n16448), .B(p_input[697]), .Z(n22306) );
  XNOR U22229 ( .A(n22327), .B(n22326), .Z(n22293) );
  XNOR U22230 ( .A(n22366), .B(n22333), .Z(n22326) );
  XNOR U22231 ( .A(n22322), .B(n22321), .Z(n22333) );
  XOR U22232 ( .A(n22367), .B(n22318), .Z(n22321) );
  XNOR U22233 ( .A(n16737), .B(p_input[683]), .Z(n22318) );
  XNOR U22234 ( .A(p_input[2060]), .B(p_input[684]), .Z(n22367) );
  XOR U22235 ( .A(p_input[2061]), .B(p_input[685]), .Z(n22322) );
  XNOR U22236 ( .A(n22332), .B(n22323), .Z(n22366) );
  XNOR U22237 ( .A(n16452), .B(p_input[674]), .Z(n22323) );
  XOR U22238 ( .A(n22368), .B(n22338), .Z(n22332) );
  XNOR U22239 ( .A(p_input[2064]), .B(p_input[688]), .Z(n22338) );
  XOR U22240 ( .A(n22329), .B(n22337), .Z(n22368) );
  XOR U22241 ( .A(n22369), .B(n22334), .Z(n22337) );
  XOR U22242 ( .A(p_input[2062]), .B(p_input[686]), .Z(n22334) );
  XNOR U22243 ( .A(p_input[2063]), .B(p_input[687]), .Z(n22369) );
  XNOR U22244 ( .A(n16740), .B(p_input[682]), .Z(n22329) );
  XNOR U22245 ( .A(n22344), .B(n22343), .Z(n22327) );
  XNOR U22246 ( .A(n22370), .B(n22349), .Z(n22343) );
  XOR U22247 ( .A(p_input[2057]), .B(p_input[681]), .Z(n22349) );
  XOR U22248 ( .A(n22340), .B(n22348), .Z(n22370) );
  XOR U22249 ( .A(n22371), .B(n22345), .Z(n22348) );
  XOR U22250 ( .A(p_input[2055]), .B(p_input[679]), .Z(n22345) );
  XNOR U22251 ( .A(p_input[2056]), .B(p_input[680]), .Z(n22371) );
  XNOR U22252 ( .A(n16459), .B(p_input[675]), .Z(n22340) );
  XNOR U22253 ( .A(n22354), .B(n22353), .Z(n22344) );
  XOR U22254 ( .A(n22372), .B(n22350), .Z(n22353) );
  XOR U22255 ( .A(p_input[2052]), .B(p_input[676]), .Z(n22350) );
  XNOR U22256 ( .A(p_input[2053]), .B(p_input[677]), .Z(n22372) );
  XOR U22257 ( .A(p_input[2054]), .B(p_input[678]), .Z(n22354) );
  XNOR U22258 ( .A(n22373), .B(n22374), .Z(n22171) );
  AND U22259 ( .A(n298), .B(n22375), .Z(n22374) );
  XNOR U22260 ( .A(n22376), .B(n22377), .Z(n298) );
  AND U22261 ( .A(n22378), .B(n22379), .Z(n22377) );
  XOR U22262 ( .A(n22376), .B(n22181), .Z(n22379) );
  XNOR U22263 ( .A(n22376), .B(n22123), .Z(n22378) );
  XOR U22264 ( .A(n22380), .B(n22381), .Z(n22376) );
  AND U22265 ( .A(n22382), .B(n22383), .Z(n22381) );
  XNOR U22266 ( .A(n22194), .B(n22380), .Z(n22383) );
  XOR U22267 ( .A(n22380), .B(n22135), .Z(n22382) );
  XOR U22268 ( .A(n22384), .B(n22385), .Z(n22380) );
  AND U22269 ( .A(n22386), .B(n22387), .Z(n22385) );
  XNOR U22270 ( .A(n22219), .B(n22384), .Z(n22387) );
  XOR U22271 ( .A(n22384), .B(n22146), .Z(n22386) );
  XOR U22272 ( .A(n22388), .B(n22389), .Z(n22384) );
  AND U22273 ( .A(n22390), .B(n22391), .Z(n22389) );
  XOR U22274 ( .A(n22388), .B(n22156), .Z(n22390) );
  XOR U22275 ( .A(n22392), .B(n22393), .Z(n22112) );
  AND U22276 ( .A(n302), .B(n22375), .Z(n22393) );
  XNOR U22277 ( .A(n22373), .B(n22392), .Z(n22375) );
  XNOR U22278 ( .A(n22394), .B(n22395), .Z(n302) );
  AND U22279 ( .A(n22396), .B(n22397), .Z(n22395) );
  XNOR U22280 ( .A(n22398), .B(n22394), .Z(n22397) );
  IV U22281 ( .A(n22181), .Z(n22398) );
  XNOR U22282 ( .A(n22399), .B(n22400), .Z(n22181) );
  AND U22283 ( .A(n305), .B(n22401), .Z(n22400) );
  XNOR U22284 ( .A(n22399), .B(n22402), .Z(n22401) );
  XNOR U22285 ( .A(n22123), .B(n22394), .Z(n22396) );
  XOR U22286 ( .A(n22403), .B(n22404), .Z(n22123) );
  AND U22287 ( .A(n313), .B(n22405), .Z(n22404) );
  XOR U22288 ( .A(n22406), .B(n22407), .Z(n22394) );
  AND U22289 ( .A(n22408), .B(n22409), .Z(n22407) );
  XNOR U22290 ( .A(n22406), .B(n22194), .Z(n22409) );
  XNOR U22291 ( .A(n22410), .B(n22411), .Z(n22194) );
  AND U22292 ( .A(n305), .B(n22412), .Z(n22411) );
  XOR U22293 ( .A(n22413), .B(n22410), .Z(n22412) );
  XNOR U22294 ( .A(n22414), .B(n22406), .Z(n22408) );
  IV U22295 ( .A(n22135), .Z(n22414) );
  XOR U22296 ( .A(n22415), .B(n22416), .Z(n22135) );
  AND U22297 ( .A(n313), .B(n22417), .Z(n22416) );
  XOR U22298 ( .A(n22418), .B(n22419), .Z(n22406) );
  AND U22299 ( .A(n22420), .B(n22421), .Z(n22419) );
  XNOR U22300 ( .A(n22418), .B(n22219), .Z(n22421) );
  XNOR U22301 ( .A(n22422), .B(n22423), .Z(n22219) );
  AND U22302 ( .A(n305), .B(n22424), .Z(n22423) );
  XNOR U22303 ( .A(n22425), .B(n22422), .Z(n22424) );
  XOR U22304 ( .A(n22146), .B(n22418), .Z(n22420) );
  XOR U22305 ( .A(n22426), .B(n22427), .Z(n22146) );
  AND U22306 ( .A(n313), .B(n22428), .Z(n22427) );
  XOR U22307 ( .A(n22388), .B(n22429), .Z(n22418) );
  AND U22308 ( .A(n22430), .B(n22391), .Z(n22429) );
  XNOR U22309 ( .A(n22265), .B(n22388), .Z(n22391) );
  XNOR U22310 ( .A(n22431), .B(n22432), .Z(n22265) );
  AND U22311 ( .A(n305), .B(n22433), .Z(n22432) );
  XOR U22312 ( .A(n22434), .B(n22431), .Z(n22433) );
  XNOR U22313 ( .A(n22435), .B(n22388), .Z(n22430) );
  IV U22314 ( .A(n22156), .Z(n22435) );
  XOR U22315 ( .A(n22436), .B(n22437), .Z(n22156) );
  AND U22316 ( .A(n313), .B(n22438), .Z(n22437) );
  XOR U22317 ( .A(n22439), .B(n22440), .Z(n22388) );
  AND U22318 ( .A(n22441), .B(n22442), .Z(n22440) );
  XNOR U22319 ( .A(n22439), .B(n22355), .Z(n22442) );
  XNOR U22320 ( .A(n22443), .B(n22444), .Z(n22355) );
  AND U22321 ( .A(n305), .B(n22445), .Z(n22444) );
  XNOR U22322 ( .A(n22446), .B(n22443), .Z(n22445) );
  XNOR U22323 ( .A(n22447), .B(n22439), .Z(n22441) );
  IV U22324 ( .A(n22168), .Z(n22447) );
  XOR U22325 ( .A(n22448), .B(n22449), .Z(n22168) );
  AND U22326 ( .A(n313), .B(n22450), .Z(n22449) );
  AND U22327 ( .A(n22392), .B(n22373), .Z(n22439) );
  XNOR U22328 ( .A(n22451), .B(n22452), .Z(n22373) );
  AND U22329 ( .A(n305), .B(n22453), .Z(n22452) );
  XNOR U22330 ( .A(n22454), .B(n22451), .Z(n22453) );
  XNOR U22331 ( .A(n22455), .B(n22456), .Z(n305) );
  AND U22332 ( .A(n22457), .B(n22458), .Z(n22456) );
  XOR U22333 ( .A(n22402), .B(n22455), .Z(n22458) );
  AND U22334 ( .A(n22459), .B(n22460), .Z(n22402) );
  XOR U22335 ( .A(n22455), .B(n22399), .Z(n22457) );
  XNOR U22336 ( .A(n22461), .B(n22462), .Z(n22399) );
  AND U22337 ( .A(n309), .B(n22405), .Z(n22462) );
  XOR U22338 ( .A(n22403), .B(n22461), .Z(n22405) );
  XOR U22339 ( .A(n22463), .B(n22464), .Z(n22455) );
  AND U22340 ( .A(n22465), .B(n22466), .Z(n22464) );
  XNOR U22341 ( .A(n22463), .B(n22459), .Z(n22466) );
  IV U22342 ( .A(n22413), .Z(n22459) );
  XOR U22343 ( .A(n22467), .B(n22468), .Z(n22413) );
  XOR U22344 ( .A(n22469), .B(n22460), .Z(n22468) );
  AND U22345 ( .A(n22425), .B(n22470), .Z(n22460) );
  AND U22346 ( .A(n22471), .B(n22472), .Z(n22469) );
  XOR U22347 ( .A(n22473), .B(n22467), .Z(n22471) );
  XNOR U22348 ( .A(n22410), .B(n22463), .Z(n22465) );
  XNOR U22349 ( .A(n22474), .B(n22475), .Z(n22410) );
  AND U22350 ( .A(n309), .B(n22417), .Z(n22475) );
  XOR U22351 ( .A(n22474), .B(n22415), .Z(n22417) );
  XOR U22352 ( .A(n22476), .B(n22477), .Z(n22463) );
  AND U22353 ( .A(n22478), .B(n22479), .Z(n22477) );
  XNOR U22354 ( .A(n22476), .B(n22425), .Z(n22479) );
  XOR U22355 ( .A(n22480), .B(n22472), .Z(n22425) );
  XNOR U22356 ( .A(n22481), .B(n22467), .Z(n22472) );
  XOR U22357 ( .A(n22482), .B(n22483), .Z(n22467) );
  AND U22358 ( .A(n22484), .B(n22485), .Z(n22483) );
  XOR U22359 ( .A(n22486), .B(n22482), .Z(n22484) );
  XNOR U22360 ( .A(n22487), .B(n22488), .Z(n22481) );
  AND U22361 ( .A(n22489), .B(n22490), .Z(n22488) );
  XOR U22362 ( .A(n22487), .B(n22491), .Z(n22489) );
  XNOR U22363 ( .A(n22473), .B(n22470), .Z(n22480) );
  AND U22364 ( .A(n22492), .B(n22493), .Z(n22470) );
  XOR U22365 ( .A(n22494), .B(n22495), .Z(n22473) );
  AND U22366 ( .A(n22496), .B(n22497), .Z(n22495) );
  XOR U22367 ( .A(n22494), .B(n22498), .Z(n22496) );
  XNOR U22368 ( .A(n22422), .B(n22476), .Z(n22478) );
  XNOR U22369 ( .A(n22499), .B(n22500), .Z(n22422) );
  AND U22370 ( .A(n309), .B(n22428), .Z(n22500) );
  XOR U22371 ( .A(n22499), .B(n22426), .Z(n22428) );
  XOR U22372 ( .A(n22501), .B(n22502), .Z(n22476) );
  AND U22373 ( .A(n22503), .B(n22504), .Z(n22502) );
  XNOR U22374 ( .A(n22501), .B(n22492), .Z(n22504) );
  IV U22375 ( .A(n22434), .Z(n22492) );
  XNOR U22376 ( .A(n22505), .B(n22485), .Z(n22434) );
  XNOR U22377 ( .A(n22506), .B(n22491), .Z(n22485) );
  XOR U22378 ( .A(n22507), .B(n22508), .Z(n22491) );
  AND U22379 ( .A(n22509), .B(n22510), .Z(n22508) );
  XOR U22380 ( .A(n22507), .B(n22511), .Z(n22509) );
  XNOR U22381 ( .A(n22490), .B(n22482), .Z(n22506) );
  XOR U22382 ( .A(n22512), .B(n22513), .Z(n22482) );
  AND U22383 ( .A(n22514), .B(n22515), .Z(n22513) );
  XNOR U22384 ( .A(n22516), .B(n22512), .Z(n22514) );
  XNOR U22385 ( .A(n22517), .B(n22487), .Z(n22490) );
  XOR U22386 ( .A(n22518), .B(n22519), .Z(n22487) );
  AND U22387 ( .A(n22520), .B(n22521), .Z(n22519) );
  XOR U22388 ( .A(n22518), .B(n22522), .Z(n22520) );
  XNOR U22389 ( .A(n22523), .B(n22524), .Z(n22517) );
  AND U22390 ( .A(n22525), .B(n22526), .Z(n22524) );
  XNOR U22391 ( .A(n22523), .B(n22527), .Z(n22525) );
  XNOR U22392 ( .A(n22486), .B(n22493), .Z(n22505) );
  AND U22393 ( .A(n22446), .B(n22528), .Z(n22493) );
  XOR U22394 ( .A(n22498), .B(n22497), .Z(n22486) );
  XNOR U22395 ( .A(n22529), .B(n22494), .Z(n22497) );
  XOR U22396 ( .A(n22530), .B(n22531), .Z(n22494) );
  AND U22397 ( .A(n22532), .B(n22533), .Z(n22531) );
  XOR U22398 ( .A(n22530), .B(n22534), .Z(n22532) );
  XNOR U22399 ( .A(n22535), .B(n22536), .Z(n22529) );
  AND U22400 ( .A(n22537), .B(n22538), .Z(n22536) );
  XOR U22401 ( .A(n22535), .B(n22539), .Z(n22537) );
  XOR U22402 ( .A(n22540), .B(n22541), .Z(n22498) );
  AND U22403 ( .A(n22542), .B(n22543), .Z(n22541) );
  XOR U22404 ( .A(n22540), .B(n22544), .Z(n22542) );
  XNOR U22405 ( .A(n22431), .B(n22501), .Z(n22503) );
  XNOR U22406 ( .A(n22545), .B(n22546), .Z(n22431) );
  AND U22407 ( .A(n309), .B(n22438), .Z(n22546) );
  XOR U22408 ( .A(n22545), .B(n22436), .Z(n22438) );
  XOR U22409 ( .A(n22547), .B(n22548), .Z(n22501) );
  AND U22410 ( .A(n22549), .B(n22550), .Z(n22548) );
  XNOR U22411 ( .A(n22547), .B(n22446), .Z(n22550) );
  XOR U22412 ( .A(n22551), .B(n22515), .Z(n22446) );
  XNOR U22413 ( .A(n22552), .B(n22522), .Z(n22515) );
  XOR U22414 ( .A(n22511), .B(n22510), .Z(n22522) );
  XNOR U22415 ( .A(n22553), .B(n22507), .Z(n22510) );
  XOR U22416 ( .A(n22554), .B(n22555), .Z(n22507) );
  AND U22417 ( .A(n22556), .B(n22557), .Z(n22555) );
  XOR U22418 ( .A(n22554), .B(n22558), .Z(n22556) );
  XNOR U22419 ( .A(n22559), .B(n22560), .Z(n22553) );
  NOR U22420 ( .A(n22561), .B(n22562), .Z(n22560) );
  XNOR U22421 ( .A(n22559), .B(n22563), .Z(n22561) );
  XOR U22422 ( .A(n22564), .B(n22565), .Z(n22511) );
  NOR U22423 ( .A(n22566), .B(n22567), .Z(n22565) );
  XNOR U22424 ( .A(n22564), .B(n22568), .Z(n22566) );
  XNOR U22425 ( .A(n22521), .B(n22512), .Z(n22552) );
  XOR U22426 ( .A(n22569), .B(n22570), .Z(n22512) );
  NOR U22427 ( .A(n22571), .B(n22572), .Z(n22570) );
  XNOR U22428 ( .A(n22569), .B(n22573), .Z(n22571) );
  XOR U22429 ( .A(n22574), .B(n22527), .Z(n22521) );
  XNOR U22430 ( .A(n22575), .B(n22576), .Z(n22527) );
  NOR U22431 ( .A(n22577), .B(n22578), .Z(n22576) );
  XNOR U22432 ( .A(n22575), .B(n22579), .Z(n22577) );
  XNOR U22433 ( .A(n22526), .B(n22518), .Z(n22574) );
  XOR U22434 ( .A(n22580), .B(n22581), .Z(n22518) );
  AND U22435 ( .A(n22582), .B(n22583), .Z(n22581) );
  XOR U22436 ( .A(n22580), .B(n22584), .Z(n22582) );
  XNOR U22437 ( .A(n22585), .B(n22523), .Z(n22526) );
  XOR U22438 ( .A(n22586), .B(n22587), .Z(n22523) );
  AND U22439 ( .A(n22588), .B(n22589), .Z(n22587) );
  XOR U22440 ( .A(n22586), .B(n22590), .Z(n22588) );
  XNOR U22441 ( .A(n22591), .B(n22592), .Z(n22585) );
  NOR U22442 ( .A(n22593), .B(n22594), .Z(n22592) );
  XOR U22443 ( .A(n22591), .B(n22595), .Z(n22593) );
  XOR U22444 ( .A(n22516), .B(n22528), .Z(n22551) );
  NOR U22445 ( .A(n22454), .B(n22596), .Z(n22528) );
  XNOR U22446 ( .A(n22534), .B(n22533), .Z(n22516) );
  XNOR U22447 ( .A(n22597), .B(n22539), .Z(n22533) );
  XOR U22448 ( .A(n22598), .B(n22599), .Z(n22539) );
  NOR U22449 ( .A(n22600), .B(n22601), .Z(n22599) );
  XNOR U22450 ( .A(n22598), .B(n22602), .Z(n22600) );
  XNOR U22451 ( .A(n22538), .B(n22530), .Z(n22597) );
  XOR U22452 ( .A(n22603), .B(n22604), .Z(n22530) );
  AND U22453 ( .A(n22605), .B(n22606), .Z(n22604) );
  XNOR U22454 ( .A(n22603), .B(n22607), .Z(n22605) );
  XNOR U22455 ( .A(n22608), .B(n22535), .Z(n22538) );
  XOR U22456 ( .A(n22609), .B(n22610), .Z(n22535) );
  AND U22457 ( .A(n22611), .B(n22612), .Z(n22610) );
  XOR U22458 ( .A(n22609), .B(n22613), .Z(n22611) );
  XNOR U22459 ( .A(n22614), .B(n22615), .Z(n22608) );
  NOR U22460 ( .A(n22616), .B(n22617), .Z(n22615) );
  XOR U22461 ( .A(n22614), .B(n22618), .Z(n22616) );
  XOR U22462 ( .A(n22544), .B(n22543), .Z(n22534) );
  XNOR U22463 ( .A(n22619), .B(n22540), .Z(n22543) );
  XOR U22464 ( .A(n22620), .B(n22621), .Z(n22540) );
  AND U22465 ( .A(n22622), .B(n22623), .Z(n22621) );
  XOR U22466 ( .A(n22620), .B(n22624), .Z(n22622) );
  XNOR U22467 ( .A(n22625), .B(n22626), .Z(n22619) );
  NOR U22468 ( .A(n22627), .B(n22628), .Z(n22626) );
  XNOR U22469 ( .A(n22625), .B(n22629), .Z(n22627) );
  XOR U22470 ( .A(n22630), .B(n22631), .Z(n22544) );
  NOR U22471 ( .A(n22632), .B(n22633), .Z(n22631) );
  XNOR U22472 ( .A(n22630), .B(n22634), .Z(n22632) );
  XNOR U22473 ( .A(n22443), .B(n22547), .Z(n22549) );
  XNOR U22474 ( .A(n22635), .B(n22636), .Z(n22443) );
  AND U22475 ( .A(n309), .B(n22450), .Z(n22636) );
  XOR U22476 ( .A(n22635), .B(n22448), .Z(n22450) );
  AND U22477 ( .A(n22451), .B(n22454), .Z(n22547) );
  XOR U22478 ( .A(n22637), .B(n22596), .Z(n22454) );
  XNOR U22479 ( .A(p_input[2048]), .B(p_input[704]), .Z(n22596) );
  XOR U22480 ( .A(n22573), .B(n22572), .Z(n22637) );
  XOR U22481 ( .A(n22638), .B(n22584), .Z(n22572) );
  XOR U22482 ( .A(n22558), .B(n22557), .Z(n22584) );
  XNOR U22483 ( .A(n22639), .B(n22563), .Z(n22557) );
  XOR U22484 ( .A(p_input[2072]), .B(p_input[728]), .Z(n22563) );
  XOR U22485 ( .A(n22554), .B(n22562), .Z(n22639) );
  XOR U22486 ( .A(n22640), .B(n22559), .Z(n22562) );
  XOR U22487 ( .A(p_input[2070]), .B(p_input[726]), .Z(n22559) );
  XNOR U22488 ( .A(p_input[2071]), .B(p_input[727]), .Z(n22640) );
  XNOR U22489 ( .A(n16727), .B(p_input[722]), .Z(n22554) );
  XNOR U22490 ( .A(n22568), .B(n22567), .Z(n22558) );
  XOR U22491 ( .A(n22641), .B(n22564), .Z(n22567) );
  XOR U22492 ( .A(p_input[2067]), .B(p_input[723]), .Z(n22564) );
  XNOR U22493 ( .A(p_input[2068]), .B(p_input[724]), .Z(n22641) );
  XOR U22494 ( .A(p_input[2069]), .B(p_input[725]), .Z(n22568) );
  XNOR U22495 ( .A(n22583), .B(n22569), .Z(n22638) );
  XNOR U22496 ( .A(n16729), .B(p_input[705]), .Z(n22569) );
  XNOR U22497 ( .A(n22642), .B(n22590), .Z(n22583) );
  XNOR U22498 ( .A(n22579), .B(n22578), .Z(n22590) );
  XOR U22499 ( .A(n22643), .B(n22575), .Z(n22578) );
  XNOR U22500 ( .A(n16444), .B(p_input[730]), .Z(n22575) );
  XNOR U22501 ( .A(p_input[2075]), .B(p_input[731]), .Z(n22643) );
  XOR U22502 ( .A(p_input[2076]), .B(p_input[732]), .Z(n22579) );
  XNOR U22503 ( .A(n22589), .B(n22580), .Z(n22642) );
  XNOR U22504 ( .A(n16732), .B(p_input[721]), .Z(n22580) );
  XOR U22505 ( .A(n22644), .B(n22595), .Z(n22589) );
  XNOR U22506 ( .A(p_input[2079]), .B(p_input[735]), .Z(n22595) );
  XOR U22507 ( .A(n22586), .B(n22594), .Z(n22644) );
  XOR U22508 ( .A(n22645), .B(n22591), .Z(n22594) );
  XOR U22509 ( .A(p_input[2077]), .B(p_input[733]), .Z(n22591) );
  XNOR U22510 ( .A(p_input[2078]), .B(p_input[734]), .Z(n22645) );
  XNOR U22511 ( .A(n16448), .B(p_input[729]), .Z(n22586) );
  XNOR U22512 ( .A(n22607), .B(n22606), .Z(n22573) );
  XNOR U22513 ( .A(n22646), .B(n22613), .Z(n22606) );
  XNOR U22514 ( .A(n22602), .B(n22601), .Z(n22613) );
  XOR U22515 ( .A(n22647), .B(n22598), .Z(n22601) );
  XNOR U22516 ( .A(n16737), .B(p_input[715]), .Z(n22598) );
  XNOR U22517 ( .A(p_input[2060]), .B(p_input[716]), .Z(n22647) );
  XOR U22518 ( .A(p_input[2061]), .B(p_input[717]), .Z(n22602) );
  XNOR U22519 ( .A(n22612), .B(n22603), .Z(n22646) );
  XNOR U22520 ( .A(n16452), .B(p_input[706]), .Z(n22603) );
  XOR U22521 ( .A(n22648), .B(n22618), .Z(n22612) );
  XNOR U22522 ( .A(p_input[2064]), .B(p_input[720]), .Z(n22618) );
  XOR U22523 ( .A(n22609), .B(n22617), .Z(n22648) );
  XOR U22524 ( .A(n22649), .B(n22614), .Z(n22617) );
  XOR U22525 ( .A(p_input[2062]), .B(p_input[718]), .Z(n22614) );
  XNOR U22526 ( .A(p_input[2063]), .B(p_input[719]), .Z(n22649) );
  XNOR U22527 ( .A(n16740), .B(p_input[714]), .Z(n22609) );
  XNOR U22528 ( .A(n22624), .B(n22623), .Z(n22607) );
  XNOR U22529 ( .A(n22650), .B(n22629), .Z(n22623) );
  XOR U22530 ( .A(p_input[2057]), .B(p_input[713]), .Z(n22629) );
  XOR U22531 ( .A(n22620), .B(n22628), .Z(n22650) );
  XOR U22532 ( .A(n22651), .B(n22625), .Z(n22628) );
  XOR U22533 ( .A(p_input[2055]), .B(p_input[711]), .Z(n22625) );
  XNOR U22534 ( .A(p_input[2056]), .B(p_input[712]), .Z(n22651) );
  XNOR U22535 ( .A(n16459), .B(p_input[707]), .Z(n22620) );
  XNOR U22536 ( .A(n22634), .B(n22633), .Z(n22624) );
  XOR U22537 ( .A(n22652), .B(n22630), .Z(n22633) );
  XOR U22538 ( .A(p_input[2052]), .B(p_input[708]), .Z(n22630) );
  XNOR U22539 ( .A(p_input[2053]), .B(p_input[709]), .Z(n22652) );
  XOR U22540 ( .A(p_input[2054]), .B(p_input[710]), .Z(n22634) );
  XNOR U22541 ( .A(n22653), .B(n22654), .Z(n22451) );
  AND U22542 ( .A(n309), .B(n22655), .Z(n22654) );
  XNOR U22543 ( .A(n22656), .B(n22657), .Z(n309) );
  AND U22544 ( .A(n22658), .B(n22659), .Z(n22657) );
  XOR U22545 ( .A(n22656), .B(n22461), .Z(n22659) );
  XNOR U22546 ( .A(n22656), .B(n22403), .Z(n22658) );
  XOR U22547 ( .A(n22660), .B(n22661), .Z(n22656) );
  AND U22548 ( .A(n22662), .B(n22663), .Z(n22661) );
  XNOR U22549 ( .A(n22474), .B(n22660), .Z(n22663) );
  XOR U22550 ( .A(n22660), .B(n22415), .Z(n22662) );
  XOR U22551 ( .A(n22664), .B(n22665), .Z(n22660) );
  AND U22552 ( .A(n22666), .B(n22667), .Z(n22665) );
  XNOR U22553 ( .A(n22499), .B(n22664), .Z(n22667) );
  XOR U22554 ( .A(n22664), .B(n22426), .Z(n22666) );
  XOR U22555 ( .A(n22668), .B(n22669), .Z(n22664) );
  AND U22556 ( .A(n22670), .B(n22671), .Z(n22669) );
  XOR U22557 ( .A(n22668), .B(n22436), .Z(n22670) );
  XOR U22558 ( .A(n22672), .B(n22673), .Z(n22392) );
  AND U22559 ( .A(n313), .B(n22655), .Z(n22673) );
  XNOR U22560 ( .A(n22653), .B(n22672), .Z(n22655) );
  XNOR U22561 ( .A(n22674), .B(n22675), .Z(n313) );
  AND U22562 ( .A(n22676), .B(n22677), .Z(n22675) );
  XNOR U22563 ( .A(n22678), .B(n22674), .Z(n22677) );
  IV U22564 ( .A(n22461), .Z(n22678) );
  XNOR U22565 ( .A(n22679), .B(n22680), .Z(n22461) );
  AND U22566 ( .A(n316), .B(n22681), .Z(n22680) );
  XNOR U22567 ( .A(n22679), .B(n22682), .Z(n22681) );
  XNOR U22568 ( .A(n22403), .B(n22674), .Z(n22676) );
  XOR U22569 ( .A(n22683), .B(n22684), .Z(n22403) );
  AND U22570 ( .A(n324), .B(n22685), .Z(n22684) );
  XOR U22571 ( .A(n22686), .B(n22687), .Z(n22674) );
  AND U22572 ( .A(n22688), .B(n22689), .Z(n22687) );
  XNOR U22573 ( .A(n22686), .B(n22474), .Z(n22689) );
  XNOR U22574 ( .A(n22690), .B(n22691), .Z(n22474) );
  AND U22575 ( .A(n316), .B(n22692), .Z(n22691) );
  XOR U22576 ( .A(n22693), .B(n22690), .Z(n22692) );
  XNOR U22577 ( .A(n22694), .B(n22686), .Z(n22688) );
  IV U22578 ( .A(n22415), .Z(n22694) );
  XOR U22579 ( .A(n22695), .B(n22696), .Z(n22415) );
  AND U22580 ( .A(n324), .B(n22697), .Z(n22696) );
  XOR U22581 ( .A(n22698), .B(n22699), .Z(n22686) );
  AND U22582 ( .A(n22700), .B(n22701), .Z(n22699) );
  XNOR U22583 ( .A(n22698), .B(n22499), .Z(n22701) );
  XNOR U22584 ( .A(n22702), .B(n22703), .Z(n22499) );
  AND U22585 ( .A(n316), .B(n22704), .Z(n22703) );
  XNOR U22586 ( .A(n22705), .B(n22702), .Z(n22704) );
  XOR U22587 ( .A(n22426), .B(n22698), .Z(n22700) );
  XOR U22588 ( .A(n22706), .B(n22707), .Z(n22426) );
  AND U22589 ( .A(n324), .B(n22708), .Z(n22707) );
  XOR U22590 ( .A(n22668), .B(n22709), .Z(n22698) );
  AND U22591 ( .A(n22710), .B(n22671), .Z(n22709) );
  XNOR U22592 ( .A(n22545), .B(n22668), .Z(n22671) );
  XNOR U22593 ( .A(n22711), .B(n22712), .Z(n22545) );
  AND U22594 ( .A(n316), .B(n22713), .Z(n22712) );
  XOR U22595 ( .A(n22714), .B(n22711), .Z(n22713) );
  XNOR U22596 ( .A(n22715), .B(n22668), .Z(n22710) );
  IV U22597 ( .A(n22436), .Z(n22715) );
  XOR U22598 ( .A(n22716), .B(n22717), .Z(n22436) );
  AND U22599 ( .A(n324), .B(n22718), .Z(n22717) );
  XOR U22600 ( .A(n22719), .B(n22720), .Z(n22668) );
  AND U22601 ( .A(n22721), .B(n22722), .Z(n22720) );
  XNOR U22602 ( .A(n22719), .B(n22635), .Z(n22722) );
  XNOR U22603 ( .A(n22723), .B(n22724), .Z(n22635) );
  AND U22604 ( .A(n316), .B(n22725), .Z(n22724) );
  XNOR U22605 ( .A(n22726), .B(n22723), .Z(n22725) );
  XNOR U22606 ( .A(n22727), .B(n22719), .Z(n22721) );
  IV U22607 ( .A(n22448), .Z(n22727) );
  XOR U22608 ( .A(n22728), .B(n22729), .Z(n22448) );
  AND U22609 ( .A(n324), .B(n22730), .Z(n22729) );
  AND U22610 ( .A(n22672), .B(n22653), .Z(n22719) );
  XNOR U22611 ( .A(n22731), .B(n22732), .Z(n22653) );
  AND U22612 ( .A(n316), .B(n22733), .Z(n22732) );
  XNOR U22613 ( .A(n22734), .B(n22731), .Z(n22733) );
  XNOR U22614 ( .A(n22735), .B(n22736), .Z(n316) );
  AND U22615 ( .A(n22737), .B(n22738), .Z(n22736) );
  XOR U22616 ( .A(n22682), .B(n22735), .Z(n22738) );
  AND U22617 ( .A(n22739), .B(n22740), .Z(n22682) );
  XOR U22618 ( .A(n22735), .B(n22679), .Z(n22737) );
  XNOR U22619 ( .A(n22741), .B(n22742), .Z(n22679) );
  AND U22620 ( .A(n320), .B(n22685), .Z(n22742) );
  XOR U22621 ( .A(n22683), .B(n22741), .Z(n22685) );
  XOR U22622 ( .A(n22743), .B(n22744), .Z(n22735) );
  AND U22623 ( .A(n22745), .B(n22746), .Z(n22744) );
  XNOR U22624 ( .A(n22743), .B(n22739), .Z(n22746) );
  IV U22625 ( .A(n22693), .Z(n22739) );
  XOR U22626 ( .A(n22747), .B(n22748), .Z(n22693) );
  XOR U22627 ( .A(n22749), .B(n22740), .Z(n22748) );
  AND U22628 ( .A(n22705), .B(n22750), .Z(n22740) );
  AND U22629 ( .A(n22751), .B(n22752), .Z(n22749) );
  XOR U22630 ( .A(n22753), .B(n22747), .Z(n22751) );
  XNOR U22631 ( .A(n22690), .B(n22743), .Z(n22745) );
  XNOR U22632 ( .A(n22754), .B(n22755), .Z(n22690) );
  AND U22633 ( .A(n320), .B(n22697), .Z(n22755) );
  XOR U22634 ( .A(n22754), .B(n22695), .Z(n22697) );
  XOR U22635 ( .A(n22756), .B(n22757), .Z(n22743) );
  AND U22636 ( .A(n22758), .B(n22759), .Z(n22757) );
  XNOR U22637 ( .A(n22756), .B(n22705), .Z(n22759) );
  XOR U22638 ( .A(n22760), .B(n22752), .Z(n22705) );
  XNOR U22639 ( .A(n22761), .B(n22747), .Z(n22752) );
  XOR U22640 ( .A(n22762), .B(n22763), .Z(n22747) );
  AND U22641 ( .A(n22764), .B(n22765), .Z(n22763) );
  XOR U22642 ( .A(n22766), .B(n22762), .Z(n22764) );
  XNOR U22643 ( .A(n22767), .B(n22768), .Z(n22761) );
  AND U22644 ( .A(n22769), .B(n22770), .Z(n22768) );
  XOR U22645 ( .A(n22767), .B(n22771), .Z(n22769) );
  XNOR U22646 ( .A(n22753), .B(n22750), .Z(n22760) );
  AND U22647 ( .A(n22772), .B(n22773), .Z(n22750) );
  XOR U22648 ( .A(n22774), .B(n22775), .Z(n22753) );
  AND U22649 ( .A(n22776), .B(n22777), .Z(n22775) );
  XOR U22650 ( .A(n22774), .B(n22778), .Z(n22776) );
  XNOR U22651 ( .A(n22702), .B(n22756), .Z(n22758) );
  XNOR U22652 ( .A(n22779), .B(n22780), .Z(n22702) );
  AND U22653 ( .A(n320), .B(n22708), .Z(n22780) );
  XOR U22654 ( .A(n22779), .B(n22706), .Z(n22708) );
  XOR U22655 ( .A(n22781), .B(n22782), .Z(n22756) );
  AND U22656 ( .A(n22783), .B(n22784), .Z(n22782) );
  XNOR U22657 ( .A(n22781), .B(n22772), .Z(n22784) );
  IV U22658 ( .A(n22714), .Z(n22772) );
  XNOR U22659 ( .A(n22785), .B(n22765), .Z(n22714) );
  XNOR U22660 ( .A(n22786), .B(n22771), .Z(n22765) );
  XOR U22661 ( .A(n22787), .B(n22788), .Z(n22771) );
  AND U22662 ( .A(n22789), .B(n22790), .Z(n22788) );
  XOR U22663 ( .A(n22787), .B(n22791), .Z(n22789) );
  XNOR U22664 ( .A(n22770), .B(n22762), .Z(n22786) );
  XOR U22665 ( .A(n22792), .B(n22793), .Z(n22762) );
  AND U22666 ( .A(n22794), .B(n22795), .Z(n22793) );
  XNOR U22667 ( .A(n22796), .B(n22792), .Z(n22794) );
  XNOR U22668 ( .A(n22797), .B(n22767), .Z(n22770) );
  XOR U22669 ( .A(n22798), .B(n22799), .Z(n22767) );
  AND U22670 ( .A(n22800), .B(n22801), .Z(n22799) );
  XOR U22671 ( .A(n22798), .B(n22802), .Z(n22800) );
  XNOR U22672 ( .A(n22803), .B(n22804), .Z(n22797) );
  AND U22673 ( .A(n22805), .B(n22806), .Z(n22804) );
  XNOR U22674 ( .A(n22803), .B(n22807), .Z(n22805) );
  XNOR U22675 ( .A(n22766), .B(n22773), .Z(n22785) );
  AND U22676 ( .A(n22726), .B(n22808), .Z(n22773) );
  XOR U22677 ( .A(n22778), .B(n22777), .Z(n22766) );
  XNOR U22678 ( .A(n22809), .B(n22774), .Z(n22777) );
  XOR U22679 ( .A(n22810), .B(n22811), .Z(n22774) );
  AND U22680 ( .A(n22812), .B(n22813), .Z(n22811) );
  XOR U22681 ( .A(n22810), .B(n22814), .Z(n22812) );
  XNOR U22682 ( .A(n22815), .B(n22816), .Z(n22809) );
  AND U22683 ( .A(n22817), .B(n22818), .Z(n22816) );
  XOR U22684 ( .A(n22815), .B(n22819), .Z(n22817) );
  XOR U22685 ( .A(n22820), .B(n22821), .Z(n22778) );
  AND U22686 ( .A(n22822), .B(n22823), .Z(n22821) );
  XOR U22687 ( .A(n22820), .B(n22824), .Z(n22822) );
  XNOR U22688 ( .A(n22711), .B(n22781), .Z(n22783) );
  XNOR U22689 ( .A(n22825), .B(n22826), .Z(n22711) );
  AND U22690 ( .A(n320), .B(n22718), .Z(n22826) );
  XOR U22691 ( .A(n22825), .B(n22716), .Z(n22718) );
  XOR U22692 ( .A(n22827), .B(n22828), .Z(n22781) );
  AND U22693 ( .A(n22829), .B(n22830), .Z(n22828) );
  XNOR U22694 ( .A(n22827), .B(n22726), .Z(n22830) );
  XOR U22695 ( .A(n22831), .B(n22795), .Z(n22726) );
  XNOR U22696 ( .A(n22832), .B(n22802), .Z(n22795) );
  XOR U22697 ( .A(n22791), .B(n22790), .Z(n22802) );
  XNOR U22698 ( .A(n22833), .B(n22787), .Z(n22790) );
  XOR U22699 ( .A(n22834), .B(n22835), .Z(n22787) );
  AND U22700 ( .A(n22836), .B(n22837), .Z(n22835) );
  XOR U22701 ( .A(n22834), .B(n22838), .Z(n22836) );
  XNOR U22702 ( .A(n22839), .B(n22840), .Z(n22833) );
  NOR U22703 ( .A(n22841), .B(n22842), .Z(n22840) );
  XNOR U22704 ( .A(n22839), .B(n22843), .Z(n22841) );
  XOR U22705 ( .A(n22844), .B(n22845), .Z(n22791) );
  NOR U22706 ( .A(n22846), .B(n22847), .Z(n22845) );
  XNOR U22707 ( .A(n22844), .B(n22848), .Z(n22846) );
  XNOR U22708 ( .A(n22801), .B(n22792), .Z(n22832) );
  XOR U22709 ( .A(n22849), .B(n22850), .Z(n22792) );
  NOR U22710 ( .A(n22851), .B(n22852), .Z(n22850) );
  XNOR U22711 ( .A(n22849), .B(n22853), .Z(n22851) );
  XOR U22712 ( .A(n22854), .B(n22807), .Z(n22801) );
  XNOR U22713 ( .A(n22855), .B(n22856), .Z(n22807) );
  NOR U22714 ( .A(n22857), .B(n22858), .Z(n22856) );
  XNOR U22715 ( .A(n22855), .B(n22859), .Z(n22857) );
  XNOR U22716 ( .A(n22806), .B(n22798), .Z(n22854) );
  XOR U22717 ( .A(n22860), .B(n22861), .Z(n22798) );
  AND U22718 ( .A(n22862), .B(n22863), .Z(n22861) );
  XOR U22719 ( .A(n22860), .B(n22864), .Z(n22862) );
  XNOR U22720 ( .A(n22865), .B(n22803), .Z(n22806) );
  XOR U22721 ( .A(n22866), .B(n22867), .Z(n22803) );
  AND U22722 ( .A(n22868), .B(n22869), .Z(n22867) );
  XOR U22723 ( .A(n22866), .B(n22870), .Z(n22868) );
  XNOR U22724 ( .A(n22871), .B(n22872), .Z(n22865) );
  NOR U22725 ( .A(n22873), .B(n22874), .Z(n22872) );
  XOR U22726 ( .A(n22871), .B(n22875), .Z(n22873) );
  XOR U22727 ( .A(n22796), .B(n22808), .Z(n22831) );
  NOR U22728 ( .A(n22734), .B(n22876), .Z(n22808) );
  XNOR U22729 ( .A(n22814), .B(n22813), .Z(n22796) );
  XNOR U22730 ( .A(n22877), .B(n22819), .Z(n22813) );
  XOR U22731 ( .A(n22878), .B(n22879), .Z(n22819) );
  NOR U22732 ( .A(n22880), .B(n22881), .Z(n22879) );
  XNOR U22733 ( .A(n22878), .B(n22882), .Z(n22880) );
  XNOR U22734 ( .A(n22818), .B(n22810), .Z(n22877) );
  XOR U22735 ( .A(n22883), .B(n22884), .Z(n22810) );
  AND U22736 ( .A(n22885), .B(n22886), .Z(n22884) );
  XNOR U22737 ( .A(n22883), .B(n22887), .Z(n22885) );
  XNOR U22738 ( .A(n22888), .B(n22815), .Z(n22818) );
  XOR U22739 ( .A(n22889), .B(n22890), .Z(n22815) );
  AND U22740 ( .A(n22891), .B(n22892), .Z(n22890) );
  XOR U22741 ( .A(n22889), .B(n22893), .Z(n22891) );
  XNOR U22742 ( .A(n22894), .B(n22895), .Z(n22888) );
  NOR U22743 ( .A(n22896), .B(n22897), .Z(n22895) );
  XOR U22744 ( .A(n22894), .B(n22898), .Z(n22896) );
  XOR U22745 ( .A(n22824), .B(n22823), .Z(n22814) );
  XNOR U22746 ( .A(n22899), .B(n22820), .Z(n22823) );
  XOR U22747 ( .A(n22900), .B(n22901), .Z(n22820) );
  AND U22748 ( .A(n22902), .B(n22903), .Z(n22901) );
  XOR U22749 ( .A(n22900), .B(n22904), .Z(n22902) );
  XNOR U22750 ( .A(n22905), .B(n22906), .Z(n22899) );
  NOR U22751 ( .A(n22907), .B(n22908), .Z(n22906) );
  XNOR U22752 ( .A(n22905), .B(n22909), .Z(n22907) );
  XOR U22753 ( .A(n22910), .B(n22911), .Z(n22824) );
  NOR U22754 ( .A(n22912), .B(n22913), .Z(n22911) );
  XNOR U22755 ( .A(n22910), .B(n22914), .Z(n22912) );
  XNOR U22756 ( .A(n22723), .B(n22827), .Z(n22829) );
  XNOR U22757 ( .A(n22915), .B(n22916), .Z(n22723) );
  AND U22758 ( .A(n320), .B(n22730), .Z(n22916) );
  XOR U22759 ( .A(n22915), .B(n22728), .Z(n22730) );
  AND U22760 ( .A(n22731), .B(n22734), .Z(n22827) );
  XOR U22761 ( .A(n22917), .B(n22876), .Z(n22734) );
  XNOR U22762 ( .A(p_input[2048]), .B(p_input[736]), .Z(n22876) );
  XOR U22763 ( .A(n22853), .B(n22852), .Z(n22917) );
  XOR U22764 ( .A(n22918), .B(n22864), .Z(n22852) );
  XOR U22765 ( .A(n22838), .B(n22837), .Z(n22864) );
  XNOR U22766 ( .A(n22919), .B(n22843), .Z(n22837) );
  XOR U22767 ( .A(p_input[2072]), .B(p_input[760]), .Z(n22843) );
  XOR U22768 ( .A(n22834), .B(n22842), .Z(n22919) );
  XOR U22769 ( .A(n22920), .B(n22839), .Z(n22842) );
  XOR U22770 ( .A(p_input[2070]), .B(p_input[758]), .Z(n22839) );
  XNOR U22771 ( .A(p_input[2071]), .B(p_input[759]), .Z(n22920) );
  XNOR U22772 ( .A(n16727), .B(p_input[754]), .Z(n22834) );
  XNOR U22773 ( .A(n22848), .B(n22847), .Z(n22838) );
  XOR U22774 ( .A(n22921), .B(n22844), .Z(n22847) );
  XOR U22775 ( .A(p_input[2067]), .B(p_input[755]), .Z(n22844) );
  XNOR U22776 ( .A(p_input[2068]), .B(p_input[756]), .Z(n22921) );
  XOR U22777 ( .A(p_input[2069]), .B(p_input[757]), .Z(n22848) );
  XNOR U22778 ( .A(n22863), .B(n22849), .Z(n22918) );
  XNOR U22779 ( .A(n16729), .B(p_input[737]), .Z(n22849) );
  XNOR U22780 ( .A(n22922), .B(n22870), .Z(n22863) );
  XNOR U22781 ( .A(n22859), .B(n22858), .Z(n22870) );
  XOR U22782 ( .A(n22923), .B(n22855), .Z(n22858) );
  XNOR U22783 ( .A(n16444), .B(p_input[762]), .Z(n22855) );
  XNOR U22784 ( .A(p_input[2075]), .B(p_input[763]), .Z(n22923) );
  XOR U22785 ( .A(p_input[2076]), .B(p_input[764]), .Z(n22859) );
  XNOR U22786 ( .A(n22869), .B(n22860), .Z(n22922) );
  XNOR U22787 ( .A(n16732), .B(p_input[753]), .Z(n22860) );
  XOR U22788 ( .A(n22924), .B(n22875), .Z(n22869) );
  XNOR U22789 ( .A(p_input[2079]), .B(p_input[767]), .Z(n22875) );
  XOR U22790 ( .A(n22866), .B(n22874), .Z(n22924) );
  XOR U22791 ( .A(n22925), .B(n22871), .Z(n22874) );
  XOR U22792 ( .A(p_input[2077]), .B(p_input[765]), .Z(n22871) );
  XNOR U22793 ( .A(p_input[2078]), .B(p_input[766]), .Z(n22925) );
  XNOR U22794 ( .A(n16448), .B(p_input[761]), .Z(n22866) );
  XNOR U22795 ( .A(n22887), .B(n22886), .Z(n22853) );
  XNOR U22796 ( .A(n22926), .B(n22893), .Z(n22886) );
  XNOR U22797 ( .A(n22882), .B(n22881), .Z(n22893) );
  XOR U22798 ( .A(n22927), .B(n22878), .Z(n22881) );
  XNOR U22799 ( .A(n16737), .B(p_input[747]), .Z(n22878) );
  XNOR U22800 ( .A(p_input[2060]), .B(p_input[748]), .Z(n22927) );
  XOR U22801 ( .A(p_input[2061]), .B(p_input[749]), .Z(n22882) );
  XNOR U22802 ( .A(n22892), .B(n22883), .Z(n22926) );
  XNOR U22803 ( .A(n16452), .B(p_input[738]), .Z(n22883) );
  XOR U22804 ( .A(n22928), .B(n22898), .Z(n22892) );
  XNOR U22805 ( .A(p_input[2064]), .B(p_input[752]), .Z(n22898) );
  XOR U22806 ( .A(n22889), .B(n22897), .Z(n22928) );
  XOR U22807 ( .A(n22929), .B(n22894), .Z(n22897) );
  XOR U22808 ( .A(p_input[2062]), .B(p_input[750]), .Z(n22894) );
  XNOR U22809 ( .A(p_input[2063]), .B(p_input[751]), .Z(n22929) );
  XNOR U22810 ( .A(n16740), .B(p_input[746]), .Z(n22889) );
  XNOR U22811 ( .A(n22904), .B(n22903), .Z(n22887) );
  XNOR U22812 ( .A(n22930), .B(n22909), .Z(n22903) );
  XOR U22813 ( .A(p_input[2057]), .B(p_input[745]), .Z(n22909) );
  XOR U22814 ( .A(n22900), .B(n22908), .Z(n22930) );
  XOR U22815 ( .A(n22931), .B(n22905), .Z(n22908) );
  XOR U22816 ( .A(p_input[2055]), .B(p_input[743]), .Z(n22905) );
  XNOR U22817 ( .A(p_input[2056]), .B(p_input[744]), .Z(n22931) );
  XNOR U22818 ( .A(n16459), .B(p_input[739]), .Z(n22900) );
  XNOR U22819 ( .A(n22914), .B(n22913), .Z(n22904) );
  XOR U22820 ( .A(n22932), .B(n22910), .Z(n22913) );
  XOR U22821 ( .A(p_input[2052]), .B(p_input[740]), .Z(n22910) );
  XNOR U22822 ( .A(p_input[2053]), .B(p_input[741]), .Z(n22932) );
  XOR U22823 ( .A(p_input[2054]), .B(p_input[742]), .Z(n22914) );
  XNOR U22824 ( .A(n22933), .B(n22934), .Z(n22731) );
  AND U22825 ( .A(n320), .B(n22935), .Z(n22934) );
  XNOR U22826 ( .A(n22936), .B(n22937), .Z(n320) );
  AND U22827 ( .A(n22938), .B(n22939), .Z(n22937) );
  XOR U22828 ( .A(n22936), .B(n22741), .Z(n22939) );
  XNOR U22829 ( .A(n22936), .B(n22683), .Z(n22938) );
  XOR U22830 ( .A(n22940), .B(n22941), .Z(n22936) );
  AND U22831 ( .A(n22942), .B(n22943), .Z(n22941) );
  XNOR U22832 ( .A(n22754), .B(n22940), .Z(n22943) );
  XOR U22833 ( .A(n22940), .B(n22695), .Z(n22942) );
  XOR U22834 ( .A(n22944), .B(n22945), .Z(n22940) );
  AND U22835 ( .A(n22946), .B(n22947), .Z(n22945) );
  XNOR U22836 ( .A(n22779), .B(n22944), .Z(n22947) );
  XOR U22837 ( .A(n22944), .B(n22706), .Z(n22946) );
  XOR U22838 ( .A(n22948), .B(n22949), .Z(n22944) );
  AND U22839 ( .A(n22950), .B(n22951), .Z(n22949) );
  XOR U22840 ( .A(n22948), .B(n22716), .Z(n22950) );
  XOR U22841 ( .A(n22952), .B(n22953), .Z(n22672) );
  AND U22842 ( .A(n324), .B(n22935), .Z(n22953) );
  XNOR U22843 ( .A(n22933), .B(n22952), .Z(n22935) );
  XNOR U22844 ( .A(n22954), .B(n22955), .Z(n324) );
  AND U22845 ( .A(n22956), .B(n22957), .Z(n22955) );
  XNOR U22846 ( .A(n22958), .B(n22954), .Z(n22957) );
  IV U22847 ( .A(n22741), .Z(n22958) );
  XNOR U22848 ( .A(n22959), .B(n22960), .Z(n22741) );
  AND U22849 ( .A(n327), .B(n22961), .Z(n22960) );
  XNOR U22850 ( .A(n22959), .B(n22962), .Z(n22961) );
  XNOR U22851 ( .A(n22683), .B(n22954), .Z(n22956) );
  XOR U22852 ( .A(n22963), .B(n22964), .Z(n22683) );
  AND U22853 ( .A(n335), .B(n22965), .Z(n22964) );
  XOR U22854 ( .A(n22966), .B(n22967), .Z(n22954) );
  AND U22855 ( .A(n22968), .B(n22969), .Z(n22967) );
  XNOR U22856 ( .A(n22966), .B(n22754), .Z(n22969) );
  XNOR U22857 ( .A(n22970), .B(n22971), .Z(n22754) );
  AND U22858 ( .A(n327), .B(n22972), .Z(n22971) );
  XOR U22859 ( .A(n22973), .B(n22970), .Z(n22972) );
  XNOR U22860 ( .A(n22974), .B(n22966), .Z(n22968) );
  IV U22861 ( .A(n22695), .Z(n22974) );
  XOR U22862 ( .A(n22975), .B(n22976), .Z(n22695) );
  AND U22863 ( .A(n335), .B(n22977), .Z(n22976) );
  XOR U22864 ( .A(n22978), .B(n22979), .Z(n22966) );
  AND U22865 ( .A(n22980), .B(n22981), .Z(n22979) );
  XNOR U22866 ( .A(n22978), .B(n22779), .Z(n22981) );
  XNOR U22867 ( .A(n22982), .B(n22983), .Z(n22779) );
  AND U22868 ( .A(n327), .B(n22984), .Z(n22983) );
  XNOR U22869 ( .A(n22985), .B(n22982), .Z(n22984) );
  XOR U22870 ( .A(n22706), .B(n22978), .Z(n22980) );
  XOR U22871 ( .A(n22986), .B(n22987), .Z(n22706) );
  AND U22872 ( .A(n335), .B(n22988), .Z(n22987) );
  XOR U22873 ( .A(n22948), .B(n22989), .Z(n22978) );
  AND U22874 ( .A(n22990), .B(n22951), .Z(n22989) );
  XNOR U22875 ( .A(n22825), .B(n22948), .Z(n22951) );
  XNOR U22876 ( .A(n22991), .B(n22992), .Z(n22825) );
  AND U22877 ( .A(n327), .B(n22993), .Z(n22992) );
  XOR U22878 ( .A(n22994), .B(n22991), .Z(n22993) );
  XNOR U22879 ( .A(n22995), .B(n22948), .Z(n22990) );
  IV U22880 ( .A(n22716), .Z(n22995) );
  XOR U22881 ( .A(n22996), .B(n22997), .Z(n22716) );
  AND U22882 ( .A(n335), .B(n22998), .Z(n22997) );
  XOR U22883 ( .A(n22999), .B(n23000), .Z(n22948) );
  AND U22884 ( .A(n23001), .B(n23002), .Z(n23000) );
  XNOR U22885 ( .A(n22999), .B(n22915), .Z(n23002) );
  XNOR U22886 ( .A(n23003), .B(n23004), .Z(n22915) );
  AND U22887 ( .A(n327), .B(n23005), .Z(n23004) );
  XNOR U22888 ( .A(n23006), .B(n23003), .Z(n23005) );
  XNOR U22889 ( .A(n23007), .B(n22999), .Z(n23001) );
  IV U22890 ( .A(n22728), .Z(n23007) );
  XOR U22891 ( .A(n23008), .B(n23009), .Z(n22728) );
  AND U22892 ( .A(n335), .B(n23010), .Z(n23009) );
  AND U22893 ( .A(n22952), .B(n22933), .Z(n22999) );
  XNOR U22894 ( .A(n23011), .B(n23012), .Z(n22933) );
  AND U22895 ( .A(n327), .B(n23013), .Z(n23012) );
  XNOR U22896 ( .A(n23014), .B(n23011), .Z(n23013) );
  XNOR U22897 ( .A(n23015), .B(n23016), .Z(n327) );
  AND U22898 ( .A(n23017), .B(n23018), .Z(n23016) );
  XOR U22899 ( .A(n22962), .B(n23015), .Z(n23018) );
  AND U22900 ( .A(n23019), .B(n23020), .Z(n22962) );
  XOR U22901 ( .A(n23015), .B(n22959), .Z(n23017) );
  XNOR U22902 ( .A(n23021), .B(n23022), .Z(n22959) );
  AND U22903 ( .A(n331), .B(n22965), .Z(n23022) );
  XOR U22904 ( .A(n22963), .B(n23021), .Z(n22965) );
  XOR U22905 ( .A(n23023), .B(n23024), .Z(n23015) );
  AND U22906 ( .A(n23025), .B(n23026), .Z(n23024) );
  XNOR U22907 ( .A(n23023), .B(n23019), .Z(n23026) );
  IV U22908 ( .A(n22973), .Z(n23019) );
  XOR U22909 ( .A(n23027), .B(n23028), .Z(n22973) );
  XOR U22910 ( .A(n23029), .B(n23020), .Z(n23028) );
  AND U22911 ( .A(n22985), .B(n23030), .Z(n23020) );
  AND U22912 ( .A(n23031), .B(n23032), .Z(n23029) );
  XOR U22913 ( .A(n23033), .B(n23027), .Z(n23031) );
  XNOR U22914 ( .A(n22970), .B(n23023), .Z(n23025) );
  XNOR U22915 ( .A(n23034), .B(n23035), .Z(n22970) );
  AND U22916 ( .A(n331), .B(n22977), .Z(n23035) );
  XOR U22917 ( .A(n23034), .B(n22975), .Z(n22977) );
  XOR U22918 ( .A(n23036), .B(n23037), .Z(n23023) );
  AND U22919 ( .A(n23038), .B(n23039), .Z(n23037) );
  XNOR U22920 ( .A(n23036), .B(n22985), .Z(n23039) );
  XOR U22921 ( .A(n23040), .B(n23032), .Z(n22985) );
  XNOR U22922 ( .A(n23041), .B(n23027), .Z(n23032) );
  XOR U22923 ( .A(n23042), .B(n23043), .Z(n23027) );
  AND U22924 ( .A(n23044), .B(n23045), .Z(n23043) );
  XOR U22925 ( .A(n23046), .B(n23042), .Z(n23044) );
  XNOR U22926 ( .A(n23047), .B(n23048), .Z(n23041) );
  AND U22927 ( .A(n23049), .B(n23050), .Z(n23048) );
  XOR U22928 ( .A(n23047), .B(n23051), .Z(n23049) );
  XNOR U22929 ( .A(n23033), .B(n23030), .Z(n23040) );
  AND U22930 ( .A(n23052), .B(n23053), .Z(n23030) );
  XOR U22931 ( .A(n23054), .B(n23055), .Z(n23033) );
  AND U22932 ( .A(n23056), .B(n23057), .Z(n23055) );
  XOR U22933 ( .A(n23054), .B(n23058), .Z(n23056) );
  XNOR U22934 ( .A(n22982), .B(n23036), .Z(n23038) );
  XNOR U22935 ( .A(n23059), .B(n23060), .Z(n22982) );
  AND U22936 ( .A(n331), .B(n22988), .Z(n23060) );
  XOR U22937 ( .A(n23059), .B(n22986), .Z(n22988) );
  XOR U22938 ( .A(n23061), .B(n23062), .Z(n23036) );
  AND U22939 ( .A(n23063), .B(n23064), .Z(n23062) );
  XNOR U22940 ( .A(n23061), .B(n23052), .Z(n23064) );
  IV U22941 ( .A(n22994), .Z(n23052) );
  XNOR U22942 ( .A(n23065), .B(n23045), .Z(n22994) );
  XNOR U22943 ( .A(n23066), .B(n23051), .Z(n23045) );
  XOR U22944 ( .A(n23067), .B(n23068), .Z(n23051) );
  AND U22945 ( .A(n23069), .B(n23070), .Z(n23068) );
  XOR U22946 ( .A(n23067), .B(n23071), .Z(n23069) );
  XNOR U22947 ( .A(n23050), .B(n23042), .Z(n23066) );
  XOR U22948 ( .A(n23072), .B(n23073), .Z(n23042) );
  AND U22949 ( .A(n23074), .B(n23075), .Z(n23073) );
  XNOR U22950 ( .A(n23076), .B(n23072), .Z(n23074) );
  XNOR U22951 ( .A(n23077), .B(n23047), .Z(n23050) );
  XOR U22952 ( .A(n23078), .B(n23079), .Z(n23047) );
  AND U22953 ( .A(n23080), .B(n23081), .Z(n23079) );
  XOR U22954 ( .A(n23078), .B(n23082), .Z(n23080) );
  XNOR U22955 ( .A(n23083), .B(n23084), .Z(n23077) );
  AND U22956 ( .A(n23085), .B(n23086), .Z(n23084) );
  XNOR U22957 ( .A(n23083), .B(n23087), .Z(n23085) );
  XNOR U22958 ( .A(n23046), .B(n23053), .Z(n23065) );
  AND U22959 ( .A(n23006), .B(n23088), .Z(n23053) );
  XOR U22960 ( .A(n23058), .B(n23057), .Z(n23046) );
  XNOR U22961 ( .A(n23089), .B(n23054), .Z(n23057) );
  XOR U22962 ( .A(n23090), .B(n23091), .Z(n23054) );
  AND U22963 ( .A(n23092), .B(n23093), .Z(n23091) );
  XOR U22964 ( .A(n23090), .B(n23094), .Z(n23092) );
  XNOR U22965 ( .A(n23095), .B(n23096), .Z(n23089) );
  AND U22966 ( .A(n23097), .B(n23098), .Z(n23096) );
  XOR U22967 ( .A(n23095), .B(n23099), .Z(n23097) );
  XOR U22968 ( .A(n23100), .B(n23101), .Z(n23058) );
  AND U22969 ( .A(n23102), .B(n23103), .Z(n23101) );
  XOR U22970 ( .A(n23100), .B(n23104), .Z(n23102) );
  XNOR U22971 ( .A(n22991), .B(n23061), .Z(n23063) );
  XNOR U22972 ( .A(n23105), .B(n23106), .Z(n22991) );
  AND U22973 ( .A(n331), .B(n22998), .Z(n23106) );
  XOR U22974 ( .A(n23105), .B(n22996), .Z(n22998) );
  XOR U22975 ( .A(n23107), .B(n23108), .Z(n23061) );
  AND U22976 ( .A(n23109), .B(n23110), .Z(n23108) );
  XNOR U22977 ( .A(n23107), .B(n23006), .Z(n23110) );
  XOR U22978 ( .A(n23111), .B(n23075), .Z(n23006) );
  XNOR U22979 ( .A(n23112), .B(n23082), .Z(n23075) );
  XOR U22980 ( .A(n23071), .B(n23070), .Z(n23082) );
  XNOR U22981 ( .A(n23113), .B(n23067), .Z(n23070) );
  XOR U22982 ( .A(n23114), .B(n23115), .Z(n23067) );
  AND U22983 ( .A(n23116), .B(n23117), .Z(n23115) );
  XOR U22984 ( .A(n23114), .B(n23118), .Z(n23116) );
  XNOR U22985 ( .A(n23119), .B(n23120), .Z(n23113) );
  NOR U22986 ( .A(n23121), .B(n23122), .Z(n23120) );
  XNOR U22987 ( .A(n23119), .B(n23123), .Z(n23121) );
  XOR U22988 ( .A(n23124), .B(n23125), .Z(n23071) );
  NOR U22989 ( .A(n23126), .B(n23127), .Z(n23125) );
  XNOR U22990 ( .A(n23124), .B(n23128), .Z(n23126) );
  XNOR U22991 ( .A(n23081), .B(n23072), .Z(n23112) );
  XOR U22992 ( .A(n23129), .B(n23130), .Z(n23072) );
  NOR U22993 ( .A(n23131), .B(n23132), .Z(n23130) );
  XNOR U22994 ( .A(n23129), .B(n23133), .Z(n23131) );
  XOR U22995 ( .A(n23134), .B(n23087), .Z(n23081) );
  XNOR U22996 ( .A(n23135), .B(n23136), .Z(n23087) );
  NOR U22997 ( .A(n23137), .B(n23138), .Z(n23136) );
  XNOR U22998 ( .A(n23135), .B(n23139), .Z(n23137) );
  XNOR U22999 ( .A(n23086), .B(n23078), .Z(n23134) );
  XOR U23000 ( .A(n23140), .B(n23141), .Z(n23078) );
  AND U23001 ( .A(n23142), .B(n23143), .Z(n23141) );
  XOR U23002 ( .A(n23140), .B(n23144), .Z(n23142) );
  XNOR U23003 ( .A(n23145), .B(n23083), .Z(n23086) );
  XOR U23004 ( .A(n23146), .B(n23147), .Z(n23083) );
  AND U23005 ( .A(n23148), .B(n23149), .Z(n23147) );
  XOR U23006 ( .A(n23146), .B(n23150), .Z(n23148) );
  XNOR U23007 ( .A(n23151), .B(n23152), .Z(n23145) );
  NOR U23008 ( .A(n23153), .B(n23154), .Z(n23152) );
  XOR U23009 ( .A(n23151), .B(n23155), .Z(n23153) );
  XOR U23010 ( .A(n23076), .B(n23088), .Z(n23111) );
  NOR U23011 ( .A(n23014), .B(n23156), .Z(n23088) );
  XNOR U23012 ( .A(n23094), .B(n23093), .Z(n23076) );
  XNOR U23013 ( .A(n23157), .B(n23099), .Z(n23093) );
  XOR U23014 ( .A(n23158), .B(n23159), .Z(n23099) );
  NOR U23015 ( .A(n23160), .B(n23161), .Z(n23159) );
  XNOR U23016 ( .A(n23158), .B(n23162), .Z(n23160) );
  XNOR U23017 ( .A(n23098), .B(n23090), .Z(n23157) );
  XOR U23018 ( .A(n23163), .B(n23164), .Z(n23090) );
  AND U23019 ( .A(n23165), .B(n23166), .Z(n23164) );
  XNOR U23020 ( .A(n23163), .B(n23167), .Z(n23165) );
  XNOR U23021 ( .A(n23168), .B(n23095), .Z(n23098) );
  XOR U23022 ( .A(n23169), .B(n23170), .Z(n23095) );
  AND U23023 ( .A(n23171), .B(n23172), .Z(n23170) );
  XOR U23024 ( .A(n23169), .B(n23173), .Z(n23171) );
  XNOR U23025 ( .A(n23174), .B(n23175), .Z(n23168) );
  NOR U23026 ( .A(n23176), .B(n23177), .Z(n23175) );
  XOR U23027 ( .A(n23174), .B(n23178), .Z(n23176) );
  XOR U23028 ( .A(n23104), .B(n23103), .Z(n23094) );
  XNOR U23029 ( .A(n23179), .B(n23100), .Z(n23103) );
  XOR U23030 ( .A(n23180), .B(n23181), .Z(n23100) );
  AND U23031 ( .A(n23182), .B(n23183), .Z(n23181) );
  XOR U23032 ( .A(n23180), .B(n23184), .Z(n23182) );
  XNOR U23033 ( .A(n23185), .B(n23186), .Z(n23179) );
  NOR U23034 ( .A(n23187), .B(n23188), .Z(n23186) );
  XNOR U23035 ( .A(n23185), .B(n23189), .Z(n23187) );
  XOR U23036 ( .A(n23190), .B(n23191), .Z(n23104) );
  NOR U23037 ( .A(n23192), .B(n23193), .Z(n23191) );
  XNOR U23038 ( .A(n23190), .B(n23194), .Z(n23192) );
  XNOR U23039 ( .A(n23003), .B(n23107), .Z(n23109) );
  XNOR U23040 ( .A(n23195), .B(n23196), .Z(n23003) );
  AND U23041 ( .A(n331), .B(n23010), .Z(n23196) );
  XOR U23042 ( .A(n23195), .B(n23008), .Z(n23010) );
  AND U23043 ( .A(n23011), .B(n23014), .Z(n23107) );
  XOR U23044 ( .A(n23197), .B(n23156), .Z(n23014) );
  XNOR U23045 ( .A(p_input[2048]), .B(p_input[768]), .Z(n23156) );
  XOR U23046 ( .A(n23133), .B(n23132), .Z(n23197) );
  XOR U23047 ( .A(n23198), .B(n23144), .Z(n23132) );
  XOR U23048 ( .A(n23118), .B(n23117), .Z(n23144) );
  XNOR U23049 ( .A(n23199), .B(n23123), .Z(n23117) );
  XOR U23050 ( .A(p_input[2072]), .B(p_input[792]), .Z(n23123) );
  XOR U23051 ( .A(n23114), .B(n23122), .Z(n23199) );
  XOR U23052 ( .A(n23200), .B(n23119), .Z(n23122) );
  XOR U23053 ( .A(p_input[2070]), .B(p_input[790]), .Z(n23119) );
  XNOR U23054 ( .A(p_input[2071]), .B(p_input[791]), .Z(n23200) );
  XNOR U23055 ( .A(n16727), .B(p_input[786]), .Z(n23114) );
  XNOR U23056 ( .A(n23128), .B(n23127), .Z(n23118) );
  XOR U23057 ( .A(n23201), .B(n23124), .Z(n23127) );
  XOR U23058 ( .A(p_input[2067]), .B(p_input[787]), .Z(n23124) );
  XNOR U23059 ( .A(p_input[2068]), .B(p_input[788]), .Z(n23201) );
  XOR U23060 ( .A(p_input[2069]), .B(p_input[789]), .Z(n23128) );
  XNOR U23061 ( .A(n23143), .B(n23129), .Z(n23198) );
  XNOR U23062 ( .A(n16729), .B(p_input[769]), .Z(n23129) );
  XNOR U23063 ( .A(n23202), .B(n23150), .Z(n23143) );
  XNOR U23064 ( .A(n23139), .B(n23138), .Z(n23150) );
  XOR U23065 ( .A(n23203), .B(n23135), .Z(n23138) );
  XNOR U23066 ( .A(n16444), .B(p_input[794]), .Z(n23135) );
  XNOR U23067 ( .A(p_input[2075]), .B(p_input[795]), .Z(n23203) );
  XOR U23068 ( .A(p_input[2076]), .B(p_input[796]), .Z(n23139) );
  XNOR U23069 ( .A(n23149), .B(n23140), .Z(n23202) );
  XNOR U23070 ( .A(n16732), .B(p_input[785]), .Z(n23140) );
  XOR U23071 ( .A(n23204), .B(n23155), .Z(n23149) );
  XNOR U23072 ( .A(p_input[2079]), .B(p_input[799]), .Z(n23155) );
  XOR U23073 ( .A(n23146), .B(n23154), .Z(n23204) );
  XOR U23074 ( .A(n23205), .B(n23151), .Z(n23154) );
  XOR U23075 ( .A(p_input[2077]), .B(p_input[797]), .Z(n23151) );
  XNOR U23076 ( .A(p_input[2078]), .B(p_input[798]), .Z(n23205) );
  XNOR U23077 ( .A(n16448), .B(p_input[793]), .Z(n23146) );
  XNOR U23078 ( .A(n23167), .B(n23166), .Z(n23133) );
  XNOR U23079 ( .A(n23206), .B(n23173), .Z(n23166) );
  XNOR U23080 ( .A(n23162), .B(n23161), .Z(n23173) );
  XOR U23081 ( .A(n23207), .B(n23158), .Z(n23161) );
  XNOR U23082 ( .A(n16737), .B(p_input[779]), .Z(n23158) );
  XNOR U23083 ( .A(p_input[2060]), .B(p_input[780]), .Z(n23207) );
  XOR U23084 ( .A(p_input[2061]), .B(p_input[781]), .Z(n23162) );
  XNOR U23085 ( .A(n23172), .B(n23163), .Z(n23206) );
  XNOR U23086 ( .A(n16452), .B(p_input[770]), .Z(n23163) );
  XOR U23087 ( .A(n23208), .B(n23178), .Z(n23172) );
  XNOR U23088 ( .A(p_input[2064]), .B(p_input[784]), .Z(n23178) );
  XOR U23089 ( .A(n23169), .B(n23177), .Z(n23208) );
  XOR U23090 ( .A(n23209), .B(n23174), .Z(n23177) );
  XOR U23091 ( .A(p_input[2062]), .B(p_input[782]), .Z(n23174) );
  XNOR U23092 ( .A(p_input[2063]), .B(p_input[783]), .Z(n23209) );
  XNOR U23093 ( .A(n16740), .B(p_input[778]), .Z(n23169) );
  XNOR U23094 ( .A(n23184), .B(n23183), .Z(n23167) );
  XNOR U23095 ( .A(n23210), .B(n23189), .Z(n23183) );
  XOR U23096 ( .A(p_input[2057]), .B(p_input[777]), .Z(n23189) );
  XOR U23097 ( .A(n23180), .B(n23188), .Z(n23210) );
  XOR U23098 ( .A(n23211), .B(n23185), .Z(n23188) );
  XOR U23099 ( .A(p_input[2055]), .B(p_input[775]), .Z(n23185) );
  XNOR U23100 ( .A(p_input[2056]), .B(p_input[776]), .Z(n23211) );
  XNOR U23101 ( .A(n16459), .B(p_input[771]), .Z(n23180) );
  XNOR U23102 ( .A(n23194), .B(n23193), .Z(n23184) );
  XOR U23103 ( .A(n23212), .B(n23190), .Z(n23193) );
  XOR U23104 ( .A(p_input[2052]), .B(p_input[772]), .Z(n23190) );
  XNOR U23105 ( .A(p_input[2053]), .B(p_input[773]), .Z(n23212) );
  XOR U23106 ( .A(p_input[2054]), .B(p_input[774]), .Z(n23194) );
  XNOR U23107 ( .A(n23213), .B(n23214), .Z(n23011) );
  AND U23108 ( .A(n331), .B(n23215), .Z(n23214) );
  XNOR U23109 ( .A(n23216), .B(n23217), .Z(n331) );
  AND U23110 ( .A(n23218), .B(n23219), .Z(n23217) );
  XOR U23111 ( .A(n23216), .B(n23021), .Z(n23219) );
  XNOR U23112 ( .A(n23216), .B(n22963), .Z(n23218) );
  XOR U23113 ( .A(n23220), .B(n23221), .Z(n23216) );
  AND U23114 ( .A(n23222), .B(n23223), .Z(n23221) );
  XNOR U23115 ( .A(n23034), .B(n23220), .Z(n23223) );
  XOR U23116 ( .A(n23220), .B(n22975), .Z(n23222) );
  XOR U23117 ( .A(n23224), .B(n23225), .Z(n23220) );
  AND U23118 ( .A(n23226), .B(n23227), .Z(n23225) );
  XNOR U23119 ( .A(n23059), .B(n23224), .Z(n23227) );
  XOR U23120 ( .A(n23224), .B(n22986), .Z(n23226) );
  XOR U23121 ( .A(n23228), .B(n23229), .Z(n23224) );
  AND U23122 ( .A(n23230), .B(n23231), .Z(n23229) );
  XOR U23123 ( .A(n23228), .B(n22996), .Z(n23230) );
  XOR U23124 ( .A(n23232), .B(n23233), .Z(n22952) );
  AND U23125 ( .A(n335), .B(n23215), .Z(n23233) );
  XNOR U23126 ( .A(n23213), .B(n23232), .Z(n23215) );
  XNOR U23127 ( .A(n23234), .B(n23235), .Z(n335) );
  AND U23128 ( .A(n23236), .B(n23237), .Z(n23235) );
  XNOR U23129 ( .A(n23238), .B(n23234), .Z(n23237) );
  IV U23130 ( .A(n23021), .Z(n23238) );
  XNOR U23131 ( .A(n23239), .B(n23240), .Z(n23021) );
  AND U23132 ( .A(n338), .B(n23241), .Z(n23240) );
  XNOR U23133 ( .A(n23239), .B(n23242), .Z(n23241) );
  XNOR U23134 ( .A(n22963), .B(n23234), .Z(n23236) );
  XOR U23135 ( .A(n23243), .B(n23244), .Z(n22963) );
  AND U23136 ( .A(n346), .B(n23245), .Z(n23244) );
  XOR U23137 ( .A(n23246), .B(n23247), .Z(n23234) );
  AND U23138 ( .A(n23248), .B(n23249), .Z(n23247) );
  XNOR U23139 ( .A(n23246), .B(n23034), .Z(n23249) );
  XNOR U23140 ( .A(n23250), .B(n23251), .Z(n23034) );
  AND U23141 ( .A(n338), .B(n23252), .Z(n23251) );
  XOR U23142 ( .A(n23253), .B(n23250), .Z(n23252) );
  XNOR U23143 ( .A(n23254), .B(n23246), .Z(n23248) );
  IV U23144 ( .A(n22975), .Z(n23254) );
  XOR U23145 ( .A(n23255), .B(n23256), .Z(n22975) );
  AND U23146 ( .A(n346), .B(n23257), .Z(n23256) );
  XOR U23147 ( .A(n23258), .B(n23259), .Z(n23246) );
  AND U23148 ( .A(n23260), .B(n23261), .Z(n23259) );
  XNOR U23149 ( .A(n23258), .B(n23059), .Z(n23261) );
  XNOR U23150 ( .A(n23262), .B(n23263), .Z(n23059) );
  AND U23151 ( .A(n338), .B(n23264), .Z(n23263) );
  XNOR U23152 ( .A(n23265), .B(n23262), .Z(n23264) );
  XOR U23153 ( .A(n22986), .B(n23258), .Z(n23260) );
  XOR U23154 ( .A(n23266), .B(n23267), .Z(n22986) );
  AND U23155 ( .A(n346), .B(n23268), .Z(n23267) );
  XOR U23156 ( .A(n23228), .B(n23269), .Z(n23258) );
  AND U23157 ( .A(n23270), .B(n23231), .Z(n23269) );
  XNOR U23158 ( .A(n23105), .B(n23228), .Z(n23231) );
  XNOR U23159 ( .A(n23271), .B(n23272), .Z(n23105) );
  AND U23160 ( .A(n338), .B(n23273), .Z(n23272) );
  XOR U23161 ( .A(n23274), .B(n23271), .Z(n23273) );
  XNOR U23162 ( .A(n23275), .B(n23228), .Z(n23270) );
  IV U23163 ( .A(n22996), .Z(n23275) );
  XOR U23164 ( .A(n23276), .B(n23277), .Z(n22996) );
  AND U23165 ( .A(n346), .B(n23278), .Z(n23277) );
  XOR U23166 ( .A(n23279), .B(n23280), .Z(n23228) );
  AND U23167 ( .A(n23281), .B(n23282), .Z(n23280) );
  XNOR U23168 ( .A(n23279), .B(n23195), .Z(n23282) );
  XNOR U23169 ( .A(n23283), .B(n23284), .Z(n23195) );
  AND U23170 ( .A(n338), .B(n23285), .Z(n23284) );
  XNOR U23171 ( .A(n23286), .B(n23283), .Z(n23285) );
  XNOR U23172 ( .A(n23287), .B(n23279), .Z(n23281) );
  IV U23173 ( .A(n23008), .Z(n23287) );
  XOR U23174 ( .A(n23288), .B(n23289), .Z(n23008) );
  AND U23175 ( .A(n346), .B(n23290), .Z(n23289) );
  AND U23176 ( .A(n23232), .B(n23213), .Z(n23279) );
  XNOR U23177 ( .A(n23291), .B(n23292), .Z(n23213) );
  AND U23178 ( .A(n338), .B(n23293), .Z(n23292) );
  XNOR U23179 ( .A(n23294), .B(n23291), .Z(n23293) );
  XNOR U23180 ( .A(n23295), .B(n23296), .Z(n338) );
  AND U23181 ( .A(n23297), .B(n23298), .Z(n23296) );
  XOR U23182 ( .A(n23242), .B(n23295), .Z(n23298) );
  AND U23183 ( .A(n23299), .B(n23300), .Z(n23242) );
  XOR U23184 ( .A(n23295), .B(n23239), .Z(n23297) );
  XNOR U23185 ( .A(n23301), .B(n23302), .Z(n23239) );
  AND U23186 ( .A(n342), .B(n23245), .Z(n23302) );
  XOR U23187 ( .A(n23243), .B(n23301), .Z(n23245) );
  XOR U23188 ( .A(n23303), .B(n23304), .Z(n23295) );
  AND U23189 ( .A(n23305), .B(n23306), .Z(n23304) );
  XNOR U23190 ( .A(n23303), .B(n23299), .Z(n23306) );
  IV U23191 ( .A(n23253), .Z(n23299) );
  XOR U23192 ( .A(n23307), .B(n23308), .Z(n23253) );
  XOR U23193 ( .A(n23309), .B(n23300), .Z(n23308) );
  AND U23194 ( .A(n23265), .B(n23310), .Z(n23300) );
  AND U23195 ( .A(n23311), .B(n23312), .Z(n23309) );
  XOR U23196 ( .A(n23313), .B(n23307), .Z(n23311) );
  XNOR U23197 ( .A(n23250), .B(n23303), .Z(n23305) );
  XNOR U23198 ( .A(n23314), .B(n23315), .Z(n23250) );
  AND U23199 ( .A(n342), .B(n23257), .Z(n23315) );
  XOR U23200 ( .A(n23314), .B(n23255), .Z(n23257) );
  XOR U23201 ( .A(n23316), .B(n23317), .Z(n23303) );
  AND U23202 ( .A(n23318), .B(n23319), .Z(n23317) );
  XNOR U23203 ( .A(n23316), .B(n23265), .Z(n23319) );
  XOR U23204 ( .A(n23320), .B(n23312), .Z(n23265) );
  XNOR U23205 ( .A(n23321), .B(n23307), .Z(n23312) );
  XOR U23206 ( .A(n23322), .B(n23323), .Z(n23307) );
  AND U23207 ( .A(n23324), .B(n23325), .Z(n23323) );
  XOR U23208 ( .A(n23326), .B(n23322), .Z(n23324) );
  XNOR U23209 ( .A(n23327), .B(n23328), .Z(n23321) );
  AND U23210 ( .A(n23329), .B(n23330), .Z(n23328) );
  XOR U23211 ( .A(n23327), .B(n23331), .Z(n23329) );
  XNOR U23212 ( .A(n23313), .B(n23310), .Z(n23320) );
  AND U23213 ( .A(n23332), .B(n23333), .Z(n23310) );
  XOR U23214 ( .A(n23334), .B(n23335), .Z(n23313) );
  AND U23215 ( .A(n23336), .B(n23337), .Z(n23335) );
  XOR U23216 ( .A(n23334), .B(n23338), .Z(n23336) );
  XNOR U23217 ( .A(n23262), .B(n23316), .Z(n23318) );
  XNOR U23218 ( .A(n23339), .B(n23340), .Z(n23262) );
  AND U23219 ( .A(n342), .B(n23268), .Z(n23340) );
  XOR U23220 ( .A(n23339), .B(n23266), .Z(n23268) );
  XOR U23221 ( .A(n23341), .B(n23342), .Z(n23316) );
  AND U23222 ( .A(n23343), .B(n23344), .Z(n23342) );
  XNOR U23223 ( .A(n23341), .B(n23332), .Z(n23344) );
  IV U23224 ( .A(n23274), .Z(n23332) );
  XNOR U23225 ( .A(n23345), .B(n23325), .Z(n23274) );
  XNOR U23226 ( .A(n23346), .B(n23331), .Z(n23325) );
  XOR U23227 ( .A(n23347), .B(n23348), .Z(n23331) );
  AND U23228 ( .A(n23349), .B(n23350), .Z(n23348) );
  XOR U23229 ( .A(n23347), .B(n23351), .Z(n23349) );
  XNOR U23230 ( .A(n23330), .B(n23322), .Z(n23346) );
  XOR U23231 ( .A(n23352), .B(n23353), .Z(n23322) );
  AND U23232 ( .A(n23354), .B(n23355), .Z(n23353) );
  XNOR U23233 ( .A(n23356), .B(n23352), .Z(n23354) );
  XNOR U23234 ( .A(n23357), .B(n23327), .Z(n23330) );
  XOR U23235 ( .A(n23358), .B(n23359), .Z(n23327) );
  AND U23236 ( .A(n23360), .B(n23361), .Z(n23359) );
  XOR U23237 ( .A(n23358), .B(n23362), .Z(n23360) );
  XNOR U23238 ( .A(n23363), .B(n23364), .Z(n23357) );
  AND U23239 ( .A(n23365), .B(n23366), .Z(n23364) );
  XNOR U23240 ( .A(n23363), .B(n23367), .Z(n23365) );
  XNOR U23241 ( .A(n23326), .B(n23333), .Z(n23345) );
  AND U23242 ( .A(n23286), .B(n23368), .Z(n23333) );
  XOR U23243 ( .A(n23338), .B(n23337), .Z(n23326) );
  XNOR U23244 ( .A(n23369), .B(n23334), .Z(n23337) );
  XOR U23245 ( .A(n23370), .B(n23371), .Z(n23334) );
  AND U23246 ( .A(n23372), .B(n23373), .Z(n23371) );
  XOR U23247 ( .A(n23370), .B(n23374), .Z(n23372) );
  XNOR U23248 ( .A(n23375), .B(n23376), .Z(n23369) );
  AND U23249 ( .A(n23377), .B(n23378), .Z(n23376) );
  XOR U23250 ( .A(n23375), .B(n23379), .Z(n23377) );
  XOR U23251 ( .A(n23380), .B(n23381), .Z(n23338) );
  AND U23252 ( .A(n23382), .B(n23383), .Z(n23381) );
  XOR U23253 ( .A(n23380), .B(n23384), .Z(n23382) );
  XNOR U23254 ( .A(n23271), .B(n23341), .Z(n23343) );
  XNOR U23255 ( .A(n23385), .B(n23386), .Z(n23271) );
  AND U23256 ( .A(n342), .B(n23278), .Z(n23386) );
  XOR U23257 ( .A(n23385), .B(n23276), .Z(n23278) );
  XOR U23258 ( .A(n23387), .B(n23388), .Z(n23341) );
  AND U23259 ( .A(n23389), .B(n23390), .Z(n23388) );
  XNOR U23260 ( .A(n23387), .B(n23286), .Z(n23390) );
  XOR U23261 ( .A(n23391), .B(n23355), .Z(n23286) );
  XNOR U23262 ( .A(n23392), .B(n23362), .Z(n23355) );
  XOR U23263 ( .A(n23351), .B(n23350), .Z(n23362) );
  XNOR U23264 ( .A(n23393), .B(n23347), .Z(n23350) );
  XOR U23265 ( .A(n23394), .B(n23395), .Z(n23347) );
  AND U23266 ( .A(n23396), .B(n23397), .Z(n23395) );
  XOR U23267 ( .A(n23394), .B(n23398), .Z(n23396) );
  XNOR U23268 ( .A(n23399), .B(n23400), .Z(n23393) );
  NOR U23269 ( .A(n23401), .B(n23402), .Z(n23400) );
  XNOR U23270 ( .A(n23399), .B(n23403), .Z(n23401) );
  XOR U23271 ( .A(n23404), .B(n23405), .Z(n23351) );
  NOR U23272 ( .A(n23406), .B(n23407), .Z(n23405) );
  XNOR U23273 ( .A(n23404), .B(n23408), .Z(n23406) );
  XNOR U23274 ( .A(n23361), .B(n23352), .Z(n23392) );
  XOR U23275 ( .A(n23409), .B(n23410), .Z(n23352) );
  NOR U23276 ( .A(n23411), .B(n23412), .Z(n23410) );
  XNOR U23277 ( .A(n23409), .B(n23413), .Z(n23411) );
  XOR U23278 ( .A(n23414), .B(n23367), .Z(n23361) );
  XNOR U23279 ( .A(n23415), .B(n23416), .Z(n23367) );
  NOR U23280 ( .A(n23417), .B(n23418), .Z(n23416) );
  XNOR U23281 ( .A(n23415), .B(n23419), .Z(n23417) );
  XNOR U23282 ( .A(n23366), .B(n23358), .Z(n23414) );
  XOR U23283 ( .A(n23420), .B(n23421), .Z(n23358) );
  AND U23284 ( .A(n23422), .B(n23423), .Z(n23421) );
  XOR U23285 ( .A(n23420), .B(n23424), .Z(n23422) );
  XNOR U23286 ( .A(n23425), .B(n23363), .Z(n23366) );
  XOR U23287 ( .A(n23426), .B(n23427), .Z(n23363) );
  AND U23288 ( .A(n23428), .B(n23429), .Z(n23427) );
  XOR U23289 ( .A(n23426), .B(n23430), .Z(n23428) );
  XNOR U23290 ( .A(n23431), .B(n23432), .Z(n23425) );
  NOR U23291 ( .A(n23433), .B(n23434), .Z(n23432) );
  XOR U23292 ( .A(n23431), .B(n23435), .Z(n23433) );
  XOR U23293 ( .A(n23356), .B(n23368), .Z(n23391) );
  NOR U23294 ( .A(n23294), .B(n23436), .Z(n23368) );
  XNOR U23295 ( .A(n23374), .B(n23373), .Z(n23356) );
  XNOR U23296 ( .A(n23437), .B(n23379), .Z(n23373) );
  XOR U23297 ( .A(n23438), .B(n23439), .Z(n23379) );
  NOR U23298 ( .A(n23440), .B(n23441), .Z(n23439) );
  XNOR U23299 ( .A(n23438), .B(n23442), .Z(n23440) );
  XNOR U23300 ( .A(n23378), .B(n23370), .Z(n23437) );
  XOR U23301 ( .A(n23443), .B(n23444), .Z(n23370) );
  AND U23302 ( .A(n23445), .B(n23446), .Z(n23444) );
  XNOR U23303 ( .A(n23443), .B(n23447), .Z(n23445) );
  XNOR U23304 ( .A(n23448), .B(n23375), .Z(n23378) );
  XOR U23305 ( .A(n23449), .B(n23450), .Z(n23375) );
  AND U23306 ( .A(n23451), .B(n23452), .Z(n23450) );
  XOR U23307 ( .A(n23449), .B(n23453), .Z(n23451) );
  XNOR U23308 ( .A(n23454), .B(n23455), .Z(n23448) );
  NOR U23309 ( .A(n23456), .B(n23457), .Z(n23455) );
  XOR U23310 ( .A(n23454), .B(n23458), .Z(n23456) );
  XOR U23311 ( .A(n23384), .B(n23383), .Z(n23374) );
  XNOR U23312 ( .A(n23459), .B(n23380), .Z(n23383) );
  XOR U23313 ( .A(n23460), .B(n23461), .Z(n23380) );
  AND U23314 ( .A(n23462), .B(n23463), .Z(n23461) );
  XOR U23315 ( .A(n23460), .B(n23464), .Z(n23462) );
  XNOR U23316 ( .A(n23465), .B(n23466), .Z(n23459) );
  NOR U23317 ( .A(n23467), .B(n23468), .Z(n23466) );
  XNOR U23318 ( .A(n23465), .B(n23469), .Z(n23467) );
  XOR U23319 ( .A(n23470), .B(n23471), .Z(n23384) );
  NOR U23320 ( .A(n23472), .B(n23473), .Z(n23471) );
  XNOR U23321 ( .A(n23470), .B(n23474), .Z(n23472) );
  XNOR U23322 ( .A(n23283), .B(n23387), .Z(n23389) );
  XNOR U23323 ( .A(n23475), .B(n23476), .Z(n23283) );
  AND U23324 ( .A(n342), .B(n23290), .Z(n23476) );
  XOR U23325 ( .A(n23475), .B(n23288), .Z(n23290) );
  AND U23326 ( .A(n23291), .B(n23294), .Z(n23387) );
  XOR U23327 ( .A(n23477), .B(n23436), .Z(n23294) );
  XNOR U23328 ( .A(p_input[2048]), .B(p_input[800]), .Z(n23436) );
  XOR U23329 ( .A(n23413), .B(n23412), .Z(n23477) );
  XOR U23330 ( .A(n23478), .B(n23424), .Z(n23412) );
  XOR U23331 ( .A(n23398), .B(n23397), .Z(n23424) );
  XNOR U23332 ( .A(n23479), .B(n23403), .Z(n23397) );
  XOR U23333 ( .A(p_input[2072]), .B(p_input[824]), .Z(n23403) );
  XOR U23334 ( .A(n23394), .B(n23402), .Z(n23479) );
  XOR U23335 ( .A(n23480), .B(n23399), .Z(n23402) );
  XOR U23336 ( .A(p_input[2070]), .B(p_input[822]), .Z(n23399) );
  XNOR U23337 ( .A(p_input[2071]), .B(p_input[823]), .Z(n23480) );
  XNOR U23338 ( .A(n16727), .B(p_input[818]), .Z(n23394) );
  XNOR U23339 ( .A(n23408), .B(n23407), .Z(n23398) );
  XOR U23340 ( .A(n23481), .B(n23404), .Z(n23407) );
  XOR U23341 ( .A(p_input[2067]), .B(p_input[819]), .Z(n23404) );
  XNOR U23342 ( .A(p_input[2068]), .B(p_input[820]), .Z(n23481) );
  XOR U23343 ( .A(p_input[2069]), .B(p_input[821]), .Z(n23408) );
  XNOR U23344 ( .A(n23423), .B(n23409), .Z(n23478) );
  XNOR U23345 ( .A(n16729), .B(p_input[801]), .Z(n23409) );
  XNOR U23346 ( .A(n23482), .B(n23430), .Z(n23423) );
  XNOR U23347 ( .A(n23419), .B(n23418), .Z(n23430) );
  XOR U23348 ( .A(n23483), .B(n23415), .Z(n23418) );
  XNOR U23349 ( .A(n16444), .B(p_input[826]), .Z(n23415) );
  XNOR U23350 ( .A(p_input[2075]), .B(p_input[827]), .Z(n23483) );
  XOR U23351 ( .A(p_input[2076]), .B(p_input[828]), .Z(n23419) );
  XNOR U23352 ( .A(n23429), .B(n23420), .Z(n23482) );
  XNOR U23353 ( .A(n16732), .B(p_input[817]), .Z(n23420) );
  XOR U23354 ( .A(n23484), .B(n23435), .Z(n23429) );
  XNOR U23355 ( .A(p_input[2079]), .B(p_input[831]), .Z(n23435) );
  XOR U23356 ( .A(n23426), .B(n23434), .Z(n23484) );
  XOR U23357 ( .A(n23485), .B(n23431), .Z(n23434) );
  XOR U23358 ( .A(p_input[2077]), .B(p_input[829]), .Z(n23431) );
  XNOR U23359 ( .A(p_input[2078]), .B(p_input[830]), .Z(n23485) );
  XNOR U23360 ( .A(n16448), .B(p_input[825]), .Z(n23426) );
  XNOR U23361 ( .A(n23447), .B(n23446), .Z(n23413) );
  XNOR U23362 ( .A(n23486), .B(n23453), .Z(n23446) );
  XNOR U23363 ( .A(n23442), .B(n23441), .Z(n23453) );
  XOR U23364 ( .A(n23487), .B(n23438), .Z(n23441) );
  XNOR U23365 ( .A(n16737), .B(p_input[811]), .Z(n23438) );
  XNOR U23366 ( .A(p_input[2060]), .B(p_input[812]), .Z(n23487) );
  XOR U23367 ( .A(p_input[2061]), .B(p_input[813]), .Z(n23442) );
  XNOR U23368 ( .A(n23452), .B(n23443), .Z(n23486) );
  XNOR U23369 ( .A(n16452), .B(p_input[802]), .Z(n23443) );
  XOR U23370 ( .A(n23488), .B(n23458), .Z(n23452) );
  XNOR U23371 ( .A(p_input[2064]), .B(p_input[816]), .Z(n23458) );
  XOR U23372 ( .A(n23449), .B(n23457), .Z(n23488) );
  XOR U23373 ( .A(n23489), .B(n23454), .Z(n23457) );
  XOR U23374 ( .A(p_input[2062]), .B(p_input[814]), .Z(n23454) );
  XNOR U23375 ( .A(p_input[2063]), .B(p_input[815]), .Z(n23489) );
  XNOR U23376 ( .A(n16740), .B(p_input[810]), .Z(n23449) );
  XNOR U23377 ( .A(n23464), .B(n23463), .Z(n23447) );
  XNOR U23378 ( .A(n23490), .B(n23469), .Z(n23463) );
  XOR U23379 ( .A(p_input[2057]), .B(p_input[809]), .Z(n23469) );
  XOR U23380 ( .A(n23460), .B(n23468), .Z(n23490) );
  XOR U23381 ( .A(n23491), .B(n23465), .Z(n23468) );
  XOR U23382 ( .A(p_input[2055]), .B(p_input[807]), .Z(n23465) );
  XNOR U23383 ( .A(p_input[2056]), .B(p_input[808]), .Z(n23491) );
  XNOR U23384 ( .A(n16459), .B(p_input[803]), .Z(n23460) );
  XNOR U23385 ( .A(n23474), .B(n23473), .Z(n23464) );
  XOR U23386 ( .A(n23492), .B(n23470), .Z(n23473) );
  XOR U23387 ( .A(p_input[2052]), .B(p_input[804]), .Z(n23470) );
  XNOR U23388 ( .A(p_input[2053]), .B(p_input[805]), .Z(n23492) );
  XOR U23389 ( .A(p_input[2054]), .B(p_input[806]), .Z(n23474) );
  XNOR U23390 ( .A(n23493), .B(n23494), .Z(n23291) );
  AND U23391 ( .A(n342), .B(n23495), .Z(n23494) );
  XNOR U23392 ( .A(n23496), .B(n23497), .Z(n342) );
  AND U23393 ( .A(n23498), .B(n23499), .Z(n23497) );
  XOR U23394 ( .A(n23496), .B(n23301), .Z(n23499) );
  XNOR U23395 ( .A(n23496), .B(n23243), .Z(n23498) );
  XOR U23396 ( .A(n23500), .B(n23501), .Z(n23496) );
  AND U23397 ( .A(n23502), .B(n23503), .Z(n23501) );
  XNOR U23398 ( .A(n23314), .B(n23500), .Z(n23503) );
  XOR U23399 ( .A(n23500), .B(n23255), .Z(n23502) );
  XOR U23400 ( .A(n23504), .B(n23505), .Z(n23500) );
  AND U23401 ( .A(n23506), .B(n23507), .Z(n23505) );
  XNOR U23402 ( .A(n23339), .B(n23504), .Z(n23507) );
  XOR U23403 ( .A(n23504), .B(n23266), .Z(n23506) );
  XOR U23404 ( .A(n23508), .B(n23509), .Z(n23504) );
  AND U23405 ( .A(n23510), .B(n23511), .Z(n23509) );
  XOR U23406 ( .A(n23508), .B(n23276), .Z(n23510) );
  XOR U23407 ( .A(n23512), .B(n23513), .Z(n23232) );
  AND U23408 ( .A(n346), .B(n23495), .Z(n23513) );
  XNOR U23409 ( .A(n23493), .B(n23512), .Z(n23495) );
  XNOR U23410 ( .A(n23514), .B(n23515), .Z(n346) );
  AND U23411 ( .A(n23516), .B(n23517), .Z(n23515) );
  XNOR U23412 ( .A(n23518), .B(n23514), .Z(n23517) );
  IV U23413 ( .A(n23301), .Z(n23518) );
  XNOR U23414 ( .A(n23519), .B(n23520), .Z(n23301) );
  AND U23415 ( .A(n349), .B(n23521), .Z(n23520) );
  XNOR U23416 ( .A(n23519), .B(n23522), .Z(n23521) );
  XNOR U23417 ( .A(n23243), .B(n23514), .Z(n23516) );
  XOR U23418 ( .A(n23523), .B(n23524), .Z(n23243) );
  AND U23419 ( .A(n357), .B(n23525), .Z(n23524) );
  XOR U23420 ( .A(n23526), .B(n23527), .Z(n23514) );
  AND U23421 ( .A(n23528), .B(n23529), .Z(n23527) );
  XNOR U23422 ( .A(n23526), .B(n23314), .Z(n23529) );
  XNOR U23423 ( .A(n23530), .B(n23531), .Z(n23314) );
  AND U23424 ( .A(n349), .B(n23532), .Z(n23531) );
  XOR U23425 ( .A(n23533), .B(n23530), .Z(n23532) );
  XNOR U23426 ( .A(n23534), .B(n23526), .Z(n23528) );
  IV U23427 ( .A(n23255), .Z(n23534) );
  XOR U23428 ( .A(n23535), .B(n23536), .Z(n23255) );
  AND U23429 ( .A(n357), .B(n23537), .Z(n23536) );
  XOR U23430 ( .A(n23538), .B(n23539), .Z(n23526) );
  AND U23431 ( .A(n23540), .B(n23541), .Z(n23539) );
  XNOR U23432 ( .A(n23538), .B(n23339), .Z(n23541) );
  XNOR U23433 ( .A(n23542), .B(n23543), .Z(n23339) );
  AND U23434 ( .A(n349), .B(n23544), .Z(n23543) );
  XNOR U23435 ( .A(n23545), .B(n23542), .Z(n23544) );
  XOR U23436 ( .A(n23266), .B(n23538), .Z(n23540) );
  XOR U23437 ( .A(n23546), .B(n23547), .Z(n23266) );
  AND U23438 ( .A(n357), .B(n23548), .Z(n23547) );
  XOR U23439 ( .A(n23508), .B(n23549), .Z(n23538) );
  AND U23440 ( .A(n23550), .B(n23511), .Z(n23549) );
  XNOR U23441 ( .A(n23385), .B(n23508), .Z(n23511) );
  XNOR U23442 ( .A(n23551), .B(n23552), .Z(n23385) );
  AND U23443 ( .A(n349), .B(n23553), .Z(n23552) );
  XOR U23444 ( .A(n23554), .B(n23551), .Z(n23553) );
  XNOR U23445 ( .A(n23555), .B(n23508), .Z(n23550) );
  IV U23446 ( .A(n23276), .Z(n23555) );
  XOR U23447 ( .A(n23556), .B(n23557), .Z(n23276) );
  AND U23448 ( .A(n357), .B(n23558), .Z(n23557) );
  XOR U23449 ( .A(n23559), .B(n23560), .Z(n23508) );
  AND U23450 ( .A(n23561), .B(n23562), .Z(n23560) );
  XNOR U23451 ( .A(n23559), .B(n23475), .Z(n23562) );
  XNOR U23452 ( .A(n23563), .B(n23564), .Z(n23475) );
  AND U23453 ( .A(n349), .B(n23565), .Z(n23564) );
  XNOR U23454 ( .A(n23566), .B(n23563), .Z(n23565) );
  XNOR U23455 ( .A(n23567), .B(n23559), .Z(n23561) );
  IV U23456 ( .A(n23288), .Z(n23567) );
  XOR U23457 ( .A(n23568), .B(n23569), .Z(n23288) );
  AND U23458 ( .A(n357), .B(n23570), .Z(n23569) );
  AND U23459 ( .A(n23512), .B(n23493), .Z(n23559) );
  XNOR U23460 ( .A(n23571), .B(n23572), .Z(n23493) );
  AND U23461 ( .A(n349), .B(n23573), .Z(n23572) );
  XNOR U23462 ( .A(n23574), .B(n23571), .Z(n23573) );
  XNOR U23463 ( .A(n23575), .B(n23576), .Z(n349) );
  AND U23464 ( .A(n23577), .B(n23578), .Z(n23576) );
  XOR U23465 ( .A(n23522), .B(n23575), .Z(n23578) );
  AND U23466 ( .A(n23579), .B(n23580), .Z(n23522) );
  XOR U23467 ( .A(n23575), .B(n23519), .Z(n23577) );
  XNOR U23468 ( .A(n23581), .B(n23582), .Z(n23519) );
  AND U23469 ( .A(n353), .B(n23525), .Z(n23582) );
  XOR U23470 ( .A(n23523), .B(n23581), .Z(n23525) );
  XOR U23471 ( .A(n23583), .B(n23584), .Z(n23575) );
  AND U23472 ( .A(n23585), .B(n23586), .Z(n23584) );
  XNOR U23473 ( .A(n23583), .B(n23579), .Z(n23586) );
  IV U23474 ( .A(n23533), .Z(n23579) );
  XOR U23475 ( .A(n23587), .B(n23588), .Z(n23533) );
  XOR U23476 ( .A(n23589), .B(n23580), .Z(n23588) );
  AND U23477 ( .A(n23545), .B(n23590), .Z(n23580) );
  AND U23478 ( .A(n23591), .B(n23592), .Z(n23589) );
  XOR U23479 ( .A(n23593), .B(n23587), .Z(n23591) );
  XNOR U23480 ( .A(n23530), .B(n23583), .Z(n23585) );
  XNOR U23481 ( .A(n23594), .B(n23595), .Z(n23530) );
  AND U23482 ( .A(n353), .B(n23537), .Z(n23595) );
  XOR U23483 ( .A(n23594), .B(n23535), .Z(n23537) );
  XOR U23484 ( .A(n23596), .B(n23597), .Z(n23583) );
  AND U23485 ( .A(n23598), .B(n23599), .Z(n23597) );
  XNOR U23486 ( .A(n23596), .B(n23545), .Z(n23599) );
  XOR U23487 ( .A(n23600), .B(n23592), .Z(n23545) );
  XNOR U23488 ( .A(n23601), .B(n23587), .Z(n23592) );
  XOR U23489 ( .A(n23602), .B(n23603), .Z(n23587) );
  AND U23490 ( .A(n23604), .B(n23605), .Z(n23603) );
  XOR U23491 ( .A(n23606), .B(n23602), .Z(n23604) );
  XNOR U23492 ( .A(n23607), .B(n23608), .Z(n23601) );
  AND U23493 ( .A(n23609), .B(n23610), .Z(n23608) );
  XOR U23494 ( .A(n23607), .B(n23611), .Z(n23609) );
  XNOR U23495 ( .A(n23593), .B(n23590), .Z(n23600) );
  AND U23496 ( .A(n23612), .B(n23613), .Z(n23590) );
  XOR U23497 ( .A(n23614), .B(n23615), .Z(n23593) );
  AND U23498 ( .A(n23616), .B(n23617), .Z(n23615) );
  XOR U23499 ( .A(n23614), .B(n23618), .Z(n23616) );
  XNOR U23500 ( .A(n23542), .B(n23596), .Z(n23598) );
  XNOR U23501 ( .A(n23619), .B(n23620), .Z(n23542) );
  AND U23502 ( .A(n353), .B(n23548), .Z(n23620) );
  XOR U23503 ( .A(n23619), .B(n23546), .Z(n23548) );
  XOR U23504 ( .A(n23621), .B(n23622), .Z(n23596) );
  AND U23505 ( .A(n23623), .B(n23624), .Z(n23622) );
  XNOR U23506 ( .A(n23621), .B(n23612), .Z(n23624) );
  IV U23507 ( .A(n23554), .Z(n23612) );
  XNOR U23508 ( .A(n23625), .B(n23605), .Z(n23554) );
  XNOR U23509 ( .A(n23626), .B(n23611), .Z(n23605) );
  XOR U23510 ( .A(n23627), .B(n23628), .Z(n23611) );
  AND U23511 ( .A(n23629), .B(n23630), .Z(n23628) );
  XOR U23512 ( .A(n23627), .B(n23631), .Z(n23629) );
  XNOR U23513 ( .A(n23610), .B(n23602), .Z(n23626) );
  XOR U23514 ( .A(n23632), .B(n23633), .Z(n23602) );
  AND U23515 ( .A(n23634), .B(n23635), .Z(n23633) );
  XNOR U23516 ( .A(n23636), .B(n23632), .Z(n23634) );
  XNOR U23517 ( .A(n23637), .B(n23607), .Z(n23610) );
  XOR U23518 ( .A(n23638), .B(n23639), .Z(n23607) );
  AND U23519 ( .A(n23640), .B(n23641), .Z(n23639) );
  XOR U23520 ( .A(n23638), .B(n23642), .Z(n23640) );
  XNOR U23521 ( .A(n23643), .B(n23644), .Z(n23637) );
  AND U23522 ( .A(n23645), .B(n23646), .Z(n23644) );
  XNOR U23523 ( .A(n23643), .B(n23647), .Z(n23645) );
  XNOR U23524 ( .A(n23606), .B(n23613), .Z(n23625) );
  AND U23525 ( .A(n23566), .B(n23648), .Z(n23613) );
  XOR U23526 ( .A(n23618), .B(n23617), .Z(n23606) );
  XNOR U23527 ( .A(n23649), .B(n23614), .Z(n23617) );
  XOR U23528 ( .A(n23650), .B(n23651), .Z(n23614) );
  AND U23529 ( .A(n23652), .B(n23653), .Z(n23651) );
  XOR U23530 ( .A(n23650), .B(n23654), .Z(n23652) );
  XNOR U23531 ( .A(n23655), .B(n23656), .Z(n23649) );
  AND U23532 ( .A(n23657), .B(n23658), .Z(n23656) );
  XOR U23533 ( .A(n23655), .B(n23659), .Z(n23657) );
  XOR U23534 ( .A(n23660), .B(n23661), .Z(n23618) );
  AND U23535 ( .A(n23662), .B(n23663), .Z(n23661) );
  XOR U23536 ( .A(n23660), .B(n23664), .Z(n23662) );
  XNOR U23537 ( .A(n23551), .B(n23621), .Z(n23623) );
  XNOR U23538 ( .A(n23665), .B(n23666), .Z(n23551) );
  AND U23539 ( .A(n353), .B(n23558), .Z(n23666) );
  XOR U23540 ( .A(n23665), .B(n23556), .Z(n23558) );
  XOR U23541 ( .A(n23667), .B(n23668), .Z(n23621) );
  AND U23542 ( .A(n23669), .B(n23670), .Z(n23668) );
  XNOR U23543 ( .A(n23667), .B(n23566), .Z(n23670) );
  XOR U23544 ( .A(n23671), .B(n23635), .Z(n23566) );
  XNOR U23545 ( .A(n23672), .B(n23642), .Z(n23635) );
  XOR U23546 ( .A(n23631), .B(n23630), .Z(n23642) );
  XNOR U23547 ( .A(n23673), .B(n23627), .Z(n23630) );
  XOR U23548 ( .A(n23674), .B(n23675), .Z(n23627) );
  AND U23549 ( .A(n23676), .B(n23677), .Z(n23675) );
  XOR U23550 ( .A(n23674), .B(n23678), .Z(n23676) );
  XNOR U23551 ( .A(n23679), .B(n23680), .Z(n23673) );
  NOR U23552 ( .A(n23681), .B(n23682), .Z(n23680) );
  XNOR U23553 ( .A(n23679), .B(n23683), .Z(n23681) );
  XOR U23554 ( .A(n23684), .B(n23685), .Z(n23631) );
  NOR U23555 ( .A(n23686), .B(n23687), .Z(n23685) );
  XNOR U23556 ( .A(n23684), .B(n23688), .Z(n23686) );
  XNOR U23557 ( .A(n23641), .B(n23632), .Z(n23672) );
  XOR U23558 ( .A(n23689), .B(n23690), .Z(n23632) );
  NOR U23559 ( .A(n23691), .B(n23692), .Z(n23690) );
  XNOR U23560 ( .A(n23689), .B(n23693), .Z(n23691) );
  XOR U23561 ( .A(n23694), .B(n23647), .Z(n23641) );
  XNOR U23562 ( .A(n23695), .B(n23696), .Z(n23647) );
  NOR U23563 ( .A(n23697), .B(n23698), .Z(n23696) );
  XNOR U23564 ( .A(n23695), .B(n23699), .Z(n23697) );
  XNOR U23565 ( .A(n23646), .B(n23638), .Z(n23694) );
  XOR U23566 ( .A(n23700), .B(n23701), .Z(n23638) );
  AND U23567 ( .A(n23702), .B(n23703), .Z(n23701) );
  XOR U23568 ( .A(n23700), .B(n23704), .Z(n23702) );
  XNOR U23569 ( .A(n23705), .B(n23643), .Z(n23646) );
  XOR U23570 ( .A(n23706), .B(n23707), .Z(n23643) );
  AND U23571 ( .A(n23708), .B(n23709), .Z(n23707) );
  XOR U23572 ( .A(n23706), .B(n23710), .Z(n23708) );
  XNOR U23573 ( .A(n23711), .B(n23712), .Z(n23705) );
  NOR U23574 ( .A(n23713), .B(n23714), .Z(n23712) );
  XOR U23575 ( .A(n23711), .B(n23715), .Z(n23713) );
  XOR U23576 ( .A(n23636), .B(n23648), .Z(n23671) );
  NOR U23577 ( .A(n23574), .B(n23716), .Z(n23648) );
  XNOR U23578 ( .A(n23654), .B(n23653), .Z(n23636) );
  XNOR U23579 ( .A(n23717), .B(n23659), .Z(n23653) );
  XOR U23580 ( .A(n23718), .B(n23719), .Z(n23659) );
  NOR U23581 ( .A(n23720), .B(n23721), .Z(n23719) );
  XNOR U23582 ( .A(n23718), .B(n23722), .Z(n23720) );
  XNOR U23583 ( .A(n23658), .B(n23650), .Z(n23717) );
  XOR U23584 ( .A(n23723), .B(n23724), .Z(n23650) );
  AND U23585 ( .A(n23725), .B(n23726), .Z(n23724) );
  XNOR U23586 ( .A(n23723), .B(n23727), .Z(n23725) );
  XNOR U23587 ( .A(n23728), .B(n23655), .Z(n23658) );
  XOR U23588 ( .A(n23729), .B(n23730), .Z(n23655) );
  AND U23589 ( .A(n23731), .B(n23732), .Z(n23730) );
  XOR U23590 ( .A(n23729), .B(n23733), .Z(n23731) );
  XNOR U23591 ( .A(n23734), .B(n23735), .Z(n23728) );
  NOR U23592 ( .A(n23736), .B(n23737), .Z(n23735) );
  XOR U23593 ( .A(n23734), .B(n23738), .Z(n23736) );
  XOR U23594 ( .A(n23664), .B(n23663), .Z(n23654) );
  XNOR U23595 ( .A(n23739), .B(n23660), .Z(n23663) );
  XOR U23596 ( .A(n23740), .B(n23741), .Z(n23660) );
  AND U23597 ( .A(n23742), .B(n23743), .Z(n23741) );
  XOR U23598 ( .A(n23740), .B(n23744), .Z(n23742) );
  XNOR U23599 ( .A(n23745), .B(n23746), .Z(n23739) );
  NOR U23600 ( .A(n23747), .B(n23748), .Z(n23746) );
  XNOR U23601 ( .A(n23745), .B(n23749), .Z(n23747) );
  XOR U23602 ( .A(n23750), .B(n23751), .Z(n23664) );
  NOR U23603 ( .A(n23752), .B(n23753), .Z(n23751) );
  XNOR U23604 ( .A(n23750), .B(n23754), .Z(n23752) );
  XNOR U23605 ( .A(n23563), .B(n23667), .Z(n23669) );
  XNOR U23606 ( .A(n23755), .B(n23756), .Z(n23563) );
  AND U23607 ( .A(n353), .B(n23570), .Z(n23756) );
  XOR U23608 ( .A(n23755), .B(n23568), .Z(n23570) );
  AND U23609 ( .A(n23571), .B(n23574), .Z(n23667) );
  XOR U23610 ( .A(n23757), .B(n23716), .Z(n23574) );
  XNOR U23611 ( .A(p_input[2048]), .B(p_input[832]), .Z(n23716) );
  XOR U23612 ( .A(n23693), .B(n23692), .Z(n23757) );
  XOR U23613 ( .A(n23758), .B(n23704), .Z(n23692) );
  XOR U23614 ( .A(n23678), .B(n23677), .Z(n23704) );
  XNOR U23615 ( .A(n23759), .B(n23683), .Z(n23677) );
  XOR U23616 ( .A(p_input[2072]), .B(p_input[856]), .Z(n23683) );
  XOR U23617 ( .A(n23674), .B(n23682), .Z(n23759) );
  XOR U23618 ( .A(n23760), .B(n23679), .Z(n23682) );
  XOR U23619 ( .A(p_input[2070]), .B(p_input[854]), .Z(n23679) );
  XNOR U23620 ( .A(p_input[2071]), .B(p_input[855]), .Z(n23760) );
  XNOR U23621 ( .A(n16727), .B(p_input[850]), .Z(n23674) );
  XNOR U23622 ( .A(n23688), .B(n23687), .Z(n23678) );
  XOR U23623 ( .A(n23761), .B(n23684), .Z(n23687) );
  XOR U23624 ( .A(p_input[2067]), .B(p_input[851]), .Z(n23684) );
  XNOR U23625 ( .A(p_input[2068]), .B(p_input[852]), .Z(n23761) );
  XOR U23626 ( .A(p_input[2069]), .B(p_input[853]), .Z(n23688) );
  XNOR U23627 ( .A(n23703), .B(n23689), .Z(n23758) );
  XNOR U23628 ( .A(n16729), .B(p_input[833]), .Z(n23689) );
  XNOR U23629 ( .A(n23762), .B(n23710), .Z(n23703) );
  XNOR U23630 ( .A(n23699), .B(n23698), .Z(n23710) );
  XOR U23631 ( .A(n23763), .B(n23695), .Z(n23698) );
  XNOR U23632 ( .A(n16444), .B(p_input[858]), .Z(n23695) );
  XNOR U23633 ( .A(p_input[2075]), .B(p_input[859]), .Z(n23763) );
  XOR U23634 ( .A(p_input[2076]), .B(p_input[860]), .Z(n23699) );
  XNOR U23635 ( .A(n23709), .B(n23700), .Z(n23762) );
  XNOR U23636 ( .A(n16732), .B(p_input[849]), .Z(n23700) );
  XOR U23637 ( .A(n23764), .B(n23715), .Z(n23709) );
  XNOR U23638 ( .A(p_input[2079]), .B(p_input[863]), .Z(n23715) );
  XOR U23639 ( .A(n23706), .B(n23714), .Z(n23764) );
  XOR U23640 ( .A(n23765), .B(n23711), .Z(n23714) );
  XOR U23641 ( .A(p_input[2077]), .B(p_input[861]), .Z(n23711) );
  XNOR U23642 ( .A(p_input[2078]), .B(p_input[862]), .Z(n23765) );
  XNOR U23643 ( .A(n16448), .B(p_input[857]), .Z(n23706) );
  XNOR U23644 ( .A(n23727), .B(n23726), .Z(n23693) );
  XNOR U23645 ( .A(n23766), .B(n23733), .Z(n23726) );
  XNOR U23646 ( .A(n23722), .B(n23721), .Z(n23733) );
  XOR U23647 ( .A(n23767), .B(n23718), .Z(n23721) );
  XNOR U23648 ( .A(n16737), .B(p_input[843]), .Z(n23718) );
  XNOR U23649 ( .A(p_input[2060]), .B(p_input[844]), .Z(n23767) );
  XOR U23650 ( .A(p_input[2061]), .B(p_input[845]), .Z(n23722) );
  XNOR U23651 ( .A(n23732), .B(n23723), .Z(n23766) );
  XNOR U23652 ( .A(n16452), .B(p_input[834]), .Z(n23723) );
  XOR U23653 ( .A(n23768), .B(n23738), .Z(n23732) );
  XNOR U23654 ( .A(p_input[2064]), .B(p_input[848]), .Z(n23738) );
  XOR U23655 ( .A(n23729), .B(n23737), .Z(n23768) );
  XOR U23656 ( .A(n23769), .B(n23734), .Z(n23737) );
  XOR U23657 ( .A(p_input[2062]), .B(p_input[846]), .Z(n23734) );
  XNOR U23658 ( .A(p_input[2063]), .B(p_input[847]), .Z(n23769) );
  XNOR U23659 ( .A(n16740), .B(p_input[842]), .Z(n23729) );
  XNOR U23660 ( .A(n23744), .B(n23743), .Z(n23727) );
  XNOR U23661 ( .A(n23770), .B(n23749), .Z(n23743) );
  XOR U23662 ( .A(p_input[2057]), .B(p_input[841]), .Z(n23749) );
  XOR U23663 ( .A(n23740), .B(n23748), .Z(n23770) );
  XOR U23664 ( .A(n23771), .B(n23745), .Z(n23748) );
  XOR U23665 ( .A(p_input[2055]), .B(p_input[839]), .Z(n23745) );
  XNOR U23666 ( .A(p_input[2056]), .B(p_input[840]), .Z(n23771) );
  XNOR U23667 ( .A(n16459), .B(p_input[835]), .Z(n23740) );
  XNOR U23668 ( .A(n23754), .B(n23753), .Z(n23744) );
  XOR U23669 ( .A(n23772), .B(n23750), .Z(n23753) );
  XOR U23670 ( .A(p_input[2052]), .B(p_input[836]), .Z(n23750) );
  XNOR U23671 ( .A(p_input[2053]), .B(p_input[837]), .Z(n23772) );
  XOR U23672 ( .A(p_input[2054]), .B(p_input[838]), .Z(n23754) );
  XNOR U23673 ( .A(n23773), .B(n23774), .Z(n23571) );
  AND U23674 ( .A(n353), .B(n23775), .Z(n23774) );
  XNOR U23675 ( .A(n23776), .B(n23777), .Z(n353) );
  AND U23676 ( .A(n23778), .B(n23779), .Z(n23777) );
  XOR U23677 ( .A(n23776), .B(n23581), .Z(n23779) );
  XNOR U23678 ( .A(n23776), .B(n23523), .Z(n23778) );
  XOR U23679 ( .A(n23780), .B(n23781), .Z(n23776) );
  AND U23680 ( .A(n23782), .B(n23783), .Z(n23781) );
  XNOR U23681 ( .A(n23594), .B(n23780), .Z(n23783) );
  XOR U23682 ( .A(n23780), .B(n23535), .Z(n23782) );
  XOR U23683 ( .A(n23784), .B(n23785), .Z(n23780) );
  AND U23684 ( .A(n23786), .B(n23787), .Z(n23785) );
  XNOR U23685 ( .A(n23619), .B(n23784), .Z(n23787) );
  XOR U23686 ( .A(n23784), .B(n23546), .Z(n23786) );
  XOR U23687 ( .A(n23788), .B(n23789), .Z(n23784) );
  AND U23688 ( .A(n23790), .B(n23791), .Z(n23789) );
  XOR U23689 ( .A(n23788), .B(n23556), .Z(n23790) );
  XOR U23690 ( .A(n23792), .B(n23793), .Z(n23512) );
  AND U23691 ( .A(n357), .B(n23775), .Z(n23793) );
  XNOR U23692 ( .A(n23773), .B(n23792), .Z(n23775) );
  XNOR U23693 ( .A(n23794), .B(n23795), .Z(n357) );
  AND U23694 ( .A(n23796), .B(n23797), .Z(n23795) );
  XNOR U23695 ( .A(n23798), .B(n23794), .Z(n23797) );
  IV U23696 ( .A(n23581), .Z(n23798) );
  XNOR U23697 ( .A(n23799), .B(n23800), .Z(n23581) );
  AND U23698 ( .A(n360), .B(n23801), .Z(n23800) );
  XNOR U23699 ( .A(n23799), .B(n23802), .Z(n23801) );
  XNOR U23700 ( .A(n23523), .B(n23794), .Z(n23796) );
  XOR U23701 ( .A(n23803), .B(n23804), .Z(n23523) );
  AND U23702 ( .A(n368), .B(n23805), .Z(n23804) );
  XOR U23703 ( .A(n23806), .B(n23807), .Z(n23794) );
  AND U23704 ( .A(n23808), .B(n23809), .Z(n23807) );
  XNOR U23705 ( .A(n23806), .B(n23594), .Z(n23809) );
  XNOR U23706 ( .A(n23810), .B(n23811), .Z(n23594) );
  AND U23707 ( .A(n360), .B(n23812), .Z(n23811) );
  XOR U23708 ( .A(n23813), .B(n23810), .Z(n23812) );
  XNOR U23709 ( .A(n23814), .B(n23806), .Z(n23808) );
  IV U23710 ( .A(n23535), .Z(n23814) );
  XOR U23711 ( .A(n23815), .B(n23816), .Z(n23535) );
  AND U23712 ( .A(n368), .B(n23817), .Z(n23816) );
  XOR U23713 ( .A(n23818), .B(n23819), .Z(n23806) );
  AND U23714 ( .A(n23820), .B(n23821), .Z(n23819) );
  XNOR U23715 ( .A(n23818), .B(n23619), .Z(n23821) );
  XNOR U23716 ( .A(n23822), .B(n23823), .Z(n23619) );
  AND U23717 ( .A(n360), .B(n23824), .Z(n23823) );
  XNOR U23718 ( .A(n23825), .B(n23822), .Z(n23824) );
  XOR U23719 ( .A(n23546), .B(n23818), .Z(n23820) );
  XOR U23720 ( .A(n23826), .B(n23827), .Z(n23546) );
  AND U23721 ( .A(n368), .B(n23828), .Z(n23827) );
  XOR U23722 ( .A(n23788), .B(n23829), .Z(n23818) );
  AND U23723 ( .A(n23830), .B(n23791), .Z(n23829) );
  XNOR U23724 ( .A(n23665), .B(n23788), .Z(n23791) );
  XNOR U23725 ( .A(n23831), .B(n23832), .Z(n23665) );
  AND U23726 ( .A(n360), .B(n23833), .Z(n23832) );
  XOR U23727 ( .A(n23834), .B(n23831), .Z(n23833) );
  XNOR U23728 ( .A(n23835), .B(n23788), .Z(n23830) );
  IV U23729 ( .A(n23556), .Z(n23835) );
  XOR U23730 ( .A(n23836), .B(n23837), .Z(n23556) );
  AND U23731 ( .A(n368), .B(n23838), .Z(n23837) );
  XOR U23732 ( .A(n23839), .B(n23840), .Z(n23788) );
  AND U23733 ( .A(n23841), .B(n23842), .Z(n23840) );
  XNOR U23734 ( .A(n23839), .B(n23755), .Z(n23842) );
  XNOR U23735 ( .A(n23843), .B(n23844), .Z(n23755) );
  AND U23736 ( .A(n360), .B(n23845), .Z(n23844) );
  XNOR U23737 ( .A(n23846), .B(n23843), .Z(n23845) );
  XNOR U23738 ( .A(n23847), .B(n23839), .Z(n23841) );
  IV U23739 ( .A(n23568), .Z(n23847) );
  XOR U23740 ( .A(n23848), .B(n23849), .Z(n23568) );
  AND U23741 ( .A(n368), .B(n23850), .Z(n23849) );
  AND U23742 ( .A(n23792), .B(n23773), .Z(n23839) );
  XNOR U23743 ( .A(n23851), .B(n23852), .Z(n23773) );
  AND U23744 ( .A(n360), .B(n23853), .Z(n23852) );
  XNOR U23745 ( .A(n23854), .B(n23851), .Z(n23853) );
  XNOR U23746 ( .A(n23855), .B(n23856), .Z(n360) );
  AND U23747 ( .A(n23857), .B(n23858), .Z(n23856) );
  XOR U23748 ( .A(n23802), .B(n23855), .Z(n23858) );
  AND U23749 ( .A(n23859), .B(n23860), .Z(n23802) );
  XOR U23750 ( .A(n23855), .B(n23799), .Z(n23857) );
  XNOR U23751 ( .A(n23861), .B(n23862), .Z(n23799) );
  AND U23752 ( .A(n364), .B(n23805), .Z(n23862) );
  XOR U23753 ( .A(n23803), .B(n23861), .Z(n23805) );
  XOR U23754 ( .A(n23863), .B(n23864), .Z(n23855) );
  AND U23755 ( .A(n23865), .B(n23866), .Z(n23864) );
  XNOR U23756 ( .A(n23863), .B(n23859), .Z(n23866) );
  IV U23757 ( .A(n23813), .Z(n23859) );
  XOR U23758 ( .A(n23867), .B(n23868), .Z(n23813) );
  XOR U23759 ( .A(n23869), .B(n23860), .Z(n23868) );
  AND U23760 ( .A(n23825), .B(n23870), .Z(n23860) );
  AND U23761 ( .A(n23871), .B(n23872), .Z(n23869) );
  XOR U23762 ( .A(n23873), .B(n23867), .Z(n23871) );
  XNOR U23763 ( .A(n23810), .B(n23863), .Z(n23865) );
  XNOR U23764 ( .A(n23874), .B(n23875), .Z(n23810) );
  AND U23765 ( .A(n364), .B(n23817), .Z(n23875) );
  XOR U23766 ( .A(n23874), .B(n23815), .Z(n23817) );
  XOR U23767 ( .A(n23876), .B(n23877), .Z(n23863) );
  AND U23768 ( .A(n23878), .B(n23879), .Z(n23877) );
  XNOR U23769 ( .A(n23876), .B(n23825), .Z(n23879) );
  XOR U23770 ( .A(n23880), .B(n23872), .Z(n23825) );
  XNOR U23771 ( .A(n23881), .B(n23867), .Z(n23872) );
  XOR U23772 ( .A(n23882), .B(n23883), .Z(n23867) );
  AND U23773 ( .A(n23884), .B(n23885), .Z(n23883) );
  XOR U23774 ( .A(n23886), .B(n23882), .Z(n23884) );
  XNOR U23775 ( .A(n23887), .B(n23888), .Z(n23881) );
  AND U23776 ( .A(n23889), .B(n23890), .Z(n23888) );
  XOR U23777 ( .A(n23887), .B(n23891), .Z(n23889) );
  XNOR U23778 ( .A(n23873), .B(n23870), .Z(n23880) );
  AND U23779 ( .A(n23892), .B(n23893), .Z(n23870) );
  XOR U23780 ( .A(n23894), .B(n23895), .Z(n23873) );
  AND U23781 ( .A(n23896), .B(n23897), .Z(n23895) );
  XOR U23782 ( .A(n23894), .B(n23898), .Z(n23896) );
  XNOR U23783 ( .A(n23822), .B(n23876), .Z(n23878) );
  XNOR U23784 ( .A(n23899), .B(n23900), .Z(n23822) );
  AND U23785 ( .A(n364), .B(n23828), .Z(n23900) );
  XOR U23786 ( .A(n23899), .B(n23826), .Z(n23828) );
  XOR U23787 ( .A(n23901), .B(n23902), .Z(n23876) );
  AND U23788 ( .A(n23903), .B(n23904), .Z(n23902) );
  XNOR U23789 ( .A(n23901), .B(n23892), .Z(n23904) );
  IV U23790 ( .A(n23834), .Z(n23892) );
  XNOR U23791 ( .A(n23905), .B(n23885), .Z(n23834) );
  XNOR U23792 ( .A(n23906), .B(n23891), .Z(n23885) );
  XOR U23793 ( .A(n23907), .B(n23908), .Z(n23891) );
  AND U23794 ( .A(n23909), .B(n23910), .Z(n23908) );
  XOR U23795 ( .A(n23907), .B(n23911), .Z(n23909) );
  XNOR U23796 ( .A(n23890), .B(n23882), .Z(n23906) );
  XOR U23797 ( .A(n23912), .B(n23913), .Z(n23882) );
  AND U23798 ( .A(n23914), .B(n23915), .Z(n23913) );
  XNOR U23799 ( .A(n23916), .B(n23912), .Z(n23914) );
  XNOR U23800 ( .A(n23917), .B(n23887), .Z(n23890) );
  XOR U23801 ( .A(n23918), .B(n23919), .Z(n23887) );
  AND U23802 ( .A(n23920), .B(n23921), .Z(n23919) );
  XOR U23803 ( .A(n23918), .B(n23922), .Z(n23920) );
  XNOR U23804 ( .A(n23923), .B(n23924), .Z(n23917) );
  AND U23805 ( .A(n23925), .B(n23926), .Z(n23924) );
  XNOR U23806 ( .A(n23923), .B(n23927), .Z(n23925) );
  XNOR U23807 ( .A(n23886), .B(n23893), .Z(n23905) );
  AND U23808 ( .A(n23846), .B(n23928), .Z(n23893) );
  XOR U23809 ( .A(n23898), .B(n23897), .Z(n23886) );
  XNOR U23810 ( .A(n23929), .B(n23894), .Z(n23897) );
  XOR U23811 ( .A(n23930), .B(n23931), .Z(n23894) );
  AND U23812 ( .A(n23932), .B(n23933), .Z(n23931) );
  XOR U23813 ( .A(n23930), .B(n23934), .Z(n23932) );
  XNOR U23814 ( .A(n23935), .B(n23936), .Z(n23929) );
  AND U23815 ( .A(n23937), .B(n23938), .Z(n23936) );
  XOR U23816 ( .A(n23935), .B(n23939), .Z(n23937) );
  XOR U23817 ( .A(n23940), .B(n23941), .Z(n23898) );
  AND U23818 ( .A(n23942), .B(n23943), .Z(n23941) );
  XOR U23819 ( .A(n23940), .B(n23944), .Z(n23942) );
  XNOR U23820 ( .A(n23831), .B(n23901), .Z(n23903) );
  XNOR U23821 ( .A(n23945), .B(n23946), .Z(n23831) );
  AND U23822 ( .A(n364), .B(n23838), .Z(n23946) );
  XOR U23823 ( .A(n23945), .B(n23836), .Z(n23838) );
  XOR U23824 ( .A(n23947), .B(n23948), .Z(n23901) );
  AND U23825 ( .A(n23949), .B(n23950), .Z(n23948) );
  XNOR U23826 ( .A(n23947), .B(n23846), .Z(n23950) );
  XOR U23827 ( .A(n23951), .B(n23915), .Z(n23846) );
  XNOR U23828 ( .A(n23952), .B(n23922), .Z(n23915) );
  XOR U23829 ( .A(n23911), .B(n23910), .Z(n23922) );
  XNOR U23830 ( .A(n23953), .B(n23907), .Z(n23910) );
  XOR U23831 ( .A(n23954), .B(n23955), .Z(n23907) );
  AND U23832 ( .A(n23956), .B(n23957), .Z(n23955) );
  XOR U23833 ( .A(n23954), .B(n23958), .Z(n23956) );
  XNOR U23834 ( .A(n23959), .B(n23960), .Z(n23953) );
  NOR U23835 ( .A(n23961), .B(n23962), .Z(n23960) );
  XNOR U23836 ( .A(n23959), .B(n23963), .Z(n23961) );
  XOR U23837 ( .A(n23964), .B(n23965), .Z(n23911) );
  NOR U23838 ( .A(n23966), .B(n23967), .Z(n23965) );
  XNOR U23839 ( .A(n23964), .B(n23968), .Z(n23966) );
  XNOR U23840 ( .A(n23921), .B(n23912), .Z(n23952) );
  XOR U23841 ( .A(n23969), .B(n23970), .Z(n23912) );
  NOR U23842 ( .A(n23971), .B(n23972), .Z(n23970) );
  XNOR U23843 ( .A(n23969), .B(n23973), .Z(n23971) );
  XOR U23844 ( .A(n23974), .B(n23927), .Z(n23921) );
  XNOR U23845 ( .A(n23975), .B(n23976), .Z(n23927) );
  NOR U23846 ( .A(n23977), .B(n23978), .Z(n23976) );
  XNOR U23847 ( .A(n23975), .B(n23979), .Z(n23977) );
  XNOR U23848 ( .A(n23926), .B(n23918), .Z(n23974) );
  XOR U23849 ( .A(n23980), .B(n23981), .Z(n23918) );
  AND U23850 ( .A(n23982), .B(n23983), .Z(n23981) );
  XOR U23851 ( .A(n23980), .B(n23984), .Z(n23982) );
  XNOR U23852 ( .A(n23985), .B(n23923), .Z(n23926) );
  XOR U23853 ( .A(n23986), .B(n23987), .Z(n23923) );
  AND U23854 ( .A(n23988), .B(n23989), .Z(n23987) );
  XOR U23855 ( .A(n23986), .B(n23990), .Z(n23988) );
  XNOR U23856 ( .A(n23991), .B(n23992), .Z(n23985) );
  NOR U23857 ( .A(n23993), .B(n23994), .Z(n23992) );
  XOR U23858 ( .A(n23991), .B(n23995), .Z(n23993) );
  XOR U23859 ( .A(n23916), .B(n23928), .Z(n23951) );
  NOR U23860 ( .A(n23854), .B(n23996), .Z(n23928) );
  XNOR U23861 ( .A(n23934), .B(n23933), .Z(n23916) );
  XNOR U23862 ( .A(n23997), .B(n23939), .Z(n23933) );
  XOR U23863 ( .A(n23998), .B(n23999), .Z(n23939) );
  NOR U23864 ( .A(n24000), .B(n24001), .Z(n23999) );
  XNOR U23865 ( .A(n23998), .B(n24002), .Z(n24000) );
  XNOR U23866 ( .A(n23938), .B(n23930), .Z(n23997) );
  XOR U23867 ( .A(n24003), .B(n24004), .Z(n23930) );
  AND U23868 ( .A(n24005), .B(n24006), .Z(n24004) );
  XNOR U23869 ( .A(n24003), .B(n24007), .Z(n24005) );
  XNOR U23870 ( .A(n24008), .B(n23935), .Z(n23938) );
  XOR U23871 ( .A(n24009), .B(n24010), .Z(n23935) );
  AND U23872 ( .A(n24011), .B(n24012), .Z(n24010) );
  XOR U23873 ( .A(n24009), .B(n24013), .Z(n24011) );
  XNOR U23874 ( .A(n24014), .B(n24015), .Z(n24008) );
  NOR U23875 ( .A(n24016), .B(n24017), .Z(n24015) );
  XOR U23876 ( .A(n24014), .B(n24018), .Z(n24016) );
  XOR U23877 ( .A(n23944), .B(n23943), .Z(n23934) );
  XNOR U23878 ( .A(n24019), .B(n23940), .Z(n23943) );
  XOR U23879 ( .A(n24020), .B(n24021), .Z(n23940) );
  AND U23880 ( .A(n24022), .B(n24023), .Z(n24021) );
  XOR U23881 ( .A(n24020), .B(n24024), .Z(n24022) );
  XNOR U23882 ( .A(n24025), .B(n24026), .Z(n24019) );
  NOR U23883 ( .A(n24027), .B(n24028), .Z(n24026) );
  XNOR U23884 ( .A(n24025), .B(n24029), .Z(n24027) );
  XOR U23885 ( .A(n24030), .B(n24031), .Z(n23944) );
  NOR U23886 ( .A(n24032), .B(n24033), .Z(n24031) );
  XNOR U23887 ( .A(n24030), .B(n24034), .Z(n24032) );
  XNOR U23888 ( .A(n23843), .B(n23947), .Z(n23949) );
  XNOR U23889 ( .A(n24035), .B(n24036), .Z(n23843) );
  AND U23890 ( .A(n364), .B(n23850), .Z(n24036) );
  XOR U23891 ( .A(n24035), .B(n23848), .Z(n23850) );
  AND U23892 ( .A(n23851), .B(n23854), .Z(n23947) );
  XOR U23893 ( .A(n24037), .B(n23996), .Z(n23854) );
  XNOR U23894 ( .A(p_input[2048]), .B(p_input[864]), .Z(n23996) );
  XOR U23895 ( .A(n23973), .B(n23972), .Z(n24037) );
  XOR U23896 ( .A(n24038), .B(n23984), .Z(n23972) );
  XOR U23897 ( .A(n23958), .B(n23957), .Z(n23984) );
  XNOR U23898 ( .A(n24039), .B(n23963), .Z(n23957) );
  XOR U23899 ( .A(p_input[2072]), .B(p_input[888]), .Z(n23963) );
  XOR U23900 ( .A(n23954), .B(n23962), .Z(n24039) );
  XOR U23901 ( .A(n24040), .B(n23959), .Z(n23962) );
  XOR U23902 ( .A(p_input[2070]), .B(p_input[886]), .Z(n23959) );
  XNOR U23903 ( .A(p_input[2071]), .B(p_input[887]), .Z(n24040) );
  XNOR U23904 ( .A(n16727), .B(p_input[882]), .Z(n23954) );
  XNOR U23905 ( .A(n23968), .B(n23967), .Z(n23958) );
  XOR U23906 ( .A(n24041), .B(n23964), .Z(n23967) );
  XOR U23907 ( .A(p_input[2067]), .B(p_input[883]), .Z(n23964) );
  XNOR U23908 ( .A(p_input[2068]), .B(p_input[884]), .Z(n24041) );
  XOR U23909 ( .A(p_input[2069]), .B(p_input[885]), .Z(n23968) );
  XNOR U23910 ( .A(n23983), .B(n23969), .Z(n24038) );
  XNOR U23911 ( .A(n16729), .B(p_input[865]), .Z(n23969) );
  XNOR U23912 ( .A(n24042), .B(n23990), .Z(n23983) );
  XNOR U23913 ( .A(n23979), .B(n23978), .Z(n23990) );
  XOR U23914 ( .A(n24043), .B(n23975), .Z(n23978) );
  XNOR U23915 ( .A(n16444), .B(p_input[890]), .Z(n23975) );
  XNOR U23916 ( .A(p_input[2075]), .B(p_input[891]), .Z(n24043) );
  XOR U23917 ( .A(p_input[2076]), .B(p_input[892]), .Z(n23979) );
  XNOR U23918 ( .A(n23989), .B(n23980), .Z(n24042) );
  XNOR U23919 ( .A(n16732), .B(p_input[881]), .Z(n23980) );
  XOR U23920 ( .A(n24044), .B(n23995), .Z(n23989) );
  XNOR U23921 ( .A(p_input[2079]), .B(p_input[895]), .Z(n23995) );
  XOR U23922 ( .A(n23986), .B(n23994), .Z(n24044) );
  XOR U23923 ( .A(n24045), .B(n23991), .Z(n23994) );
  XOR U23924 ( .A(p_input[2077]), .B(p_input[893]), .Z(n23991) );
  XNOR U23925 ( .A(p_input[2078]), .B(p_input[894]), .Z(n24045) );
  XNOR U23926 ( .A(n16448), .B(p_input[889]), .Z(n23986) );
  XNOR U23927 ( .A(n24007), .B(n24006), .Z(n23973) );
  XNOR U23928 ( .A(n24046), .B(n24013), .Z(n24006) );
  XNOR U23929 ( .A(n24002), .B(n24001), .Z(n24013) );
  XOR U23930 ( .A(n24047), .B(n23998), .Z(n24001) );
  XNOR U23931 ( .A(n16737), .B(p_input[875]), .Z(n23998) );
  XNOR U23932 ( .A(p_input[2060]), .B(p_input[876]), .Z(n24047) );
  XOR U23933 ( .A(p_input[2061]), .B(p_input[877]), .Z(n24002) );
  XNOR U23934 ( .A(n24012), .B(n24003), .Z(n24046) );
  XNOR U23935 ( .A(n16452), .B(p_input[866]), .Z(n24003) );
  XOR U23936 ( .A(n24048), .B(n24018), .Z(n24012) );
  XNOR U23937 ( .A(p_input[2064]), .B(p_input[880]), .Z(n24018) );
  XOR U23938 ( .A(n24009), .B(n24017), .Z(n24048) );
  XOR U23939 ( .A(n24049), .B(n24014), .Z(n24017) );
  XOR U23940 ( .A(p_input[2062]), .B(p_input[878]), .Z(n24014) );
  XNOR U23941 ( .A(p_input[2063]), .B(p_input[879]), .Z(n24049) );
  XNOR U23942 ( .A(n16740), .B(p_input[874]), .Z(n24009) );
  XNOR U23943 ( .A(n24024), .B(n24023), .Z(n24007) );
  XNOR U23944 ( .A(n24050), .B(n24029), .Z(n24023) );
  XOR U23945 ( .A(p_input[2057]), .B(p_input[873]), .Z(n24029) );
  XOR U23946 ( .A(n24020), .B(n24028), .Z(n24050) );
  XOR U23947 ( .A(n24051), .B(n24025), .Z(n24028) );
  XOR U23948 ( .A(p_input[2055]), .B(p_input[871]), .Z(n24025) );
  XNOR U23949 ( .A(p_input[2056]), .B(p_input[872]), .Z(n24051) );
  XNOR U23950 ( .A(n16459), .B(p_input[867]), .Z(n24020) );
  XNOR U23951 ( .A(n24034), .B(n24033), .Z(n24024) );
  XOR U23952 ( .A(n24052), .B(n24030), .Z(n24033) );
  XOR U23953 ( .A(p_input[2052]), .B(p_input[868]), .Z(n24030) );
  XNOR U23954 ( .A(p_input[2053]), .B(p_input[869]), .Z(n24052) );
  XOR U23955 ( .A(p_input[2054]), .B(p_input[870]), .Z(n24034) );
  XNOR U23956 ( .A(n24053), .B(n24054), .Z(n23851) );
  AND U23957 ( .A(n364), .B(n24055), .Z(n24054) );
  XNOR U23958 ( .A(n24056), .B(n24057), .Z(n364) );
  AND U23959 ( .A(n24058), .B(n24059), .Z(n24057) );
  XOR U23960 ( .A(n24056), .B(n23861), .Z(n24059) );
  XNOR U23961 ( .A(n24056), .B(n23803), .Z(n24058) );
  XOR U23962 ( .A(n24060), .B(n24061), .Z(n24056) );
  AND U23963 ( .A(n24062), .B(n24063), .Z(n24061) );
  XNOR U23964 ( .A(n23874), .B(n24060), .Z(n24063) );
  XOR U23965 ( .A(n24060), .B(n23815), .Z(n24062) );
  XOR U23966 ( .A(n24064), .B(n24065), .Z(n24060) );
  AND U23967 ( .A(n24066), .B(n24067), .Z(n24065) );
  XNOR U23968 ( .A(n23899), .B(n24064), .Z(n24067) );
  XOR U23969 ( .A(n24064), .B(n23826), .Z(n24066) );
  XOR U23970 ( .A(n24068), .B(n24069), .Z(n24064) );
  AND U23971 ( .A(n24070), .B(n24071), .Z(n24069) );
  XOR U23972 ( .A(n24068), .B(n23836), .Z(n24070) );
  XOR U23973 ( .A(n24072), .B(n24073), .Z(n23792) );
  AND U23974 ( .A(n368), .B(n24055), .Z(n24073) );
  XNOR U23975 ( .A(n24053), .B(n24072), .Z(n24055) );
  XNOR U23976 ( .A(n24074), .B(n24075), .Z(n368) );
  AND U23977 ( .A(n24076), .B(n24077), .Z(n24075) );
  XNOR U23978 ( .A(n24078), .B(n24074), .Z(n24077) );
  IV U23979 ( .A(n23861), .Z(n24078) );
  XNOR U23980 ( .A(n24079), .B(n24080), .Z(n23861) );
  AND U23981 ( .A(n371), .B(n24081), .Z(n24080) );
  XNOR U23982 ( .A(n24079), .B(n24082), .Z(n24081) );
  XNOR U23983 ( .A(n23803), .B(n24074), .Z(n24076) );
  XOR U23984 ( .A(n24083), .B(n24084), .Z(n23803) );
  AND U23985 ( .A(n379), .B(n24085), .Z(n24084) );
  XOR U23986 ( .A(n24086), .B(n24087), .Z(n24074) );
  AND U23987 ( .A(n24088), .B(n24089), .Z(n24087) );
  XNOR U23988 ( .A(n24086), .B(n23874), .Z(n24089) );
  XNOR U23989 ( .A(n24090), .B(n24091), .Z(n23874) );
  AND U23990 ( .A(n371), .B(n24092), .Z(n24091) );
  XOR U23991 ( .A(n24093), .B(n24090), .Z(n24092) );
  XNOR U23992 ( .A(n24094), .B(n24086), .Z(n24088) );
  IV U23993 ( .A(n23815), .Z(n24094) );
  XOR U23994 ( .A(n24095), .B(n24096), .Z(n23815) );
  AND U23995 ( .A(n379), .B(n24097), .Z(n24096) );
  XOR U23996 ( .A(n24098), .B(n24099), .Z(n24086) );
  AND U23997 ( .A(n24100), .B(n24101), .Z(n24099) );
  XNOR U23998 ( .A(n24098), .B(n23899), .Z(n24101) );
  XNOR U23999 ( .A(n24102), .B(n24103), .Z(n23899) );
  AND U24000 ( .A(n371), .B(n24104), .Z(n24103) );
  XNOR U24001 ( .A(n24105), .B(n24102), .Z(n24104) );
  XOR U24002 ( .A(n23826), .B(n24098), .Z(n24100) );
  XOR U24003 ( .A(n24106), .B(n24107), .Z(n23826) );
  AND U24004 ( .A(n379), .B(n24108), .Z(n24107) );
  XOR U24005 ( .A(n24068), .B(n24109), .Z(n24098) );
  AND U24006 ( .A(n24110), .B(n24071), .Z(n24109) );
  XNOR U24007 ( .A(n23945), .B(n24068), .Z(n24071) );
  XNOR U24008 ( .A(n24111), .B(n24112), .Z(n23945) );
  AND U24009 ( .A(n371), .B(n24113), .Z(n24112) );
  XOR U24010 ( .A(n24114), .B(n24111), .Z(n24113) );
  XNOR U24011 ( .A(n24115), .B(n24068), .Z(n24110) );
  IV U24012 ( .A(n23836), .Z(n24115) );
  XOR U24013 ( .A(n24116), .B(n24117), .Z(n23836) );
  AND U24014 ( .A(n379), .B(n24118), .Z(n24117) );
  XOR U24015 ( .A(n24119), .B(n24120), .Z(n24068) );
  AND U24016 ( .A(n24121), .B(n24122), .Z(n24120) );
  XNOR U24017 ( .A(n24119), .B(n24035), .Z(n24122) );
  XNOR U24018 ( .A(n24123), .B(n24124), .Z(n24035) );
  AND U24019 ( .A(n371), .B(n24125), .Z(n24124) );
  XNOR U24020 ( .A(n24126), .B(n24123), .Z(n24125) );
  XNOR U24021 ( .A(n24127), .B(n24119), .Z(n24121) );
  IV U24022 ( .A(n23848), .Z(n24127) );
  XOR U24023 ( .A(n24128), .B(n24129), .Z(n23848) );
  AND U24024 ( .A(n379), .B(n24130), .Z(n24129) );
  AND U24025 ( .A(n24072), .B(n24053), .Z(n24119) );
  XNOR U24026 ( .A(n24131), .B(n24132), .Z(n24053) );
  AND U24027 ( .A(n371), .B(n24133), .Z(n24132) );
  XNOR U24028 ( .A(n24134), .B(n24131), .Z(n24133) );
  XNOR U24029 ( .A(n24135), .B(n24136), .Z(n371) );
  AND U24030 ( .A(n24137), .B(n24138), .Z(n24136) );
  XOR U24031 ( .A(n24082), .B(n24135), .Z(n24138) );
  AND U24032 ( .A(n24139), .B(n24140), .Z(n24082) );
  XOR U24033 ( .A(n24135), .B(n24079), .Z(n24137) );
  XNOR U24034 ( .A(n24141), .B(n24142), .Z(n24079) );
  AND U24035 ( .A(n375), .B(n24085), .Z(n24142) );
  XOR U24036 ( .A(n24083), .B(n24141), .Z(n24085) );
  XOR U24037 ( .A(n24143), .B(n24144), .Z(n24135) );
  AND U24038 ( .A(n24145), .B(n24146), .Z(n24144) );
  XNOR U24039 ( .A(n24143), .B(n24139), .Z(n24146) );
  IV U24040 ( .A(n24093), .Z(n24139) );
  XOR U24041 ( .A(n24147), .B(n24148), .Z(n24093) );
  XOR U24042 ( .A(n24149), .B(n24140), .Z(n24148) );
  AND U24043 ( .A(n24105), .B(n24150), .Z(n24140) );
  AND U24044 ( .A(n24151), .B(n24152), .Z(n24149) );
  XOR U24045 ( .A(n24153), .B(n24147), .Z(n24151) );
  XNOR U24046 ( .A(n24090), .B(n24143), .Z(n24145) );
  XNOR U24047 ( .A(n24154), .B(n24155), .Z(n24090) );
  AND U24048 ( .A(n375), .B(n24097), .Z(n24155) );
  XOR U24049 ( .A(n24154), .B(n24095), .Z(n24097) );
  XOR U24050 ( .A(n24156), .B(n24157), .Z(n24143) );
  AND U24051 ( .A(n24158), .B(n24159), .Z(n24157) );
  XNOR U24052 ( .A(n24156), .B(n24105), .Z(n24159) );
  XOR U24053 ( .A(n24160), .B(n24152), .Z(n24105) );
  XNOR U24054 ( .A(n24161), .B(n24147), .Z(n24152) );
  XOR U24055 ( .A(n24162), .B(n24163), .Z(n24147) );
  AND U24056 ( .A(n24164), .B(n24165), .Z(n24163) );
  XOR U24057 ( .A(n24166), .B(n24162), .Z(n24164) );
  XNOR U24058 ( .A(n24167), .B(n24168), .Z(n24161) );
  AND U24059 ( .A(n24169), .B(n24170), .Z(n24168) );
  XOR U24060 ( .A(n24167), .B(n24171), .Z(n24169) );
  XNOR U24061 ( .A(n24153), .B(n24150), .Z(n24160) );
  AND U24062 ( .A(n24172), .B(n24173), .Z(n24150) );
  XOR U24063 ( .A(n24174), .B(n24175), .Z(n24153) );
  AND U24064 ( .A(n24176), .B(n24177), .Z(n24175) );
  XOR U24065 ( .A(n24174), .B(n24178), .Z(n24176) );
  XNOR U24066 ( .A(n24102), .B(n24156), .Z(n24158) );
  XNOR U24067 ( .A(n24179), .B(n24180), .Z(n24102) );
  AND U24068 ( .A(n375), .B(n24108), .Z(n24180) );
  XOR U24069 ( .A(n24179), .B(n24106), .Z(n24108) );
  XOR U24070 ( .A(n24181), .B(n24182), .Z(n24156) );
  AND U24071 ( .A(n24183), .B(n24184), .Z(n24182) );
  XNOR U24072 ( .A(n24181), .B(n24172), .Z(n24184) );
  IV U24073 ( .A(n24114), .Z(n24172) );
  XNOR U24074 ( .A(n24185), .B(n24165), .Z(n24114) );
  XNOR U24075 ( .A(n24186), .B(n24171), .Z(n24165) );
  XOR U24076 ( .A(n24187), .B(n24188), .Z(n24171) );
  AND U24077 ( .A(n24189), .B(n24190), .Z(n24188) );
  XOR U24078 ( .A(n24187), .B(n24191), .Z(n24189) );
  XNOR U24079 ( .A(n24170), .B(n24162), .Z(n24186) );
  XOR U24080 ( .A(n24192), .B(n24193), .Z(n24162) );
  AND U24081 ( .A(n24194), .B(n24195), .Z(n24193) );
  XNOR U24082 ( .A(n24196), .B(n24192), .Z(n24194) );
  XNOR U24083 ( .A(n24197), .B(n24167), .Z(n24170) );
  XOR U24084 ( .A(n24198), .B(n24199), .Z(n24167) );
  AND U24085 ( .A(n24200), .B(n24201), .Z(n24199) );
  XOR U24086 ( .A(n24198), .B(n24202), .Z(n24200) );
  XNOR U24087 ( .A(n24203), .B(n24204), .Z(n24197) );
  AND U24088 ( .A(n24205), .B(n24206), .Z(n24204) );
  XNOR U24089 ( .A(n24203), .B(n24207), .Z(n24205) );
  XNOR U24090 ( .A(n24166), .B(n24173), .Z(n24185) );
  AND U24091 ( .A(n24126), .B(n24208), .Z(n24173) );
  XOR U24092 ( .A(n24178), .B(n24177), .Z(n24166) );
  XNOR U24093 ( .A(n24209), .B(n24174), .Z(n24177) );
  XOR U24094 ( .A(n24210), .B(n24211), .Z(n24174) );
  AND U24095 ( .A(n24212), .B(n24213), .Z(n24211) );
  XOR U24096 ( .A(n24210), .B(n24214), .Z(n24212) );
  XNOR U24097 ( .A(n24215), .B(n24216), .Z(n24209) );
  AND U24098 ( .A(n24217), .B(n24218), .Z(n24216) );
  XOR U24099 ( .A(n24215), .B(n24219), .Z(n24217) );
  XOR U24100 ( .A(n24220), .B(n24221), .Z(n24178) );
  AND U24101 ( .A(n24222), .B(n24223), .Z(n24221) );
  XOR U24102 ( .A(n24220), .B(n24224), .Z(n24222) );
  XNOR U24103 ( .A(n24111), .B(n24181), .Z(n24183) );
  XNOR U24104 ( .A(n24225), .B(n24226), .Z(n24111) );
  AND U24105 ( .A(n375), .B(n24118), .Z(n24226) );
  XOR U24106 ( .A(n24225), .B(n24116), .Z(n24118) );
  XOR U24107 ( .A(n24227), .B(n24228), .Z(n24181) );
  AND U24108 ( .A(n24229), .B(n24230), .Z(n24228) );
  XNOR U24109 ( .A(n24227), .B(n24126), .Z(n24230) );
  XOR U24110 ( .A(n24231), .B(n24195), .Z(n24126) );
  XNOR U24111 ( .A(n24232), .B(n24202), .Z(n24195) );
  XOR U24112 ( .A(n24191), .B(n24190), .Z(n24202) );
  XNOR U24113 ( .A(n24233), .B(n24187), .Z(n24190) );
  XOR U24114 ( .A(n24234), .B(n24235), .Z(n24187) );
  AND U24115 ( .A(n24236), .B(n24237), .Z(n24235) );
  XOR U24116 ( .A(n24234), .B(n24238), .Z(n24236) );
  XNOR U24117 ( .A(n24239), .B(n24240), .Z(n24233) );
  NOR U24118 ( .A(n24241), .B(n24242), .Z(n24240) );
  XNOR U24119 ( .A(n24239), .B(n24243), .Z(n24241) );
  XOR U24120 ( .A(n24244), .B(n24245), .Z(n24191) );
  NOR U24121 ( .A(n24246), .B(n24247), .Z(n24245) );
  XNOR U24122 ( .A(n24244), .B(n24248), .Z(n24246) );
  XNOR U24123 ( .A(n24201), .B(n24192), .Z(n24232) );
  XOR U24124 ( .A(n24249), .B(n24250), .Z(n24192) );
  NOR U24125 ( .A(n24251), .B(n24252), .Z(n24250) );
  XNOR U24126 ( .A(n24249), .B(n24253), .Z(n24251) );
  XOR U24127 ( .A(n24254), .B(n24207), .Z(n24201) );
  XNOR U24128 ( .A(n24255), .B(n24256), .Z(n24207) );
  NOR U24129 ( .A(n24257), .B(n24258), .Z(n24256) );
  XNOR U24130 ( .A(n24255), .B(n24259), .Z(n24257) );
  XNOR U24131 ( .A(n24206), .B(n24198), .Z(n24254) );
  XOR U24132 ( .A(n24260), .B(n24261), .Z(n24198) );
  AND U24133 ( .A(n24262), .B(n24263), .Z(n24261) );
  XOR U24134 ( .A(n24260), .B(n24264), .Z(n24262) );
  XNOR U24135 ( .A(n24265), .B(n24203), .Z(n24206) );
  XOR U24136 ( .A(n24266), .B(n24267), .Z(n24203) );
  AND U24137 ( .A(n24268), .B(n24269), .Z(n24267) );
  XOR U24138 ( .A(n24266), .B(n24270), .Z(n24268) );
  XNOR U24139 ( .A(n24271), .B(n24272), .Z(n24265) );
  NOR U24140 ( .A(n24273), .B(n24274), .Z(n24272) );
  XOR U24141 ( .A(n24271), .B(n24275), .Z(n24273) );
  XOR U24142 ( .A(n24196), .B(n24208), .Z(n24231) );
  NOR U24143 ( .A(n24134), .B(n24276), .Z(n24208) );
  XNOR U24144 ( .A(n24214), .B(n24213), .Z(n24196) );
  XNOR U24145 ( .A(n24277), .B(n24219), .Z(n24213) );
  XOR U24146 ( .A(n24278), .B(n24279), .Z(n24219) );
  NOR U24147 ( .A(n24280), .B(n24281), .Z(n24279) );
  XNOR U24148 ( .A(n24278), .B(n24282), .Z(n24280) );
  XNOR U24149 ( .A(n24218), .B(n24210), .Z(n24277) );
  XOR U24150 ( .A(n24283), .B(n24284), .Z(n24210) );
  AND U24151 ( .A(n24285), .B(n24286), .Z(n24284) );
  XNOR U24152 ( .A(n24283), .B(n24287), .Z(n24285) );
  XNOR U24153 ( .A(n24288), .B(n24215), .Z(n24218) );
  XOR U24154 ( .A(n24289), .B(n24290), .Z(n24215) );
  AND U24155 ( .A(n24291), .B(n24292), .Z(n24290) );
  XOR U24156 ( .A(n24289), .B(n24293), .Z(n24291) );
  XNOR U24157 ( .A(n24294), .B(n24295), .Z(n24288) );
  NOR U24158 ( .A(n24296), .B(n24297), .Z(n24295) );
  XOR U24159 ( .A(n24294), .B(n24298), .Z(n24296) );
  XOR U24160 ( .A(n24224), .B(n24223), .Z(n24214) );
  XNOR U24161 ( .A(n24299), .B(n24220), .Z(n24223) );
  XOR U24162 ( .A(n24300), .B(n24301), .Z(n24220) );
  AND U24163 ( .A(n24302), .B(n24303), .Z(n24301) );
  XOR U24164 ( .A(n24300), .B(n24304), .Z(n24302) );
  XNOR U24165 ( .A(n24305), .B(n24306), .Z(n24299) );
  NOR U24166 ( .A(n24307), .B(n24308), .Z(n24306) );
  XNOR U24167 ( .A(n24305), .B(n24309), .Z(n24307) );
  XOR U24168 ( .A(n24310), .B(n24311), .Z(n24224) );
  NOR U24169 ( .A(n24312), .B(n24313), .Z(n24311) );
  XNOR U24170 ( .A(n24310), .B(n24314), .Z(n24312) );
  XNOR U24171 ( .A(n24123), .B(n24227), .Z(n24229) );
  XNOR U24172 ( .A(n24315), .B(n24316), .Z(n24123) );
  AND U24173 ( .A(n375), .B(n24130), .Z(n24316) );
  XOR U24174 ( .A(n24315), .B(n24128), .Z(n24130) );
  AND U24175 ( .A(n24131), .B(n24134), .Z(n24227) );
  XOR U24176 ( .A(n24317), .B(n24276), .Z(n24134) );
  XNOR U24177 ( .A(p_input[2048]), .B(p_input[896]), .Z(n24276) );
  XOR U24178 ( .A(n24253), .B(n24252), .Z(n24317) );
  XOR U24179 ( .A(n24318), .B(n24264), .Z(n24252) );
  XOR U24180 ( .A(n24238), .B(n24237), .Z(n24264) );
  XNOR U24181 ( .A(n24319), .B(n24243), .Z(n24237) );
  XOR U24182 ( .A(p_input[2072]), .B(p_input[920]), .Z(n24243) );
  XOR U24183 ( .A(n24234), .B(n24242), .Z(n24319) );
  XOR U24184 ( .A(n24320), .B(n24239), .Z(n24242) );
  XOR U24185 ( .A(p_input[2070]), .B(p_input[918]), .Z(n24239) );
  XNOR U24186 ( .A(p_input[2071]), .B(p_input[919]), .Z(n24320) );
  XNOR U24187 ( .A(n16727), .B(p_input[914]), .Z(n24234) );
  XNOR U24188 ( .A(n24248), .B(n24247), .Z(n24238) );
  XOR U24189 ( .A(n24321), .B(n24244), .Z(n24247) );
  XOR U24190 ( .A(p_input[2067]), .B(p_input[915]), .Z(n24244) );
  XNOR U24191 ( .A(p_input[2068]), .B(p_input[916]), .Z(n24321) );
  XOR U24192 ( .A(p_input[2069]), .B(p_input[917]), .Z(n24248) );
  XNOR U24193 ( .A(n24263), .B(n24249), .Z(n24318) );
  XNOR U24194 ( .A(n16729), .B(p_input[897]), .Z(n24249) );
  XNOR U24195 ( .A(n24322), .B(n24270), .Z(n24263) );
  XNOR U24196 ( .A(n24259), .B(n24258), .Z(n24270) );
  XOR U24197 ( .A(n24323), .B(n24255), .Z(n24258) );
  XNOR U24198 ( .A(n16444), .B(p_input[922]), .Z(n24255) );
  XNOR U24199 ( .A(p_input[2075]), .B(p_input[923]), .Z(n24323) );
  XOR U24200 ( .A(p_input[2076]), .B(p_input[924]), .Z(n24259) );
  XNOR U24201 ( .A(n24269), .B(n24260), .Z(n24322) );
  XNOR U24202 ( .A(n16732), .B(p_input[913]), .Z(n24260) );
  XOR U24203 ( .A(n24324), .B(n24275), .Z(n24269) );
  XNOR U24204 ( .A(p_input[2079]), .B(p_input[927]), .Z(n24275) );
  XOR U24205 ( .A(n24266), .B(n24274), .Z(n24324) );
  XOR U24206 ( .A(n24325), .B(n24271), .Z(n24274) );
  XOR U24207 ( .A(p_input[2077]), .B(p_input[925]), .Z(n24271) );
  XNOR U24208 ( .A(p_input[2078]), .B(p_input[926]), .Z(n24325) );
  XNOR U24209 ( .A(n16448), .B(p_input[921]), .Z(n24266) );
  XNOR U24210 ( .A(n24287), .B(n24286), .Z(n24253) );
  XNOR U24211 ( .A(n24326), .B(n24293), .Z(n24286) );
  XNOR U24212 ( .A(n24282), .B(n24281), .Z(n24293) );
  XOR U24213 ( .A(n24327), .B(n24278), .Z(n24281) );
  XNOR U24214 ( .A(n16737), .B(p_input[907]), .Z(n24278) );
  XNOR U24215 ( .A(p_input[2060]), .B(p_input[908]), .Z(n24327) );
  XOR U24216 ( .A(p_input[2061]), .B(p_input[909]), .Z(n24282) );
  XNOR U24217 ( .A(n24292), .B(n24283), .Z(n24326) );
  XNOR U24218 ( .A(n16452), .B(p_input[898]), .Z(n24283) );
  XOR U24219 ( .A(n24328), .B(n24298), .Z(n24292) );
  XNOR U24220 ( .A(p_input[2064]), .B(p_input[912]), .Z(n24298) );
  XOR U24221 ( .A(n24289), .B(n24297), .Z(n24328) );
  XOR U24222 ( .A(n24329), .B(n24294), .Z(n24297) );
  XOR U24223 ( .A(p_input[2062]), .B(p_input[910]), .Z(n24294) );
  XNOR U24224 ( .A(p_input[2063]), .B(p_input[911]), .Z(n24329) );
  XNOR U24225 ( .A(n16740), .B(p_input[906]), .Z(n24289) );
  XNOR U24226 ( .A(n24304), .B(n24303), .Z(n24287) );
  XNOR U24227 ( .A(n24330), .B(n24309), .Z(n24303) );
  XOR U24228 ( .A(p_input[2057]), .B(p_input[905]), .Z(n24309) );
  XOR U24229 ( .A(n24300), .B(n24308), .Z(n24330) );
  XOR U24230 ( .A(n24331), .B(n24305), .Z(n24308) );
  XOR U24231 ( .A(p_input[2055]), .B(p_input[903]), .Z(n24305) );
  XNOR U24232 ( .A(p_input[2056]), .B(p_input[904]), .Z(n24331) );
  XNOR U24233 ( .A(n16459), .B(p_input[899]), .Z(n24300) );
  XNOR U24234 ( .A(n24314), .B(n24313), .Z(n24304) );
  XOR U24235 ( .A(n24332), .B(n24310), .Z(n24313) );
  XOR U24236 ( .A(p_input[2052]), .B(p_input[900]), .Z(n24310) );
  XNOR U24237 ( .A(p_input[2053]), .B(p_input[901]), .Z(n24332) );
  XOR U24238 ( .A(p_input[2054]), .B(p_input[902]), .Z(n24314) );
  XNOR U24239 ( .A(n24333), .B(n24334), .Z(n24131) );
  AND U24240 ( .A(n375), .B(n24335), .Z(n24334) );
  XNOR U24241 ( .A(n24336), .B(n24337), .Z(n375) );
  AND U24242 ( .A(n24338), .B(n24339), .Z(n24337) );
  XOR U24243 ( .A(n24336), .B(n24141), .Z(n24339) );
  XNOR U24244 ( .A(n24336), .B(n24083), .Z(n24338) );
  XOR U24245 ( .A(n24340), .B(n24341), .Z(n24336) );
  AND U24246 ( .A(n24342), .B(n24343), .Z(n24341) );
  XNOR U24247 ( .A(n24154), .B(n24340), .Z(n24343) );
  XOR U24248 ( .A(n24340), .B(n24095), .Z(n24342) );
  XOR U24249 ( .A(n24344), .B(n24345), .Z(n24340) );
  AND U24250 ( .A(n24346), .B(n24347), .Z(n24345) );
  XNOR U24251 ( .A(n24179), .B(n24344), .Z(n24347) );
  XOR U24252 ( .A(n24344), .B(n24106), .Z(n24346) );
  XOR U24253 ( .A(n24348), .B(n24349), .Z(n24344) );
  AND U24254 ( .A(n24350), .B(n24351), .Z(n24349) );
  XOR U24255 ( .A(n24348), .B(n24116), .Z(n24350) );
  XOR U24256 ( .A(n24352), .B(n24353), .Z(n24072) );
  AND U24257 ( .A(n379), .B(n24335), .Z(n24353) );
  XNOR U24258 ( .A(n24333), .B(n24352), .Z(n24335) );
  XNOR U24259 ( .A(n24354), .B(n24355), .Z(n379) );
  AND U24260 ( .A(n24356), .B(n24357), .Z(n24355) );
  XNOR U24261 ( .A(n24358), .B(n24354), .Z(n24357) );
  IV U24262 ( .A(n24141), .Z(n24358) );
  XNOR U24263 ( .A(n24359), .B(n24360), .Z(n24141) );
  AND U24264 ( .A(n382), .B(n24361), .Z(n24360) );
  XNOR U24265 ( .A(n24359), .B(n24362), .Z(n24361) );
  XNOR U24266 ( .A(n24083), .B(n24354), .Z(n24356) );
  XOR U24267 ( .A(n24363), .B(n24364), .Z(n24083) );
  AND U24268 ( .A(n390), .B(n24365), .Z(n24364) );
  XOR U24269 ( .A(n24366), .B(n24367), .Z(n24354) );
  AND U24270 ( .A(n24368), .B(n24369), .Z(n24367) );
  XNOR U24271 ( .A(n24366), .B(n24154), .Z(n24369) );
  XNOR U24272 ( .A(n24370), .B(n24371), .Z(n24154) );
  AND U24273 ( .A(n382), .B(n24372), .Z(n24371) );
  XOR U24274 ( .A(n24373), .B(n24370), .Z(n24372) );
  XNOR U24275 ( .A(n24374), .B(n24366), .Z(n24368) );
  IV U24276 ( .A(n24095), .Z(n24374) );
  XOR U24277 ( .A(n24375), .B(n24376), .Z(n24095) );
  AND U24278 ( .A(n390), .B(n24377), .Z(n24376) );
  XOR U24279 ( .A(n24378), .B(n24379), .Z(n24366) );
  AND U24280 ( .A(n24380), .B(n24381), .Z(n24379) );
  XNOR U24281 ( .A(n24378), .B(n24179), .Z(n24381) );
  XNOR U24282 ( .A(n24382), .B(n24383), .Z(n24179) );
  AND U24283 ( .A(n382), .B(n24384), .Z(n24383) );
  XNOR U24284 ( .A(n24385), .B(n24382), .Z(n24384) );
  XOR U24285 ( .A(n24106), .B(n24378), .Z(n24380) );
  XOR U24286 ( .A(n24386), .B(n24387), .Z(n24106) );
  AND U24287 ( .A(n390), .B(n24388), .Z(n24387) );
  XOR U24288 ( .A(n24348), .B(n24389), .Z(n24378) );
  AND U24289 ( .A(n24390), .B(n24351), .Z(n24389) );
  XNOR U24290 ( .A(n24225), .B(n24348), .Z(n24351) );
  XNOR U24291 ( .A(n24391), .B(n24392), .Z(n24225) );
  AND U24292 ( .A(n382), .B(n24393), .Z(n24392) );
  XOR U24293 ( .A(n24394), .B(n24391), .Z(n24393) );
  XNOR U24294 ( .A(n24395), .B(n24348), .Z(n24390) );
  IV U24295 ( .A(n24116), .Z(n24395) );
  XOR U24296 ( .A(n24396), .B(n24397), .Z(n24116) );
  AND U24297 ( .A(n390), .B(n24398), .Z(n24397) );
  XOR U24298 ( .A(n24399), .B(n24400), .Z(n24348) );
  AND U24299 ( .A(n24401), .B(n24402), .Z(n24400) );
  XNOR U24300 ( .A(n24399), .B(n24315), .Z(n24402) );
  XNOR U24301 ( .A(n24403), .B(n24404), .Z(n24315) );
  AND U24302 ( .A(n382), .B(n24405), .Z(n24404) );
  XNOR U24303 ( .A(n24406), .B(n24403), .Z(n24405) );
  XNOR U24304 ( .A(n24407), .B(n24399), .Z(n24401) );
  IV U24305 ( .A(n24128), .Z(n24407) );
  XOR U24306 ( .A(n24408), .B(n24409), .Z(n24128) );
  AND U24307 ( .A(n390), .B(n24410), .Z(n24409) );
  AND U24308 ( .A(n24352), .B(n24333), .Z(n24399) );
  XNOR U24309 ( .A(n24411), .B(n24412), .Z(n24333) );
  AND U24310 ( .A(n382), .B(n24413), .Z(n24412) );
  XNOR U24311 ( .A(n24414), .B(n24411), .Z(n24413) );
  XNOR U24312 ( .A(n24415), .B(n24416), .Z(n382) );
  AND U24313 ( .A(n24417), .B(n24418), .Z(n24416) );
  XOR U24314 ( .A(n24362), .B(n24415), .Z(n24418) );
  AND U24315 ( .A(n24419), .B(n24420), .Z(n24362) );
  XOR U24316 ( .A(n24415), .B(n24359), .Z(n24417) );
  XNOR U24317 ( .A(n24421), .B(n24422), .Z(n24359) );
  AND U24318 ( .A(n386), .B(n24365), .Z(n24422) );
  XOR U24319 ( .A(n24363), .B(n24421), .Z(n24365) );
  XOR U24320 ( .A(n24423), .B(n24424), .Z(n24415) );
  AND U24321 ( .A(n24425), .B(n24426), .Z(n24424) );
  XNOR U24322 ( .A(n24423), .B(n24419), .Z(n24426) );
  IV U24323 ( .A(n24373), .Z(n24419) );
  XOR U24324 ( .A(n24427), .B(n24428), .Z(n24373) );
  XOR U24325 ( .A(n24429), .B(n24420), .Z(n24428) );
  AND U24326 ( .A(n24385), .B(n24430), .Z(n24420) );
  AND U24327 ( .A(n24431), .B(n24432), .Z(n24429) );
  XOR U24328 ( .A(n24433), .B(n24427), .Z(n24431) );
  XNOR U24329 ( .A(n24370), .B(n24423), .Z(n24425) );
  XNOR U24330 ( .A(n24434), .B(n24435), .Z(n24370) );
  AND U24331 ( .A(n386), .B(n24377), .Z(n24435) );
  XOR U24332 ( .A(n24434), .B(n24375), .Z(n24377) );
  XOR U24333 ( .A(n24436), .B(n24437), .Z(n24423) );
  AND U24334 ( .A(n24438), .B(n24439), .Z(n24437) );
  XNOR U24335 ( .A(n24436), .B(n24385), .Z(n24439) );
  XOR U24336 ( .A(n24440), .B(n24432), .Z(n24385) );
  XNOR U24337 ( .A(n24441), .B(n24427), .Z(n24432) );
  XOR U24338 ( .A(n24442), .B(n24443), .Z(n24427) );
  AND U24339 ( .A(n24444), .B(n24445), .Z(n24443) );
  XOR U24340 ( .A(n24446), .B(n24442), .Z(n24444) );
  XNOR U24341 ( .A(n24447), .B(n24448), .Z(n24441) );
  AND U24342 ( .A(n24449), .B(n24450), .Z(n24448) );
  XOR U24343 ( .A(n24447), .B(n24451), .Z(n24449) );
  XNOR U24344 ( .A(n24433), .B(n24430), .Z(n24440) );
  AND U24345 ( .A(n24452), .B(n24453), .Z(n24430) );
  XOR U24346 ( .A(n24454), .B(n24455), .Z(n24433) );
  AND U24347 ( .A(n24456), .B(n24457), .Z(n24455) );
  XOR U24348 ( .A(n24454), .B(n24458), .Z(n24456) );
  XNOR U24349 ( .A(n24382), .B(n24436), .Z(n24438) );
  XNOR U24350 ( .A(n24459), .B(n24460), .Z(n24382) );
  AND U24351 ( .A(n386), .B(n24388), .Z(n24460) );
  XOR U24352 ( .A(n24459), .B(n24386), .Z(n24388) );
  XOR U24353 ( .A(n24461), .B(n24462), .Z(n24436) );
  AND U24354 ( .A(n24463), .B(n24464), .Z(n24462) );
  XNOR U24355 ( .A(n24461), .B(n24452), .Z(n24464) );
  IV U24356 ( .A(n24394), .Z(n24452) );
  XNOR U24357 ( .A(n24465), .B(n24445), .Z(n24394) );
  XNOR U24358 ( .A(n24466), .B(n24451), .Z(n24445) );
  XOR U24359 ( .A(n24467), .B(n24468), .Z(n24451) );
  AND U24360 ( .A(n24469), .B(n24470), .Z(n24468) );
  XOR U24361 ( .A(n24467), .B(n24471), .Z(n24469) );
  XNOR U24362 ( .A(n24450), .B(n24442), .Z(n24466) );
  XOR U24363 ( .A(n24472), .B(n24473), .Z(n24442) );
  AND U24364 ( .A(n24474), .B(n24475), .Z(n24473) );
  XNOR U24365 ( .A(n24476), .B(n24472), .Z(n24474) );
  XNOR U24366 ( .A(n24477), .B(n24447), .Z(n24450) );
  XOR U24367 ( .A(n24478), .B(n24479), .Z(n24447) );
  AND U24368 ( .A(n24480), .B(n24481), .Z(n24479) );
  XOR U24369 ( .A(n24478), .B(n24482), .Z(n24480) );
  XNOR U24370 ( .A(n24483), .B(n24484), .Z(n24477) );
  AND U24371 ( .A(n24485), .B(n24486), .Z(n24484) );
  XNOR U24372 ( .A(n24483), .B(n24487), .Z(n24485) );
  XNOR U24373 ( .A(n24446), .B(n24453), .Z(n24465) );
  AND U24374 ( .A(n24406), .B(n24488), .Z(n24453) );
  XOR U24375 ( .A(n24458), .B(n24457), .Z(n24446) );
  XNOR U24376 ( .A(n24489), .B(n24454), .Z(n24457) );
  XOR U24377 ( .A(n24490), .B(n24491), .Z(n24454) );
  AND U24378 ( .A(n24492), .B(n24493), .Z(n24491) );
  XOR U24379 ( .A(n24490), .B(n24494), .Z(n24492) );
  XNOR U24380 ( .A(n24495), .B(n24496), .Z(n24489) );
  AND U24381 ( .A(n24497), .B(n24498), .Z(n24496) );
  XOR U24382 ( .A(n24495), .B(n24499), .Z(n24497) );
  XOR U24383 ( .A(n24500), .B(n24501), .Z(n24458) );
  AND U24384 ( .A(n24502), .B(n24503), .Z(n24501) );
  XOR U24385 ( .A(n24500), .B(n24504), .Z(n24502) );
  XNOR U24386 ( .A(n24391), .B(n24461), .Z(n24463) );
  XNOR U24387 ( .A(n24505), .B(n24506), .Z(n24391) );
  AND U24388 ( .A(n386), .B(n24398), .Z(n24506) );
  XOR U24389 ( .A(n24505), .B(n24396), .Z(n24398) );
  XOR U24390 ( .A(n24507), .B(n24508), .Z(n24461) );
  AND U24391 ( .A(n24509), .B(n24510), .Z(n24508) );
  XNOR U24392 ( .A(n24507), .B(n24406), .Z(n24510) );
  XOR U24393 ( .A(n24511), .B(n24475), .Z(n24406) );
  XNOR U24394 ( .A(n24512), .B(n24482), .Z(n24475) );
  XOR U24395 ( .A(n24471), .B(n24470), .Z(n24482) );
  XNOR U24396 ( .A(n24513), .B(n24467), .Z(n24470) );
  XOR U24397 ( .A(n24514), .B(n24515), .Z(n24467) );
  AND U24398 ( .A(n24516), .B(n24517), .Z(n24515) );
  XOR U24399 ( .A(n24514), .B(n24518), .Z(n24516) );
  XNOR U24400 ( .A(n24519), .B(n24520), .Z(n24513) );
  NOR U24401 ( .A(n24521), .B(n24522), .Z(n24520) );
  XNOR U24402 ( .A(n24519), .B(n24523), .Z(n24521) );
  XOR U24403 ( .A(n24524), .B(n24525), .Z(n24471) );
  NOR U24404 ( .A(n24526), .B(n24527), .Z(n24525) );
  XNOR U24405 ( .A(n24524), .B(n24528), .Z(n24526) );
  XNOR U24406 ( .A(n24481), .B(n24472), .Z(n24512) );
  XOR U24407 ( .A(n24529), .B(n24530), .Z(n24472) );
  NOR U24408 ( .A(n24531), .B(n24532), .Z(n24530) );
  XNOR U24409 ( .A(n24529), .B(n24533), .Z(n24531) );
  XOR U24410 ( .A(n24534), .B(n24487), .Z(n24481) );
  XNOR U24411 ( .A(n24535), .B(n24536), .Z(n24487) );
  NOR U24412 ( .A(n24537), .B(n24538), .Z(n24536) );
  XNOR U24413 ( .A(n24535), .B(n24539), .Z(n24537) );
  XNOR U24414 ( .A(n24486), .B(n24478), .Z(n24534) );
  XOR U24415 ( .A(n24540), .B(n24541), .Z(n24478) );
  AND U24416 ( .A(n24542), .B(n24543), .Z(n24541) );
  XOR U24417 ( .A(n24540), .B(n24544), .Z(n24542) );
  XNOR U24418 ( .A(n24545), .B(n24483), .Z(n24486) );
  XOR U24419 ( .A(n24546), .B(n24547), .Z(n24483) );
  AND U24420 ( .A(n24548), .B(n24549), .Z(n24547) );
  XOR U24421 ( .A(n24546), .B(n24550), .Z(n24548) );
  XNOR U24422 ( .A(n24551), .B(n24552), .Z(n24545) );
  NOR U24423 ( .A(n24553), .B(n24554), .Z(n24552) );
  XOR U24424 ( .A(n24551), .B(n24555), .Z(n24553) );
  XOR U24425 ( .A(n24476), .B(n24488), .Z(n24511) );
  NOR U24426 ( .A(n24414), .B(n24556), .Z(n24488) );
  XNOR U24427 ( .A(n24494), .B(n24493), .Z(n24476) );
  XNOR U24428 ( .A(n24557), .B(n24499), .Z(n24493) );
  XOR U24429 ( .A(n24558), .B(n24559), .Z(n24499) );
  NOR U24430 ( .A(n24560), .B(n24561), .Z(n24559) );
  XNOR U24431 ( .A(n24558), .B(n24562), .Z(n24560) );
  XNOR U24432 ( .A(n24498), .B(n24490), .Z(n24557) );
  XOR U24433 ( .A(n24563), .B(n24564), .Z(n24490) );
  AND U24434 ( .A(n24565), .B(n24566), .Z(n24564) );
  XNOR U24435 ( .A(n24563), .B(n24567), .Z(n24565) );
  XNOR U24436 ( .A(n24568), .B(n24495), .Z(n24498) );
  XOR U24437 ( .A(n24569), .B(n24570), .Z(n24495) );
  AND U24438 ( .A(n24571), .B(n24572), .Z(n24570) );
  XOR U24439 ( .A(n24569), .B(n24573), .Z(n24571) );
  XNOR U24440 ( .A(n24574), .B(n24575), .Z(n24568) );
  NOR U24441 ( .A(n24576), .B(n24577), .Z(n24575) );
  XOR U24442 ( .A(n24574), .B(n24578), .Z(n24576) );
  XOR U24443 ( .A(n24504), .B(n24503), .Z(n24494) );
  XNOR U24444 ( .A(n24579), .B(n24500), .Z(n24503) );
  XOR U24445 ( .A(n24580), .B(n24581), .Z(n24500) );
  AND U24446 ( .A(n24582), .B(n24583), .Z(n24581) );
  XOR U24447 ( .A(n24580), .B(n24584), .Z(n24582) );
  XNOR U24448 ( .A(n24585), .B(n24586), .Z(n24579) );
  NOR U24449 ( .A(n24587), .B(n24588), .Z(n24586) );
  XNOR U24450 ( .A(n24585), .B(n24589), .Z(n24587) );
  XOR U24451 ( .A(n24590), .B(n24591), .Z(n24504) );
  NOR U24452 ( .A(n24592), .B(n24593), .Z(n24591) );
  XNOR U24453 ( .A(n24590), .B(n24594), .Z(n24592) );
  XNOR U24454 ( .A(n24403), .B(n24507), .Z(n24509) );
  XNOR U24455 ( .A(n24595), .B(n24596), .Z(n24403) );
  AND U24456 ( .A(n386), .B(n24410), .Z(n24596) );
  XOR U24457 ( .A(n24595), .B(n24408), .Z(n24410) );
  AND U24458 ( .A(n24411), .B(n24414), .Z(n24507) );
  XOR U24459 ( .A(n24597), .B(n24556), .Z(n24414) );
  XNOR U24460 ( .A(p_input[2048]), .B(p_input[928]), .Z(n24556) );
  XOR U24461 ( .A(n24533), .B(n24532), .Z(n24597) );
  XOR U24462 ( .A(n24598), .B(n24544), .Z(n24532) );
  XOR U24463 ( .A(n24518), .B(n24517), .Z(n24544) );
  XNOR U24464 ( .A(n24599), .B(n24523), .Z(n24517) );
  XOR U24465 ( .A(p_input[2072]), .B(p_input[952]), .Z(n24523) );
  XOR U24466 ( .A(n24514), .B(n24522), .Z(n24599) );
  XOR U24467 ( .A(n24600), .B(n24519), .Z(n24522) );
  XOR U24468 ( .A(p_input[2070]), .B(p_input[950]), .Z(n24519) );
  XNOR U24469 ( .A(p_input[2071]), .B(p_input[951]), .Z(n24600) );
  XNOR U24470 ( .A(n16727), .B(p_input[946]), .Z(n24514) );
  XNOR U24471 ( .A(n24528), .B(n24527), .Z(n24518) );
  XOR U24472 ( .A(n24601), .B(n24524), .Z(n24527) );
  XOR U24473 ( .A(p_input[2067]), .B(p_input[947]), .Z(n24524) );
  XNOR U24474 ( .A(p_input[2068]), .B(p_input[948]), .Z(n24601) );
  XOR U24475 ( .A(p_input[2069]), .B(p_input[949]), .Z(n24528) );
  XNOR U24476 ( .A(n24543), .B(n24529), .Z(n24598) );
  XNOR U24477 ( .A(n16729), .B(p_input[929]), .Z(n24529) );
  XNOR U24478 ( .A(n24602), .B(n24550), .Z(n24543) );
  XNOR U24479 ( .A(n24539), .B(n24538), .Z(n24550) );
  XOR U24480 ( .A(n24603), .B(n24535), .Z(n24538) );
  XNOR U24481 ( .A(n16444), .B(p_input[954]), .Z(n24535) );
  XNOR U24482 ( .A(p_input[2075]), .B(p_input[955]), .Z(n24603) );
  XOR U24483 ( .A(p_input[2076]), .B(p_input[956]), .Z(n24539) );
  XNOR U24484 ( .A(n24549), .B(n24540), .Z(n24602) );
  XNOR U24485 ( .A(n16732), .B(p_input[945]), .Z(n24540) );
  XOR U24486 ( .A(n24604), .B(n24555), .Z(n24549) );
  XNOR U24487 ( .A(p_input[2079]), .B(p_input[959]), .Z(n24555) );
  XOR U24488 ( .A(n24546), .B(n24554), .Z(n24604) );
  XOR U24489 ( .A(n24605), .B(n24551), .Z(n24554) );
  XOR U24490 ( .A(p_input[2077]), .B(p_input[957]), .Z(n24551) );
  XNOR U24491 ( .A(p_input[2078]), .B(p_input[958]), .Z(n24605) );
  XNOR U24492 ( .A(n16448), .B(p_input[953]), .Z(n24546) );
  XNOR U24493 ( .A(n24567), .B(n24566), .Z(n24533) );
  XNOR U24494 ( .A(n24606), .B(n24573), .Z(n24566) );
  XNOR U24495 ( .A(n24562), .B(n24561), .Z(n24573) );
  XOR U24496 ( .A(n24607), .B(n24558), .Z(n24561) );
  XNOR U24497 ( .A(n16737), .B(p_input[939]), .Z(n24558) );
  XNOR U24498 ( .A(p_input[2060]), .B(p_input[940]), .Z(n24607) );
  XOR U24499 ( .A(p_input[2061]), .B(p_input[941]), .Z(n24562) );
  XNOR U24500 ( .A(n24572), .B(n24563), .Z(n24606) );
  XNOR U24501 ( .A(n16452), .B(p_input[930]), .Z(n24563) );
  XOR U24502 ( .A(n24608), .B(n24578), .Z(n24572) );
  XNOR U24503 ( .A(p_input[2064]), .B(p_input[944]), .Z(n24578) );
  XOR U24504 ( .A(n24569), .B(n24577), .Z(n24608) );
  XOR U24505 ( .A(n24609), .B(n24574), .Z(n24577) );
  XOR U24506 ( .A(p_input[2062]), .B(p_input[942]), .Z(n24574) );
  XNOR U24507 ( .A(p_input[2063]), .B(p_input[943]), .Z(n24609) );
  XNOR U24508 ( .A(n16740), .B(p_input[938]), .Z(n24569) );
  XNOR U24509 ( .A(n24584), .B(n24583), .Z(n24567) );
  XNOR U24510 ( .A(n24610), .B(n24589), .Z(n24583) );
  XOR U24511 ( .A(p_input[2057]), .B(p_input[937]), .Z(n24589) );
  XOR U24512 ( .A(n24580), .B(n24588), .Z(n24610) );
  XOR U24513 ( .A(n24611), .B(n24585), .Z(n24588) );
  XOR U24514 ( .A(p_input[2055]), .B(p_input[935]), .Z(n24585) );
  XNOR U24515 ( .A(p_input[2056]), .B(p_input[936]), .Z(n24611) );
  XNOR U24516 ( .A(n16459), .B(p_input[931]), .Z(n24580) );
  XNOR U24517 ( .A(n24594), .B(n24593), .Z(n24584) );
  XOR U24518 ( .A(n24612), .B(n24590), .Z(n24593) );
  XOR U24519 ( .A(p_input[2052]), .B(p_input[932]), .Z(n24590) );
  XNOR U24520 ( .A(p_input[2053]), .B(p_input[933]), .Z(n24612) );
  XOR U24521 ( .A(p_input[2054]), .B(p_input[934]), .Z(n24594) );
  XNOR U24522 ( .A(n24613), .B(n24614), .Z(n24411) );
  AND U24523 ( .A(n386), .B(n24615), .Z(n24614) );
  XNOR U24524 ( .A(n24616), .B(n24617), .Z(n386) );
  AND U24525 ( .A(n24618), .B(n24619), .Z(n24617) );
  XOR U24526 ( .A(n24616), .B(n24421), .Z(n24619) );
  XNOR U24527 ( .A(n24616), .B(n24363), .Z(n24618) );
  XOR U24528 ( .A(n24620), .B(n24621), .Z(n24616) );
  AND U24529 ( .A(n24622), .B(n24623), .Z(n24621) );
  XNOR U24530 ( .A(n24434), .B(n24620), .Z(n24623) );
  XOR U24531 ( .A(n24620), .B(n24375), .Z(n24622) );
  XOR U24532 ( .A(n24624), .B(n24625), .Z(n24620) );
  AND U24533 ( .A(n24626), .B(n24627), .Z(n24625) );
  XNOR U24534 ( .A(n24459), .B(n24624), .Z(n24627) );
  XOR U24535 ( .A(n24624), .B(n24386), .Z(n24626) );
  XOR U24536 ( .A(n24628), .B(n24629), .Z(n24624) );
  AND U24537 ( .A(n24630), .B(n24631), .Z(n24629) );
  XOR U24538 ( .A(n24628), .B(n24396), .Z(n24630) );
  XOR U24539 ( .A(n24632), .B(n24633), .Z(n24352) );
  AND U24540 ( .A(n390), .B(n24615), .Z(n24633) );
  XNOR U24541 ( .A(n24613), .B(n24632), .Z(n24615) );
  XNOR U24542 ( .A(n24634), .B(n24635), .Z(n390) );
  AND U24543 ( .A(n24636), .B(n24637), .Z(n24635) );
  XNOR U24544 ( .A(n24638), .B(n24634), .Z(n24637) );
  IV U24545 ( .A(n24421), .Z(n24638) );
  XNOR U24546 ( .A(n24639), .B(n24640), .Z(n24421) );
  AND U24547 ( .A(n393), .B(n24641), .Z(n24640) );
  XNOR U24548 ( .A(n24639), .B(n24642), .Z(n24641) );
  XNOR U24549 ( .A(n24363), .B(n24634), .Z(n24636) );
  XOR U24550 ( .A(n24643), .B(n24644), .Z(n24363) );
  AND U24551 ( .A(n401), .B(n24645), .Z(n24644) );
  XOR U24552 ( .A(n24646), .B(n24647), .Z(n24634) );
  AND U24553 ( .A(n24648), .B(n24649), .Z(n24647) );
  XNOR U24554 ( .A(n24646), .B(n24434), .Z(n24649) );
  XNOR U24555 ( .A(n24650), .B(n24651), .Z(n24434) );
  AND U24556 ( .A(n393), .B(n24652), .Z(n24651) );
  XOR U24557 ( .A(n24653), .B(n24650), .Z(n24652) );
  XNOR U24558 ( .A(n24654), .B(n24646), .Z(n24648) );
  IV U24559 ( .A(n24375), .Z(n24654) );
  XOR U24560 ( .A(n24655), .B(n24656), .Z(n24375) );
  AND U24561 ( .A(n401), .B(n24657), .Z(n24656) );
  XOR U24562 ( .A(n24658), .B(n24659), .Z(n24646) );
  AND U24563 ( .A(n24660), .B(n24661), .Z(n24659) );
  XNOR U24564 ( .A(n24658), .B(n24459), .Z(n24661) );
  XNOR U24565 ( .A(n24662), .B(n24663), .Z(n24459) );
  AND U24566 ( .A(n393), .B(n24664), .Z(n24663) );
  XNOR U24567 ( .A(n24665), .B(n24662), .Z(n24664) );
  XOR U24568 ( .A(n24386), .B(n24658), .Z(n24660) );
  XOR U24569 ( .A(n24666), .B(n24667), .Z(n24386) );
  AND U24570 ( .A(n401), .B(n24668), .Z(n24667) );
  XOR U24571 ( .A(n24628), .B(n24669), .Z(n24658) );
  AND U24572 ( .A(n24670), .B(n24631), .Z(n24669) );
  XNOR U24573 ( .A(n24505), .B(n24628), .Z(n24631) );
  XNOR U24574 ( .A(n24671), .B(n24672), .Z(n24505) );
  AND U24575 ( .A(n393), .B(n24673), .Z(n24672) );
  XOR U24576 ( .A(n24674), .B(n24671), .Z(n24673) );
  XNOR U24577 ( .A(n24675), .B(n24628), .Z(n24670) );
  IV U24578 ( .A(n24396), .Z(n24675) );
  XOR U24579 ( .A(n24676), .B(n24677), .Z(n24396) );
  AND U24580 ( .A(n401), .B(n24678), .Z(n24677) );
  XOR U24581 ( .A(n24679), .B(n24680), .Z(n24628) );
  AND U24582 ( .A(n24681), .B(n24682), .Z(n24680) );
  XNOR U24583 ( .A(n24679), .B(n24595), .Z(n24682) );
  XNOR U24584 ( .A(n24683), .B(n24684), .Z(n24595) );
  AND U24585 ( .A(n393), .B(n24685), .Z(n24684) );
  XNOR U24586 ( .A(n24686), .B(n24683), .Z(n24685) );
  XNOR U24587 ( .A(n24687), .B(n24679), .Z(n24681) );
  IV U24588 ( .A(n24408), .Z(n24687) );
  XOR U24589 ( .A(n24688), .B(n24689), .Z(n24408) );
  AND U24590 ( .A(n401), .B(n24690), .Z(n24689) );
  AND U24591 ( .A(n24632), .B(n24613), .Z(n24679) );
  XNOR U24592 ( .A(n24691), .B(n24692), .Z(n24613) );
  AND U24593 ( .A(n393), .B(n24693), .Z(n24692) );
  XNOR U24594 ( .A(n24694), .B(n24691), .Z(n24693) );
  XNOR U24595 ( .A(n24695), .B(n24696), .Z(n393) );
  AND U24596 ( .A(n24697), .B(n24698), .Z(n24696) );
  XOR U24597 ( .A(n24642), .B(n24695), .Z(n24698) );
  AND U24598 ( .A(n24699), .B(n24700), .Z(n24642) );
  XOR U24599 ( .A(n24695), .B(n24639), .Z(n24697) );
  XNOR U24600 ( .A(n24701), .B(n24702), .Z(n24639) );
  AND U24601 ( .A(n397), .B(n24645), .Z(n24702) );
  XOR U24602 ( .A(n24643), .B(n24701), .Z(n24645) );
  XOR U24603 ( .A(n24703), .B(n24704), .Z(n24695) );
  AND U24604 ( .A(n24705), .B(n24706), .Z(n24704) );
  XNOR U24605 ( .A(n24703), .B(n24699), .Z(n24706) );
  IV U24606 ( .A(n24653), .Z(n24699) );
  XOR U24607 ( .A(n24707), .B(n24708), .Z(n24653) );
  XOR U24608 ( .A(n24709), .B(n24700), .Z(n24708) );
  AND U24609 ( .A(n24665), .B(n24710), .Z(n24700) );
  AND U24610 ( .A(n24711), .B(n24712), .Z(n24709) );
  XOR U24611 ( .A(n24713), .B(n24707), .Z(n24711) );
  XNOR U24612 ( .A(n24650), .B(n24703), .Z(n24705) );
  XNOR U24613 ( .A(n24714), .B(n24715), .Z(n24650) );
  AND U24614 ( .A(n397), .B(n24657), .Z(n24715) );
  XOR U24615 ( .A(n24714), .B(n24655), .Z(n24657) );
  XOR U24616 ( .A(n24716), .B(n24717), .Z(n24703) );
  AND U24617 ( .A(n24718), .B(n24719), .Z(n24717) );
  XNOR U24618 ( .A(n24716), .B(n24665), .Z(n24719) );
  XOR U24619 ( .A(n24720), .B(n24712), .Z(n24665) );
  XNOR U24620 ( .A(n24721), .B(n24707), .Z(n24712) );
  XOR U24621 ( .A(n24722), .B(n24723), .Z(n24707) );
  AND U24622 ( .A(n24724), .B(n24725), .Z(n24723) );
  XOR U24623 ( .A(n24726), .B(n24722), .Z(n24724) );
  XNOR U24624 ( .A(n24727), .B(n24728), .Z(n24721) );
  AND U24625 ( .A(n24729), .B(n24730), .Z(n24728) );
  XOR U24626 ( .A(n24727), .B(n24731), .Z(n24729) );
  XNOR U24627 ( .A(n24713), .B(n24710), .Z(n24720) );
  AND U24628 ( .A(n24732), .B(n24733), .Z(n24710) );
  XOR U24629 ( .A(n24734), .B(n24735), .Z(n24713) );
  AND U24630 ( .A(n24736), .B(n24737), .Z(n24735) );
  XOR U24631 ( .A(n24734), .B(n24738), .Z(n24736) );
  XNOR U24632 ( .A(n24662), .B(n24716), .Z(n24718) );
  XNOR U24633 ( .A(n24739), .B(n24740), .Z(n24662) );
  AND U24634 ( .A(n397), .B(n24668), .Z(n24740) );
  XOR U24635 ( .A(n24739), .B(n24666), .Z(n24668) );
  XOR U24636 ( .A(n24741), .B(n24742), .Z(n24716) );
  AND U24637 ( .A(n24743), .B(n24744), .Z(n24742) );
  XNOR U24638 ( .A(n24741), .B(n24732), .Z(n24744) );
  IV U24639 ( .A(n24674), .Z(n24732) );
  XNOR U24640 ( .A(n24745), .B(n24725), .Z(n24674) );
  XNOR U24641 ( .A(n24746), .B(n24731), .Z(n24725) );
  XOR U24642 ( .A(n24747), .B(n24748), .Z(n24731) );
  AND U24643 ( .A(n24749), .B(n24750), .Z(n24748) );
  XOR U24644 ( .A(n24747), .B(n24751), .Z(n24749) );
  XNOR U24645 ( .A(n24730), .B(n24722), .Z(n24746) );
  XOR U24646 ( .A(n24752), .B(n24753), .Z(n24722) );
  AND U24647 ( .A(n24754), .B(n24755), .Z(n24753) );
  XNOR U24648 ( .A(n24756), .B(n24752), .Z(n24754) );
  XNOR U24649 ( .A(n24757), .B(n24727), .Z(n24730) );
  XOR U24650 ( .A(n24758), .B(n24759), .Z(n24727) );
  AND U24651 ( .A(n24760), .B(n24761), .Z(n24759) );
  XOR U24652 ( .A(n24758), .B(n24762), .Z(n24760) );
  XNOR U24653 ( .A(n24763), .B(n24764), .Z(n24757) );
  AND U24654 ( .A(n24765), .B(n24766), .Z(n24764) );
  XNOR U24655 ( .A(n24763), .B(n24767), .Z(n24765) );
  XNOR U24656 ( .A(n24726), .B(n24733), .Z(n24745) );
  AND U24657 ( .A(n24686), .B(n24768), .Z(n24733) );
  XOR U24658 ( .A(n24738), .B(n24737), .Z(n24726) );
  XNOR U24659 ( .A(n24769), .B(n24734), .Z(n24737) );
  XOR U24660 ( .A(n24770), .B(n24771), .Z(n24734) );
  AND U24661 ( .A(n24772), .B(n24773), .Z(n24771) );
  XOR U24662 ( .A(n24770), .B(n24774), .Z(n24772) );
  XNOR U24663 ( .A(n24775), .B(n24776), .Z(n24769) );
  AND U24664 ( .A(n24777), .B(n24778), .Z(n24776) );
  XOR U24665 ( .A(n24775), .B(n24779), .Z(n24777) );
  XOR U24666 ( .A(n24780), .B(n24781), .Z(n24738) );
  AND U24667 ( .A(n24782), .B(n24783), .Z(n24781) );
  XOR U24668 ( .A(n24780), .B(n24784), .Z(n24782) );
  XNOR U24669 ( .A(n24671), .B(n24741), .Z(n24743) );
  XNOR U24670 ( .A(n24785), .B(n24786), .Z(n24671) );
  AND U24671 ( .A(n397), .B(n24678), .Z(n24786) );
  XOR U24672 ( .A(n24785), .B(n24676), .Z(n24678) );
  XOR U24673 ( .A(n24787), .B(n24788), .Z(n24741) );
  AND U24674 ( .A(n24789), .B(n24790), .Z(n24788) );
  XNOR U24675 ( .A(n24787), .B(n24686), .Z(n24790) );
  XOR U24676 ( .A(n24791), .B(n24755), .Z(n24686) );
  XNOR U24677 ( .A(n24792), .B(n24762), .Z(n24755) );
  XOR U24678 ( .A(n24751), .B(n24750), .Z(n24762) );
  XNOR U24679 ( .A(n24793), .B(n24747), .Z(n24750) );
  XOR U24680 ( .A(n24794), .B(n24795), .Z(n24747) );
  AND U24681 ( .A(n24796), .B(n24797), .Z(n24795) );
  XOR U24682 ( .A(n24794), .B(n24798), .Z(n24796) );
  XNOR U24683 ( .A(n24799), .B(n24800), .Z(n24793) );
  NOR U24684 ( .A(n24801), .B(n24802), .Z(n24800) );
  XNOR U24685 ( .A(n24799), .B(n24803), .Z(n24801) );
  XOR U24686 ( .A(n24804), .B(n24805), .Z(n24751) );
  NOR U24687 ( .A(n24806), .B(n24807), .Z(n24805) );
  XNOR U24688 ( .A(n24804), .B(n24808), .Z(n24806) );
  XNOR U24689 ( .A(n24761), .B(n24752), .Z(n24792) );
  XOR U24690 ( .A(n24809), .B(n24810), .Z(n24752) );
  NOR U24691 ( .A(n24811), .B(n24812), .Z(n24810) );
  XNOR U24692 ( .A(n24809), .B(n24813), .Z(n24811) );
  XOR U24693 ( .A(n24814), .B(n24767), .Z(n24761) );
  XNOR U24694 ( .A(n24815), .B(n24816), .Z(n24767) );
  NOR U24695 ( .A(n24817), .B(n24818), .Z(n24816) );
  XNOR U24696 ( .A(n24815), .B(n24819), .Z(n24817) );
  XNOR U24697 ( .A(n24766), .B(n24758), .Z(n24814) );
  XOR U24698 ( .A(n24820), .B(n24821), .Z(n24758) );
  AND U24699 ( .A(n24822), .B(n24823), .Z(n24821) );
  XOR U24700 ( .A(n24820), .B(n24824), .Z(n24822) );
  XNOR U24701 ( .A(n24825), .B(n24763), .Z(n24766) );
  XOR U24702 ( .A(n24826), .B(n24827), .Z(n24763) );
  AND U24703 ( .A(n24828), .B(n24829), .Z(n24827) );
  XOR U24704 ( .A(n24826), .B(n24830), .Z(n24828) );
  XNOR U24705 ( .A(n24831), .B(n24832), .Z(n24825) );
  NOR U24706 ( .A(n24833), .B(n24834), .Z(n24832) );
  XOR U24707 ( .A(n24831), .B(n24835), .Z(n24833) );
  XOR U24708 ( .A(n24756), .B(n24768), .Z(n24791) );
  NOR U24709 ( .A(n24694), .B(n24836), .Z(n24768) );
  XNOR U24710 ( .A(n24774), .B(n24773), .Z(n24756) );
  XNOR U24711 ( .A(n24837), .B(n24779), .Z(n24773) );
  XOR U24712 ( .A(n24838), .B(n24839), .Z(n24779) );
  NOR U24713 ( .A(n24840), .B(n24841), .Z(n24839) );
  XNOR U24714 ( .A(n24838), .B(n24842), .Z(n24840) );
  XNOR U24715 ( .A(n24778), .B(n24770), .Z(n24837) );
  XOR U24716 ( .A(n24843), .B(n24844), .Z(n24770) );
  AND U24717 ( .A(n24845), .B(n24846), .Z(n24844) );
  XNOR U24718 ( .A(n24843), .B(n24847), .Z(n24845) );
  XNOR U24719 ( .A(n24848), .B(n24775), .Z(n24778) );
  XOR U24720 ( .A(n24849), .B(n24850), .Z(n24775) );
  AND U24721 ( .A(n24851), .B(n24852), .Z(n24850) );
  XOR U24722 ( .A(n24849), .B(n24853), .Z(n24851) );
  XNOR U24723 ( .A(n24854), .B(n24855), .Z(n24848) );
  NOR U24724 ( .A(n24856), .B(n24857), .Z(n24855) );
  XOR U24725 ( .A(n24854), .B(n24858), .Z(n24856) );
  XOR U24726 ( .A(n24784), .B(n24783), .Z(n24774) );
  XNOR U24727 ( .A(n24859), .B(n24780), .Z(n24783) );
  XOR U24728 ( .A(n24860), .B(n24861), .Z(n24780) );
  AND U24729 ( .A(n24862), .B(n24863), .Z(n24861) );
  XOR U24730 ( .A(n24860), .B(n24864), .Z(n24862) );
  XNOR U24731 ( .A(n24865), .B(n24866), .Z(n24859) );
  NOR U24732 ( .A(n24867), .B(n24868), .Z(n24866) );
  XNOR U24733 ( .A(n24865), .B(n24869), .Z(n24867) );
  XOR U24734 ( .A(n24870), .B(n24871), .Z(n24784) );
  NOR U24735 ( .A(n24872), .B(n24873), .Z(n24871) );
  XNOR U24736 ( .A(n24870), .B(n24874), .Z(n24872) );
  XNOR U24737 ( .A(n24683), .B(n24787), .Z(n24789) );
  XNOR U24738 ( .A(n24875), .B(n24876), .Z(n24683) );
  AND U24739 ( .A(n397), .B(n24690), .Z(n24876) );
  XOR U24740 ( .A(n24875), .B(n24688), .Z(n24690) );
  AND U24741 ( .A(n24691), .B(n24694), .Z(n24787) );
  XOR U24742 ( .A(n24877), .B(n24836), .Z(n24694) );
  XNOR U24743 ( .A(p_input[2048]), .B(p_input[960]), .Z(n24836) );
  XOR U24744 ( .A(n24813), .B(n24812), .Z(n24877) );
  XOR U24745 ( .A(n24878), .B(n24824), .Z(n24812) );
  XOR U24746 ( .A(n24798), .B(n24797), .Z(n24824) );
  XNOR U24747 ( .A(n24879), .B(n24803), .Z(n24797) );
  XOR U24748 ( .A(p_input[2072]), .B(p_input[984]), .Z(n24803) );
  XOR U24749 ( .A(n24794), .B(n24802), .Z(n24879) );
  XOR U24750 ( .A(n24880), .B(n24799), .Z(n24802) );
  XOR U24751 ( .A(p_input[2070]), .B(p_input[982]), .Z(n24799) );
  XNOR U24752 ( .A(p_input[2071]), .B(p_input[983]), .Z(n24880) );
  XNOR U24753 ( .A(n16727), .B(p_input[978]), .Z(n24794) );
  XNOR U24754 ( .A(n24808), .B(n24807), .Z(n24798) );
  XOR U24755 ( .A(n24881), .B(n24804), .Z(n24807) );
  XOR U24756 ( .A(p_input[2067]), .B(p_input[979]), .Z(n24804) );
  XNOR U24757 ( .A(p_input[2068]), .B(p_input[980]), .Z(n24881) );
  XOR U24758 ( .A(p_input[2069]), .B(p_input[981]), .Z(n24808) );
  XNOR U24759 ( .A(n24823), .B(n24809), .Z(n24878) );
  XNOR U24760 ( .A(n16729), .B(p_input[961]), .Z(n24809) );
  XNOR U24761 ( .A(n24882), .B(n24830), .Z(n24823) );
  XNOR U24762 ( .A(n24819), .B(n24818), .Z(n24830) );
  XOR U24763 ( .A(n24883), .B(n24815), .Z(n24818) );
  XNOR U24764 ( .A(n16444), .B(p_input[986]), .Z(n24815) );
  XNOR U24765 ( .A(p_input[2075]), .B(p_input[987]), .Z(n24883) );
  XOR U24766 ( .A(p_input[2076]), .B(p_input[988]), .Z(n24819) );
  XNOR U24767 ( .A(n24829), .B(n24820), .Z(n24882) );
  XNOR U24768 ( .A(n16732), .B(p_input[977]), .Z(n24820) );
  XOR U24769 ( .A(n24884), .B(n24835), .Z(n24829) );
  XNOR U24770 ( .A(p_input[2079]), .B(p_input[991]), .Z(n24835) );
  XOR U24771 ( .A(n24826), .B(n24834), .Z(n24884) );
  XOR U24772 ( .A(n24885), .B(n24831), .Z(n24834) );
  XOR U24773 ( .A(p_input[2077]), .B(p_input[989]), .Z(n24831) );
  XNOR U24774 ( .A(p_input[2078]), .B(p_input[990]), .Z(n24885) );
  XNOR U24775 ( .A(n16448), .B(p_input[985]), .Z(n24826) );
  XNOR U24776 ( .A(n24847), .B(n24846), .Z(n24813) );
  XNOR U24777 ( .A(n24886), .B(n24853), .Z(n24846) );
  XNOR U24778 ( .A(n24842), .B(n24841), .Z(n24853) );
  XOR U24779 ( .A(n24887), .B(n24838), .Z(n24841) );
  XNOR U24780 ( .A(n16737), .B(p_input[971]), .Z(n24838) );
  XNOR U24781 ( .A(p_input[2060]), .B(p_input[972]), .Z(n24887) );
  XOR U24782 ( .A(p_input[2061]), .B(p_input[973]), .Z(n24842) );
  XNOR U24783 ( .A(n24852), .B(n24843), .Z(n24886) );
  XNOR U24784 ( .A(n16452), .B(p_input[962]), .Z(n24843) );
  XOR U24785 ( .A(n24888), .B(n24858), .Z(n24852) );
  XNOR U24786 ( .A(p_input[2064]), .B(p_input[976]), .Z(n24858) );
  XOR U24787 ( .A(n24849), .B(n24857), .Z(n24888) );
  XOR U24788 ( .A(n24889), .B(n24854), .Z(n24857) );
  XOR U24789 ( .A(p_input[2062]), .B(p_input[974]), .Z(n24854) );
  XNOR U24790 ( .A(p_input[2063]), .B(p_input[975]), .Z(n24889) );
  XNOR U24791 ( .A(n16740), .B(p_input[970]), .Z(n24849) );
  XNOR U24792 ( .A(n24864), .B(n24863), .Z(n24847) );
  XNOR U24793 ( .A(n24890), .B(n24869), .Z(n24863) );
  XOR U24794 ( .A(p_input[2057]), .B(p_input[969]), .Z(n24869) );
  XOR U24795 ( .A(n24860), .B(n24868), .Z(n24890) );
  XOR U24796 ( .A(n24891), .B(n24865), .Z(n24868) );
  XOR U24797 ( .A(p_input[2055]), .B(p_input[967]), .Z(n24865) );
  XNOR U24798 ( .A(p_input[2056]), .B(p_input[968]), .Z(n24891) );
  XNOR U24799 ( .A(n16459), .B(p_input[963]), .Z(n24860) );
  XNOR U24800 ( .A(n24874), .B(n24873), .Z(n24864) );
  XOR U24801 ( .A(n24892), .B(n24870), .Z(n24873) );
  XOR U24802 ( .A(p_input[2052]), .B(p_input[964]), .Z(n24870) );
  XNOR U24803 ( .A(p_input[2053]), .B(p_input[965]), .Z(n24892) );
  XOR U24804 ( .A(p_input[2054]), .B(p_input[966]), .Z(n24874) );
  XNOR U24805 ( .A(n24893), .B(n24894), .Z(n24691) );
  AND U24806 ( .A(n397), .B(n24895), .Z(n24894) );
  XNOR U24807 ( .A(n24896), .B(n24897), .Z(n397) );
  AND U24808 ( .A(n24898), .B(n24899), .Z(n24897) );
  XOR U24809 ( .A(n24896), .B(n24701), .Z(n24899) );
  XNOR U24810 ( .A(n24896), .B(n24643), .Z(n24898) );
  XOR U24811 ( .A(n24900), .B(n24901), .Z(n24896) );
  AND U24812 ( .A(n24902), .B(n24903), .Z(n24901) );
  XNOR U24813 ( .A(n24714), .B(n24900), .Z(n24903) );
  XOR U24814 ( .A(n24900), .B(n24655), .Z(n24902) );
  XOR U24815 ( .A(n24904), .B(n24905), .Z(n24900) );
  AND U24816 ( .A(n24906), .B(n24907), .Z(n24905) );
  XNOR U24817 ( .A(n24739), .B(n24904), .Z(n24907) );
  XOR U24818 ( .A(n24904), .B(n24666), .Z(n24906) );
  XOR U24819 ( .A(n24908), .B(n24909), .Z(n24904) );
  AND U24820 ( .A(n24910), .B(n24911), .Z(n24909) );
  XOR U24821 ( .A(n24908), .B(n24676), .Z(n24910) );
  XOR U24822 ( .A(n24912), .B(n24913), .Z(n24632) );
  AND U24823 ( .A(n401), .B(n24895), .Z(n24913) );
  XNOR U24824 ( .A(n24893), .B(n24912), .Z(n24895) );
  XNOR U24825 ( .A(n24914), .B(n24915), .Z(n401) );
  AND U24826 ( .A(n24916), .B(n24917), .Z(n24915) );
  XNOR U24827 ( .A(n24918), .B(n24914), .Z(n24917) );
  IV U24828 ( .A(n24701), .Z(n24918) );
  XNOR U24829 ( .A(n24919), .B(n24920), .Z(n24701) );
  AND U24830 ( .A(n404), .B(n24921), .Z(n24920) );
  XNOR U24831 ( .A(n24919), .B(n24922), .Z(n24921) );
  XNOR U24832 ( .A(n24643), .B(n24914), .Z(n24916) );
  XOR U24833 ( .A(n24923), .B(n24924), .Z(n24643) );
  AND U24834 ( .A(n412), .B(n24925), .Z(n24924) );
  XOR U24835 ( .A(n24926), .B(n24927), .Z(n24914) );
  AND U24836 ( .A(n24928), .B(n24929), .Z(n24927) );
  XNOR U24837 ( .A(n24926), .B(n24714), .Z(n24929) );
  XNOR U24838 ( .A(n24930), .B(n24931), .Z(n24714) );
  AND U24839 ( .A(n404), .B(n24932), .Z(n24931) );
  XOR U24840 ( .A(n24933), .B(n24930), .Z(n24932) );
  XNOR U24841 ( .A(n24934), .B(n24926), .Z(n24928) );
  IV U24842 ( .A(n24655), .Z(n24934) );
  XOR U24843 ( .A(n24935), .B(n24936), .Z(n24655) );
  AND U24844 ( .A(n412), .B(n24937), .Z(n24936) );
  XOR U24845 ( .A(n24938), .B(n24939), .Z(n24926) );
  AND U24846 ( .A(n24940), .B(n24941), .Z(n24939) );
  XNOR U24847 ( .A(n24938), .B(n24739), .Z(n24941) );
  XNOR U24848 ( .A(n24942), .B(n24943), .Z(n24739) );
  AND U24849 ( .A(n404), .B(n24944), .Z(n24943) );
  XNOR U24850 ( .A(n24945), .B(n24942), .Z(n24944) );
  XOR U24851 ( .A(n24666), .B(n24938), .Z(n24940) );
  XOR U24852 ( .A(n24946), .B(n24947), .Z(n24666) );
  AND U24853 ( .A(n412), .B(n24948), .Z(n24947) );
  XOR U24854 ( .A(n24908), .B(n24949), .Z(n24938) );
  AND U24855 ( .A(n24950), .B(n24911), .Z(n24949) );
  XNOR U24856 ( .A(n24785), .B(n24908), .Z(n24911) );
  XNOR U24857 ( .A(n24951), .B(n24952), .Z(n24785) );
  AND U24858 ( .A(n404), .B(n24953), .Z(n24952) );
  XOR U24859 ( .A(n24954), .B(n24951), .Z(n24953) );
  XNOR U24860 ( .A(n24955), .B(n24908), .Z(n24950) );
  IV U24861 ( .A(n24676), .Z(n24955) );
  XOR U24862 ( .A(n24956), .B(n24957), .Z(n24676) );
  AND U24863 ( .A(n412), .B(n24958), .Z(n24957) );
  XOR U24864 ( .A(n24959), .B(n24960), .Z(n24908) );
  AND U24865 ( .A(n24961), .B(n24962), .Z(n24960) );
  XNOR U24866 ( .A(n24959), .B(n24875), .Z(n24962) );
  XNOR U24867 ( .A(n24963), .B(n24964), .Z(n24875) );
  AND U24868 ( .A(n404), .B(n24965), .Z(n24964) );
  XNOR U24869 ( .A(n24966), .B(n24963), .Z(n24965) );
  XNOR U24870 ( .A(n24967), .B(n24959), .Z(n24961) );
  IV U24871 ( .A(n24688), .Z(n24967) );
  XOR U24872 ( .A(n24968), .B(n24969), .Z(n24688) );
  AND U24873 ( .A(n412), .B(n24970), .Z(n24969) );
  AND U24874 ( .A(n24912), .B(n24893), .Z(n24959) );
  XNOR U24875 ( .A(n24971), .B(n24972), .Z(n24893) );
  AND U24876 ( .A(n404), .B(n24973), .Z(n24972) );
  XNOR U24877 ( .A(n24974), .B(n24971), .Z(n24973) );
  XNOR U24878 ( .A(n24975), .B(n24976), .Z(n404) );
  AND U24879 ( .A(n24977), .B(n24978), .Z(n24976) );
  XOR U24880 ( .A(n24922), .B(n24975), .Z(n24978) );
  AND U24881 ( .A(n24979), .B(n24980), .Z(n24922) );
  XOR U24882 ( .A(n24975), .B(n24919), .Z(n24977) );
  XNOR U24883 ( .A(n24981), .B(n24982), .Z(n24919) );
  AND U24884 ( .A(n408), .B(n24925), .Z(n24982) );
  XOR U24885 ( .A(n24923), .B(n24981), .Z(n24925) );
  XOR U24886 ( .A(n24983), .B(n24984), .Z(n24975) );
  AND U24887 ( .A(n24985), .B(n24986), .Z(n24984) );
  XNOR U24888 ( .A(n24983), .B(n24979), .Z(n24986) );
  IV U24889 ( .A(n24933), .Z(n24979) );
  XOR U24890 ( .A(n24987), .B(n24988), .Z(n24933) );
  XOR U24891 ( .A(n24989), .B(n24980), .Z(n24988) );
  AND U24892 ( .A(n24945), .B(n24990), .Z(n24980) );
  AND U24893 ( .A(n24991), .B(n24992), .Z(n24989) );
  XOR U24894 ( .A(n24993), .B(n24987), .Z(n24991) );
  XNOR U24895 ( .A(n24930), .B(n24983), .Z(n24985) );
  XNOR U24896 ( .A(n24994), .B(n24995), .Z(n24930) );
  AND U24897 ( .A(n408), .B(n24937), .Z(n24995) );
  XOR U24898 ( .A(n24994), .B(n24935), .Z(n24937) );
  XOR U24899 ( .A(n24996), .B(n24997), .Z(n24983) );
  AND U24900 ( .A(n24998), .B(n24999), .Z(n24997) );
  XNOR U24901 ( .A(n24996), .B(n24945), .Z(n24999) );
  XOR U24902 ( .A(n25000), .B(n24992), .Z(n24945) );
  XNOR U24903 ( .A(n25001), .B(n24987), .Z(n24992) );
  XOR U24904 ( .A(n25002), .B(n25003), .Z(n24987) );
  AND U24905 ( .A(n25004), .B(n25005), .Z(n25003) );
  XOR U24906 ( .A(n25006), .B(n25002), .Z(n25004) );
  XNOR U24907 ( .A(n25007), .B(n25008), .Z(n25001) );
  AND U24908 ( .A(n25009), .B(n25010), .Z(n25008) );
  XOR U24909 ( .A(n25007), .B(n25011), .Z(n25009) );
  XNOR U24910 ( .A(n24993), .B(n24990), .Z(n25000) );
  AND U24911 ( .A(n25012), .B(n25013), .Z(n24990) );
  XOR U24912 ( .A(n25014), .B(n25015), .Z(n24993) );
  AND U24913 ( .A(n25016), .B(n25017), .Z(n25015) );
  XOR U24914 ( .A(n25014), .B(n25018), .Z(n25016) );
  XNOR U24915 ( .A(n24942), .B(n24996), .Z(n24998) );
  XNOR U24916 ( .A(n25019), .B(n25020), .Z(n24942) );
  AND U24917 ( .A(n408), .B(n24948), .Z(n25020) );
  XOR U24918 ( .A(n25019), .B(n24946), .Z(n24948) );
  XOR U24919 ( .A(n25021), .B(n25022), .Z(n24996) );
  AND U24920 ( .A(n25023), .B(n25024), .Z(n25022) );
  XNOR U24921 ( .A(n25021), .B(n25012), .Z(n25024) );
  IV U24922 ( .A(n24954), .Z(n25012) );
  XNOR U24923 ( .A(n25025), .B(n25005), .Z(n24954) );
  XNOR U24924 ( .A(n25026), .B(n25011), .Z(n25005) );
  XOR U24925 ( .A(n25027), .B(n25028), .Z(n25011) );
  AND U24926 ( .A(n25029), .B(n25030), .Z(n25028) );
  XOR U24927 ( .A(n25027), .B(n25031), .Z(n25029) );
  XNOR U24928 ( .A(n25010), .B(n25002), .Z(n25026) );
  XOR U24929 ( .A(n25032), .B(n25033), .Z(n25002) );
  AND U24930 ( .A(n25034), .B(n25035), .Z(n25033) );
  XNOR U24931 ( .A(n25036), .B(n25032), .Z(n25034) );
  XNOR U24932 ( .A(n25037), .B(n25007), .Z(n25010) );
  XOR U24933 ( .A(n25038), .B(n25039), .Z(n25007) );
  AND U24934 ( .A(n25040), .B(n25041), .Z(n25039) );
  XOR U24935 ( .A(n25038), .B(n25042), .Z(n25040) );
  XNOR U24936 ( .A(n25043), .B(n25044), .Z(n25037) );
  AND U24937 ( .A(n25045), .B(n25046), .Z(n25044) );
  XNOR U24938 ( .A(n25043), .B(n25047), .Z(n25045) );
  XNOR U24939 ( .A(n25006), .B(n25013), .Z(n25025) );
  AND U24940 ( .A(n24966), .B(n25048), .Z(n25013) );
  XOR U24941 ( .A(n25018), .B(n25017), .Z(n25006) );
  XNOR U24942 ( .A(n25049), .B(n25014), .Z(n25017) );
  XOR U24943 ( .A(n25050), .B(n25051), .Z(n25014) );
  AND U24944 ( .A(n25052), .B(n25053), .Z(n25051) );
  XOR U24945 ( .A(n25050), .B(n25054), .Z(n25052) );
  XNOR U24946 ( .A(n25055), .B(n25056), .Z(n25049) );
  AND U24947 ( .A(n25057), .B(n25058), .Z(n25056) );
  XOR U24948 ( .A(n25055), .B(n25059), .Z(n25057) );
  XOR U24949 ( .A(n25060), .B(n25061), .Z(n25018) );
  AND U24950 ( .A(n25062), .B(n25063), .Z(n25061) );
  XOR U24951 ( .A(n25060), .B(n25064), .Z(n25062) );
  XNOR U24952 ( .A(n24951), .B(n25021), .Z(n25023) );
  XNOR U24953 ( .A(n25065), .B(n25066), .Z(n24951) );
  AND U24954 ( .A(n408), .B(n24958), .Z(n25066) );
  XOR U24955 ( .A(n25065), .B(n24956), .Z(n24958) );
  XOR U24956 ( .A(n25067), .B(n25068), .Z(n25021) );
  AND U24957 ( .A(n25069), .B(n25070), .Z(n25068) );
  XNOR U24958 ( .A(n25067), .B(n24966), .Z(n25070) );
  XOR U24959 ( .A(n25071), .B(n25035), .Z(n24966) );
  XNOR U24960 ( .A(n25072), .B(n25042), .Z(n25035) );
  XOR U24961 ( .A(n25031), .B(n25030), .Z(n25042) );
  XNOR U24962 ( .A(n25073), .B(n25027), .Z(n25030) );
  XOR U24963 ( .A(n25074), .B(n25075), .Z(n25027) );
  AND U24964 ( .A(n25076), .B(n25077), .Z(n25075) );
  XNOR U24965 ( .A(n25078), .B(n25079), .Z(n25076) );
  IV U24966 ( .A(n25074), .Z(n25078) );
  XNOR U24967 ( .A(n25080), .B(n25081), .Z(n25073) );
  NOR U24968 ( .A(n25082), .B(n25083), .Z(n25081) );
  XNOR U24969 ( .A(n25080), .B(n25084), .Z(n25082) );
  XOR U24970 ( .A(n25085), .B(n25086), .Z(n25031) );
  NOR U24971 ( .A(n25087), .B(n25088), .Z(n25086) );
  XNOR U24972 ( .A(n25085), .B(n25089), .Z(n25087) );
  XNOR U24973 ( .A(n25041), .B(n25032), .Z(n25072) );
  XOR U24974 ( .A(n25090), .B(n25091), .Z(n25032) );
  AND U24975 ( .A(n25092), .B(n25093), .Z(n25091) );
  XOR U24976 ( .A(n25090), .B(n25094), .Z(n25092) );
  XOR U24977 ( .A(n25095), .B(n25047), .Z(n25041) );
  XOR U24978 ( .A(n25096), .B(n25097), .Z(n25047) );
  NOR U24979 ( .A(n25098), .B(n25099), .Z(n25097) );
  XOR U24980 ( .A(n25096), .B(n25100), .Z(n25098) );
  XNOR U24981 ( .A(n25046), .B(n25038), .Z(n25095) );
  XOR U24982 ( .A(n25101), .B(n25102), .Z(n25038) );
  AND U24983 ( .A(n25103), .B(n25104), .Z(n25102) );
  XOR U24984 ( .A(n25101), .B(n25105), .Z(n25103) );
  XNOR U24985 ( .A(n25106), .B(n25043), .Z(n25046) );
  XOR U24986 ( .A(n25107), .B(n25108), .Z(n25043) );
  AND U24987 ( .A(n25109), .B(n25110), .Z(n25108) );
  XNOR U24988 ( .A(n25111), .B(n25112), .Z(n25109) );
  IV U24989 ( .A(n25107), .Z(n25111) );
  XNOR U24990 ( .A(n25113), .B(n25114), .Z(n25106) );
  NOR U24991 ( .A(n25115), .B(n25116), .Z(n25114) );
  XNOR U24992 ( .A(n25113), .B(n25117), .Z(n25115) );
  XOR U24993 ( .A(n25036), .B(n25048), .Z(n25071) );
  NOR U24994 ( .A(n24974), .B(n25118), .Z(n25048) );
  XNOR U24995 ( .A(n25054), .B(n25053), .Z(n25036) );
  XNOR U24996 ( .A(n25119), .B(n25059), .Z(n25053) );
  XNOR U24997 ( .A(n25120), .B(n25121), .Z(n25059) );
  NOR U24998 ( .A(n25122), .B(n25123), .Z(n25121) );
  XOR U24999 ( .A(n25120), .B(n25124), .Z(n25122) );
  XNOR U25000 ( .A(n25058), .B(n25050), .Z(n25119) );
  XOR U25001 ( .A(n25125), .B(n25126), .Z(n25050) );
  AND U25002 ( .A(n25127), .B(n25128), .Z(n25126) );
  XOR U25003 ( .A(n25125), .B(n25129), .Z(n25127) );
  XNOR U25004 ( .A(n25130), .B(n25055), .Z(n25058) );
  XOR U25005 ( .A(n25131), .B(n25132), .Z(n25055) );
  AND U25006 ( .A(n25133), .B(n25134), .Z(n25132) );
  XNOR U25007 ( .A(n25135), .B(n25136), .Z(n25133) );
  IV U25008 ( .A(n25131), .Z(n25135) );
  XNOR U25009 ( .A(n25137), .B(n25138), .Z(n25130) );
  NOR U25010 ( .A(n25139), .B(n25140), .Z(n25138) );
  XNOR U25011 ( .A(n25137), .B(n25141), .Z(n25139) );
  XOR U25012 ( .A(n25064), .B(n25063), .Z(n25054) );
  XNOR U25013 ( .A(n25142), .B(n25060), .Z(n25063) );
  XOR U25014 ( .A(n25143), .B(n25144), .Z(n25060) );
  AND U25015 ( .A(n25145), .B(n25146), .Z(n25144) );
  XOR U25016 ( .A(n25143), .B(n25147), .Z(n25145) );
  XNOR U25017 ( .A(n25148), .B(n25149), .Z(n25142) );
  NOR U25018 ( .A(n25150), .B(n25151), .Z(n25149) );
  XNOR U25019 ( .A(n25148), .B(n25152), .Z(n25150) );
  XOR U25020 ( .A(n25153), .B(n25154), .Z(n25064) );
  NOR U25021 ( .A(n25155), .B(n25156), .Z(n25154) );
  XNOR U25022 ( .A(n25153), .B(n25157), .Z(n25155) );
  XNOR U25023 ( .A(n24963), .B(n25067), .Z(n25069) );
  XNOR U25024 ( .A(n25158), .B(n25159), .Z(n24963) );
  AND U25025 ( .A(n408), .B(n24970), .Z(n25159) );
  XOR U25026 ( .A(n25158), .B(n24968), .Z(n24970) );
  AND U25027 ( .A(n24971), .B(n24974), .Z(n25067) );
  XOR U25028 ( .A(n25160), .B(n25118), .Z(n24974) );
  XNOR U25029 ( .A(p_input[2048]), .B(p_input[992]), .Z(n25118) );
  XNOR U25030 ( .A(n25094), .B(n25093), .Z(n25160) );
  XNOR U25031 ( .A(n25161), .B(n25105), .Z(n25093) );
  XOR U25032 ( .A(n25079), .B(n25077), .Z(n25105) );
  XNOR U25033 ( .A(n25162), .B(n25084), .Z(n25077) );
  XOR U25034 ( .A(p_input[1016]), .B(p_input[2072]), .Z(n25084) );
  XOR U25035 ( .A(n25074), .B(n25083), .Z(n25162) );
  XOR U25036 ( .A(n25163), .B(n25080), .Z(n25083) );
  XOR U25037 ( .A(p_input[1014]), .B(p_input[2070]), .Z(n25080) );
  XOR U25038 ( .A(p_input[1015]), .B(n17295), .Z(n25163) );
  XOR U25039 ( .A(p_input[1010]), .B(p_input[2066]), .Z(n25074) );
  XNOR U25040 ( .A(n25089), .B(n25088), .Z(n25079) );
  XOR U25041 ( .A(n25164), .B(n25085), .Z(n25088) );
  XOR U25042 ( .A(p_input[1011]), .B(p_input[2067]), .Z(n25085) );
  XOR U25043 ( .A(p_input[1012]), .B(n17297), .Z(n25164) );
  XOR U25044 ( .A(p_input[1013]), .B(p_input[2069]), .Z(n25089) );
  XNOR U25045 ( .A(n25104), .B(n25090), .Z(n25161) );
  XNOR U25046 ( .A(n16729), .B(p_input[993]), .Z(n25090) );
  XNOR U25047 ( .A(n25165), .B(n25112), .Z(n25104) );
  XNOR U25048 ( .A(n25100), .B(n25099), .Z(n25112) );
  XNOR U25049 ( .A(n25166), .B(n25096), .Z(n25099) );
  XNOR U25050 ( .A(p_input[1018]), .B(p_input[2074]), .Z(n25096) );
  XOR U25051 ( .A(p_input[1019]), .B(n17300), .Z(n25166) );
  XOR U25052 ( .A(p_input[1020]), .B(p_input[2076]), .Z(n25100) );
  XOR U25053 ( .A(n25110), .B(n25167), .Z(n25165) );
  IV U25054 ( .A(n25101), .Z(n25167) );
  XOR U25055 ( .A(p_input[1009]), .B(p_input[2065]), .Z(n25101) );
  XNOR U25056 ( .A(n25168), .B(n25117), .Z(n25110) );
  XNOR U25057 ( .A(p_input[1023]), .B(n17303), .Z(n25117) );
  XOR U25058 ( .A(n25107), .B(n25116), .Z(n25168) );
  XOR U25059 ( .A(n25169), .B(n25113), .Z(n25116) );
  XOR U25060 ( .A(p_input[1021]), .B(p_input[2077]), .Z(n25113) );
  XOR U25061 ( .A(p_input[1022]), .B(n17305), .Z(n25169) );
  XOR U25062 ( .A(p_input[1017]), .B(p_input[2073]), .Z(n25107) );
  XOR U25063 ( .A(n25129), .B(n25128), .Z(n25094) );
  XNOR U25064 ( .A(n25170), .B(n25136), .Z(n25128) );
  XNOR U25065 ( .A(n25124), .B(n25123), .Z(n25136) );
  XNOR U25066 ( .A(n25171), .B(n25120), .Z(n25123) );
  XNOR U25067 ( .A(p_input[1003]), .B(p_input[2059]), .Z(n25120) );
  XOR U25068 ( .A(p_input[1004]), .B(n16451), .Z(n25171) );
  XOR U25069 ( .A(p_input[1005]), .B(p_input[2061]), .Z(n25124) );
  XNOR U25070 ( .A(n25134), .B(n25125), .Z(n25170) );
  XNOR U25071 ( .A(n16452), .B(p_input[994]), .Z(n25125) );
  XNOR U25072 ( .A(n25172), .B(n25141), .Z(n25134) );
  XNOR U25073 ( .A(p_input[1008]), .B(n16454), .Z(n25141) );
  XOR U25074 ( .A(n25131), .B(n25140), .Z(n25172) );
  XOR U25075 ( .A(n25173), .B(n25137), .Z(n25140) );
  XOR U25076 ( .A(p_input[1006]), .B(p_input[2062]), .Z(n25137) );
  XOR U25077 ( .A(p_input[1007]), .B(n16456), .Z(n25173) );
  XOR U25078 ( .A(p_input[1002]), .B(p_input[2058]), .Z(n25131) );
  XOR U25079 ( .A(n25147), .B(n25146), .Z(n25129) );
  XNOR U25080 ( .A(n25174), .B(n25152), .Z(n25146) );
  XOR U25081 ( .A(p_input[1001]), .B(p_input[2057]), .Z(n25152) );
  XOR U25082 ( .A(n25143), .B(n25151), .Z(n25174) );
  XOR U25083 ( .A(n25175), .B(n25148), .Z(n25151) );
  XOR U25084 ( .A(p_input[2055]), .B(p_input[999]), .Z(n25148) );
  XOR U25085 ( .A(p_input[1000]), .B(n17312), .Z(n25175) );
  XNOR U25086 ( .A(n16459), .B(p_input[995]), .Z(n25143) );
  IV U25087 ( .A(p_input[2051]), .Z(n16459) );
  XNOR U25088 ( .A(n25157), .B(n25156), .Z(n25147) );
  XOR U25089 ( .A(n25176), .B(n25153), .Z(n25156) );
  XOR U25090 ( .A(p_input[2052]), .B(p_input[996]), .Z(n25153) );
  XNOR U25091 ( .A(p_input[2053]), .B(p_input[997]), .Z(n25176) );
  XOR U25092 ( .A(p_input[2054]), .B(p_input[998]), .Z(n25157) );
  XNOR U25093 ( .A(n25177), .B(n25178), .Z(n24971) );
  AND U25094 ( .A(n408), .B(n25179), .Z(n25178) );
  XNOR U25095 ( .A(n25180), .B(n25181), .Z(n408) );
  AND U25096 ( .A(n25182), .B(n25183), .Z(n25181) );
  XOR U25097 ( .A(n25180), .B(n24981), .Z(n25183) );
  XNOR U25098 ( .A(n25180), .B(n24923), .Z(n25182) );
  XOR U25099 ( .A(n25184), .B(n25185), .Z(n25180) );
  AND U25100 ( .A(n25186), .B(n25187), .Z(n25185) );
  XNOR U25101 ( .A(n24994), .B(n25184), .Z(n25187) );
  XOR U25102 ( .A(n25184), .B(n24935), .Z(n25186) );
  XOR U25103 ( .A(n25188), .B(n25189), .Z(n25184) );
  AND U25104 ( .A(n25190), .B(n25191), .Z(n25189) );
  XNOR U25105 ( .A(n25019), .B(n25188), .Z(n25191) );
  XOR U25106 ( .A(n25188), .B(n24946), .Z(n25190) );
  XOR U25107 ( .A(n25192), .B(n25193), .Z(n25188) );
  AND U25108 ( .A(n25194), .B(n25195), .Z(n25193) );
  XOR U25109 ( .A(n25192), .B(n24956), .Z(n25194) );
  XOR U25110 ( .A(n25196), .B(n25197), .Z(n24912) );
  AND U25111 ( .A(n412), .B(n25179), .Z(n25197) );
  XNOR U25112 ( .A(n25177), .B(n25196), .Z(n25179) );
  XNOR U25113 ( .A(n25198), .B(n25199), .Z(n412) );
  AND U25114 ( .A(n25200), .B(n25201), .Z(n25199) );
  XNOR U25115 ( .A(n25202), .B(n25198), .Z(n25201) );
  IV U25116 ( .A(n24981), .Z(n25202) );
  XNOR U25117 ( .A(n25203), .B(n25204), .Z(n24981) );
  AND U25118 ( .A(n415), .B(n25205), .Z(n25204) );
  XNOR U25119 ( .A(n25203), .B(n25206), .Z(n25205) );
  XNOR U25120 ( .A(n24923), .B(n25198), .Z(n25200) );
  XOR U25121 ( .A(n25207), .B(n25208), .Z(n24923) );
  AND U25122 ( .A(n423), .B(n25209), .Z(n25208) );
  XOR U25123 ( .A(n25210), .B(n25211), .Z(n25198) );
  AND U25124 ( .A(n25212), .B(n25213), .Z(n25211) );
  XNOR U25125 ( .A(n25210), .B(n24994), .Z(n25213) );
  XNOR U25126 ( .A(n25214), .B(n25215), .Z(n24994) );
  AND U25127 ( .A(n415), .B(n25216), .Z(n25215) );
  XOR U25128 ( .A(n25217), .B(n25214), .Z(n25216) );
  XNOR U25129 ( .A(n25218), .B(n25210), .Z(n25212) );
  IV U25130 ( .A(n24935), .Z(n25218) );
  XOR U25131 ( .A(n25219), .B(n25220), .Z(n24935) );
  AND U25132 ( .A(n423), .B(n25221), .Z(n25220) );
  XOR U25133 ( .A(n25222), .B(n25223), .Z(n25210) );
  AND U25134 ( .A(n25224), .B(n25225), .Z(n25223) );
  XNOR U25135 ( .A(n25222), .B(n25019), .Z(n25225) );
  XNOR U25136 ( .A(n25226), .B(n25227), .Z(n25019) );
  AND U25137 ( .A(n415), .B(n25228), .Z(n25227) );
  XNOR U25138 ( .A(n25229), .B(n25226), .Z(n25228) );
  XOR U25139 ( .A(n24946), .B(n25222), .Z(n25224) );
  XOR U25140 ( .A(n25230), .B(n25231), .Z(n24946) );
  AND U25141 ( .A(n423), .B(n25232), .Z(n25231) );
  XOR U25142 ( .A(n25192), .B(n25233), .Z(n25222) );
  AND U25143 ( .A(n25234), .B(n25195), .Z(n25233) );
  XNOR U25144 ( .A(n25065), .B(n25192), .Z(n25195) );
  XNOR U25145 ( .A(n25235), .B(n25236), .Z(n25065) );
  AND U25146 ( .A(n415), .B(n25237), .Z(n25236) );
  XOR U25147 ( .A(n25238), .B(n25235), .Z(n25237) );
  XNOR U25148 ( .A(n25239), .B(n25192), .Z(n25234) );
  IV U25149 ( .A(n24956), .Z(n25239) );
  XOR U25150 ( .A(n25240), .B(n25241), .Z(n24956) );
  AND U25151 ( .A(n423), .B(n25242), .Z(n25241) );
  XOR U25152 ( .A(n25243), .B(n25244), .Z(n25192) );
  AND U25153 ( .A(n25245), .B(n25246), .Z(n25244) );
  XNOR U25154 ( .A(n25243), .B(n25158), .Z(n25246) );
  XNOR U25155 ( .A(n25247), .B(n25248), .Z(n25158) );
  AND U25156 ( .A(n415), .B(n25249), .Z(n25248) );
  XNOR U25157 ( .A(n25250), .B(n25247), .Z(n25249) );
  XNOR U25158 ( .A(n25251), .B(n25243), .Z(n25245) );
  IV U25159 ( .A(n24968), .Z(n25251) );
  XOR U25160 ( .A(n25252), .B(n25253), .Z(n24968) );
  AND U25161 ( .A(n423), .B(n25254), .Z(n25253) );
  AND U25162 ( .A(n25196), .B(n25177), .Z(n25243) );
  XNOR U25163 ( .A(n25255), .B(n25256), .Z(n25177) );
  AND U25164 ( .A(n415), .B(n25257), .Z(n25256) );
  XNOR U25165 ( .A(n25258), .B(n25255), .Z(n25257) );
  XNOR U25166 ( .A(n25259), .B(n25260), .Z(n415) );
  AND U25167 ( .A(n25261), .B(n25262), .Z(n25260) );
  XOR U25168 ( .A(n25206), .B(n25259), .Z(n25262) );
  AND U25169 ( .A(n25263), .B(n25264), .Z(n25206) );
  XOR U25170 ( .A(n25259), .B(n25203), .Z(n25261) );
  XNOR U25171 ( .A(n25265), .B(n25266), .Z(n25203) );
  AND U25172 ( .A(n419), .B(n25209), .Z(n25266) );
  XOR U25173 ( .A(n25207), .B(n25265), .Z(n25209) );
  XOR U25174 ( .A(n25267), .B(n25268), .Z(n25259) );
  AND U25175 ( .A(n25269), .B(n25270), .Z(n25268) );
  XNOR U25176 ( .A(n25267), .B(n25263), .Z(n25270) );
  IV U25177 ( .A(n25217), .Z(n25263) );
  XOR U25178 ( .A(n25271), .B(n25272), .Z(n25217) );
  XOR U25179 ( .A(n25273), .B(n25264), .Z(n25272) );
  AND U25180 ( .A(n25229), .B(n25274), .Z(n25264) );
  AND U25181 ( .A(n25275), .B(n25276), .Z(n25273) );
  XOR U25182 ( .A(n25277), .B(n25271), .Z(n25275) );
  XNOR U25183 ( .A(n25214), .B(n25267), .Z(n25269) );
  XNOR U25184 ( .A(n25278), .B(n25279), .Z(n25214) );
  AND U25185 ( .A(n419), .B(n25221), .Z(n25279) );
  XOR U25186 ( .A(n25278), .B(n25219), .Z(n25221) );
  XOR U25187 ( .A(n25280), .B(n25281), .Z(n25267) );
  AND U25188 ( .A(n25282), .B(n25283), .Z(n25281) );
  XNOR U25189 ( .A(n25280), .B(n25229), .Z(n25283) );
  XOR U25190 ( .A(n25284), .B(n25276), .Z(n25229) );
  XNOR U25191 ( .A(n25285), .B(n25271), .Z(n25276) );
  XOR U25192 ( .A(n25286), .B(n25287), .Z(n25271) );
  AND U25193 ( .A(n25288), .B(n25289), .Z(n25287) );
  XOR U25194 ( .A(n25290), .B(n25286), .Z(n25288) );
  XNOR U25195 ( .A(n25291), .B(n25292), .Z(n25285) );
  AND U25196 ( .A(n25293), .B(n25294), .Z(n25292) );
  XOR U25197 ( .A(n25291), .B(n25295), .Z(n25293) );
  XNOR U25198 ( .A(n25277), .B(n25274), .Z(n25284) );
  AND U25199 ( .A(n25296), .B(n25297), .Z(n25274) );
  XOR U25200 ( .A(n25298), .B(n25299), .Z(n25277) );
  AND U25201 ( .A(n25300), .B(n25301), .Z(n25299) );
  XOR U25202 ( .A(n25298), .B(n25302), .Z(n25300) );
  XNOR U25203 ( .A(n25226), .B(n25280), .Z(n25282) );
  XNOR U25204 ( .A(n25303), .B(n25304), .Z(n25226) );
  AND U25205 ( .A(n419), .B(n25232), .Z(n25304) );
  XOR U25206 ( .A(n25303), .B(n25230), .Z(n25232) );
  XOR U25207 ( .A(n25305), .B(n25306), .Z(n25280) );
  AND U25208 ( .A(n25307), .B(n25308), .Z(n25306) );
  XNOR U25209 ( .A(n25305), .B(n25296), .Z(n25308) );
  IV U25210 ( .A(n25238), .Z(n25296) );
  XNOR U25211 ( .A(n25309), .B(n25289), .Z(n25238) );
  XNOR U25212 ( .A(n25310), .B(n25295), .Z(n25289) );
  XOR U25213 ( .A(n25311), .B(n25312), .Z(n25295) );
  AND U25214 ( .A(n25313), .B(n25314), .Z(n25312) );
  XOR U25215 ( .A(n25311), .B(n25315), .Z(n25313) );
  XNOR U25216 ( .A(n25294), .B(n25286), .Z(n25310) );
  XOR U25217 ( .A(n25316), .B(n25317), .Z(n25286) );
  AND U25218 ( .A(n25318), .B(n25319), .Z(n25317) );
  XNOR U25219 ( .A(n25320), .B(n25316), .Z(n25318) );
  XNOR U25220 ( .A(n25321), .B(n25291), .Z(n25294) );
  XOR U25221 ( .A(n25322), .B(n25323), .Z(n25291) );
  AND U25222 ( .A(n25324), .B(n25325), .Z(n25323) );
  XOR U25223 ( .A(n25322), .B(n25326), .Z(n25324) );
  XNOR U25224 ( .A(n25327), .B(n25328), .Z(n25321) );
  AND U25225 ( .A(n25329), .B(n25330), .Z(n25328) );
  XNOR U25226 ( .A(n25327), .B(n25331), .Z(n25329) );
  XNOR U25227 ( .A(n25290), .B(n25297), .Z(n25309) );
  AND U25228 ( .A(n25250), .B(n25332), .Z(n25297) );
  XOR U25229 ( .A(n25302), .B(n25301), .Z(n25290) );
  XNOR U25230 ( .A(n25333), .B(n25298), .Z(n25301) );
  XOR U25231 ( .A(n25334), .B(n25335), .Z(n25298) );
  AND U25232 ( .A(n25336), .B(n25337), .Z(n25335) );
  XOR U25233 ( .A(n25334), .B(n25338), .Z(n25336) );
  XNOR U25234 ( .A(n25339), .B(n25340), .Z(n25333) );
  AND U25235 ( .A(n25341), .B(n25342), .Z(n25340) );
  XOR U25236 ( .A(n25339), .B(n25343), .Z(n25341) );
  XOR U25237 ( .A(n25344), .B(n25345), .Z(n25302) );
  AND U25238 ( .A(n25346), .B(n25347), .Z(n25345) );
  XOR U25239 ( .A(n25344), .B(n25348), .Z(n25346) );
  XNOR U25240 ( .A(n25235), .B(n25305), .Z(n25307) );
  XNOR U25241 ( .A(n25349), .B(n25350), .Z(n25235) );
  AND U25242 ( .A(n419), .B(n25242), .Z(n25350) );
  XOR U25243 ( .A(n25349), .B(n25240), .Z(n25242) );
  XOR U25244 ( .A(n25351), .B(n25352), .Z(n25305) );
  AND U25245 ( .A(n25353), .B(n25354), .Z(n25352) );
  XNOR U25246 ( .A(n25351), .B(n25250), .Z(n25354) );
  XOR U25247 ( .A(n25355), .B(n25319), .Z(n25250) );
  XNOR U25248 ( .A(n25356), .B(n25326), .Z(n25319) );
  XOR U25249 ( .A(n25315), .B(n25314), .Z(n25326) );
  XNOR U25250 ( .A(n25357), .B(n25311), .Z(n25314) );
  XOR U25251 ( .A(n25358), .B(n25359), .Z(n25311) );
  AND U25252 ( .A(n25360), .B(n25361), .Z(n25359) );
  XNOR U25253 ( .A(n25362), .B(n25363), .Z(n25360) );
  IV U25254 ( .A(n25358), .Z(n25362) );
  XNOR U25255 ( .A(n25364), .B(n25365), .Z(n25357) );
  NOR U25256 ( .A(n25366), .B(n25367), .Z(n25365) );
  XNOR U25257 ( .A(n25364), .B(n25368), .Z(n25366) );
  XOR U25258 ( .A(n25369), .B(n25370), .Z(n25315) );
  NOR U25259 ( .A(n25371), .B(n25372), .Z(n25370) );
  XNOR U25260 ( .A(n25369), .B(n25373), .Z(n25371) );
  XNOR U25261 ( .A(n25325), .B(n25316), .Z(n25356) );
  XOR U25262 ( .A(n25374), .B(n25375), .Z(n25316) );
  AND U25263 ( .A(n25376), .B(n25377), .Z(n25375) );
  XOR U25264 ( .A(n25374), .B(n25378), .Z(n25376) );
  XOR U25265 ( .A(n25379), .B(n25331), .Z(n25325) );
  XOR U25266 ( .A(n25380), .B(n25381), .Z(n25331) );
  NOR U25267 ( .A(n25382), .B(n25383), .Z(n25381) );
  XOR U25268 ( .A(n25380), .B(n25384), .Z(n25382) );
  XNOR U25269 ( .A(n25330), .B(n25322), .Z(n25379) );
  XOR U25270 ( .A(n25385), .B(n25386), .Z(n25322) );
  AND U25271 ( .A(n25387), .B(n25388), .Z(n25386) );
  XOR U25272 ( .A(n25385), .B(n25389), .Z(n25387) );
  XNOR U25273 ( .A(n25390), .B(n25327), .Z(n25330) );
  XOR U25274 ( .A(n25391), .B(n25392), .Z(n25327) );
  AND U25275 ( .A(n25393), .B(n25394), .Z(n25392) );
  XNOR U25276 ( .A(n25395), .B(n25396), .Z(n25393) );
  IV U25277 ( .A(n25391), .Z(n25395) );
  XNOR U25278 ( .A(n25397), .B(n25398), .Z(n25390) );
  NOR U25279 ( .A(n25399), .B(n25400), .Z(n25398) );
  XNOR U25280 ( .A(n25397), .B(n25401), .Z(n25399) );
  XOR U25281 ( .A(n25320), .B(n25332), .Z(n25355) );
  NOR U25282 ( .A(n25258), .B(n25402), .Z(n25332) );
  XNOR U25283 ( .A(n25338), .B(n25337), .Z(n25320) );
  XNOR U25284 ( .A(n25403), .B(n25343), .Z(n25337) );
  XNOR U25285 ( .A(n25404), .B(n25405), .Z(n25343) );
  NOR U25286 ( .A(n25406), .B(n25407), .Z(n25405) );
  XOR U25287 ( .A(n25404), .B(n25408), .Z(n25406) );
  XNOR U25288 ( .A(n25342), .B(n25334), .Z(n25403) );
  XOR U25289 ( .A(n25409), .B(n25410), .Z(n25334) );
  AND U25290 ( .A(n25411), .B(n25412), .Z(n25410) );
  XOR U25291 ( .A(n25409), .B(n25413), .Z(n25411) );
  XNOR U25292 ( .A(n25414), .B(n25339), .Z(n25342) );
  XOR U25293 ( .A(n25415), .B(n25416), .Z(n25339) );
  AND U25294 ( .A(n25417), .B(n25418), .Z(n25416) );
  XNOR U25295 ( .A(n25419), .B(n25420), .Z(n25417) );
  IV U25296 ( .A(n25415), .Z(n25419) );
  XNOR U25297 ( .A(n25421), .B(n25422), .Z(n25414) );
  NOR U25298 ( .A(n25423), .B(n25424), .Z(n25422) );
  XNOR U25299 ( .A(n25421), .B(n25425), .Z(n25423) );
  XOR U25300 ( .A(n25348), .B(n25347), .Z(n25338) );
  XNOR U25301 ( .A(n25426), .B(n25344), .Z(n25347) );
  XOR U25302 ( .A(n25427), .B(n25428), .Z(n25344) );
  AND U25303 ( .A(n25429), .B(n25430), .Z(n25428) );
  XNOR U25304 ( .A(n25431), .B(n25432), .Z(n25429) );
  IV U25305 ( .A(n25427), .Z(n25431) );
  XNOR U25306 ( .A(n25433), .B(n25434), .Z(n25426) );
  NOR U25307 ( .A(n25435), .B(n25436), .Z(n25434) );
  XNOR U25308 ( .A(n25433), .B(n25437), .Z(n25435) );
  XOR U25309 ( .A(n25438), .B(n25439), .Z(n25348) );
  NOR U25310 ( .A(n25440), .B(n25441), .Z(n25439) );
  XNOR U25311 ( .A(n25438), .B(n25442), .Z(n25440) );
  XNOR U25312 ( .A(n25247), .B(n25351), .Z(n25353) );
  XNOR U25313 ( .A(n25443), .B(n25444), .Z(n25247) );
  AND U25314 ( .A(n419), .B(n25254), .Z(n25444) );
  XOR U25315 ( .A(n25443), .B(n25252), .Z(n25254) );
  AND U25316 ( .A(n25255), .B(n25258), .Z(n25351) );
  XOR U25317 ( .A(n25445), .B(n25402), .Z(n25258) );
  XNOR U25318 ( .A(p_input[1024]), .B(p_input[2048]), .Z(n25402) );
  XNOR U25319 ( .A(n25378), .B(n25377), .Z(n25445) );
  XNOR U25320 ( .A(n25446), .B(n25389), .Z(n25377) );
  XOR U25321 ( .A(n25363), .B(n25361), .Z(n25389) );
  XNOR U25322 ( .A(n25447), .B(n25368), .Z(n25361) );
  XOR U25323 ( .A(p_input[1048]), .B(p_input[2072]), .Z(n25368) );
  XOR U25324 ( .A(n25358), .B(n25367), .Z(n25447) );
  XOR U25325 ( .A(n25448), .B(n25364), .Z(n25367) );
  XOR U25326 ( .A(p_input[1046]), .B(p_input[2070]), .Z(n25364) );
  XOR U25327 ( .A(p_input[1047]), .B(n17295), .Z(n25448) );
  XOR U25328 ( .A(p_input[1042]), .B(p_input[2066]), .Z(n25358) );
  XNOR U25329 ( .A(n25373), .B(n25372), .Z(n25363) );
  XOR U25330 ( .A(n25449), .B(n25369), .Z(n25372) );
  XOR U25331 ( .A(p_input[1043]), .B(p_input[2067]), .Z(n25369) );
  XOR U25332 ( .A(p_input[1044]), .B(n17297), .Z(n25449) );
  XOR U25333 ( .A(p_input[1045]), .B(p_input[2069]), .Z(n25373) );
  XOR U25334 ( .A(n25388), .B(n25450), .Z(n25446) );
  IV U25335 ( .A(n25374), .Z(n25450) );
  XOR U25336 ( .A(p_input[1025]), .B(p_input[2049]), .Z(n25374) );
  XNOR U25337 ( .A(n25451), .B(n25396), .Z(n25388) );
  XNOR U25338 ( .A(n25384), .B(n25383), .Z(n25396) );
  XNOR U25339 ( .A(n25452), .B(n25380), .Z(n25383) );
  XNOR U25340 ( .A(p_input[1050]), .B(p_input[2074]), .Z(n25380) );
  XOR U25341 ( .A(p_input[1051]), .B(n17300), .Z(n25452) );
  XOR U25342 ( .A(p_input[1052]), .B(p_input[2076]), .Z(n25384) );
  XOR U25343 ( .A(n25394), .B(n25453), .Z(n25451) );
  IV U25344 ( .A(n25385), .Z(n25453) );
  XOR U25345 ( .A(p_input[1041]), .B(p_input[2065]), .Z(n25385) );
  XNOR U25346 ( .A(n25454), .B(n25401), .Z(n25394) );
  XNOR U25347 ( .A(p_input[1055]), .B(n17303), .Z(n25401) );
  XOR U25348 ( .A(n25391), .B(n25400), .Z(n25454) );
  XOR U25349 ( .A(n25455), .B(n25397), .Z(n25400) );
  XOR U25350 ( .A(p_input[1053]), .B(p_input[2077]), .Z(n25397) );
  XOR U25351 ( .A(p_input[1054]), .B(n17305), .Z(n25455) );
  XOR U25352 ( .A(p_input[1049]), .B(p_input[2073]), .Z(n25391) );
  XOR U25353 ( .A(n25413), .B(n25412), .Z(n25378) );
  XNOR U25354 ( .A(n25456), .B(n25420), .Z(n25412) );
  XNOR U25355 ( .A(n25408), .B(n25407), .Z(n25420) );
  XNOR U25356 ( .A(n25457), .B(n25404), .Z(n25407) );
  XNOR U25357 ( .A(p_input[1035]), .B(p_input[2059]), .Z(n25404) );
  XOR U25358 ( .A(p_input[1036]), .B(n16451), .Z(n25457) );
  XOR U25359 ( .A(p_input[1037]), .B(p_input[2061]), .Z(n25408) );
  XOR U25360 ( .A(n25418), .B(n25458), .Z(n25456) );
  IV U25361 ( .A(n25409), .Z(n25458) );
  XOR U25362 ( .A(p_input[1026]), .B(p_input[2050]), .Z(n25409) );
  XNOR U25363 ( .A(n25459), .B(n25425), .Z(n25418) );
  XNOR U25364 ( .A(p_input[1040]), .B(n16454), .Z(n25425) );
  XOR U25365 ( .A(n25415), .B(n25424), .Z(n25459) );
  XOR U25366 ( .A(n25460), .B(n25421), .Z(n25424) );
  XOR U25367 ( .A(p_input[1038]), .B(p_input[2062]), .Z(n25421) );
  XOR U25368 ( .A(p_input[1039]), .B(n16456), .Z(n25460) );
  XOR U25369 ( .A(p_input[1034]), .B(p_input[2058]), .Z(n25415) );
  XOR U25370 ( .A(n25432), .B(n25430), .Z(n25413) );
  XNOR U25371 ( .A(n25461), .B(n25437), .Z(n25430) );
  XOR U25372 ( .A(p_input[1033]), .B(p_input[2057]), .Z(n25437) );
  XOR U25373 ( .A(n25427), .B(n25436), .Z(n25461) );
  XOR U25374 ( .A(n25462), .B(n25433), .Z(n25436) );
  XOR U25375 ( .A(p_input[1031]), .B(p_input[2055]), .Z(n25433) );
  XOR U25376 ( .A(p_input[1032]), .B(n17312), .Z(n25462) );
  XOR U25377 ( .A(p_input[1027]), .B(p_input[2051]), .Z(n25427) );
  XNOR U25378 ( .A(n25442), .B(n25441), .Z(n25432) );
  XOR U25379 ( .A(n25463), .B(n25438), .Z(n25441) );
  XOR U25380 ( .A(p_input[1028]), .B(p_input[2052]), .Z(n25438) );
  XOR U25381 ( .A(p_input[1029]), .B(n17314), .Z(n25463) );
  XOR U25382 ( .A(p_input[1030]), .B(p_input[2054]), .Z(n25442) );
  XNOR U25383 ( .A(n25464), .B(n25465), .Z(n25255) );
  AND U25384 ( .A(n419), .B(n25466), .Z(n25465) );
  XNOR U25385 ( .A(n25467), .B(n25468), .Z(n419) );
  AND U25386 ( .A(n25469), .B(n25470), .Z(n25468) );
  XOR U25387 ( .A(n25467), .B(n25265), .Z(n25470) );
  XNOR U25388 ( .A(n25467), .B(n25207), .Z(n25469) );
  XOR U25389 ( .A(n25471), .B(n25472), .Z(n25467) );
  AND U25390 ( .A(n25473), .B(n25474), .Z(n25472) );
  XNOR U25391 ( .A(n25278), .B(n25471), .Z(n25474) );
  XOR U25392 ( .A(n25471), .B(n25219), .Z(n25473) );
  XOR U25393 ( .A(n25475), .B(n25476), .Z(n25471) );
  AND U25394 ( .A(n25477), .B(n25478), .Z(n25476) );
  XNOR U25395 ( .A(n25303), .B(n25475), .Z(n25478) );
  XOR U25396 ( .A(n25475), .B(n25230), .Z(n25477) );
  XOR U25397 ( .A(n25479), .B(n25480), .Z(n25475) );
  AND U25398 ( .A(n25481), .B(n25482), .Z(n25480) );
  XOR U25399 ( .A(n25479), .B(n25240), .Z(n25481) );
  XOR U25400 ( .A(n25483), .B(n25484), .Z(n25196) );
  AND U25401 ( .A(n423), .B(n25466), .Z(n25484) );
  XNOR U25402 ( .A(n25464), .B(n25483), .Z(n25466) );
  XNOR U25403 ( .A(n25485), .B(n25486), .Z(n423) );
  AND U25404 ( .A(n25487), .B(n25488), .Z(n25486) );
  XNOR U25405 ( .A(n25489), .B(n25485), .Z(n25488) );
  IV U25406 ( .A(n25265), .Z(n25489) );
  XNOR U25407 ( .A(n25490), .B(n25491), .Z(n25265) );
  AND U25408 ( .A(n426), .B(n25492), .Z(n25491) );
  XNOR U25409 ( .A(n25490), .B(n25493), .Z(n25492) );
  XNOR U25410 ( .A(n25207), .B(n25485), .Z(n25487) );
  XOR U25411 ( .A(n25494), .B(n25495), .Z(n25207) );
  AND U25412 ( .A(n434), .B(n25496), .Z(n25495) );
  XOR U25413 ( .A(n25497), .B(n25498), .Z(n25485) );
  AND U25414 ( .A(n25499), .B(n25500), .Z(n25498) );
  XNOR U25415 ( .A(n25497), .B(n25278), .Z(n25500) );
  XNOR U25416 ( .A(n25501), .B(n25502), .Z(n25278) );
  AND U25417 ( .A(n426), .B(n25503), .Z(n25502) );
  XOR U25418 ( .A(n25504), .B(n25501), .Z(n25503) );
  XNOR U25419 ( .A(n25505), .B(n25497), .Z(n25499) );
  IV U25420 ( .A(n25219), .Z(n25505) );
  XOR U25421 ( .A(n25506), .B(n25507), .Z(n25219) );
  AND U25422 ( .A(n434), .B(n25508), .Z(n25507) );
  XOR U25423 ( .A(n25509), .B(n25510), .Z(n25497) );
  AND U25424 ( .A(n25511), .B(n25512), .Z(n25510) );
  XNOR U25425 ( .A(n25509), .B(n25303), .Z(n25512) );
  XNOR U25426 ( .A(n25513), .B(n25514), .Z(n25303) );
  AND U25427 ( .A(n426), .B(n25515), .Z(n25514) );
  XNOR U25428 ( .A(n25516), .B(n25513), .Z(n25515) );
  XOR U25429 ( .A(n25230), .B(n25509), .Z(n25511) );
  XOR U25430 ( .A(n25517), .B(n25518), .Z(n25230) );
  AND U25431 ( .A(n434), .B(n25519), .Z(n25518) );
  XOR U25432 ( .A(n25479), .B(n25520), .Z(n25509) );
  AND U25433 ( .A(n25521), .B(n25482), .Z(n25520) );
  XNOR U25434 ( .A(n25349), .B(n25479), .Z(n25482) );
  XNOR U25435 ( .A(n25522), .B(n25523), .Z(n25349) );
  AND U25436 ( .A(n426), .B(n25524), .Z(n25523) );
  XOR U25437 ( .A(n25525), .B(n25522), .Z(n25524) );
  XNOR U25438 ( .A(n25526), .B(n25479), .Z(n25521) );
  IV U25439 ( .A(n25240), .Z(n25526) );
  XOR U25440 ( .A(n25527), .B(n25528), .Z(n25240) );
  AND U25441 ( .A(n434), .B(n25529), .Z(n25528) );
  XOR U25442 ( .A(n25530), .B(n25531), .Z(n25479) );
  AND U25443 ( .A(n25532), .B(n25533), .Z(n25531) );
  XNOR U25444 ( .A(n25530), .B(n25443), .Z(n25533) );
  XNOR U25445 ( .A(n25534), .B(n25535), .Z(n25443) );
  AND U25446 ( .A(n426), .B(n25536), .Z(n25535) );
  XNOR U25447 ( .A(n25537), .B(n25534), .Z(n25536) );
  XNOR U25448 ( .A(n25538), .B(n25530), .Z(n25532) );
  IV U25449 ( .A(n25252), .Z(n25538) );
  XOR U25450 ( .A(n25539), .B(n25540), .Z(n25252) );
  AND U25451 ( .A(n434), .B(n25541), .Z(n25540) );
  AND U25452 ( .A(n25483), .B(n25464), .Z(n25530) );
  XNOR U25453 ( .A(n25542), .B(n25543), .Z(n25464) );
  AND U25454 ( .A(n426), .B(n25544), .Z(n25543) );
  XNOR U25455 ( .A(n25545), .B(n25542), .Z(n25544) );
  XNOR U25456 ( .A(n25546), .B(n25547), .Z(n426) );
  AND U25457 ( .A(n25548), .B(n25549), .Z(n25547) );
  XOR U25458 ( .A(n25493), .B(n25546), .Z(n25549) );
  AND U25459 ( .A(n25550), .B(n25551), .Z(n25493) );
  XOR U25460 ( .A(n25546), .B(n25490), .Z(n25548) );
  XNOR U25461 ( .A(n25552), .B(n25553), .Z(n25490) );
  AND U25462 ( .A(n430), .B(n25496), .Z(n25553) );
  XOR U25463 ( .A(n25494), .B(n25552), .Z(n25496) );
  XOR U25464 ( .A(n25554), .B(n25555), .Z(n25546) );
  AND U25465 ( .A(n25556), .B(n25557), .Z(n25555) );
  XNOR U25466 ( .A(n25554), .B(n25550), .Z(n25557) );
  IV U25467 ( .A(n25504), .Z(n25550) );
  XOR U25468 ( .A(n25558), .B(n25559), .Z(n25504) );
  XOR U25469 ( .A(n25560), .B(n25551), .Z(n25559) );
  AND U25470 ( .A(n25516), .B(n25561), .Z(n25551) );
  AND U25471 ( .A(n25562), .B(n25563), .Z(n25560) );
  XOR U25472 ( .A(n25564), .B(n25558), .Z(n25562) );
  XNOR U25473 ( .A(n25501), .B(n25554), .Z(n25556) );
  XNOR U25474 ( .A(n25565), .B(n25566), .Z(n25501) );
  AND U25475 ( .A(n430), .B(n25508), .Z(n25566) );
  XOR U25476 ( .A(n25565), .B(n25506), .Z(n25508) );
  XOR U25477 ( .A(n25567), .B(n25568), .Z(n25554) );
  AND U25478 ( .A(n25569), .B(n25570), .Z(n25568) );
  XNOR U25479 ( .A(n25567), .B(n25516), .Z(n25570) );
  XOR U25480 ( .A(n25571), .B(n25563), .Z(n25516) );
  XNOR U25481 ( .A(n25572), .B(n25558), .Z(n25563) );
  XOR U25482 ( .A(n25573), .B(n25574), .Z(n25558) );
  AND U25483 ( .A(n25575), .B(n25576), .Z(n25574) );
  XOR U25484 ( .A(n25577), .B(n25573), .Z(n25575) );
  XNOR U25485 ( .A(n25578), .B(n25579), .Z(n25572) );
  AND U25486 ( .A(n25580), .B(n25581), .Z(n25579) );
  XOR U25487 ( .A(n25578), .B(n25582), .Z(n25580) );
  XNOR U25488 ( .A(n25564), .B(n25561), .Z(n25571) );
  AND U25489 ( .A(n25583), .B(n25584), .Z(n25561) );
  XOR U25490 ( .A(n25585), .B(n25586), .Z(n25564) );
  AND U25491 ( .A(n25587), .B(n25588), .Z(n25586) );
  XOR U25492 ( .A(n25585), .B(n25589), .Z(n25587) );
  XNOR U25493 ( .A(n25513), .B(n25567), .Z(n25569) );
  XNOR U25494 ( .A(n25590), .B(n25591), .Z(n25513) );
  AND U25495 ( .A(n430), .B(n25519), .Z(n25591) );
  XOR U25496 ( .A(n25590), .B(n25517), .Z(n25519) );
  XOR U25497 ( .A(n25592), .B(n25593), .Z(n25567) );
  AND U25498 ( .A(n25594), .B(n25595), .Z(n25593) );
  XNOR U25499 ( .A(n25592), .B(n25583), .Z(n25595) );
  IV U25500 ( .A(n25525), .Z(n25583) );
  XNOR U25501 ( .A(n25596), .B(n25576), .Z(n25525) );
  XNOR U25502 ( .A(n25597), .B(n25582), .Z(n25576) );
  XOR U25503 ( .A(n25598), .B(n25599), .Z(n25582) );
  AND U25504 ( .A(n25600), .B(n25601), .Z(n25599) );
  XOR U25505 ( .A(n25598), .B(n25602), .Z(n25600) );
  XNOR U25506 ( .A(n25581), .B(n25573), .Z(n25597) );
  XOR U25507 ( .A(n25603), .B(n25604), .Z(n25573) );
  AND U25508 ( .A(n25605), .B(n25606), .Z(n25604) );
  XNOR U25509 ( .A(n25607), .B(n25603), .Z(n25605) );
  XNOR U25510 ( .A(n25608), .B(n25578), .Z(n25581) );
  XOR U25511 ( .A(n25609), .B(n25610), .Z(n25578) );
  AND U25512 ( .A(n25611), .B(n25612), .Z(n25610) );
  XOR U25513 ( .A(n25609), .B(n25613), .Z(n25611) );
  XNOR U25514 ( .A(n25614), .B(n25615), .Z(n25608) );
  AND U25515 ( .A(n25616), .B(n25617), .Z(n25615) );
  XNOR U25516 ( .A(n25614), .B(n25618), .Z(n25616) );
  XNOR U25517 ( .A(n25577), .B(n25584), .Z(n25596) );
  AND U25518 ( .A(n25537), .B(n25619), .Z(n25584) );
  XOR U25519 ( .A(n25589), .B(n25588), .Z(n25577) );
  XNOR U25520 ( .A(n25620), .B(n25585), .Z(n25588) );
  XOR U25521 ( .A(n25621), .B(n25622), .Z(n25585) );
  AND U25522 ( .A(n25623), .B(n25624), .Z(n25622) );
  XOR U25523 ( .A(n25621), .B(n25625), .Z(n25623) );
  XNOR U25524 ( .A(n25626), .B(n25627), .Z(n25620) );
  AND U25525 ( .A(n25628), .B(n25629), .Z(n25627) );
  XOR U25526 ( .A(n25626), .B(n25630), .Z(n25628) );
  XOR U25527 ( .A(n25631), .B(n25632), .Z(n25589) );
  AND U25528 ( .A(n25633), .B(n25634), .Z(n25632) );
  XOR U25529 ( .A(n25631), .B(n25635), .Z(n25633) );
  XNOR U25530 ( .A(n25522), .B(n25592), .Z(n25594) );
  XNOR U25531 ( .A(n25636), .B(n25637), .Z(n25522) );
  AND U25532 ( .A(n430), .B(n25529), .Z(n25637) );
  XOR U25533 ( .A(n25636), .B(n25527), .Z(n25529) );
  XOR U25534 ( .A(n25638), .B(n25639), .Z(n25592) );
  AND U25535 ( .A(n25640), .B(n25641), .Z(n25639) );
  XNOR U25536 ( .A(n25638), .B(n25537), .Z(n25641) );
  XOR U25537 ( .A(n25642), .B(n25606), .Z(n25537) );
  XNOR U25538 ( .A(n25643), .B(n25613), .Z(n25606) );
  XOR U25539 ( .A(n25602), .B(n25601), .Z(n25613) );
  XNOR U25540 ( .A(n25644), .B(n25598), .Z(n25601) );
  XOR U25541 ( .A(n25645), .B(n25646), .Z(n25598) );
  AND U25542 ( .A(n25647), .B(n25648), .Z(n25646) );
  XNOR U25543 ( .A(n25649), .B(n25650), .Z(n25647) );
  IV U25544 ( .A(n25645), .Z(n25649) );
  XNOR U25545 ( .A(n25651), .B(n25652), .Z(n25644) );
  NOR U25546 ( .A(n25653), .B(n25654), .Z(n25652) );
  XNOR U25547 ( .A(n25651), .B(n25655), .Z(n25653) );
  XOR U25548 ( .A(n25656), .B(n25657), .Z(n25602) );
  NOR U25549 ( .A(n25658), .B(n25659), .Z(n25657) );
  XNOR U25550 ( .A(n25656), .B(n25660), .Z(n25658) );
  XNOR U25551 ( .A(n25612), .B(n25603), .Z(n25643) );
  XOR U25552 ( .A(n25661), .B(n25662), .Z(n25603) );
  AND U25553 ( .A(n25663), .B(n25664), .Z(n25662) );
  XOR U25554 ( .A(n25661), .B(n25665), .Z(n25663) );
  XOR U25555 ( .A(n25666), .B(n25618), .Z(n25612) );
  XOR U25556 ( .A(n25667), .B(n25668), .Z(n25618) );
  NOR U25557 ( .A(n25669), .B(n25670), .Z(n25668) );
  XOR U25558 ( .A(n25667), .B(n25671), .Z(n25669) );
  XNOR U25559 ( .A(n25617), .B(n25609), .Z(n25666) );
  XOR U25560 ( .A(n25672), .B(n25673), .Z(n25609) );
  AND U25561 ( .A(n25674), .B(n25675), .Z(n25673) );
  XOR U25562 ( .A(n25672), .B(n25676), .Z(n25674) );
  XNOR U25563 ( .A(n25677), .B(n25614), .Z(n25617) );
  XOR U25564 ( .A(n25678), .B(n25679), .Z(n25614) );
  AND U25565 ( .A(n25680), .B(n25681), .Z(n25679) );
  XNOR U25566 ( .A(n25682), .B(n25683), .Z(n25680) );
  IV U25567 ( .A(n25678), .Z(n25682) );
  XNOR U25568 ( .A(n25684), .B(n25685), .Z(n25677) );
  NOR U25569 ( .A(n25686), .B(n25687), .Z(n25685) );
  XNOR U25570 ( .A(n25684), .B(n25688), .Z(n25686) );
  XOR U25571 ( .A(n25607), .B(n25619), .Z(n25642) );
  NOR U25572 ( .A(n25545), .B(n25689), .Z(n25619) );
  XNOR U25573 ( .A(n25625), .B(n25624), .Z(n25607) );
  XNOR U25574 ( .A(n25690), .B(n25630), .Z(n25624) );
  XNOR U25575 ( .A(n25691), .B(n25692), .Z(n25630) );
  NOR U25576 ( .A(n25693), .B(n25694), .Z(n25692) );
  XOR U25577 ( .A(n25691), .B(n25695), .Z(n25693) );
  XNOR U25578 ( .A(n25629), .B(n25621), .Z(n25690) );
  XOR U25579 ( .A(n25696), .B(n25697), .Z(n25621) );
  AND U25580 ( .A(n25698), .B(n25699), .Z(n25697) );
  XOR U25581 ( .A(n25696), .B(n25700), .Z(n25698) );
  XNOR U25582 ( .A(n25701), .B(n25626), .Z(n25629) );
  XOR U25583 ( .A(n25702), .B(n25703), .Z(n25626) );
  AND U25584 ( .A(n25704), .B(n25705), .Z(n25703) );
  XNOR U25585 ( .A(n25706), .B(n25707), .Z(n25704) );
  IV U25586 ( .A(n25702), .Z(n25706) );
  XNOR U25587 ( .A(n25708), .B(n25709), .Z(n25701) );
  NOR U25588 ( .A(n25710), .B(n25711), .Z(n25709) );
  XNOR U25589 ( .A(n25708), .B(n25712), .Z(n25710) );
  XOR U25590 ( .A(n25635), .B(n25634), .Z(n25625) );
  XNOR U25591 ( .A(n25713), .B(n25631), .Z(n25634) );
  XOR U25592 ( .A(n25714), .B(n25715), .Z(n25631) );
  AND U25593 ( .A(n25716), .B(n25717), .Z(n25715) );
  XNOR U25594 ( .A(n25718), .B(n25719), .Z(n25716) );
  IV U25595 ( .A(n25714), .Z(n25718) );
  XNOR U25596 ( .A(n25720), .B(n25721), .Z(n25713) );
  NOR U25597 ( .A(n25722), .B(n25723), .Z(n25721) );
  XNOR U25598 ( .A(n25720), .B(n25724), .Z(n25722) );
  XOR U25599 ( .A(n25725), .B(n25726), .Z(n25635) );
  NOR U25600 ( .A(n25727), .B(n25728), .Z(n25726) );
  XNOR U25601 ( .A(n25725), .B(n25729), .Z(n25727) );
  XNOR U25602 ( .A(n25534), .B(n25638), .Z(n25640) );
  XNOR U25603 ( .A(n25730), .B(n25731), .Z(n25534) );
  AND U25604 ( .A(n430), .B(n25541), .Z(n25731) );
  XOR U25605 ( .A(n25730), .B(n25539), .Z(n25541) );
  AND U25606 ( .A(n25542), .B(n25545), .Z(n25638) );
  XOR U25607 ( .A(n25732), .B(n25689), .Z(n25545) );
  XNOR U25608 ( .A(p_input[1056]), .B(p_input[2048]), .Z(n25689) );
  XNOR U25609 ( .A(n25665), .B(n25664), .Z(n25732) );
  XNOR U25610 ( .A(n25733), .B(n25676), .Z(n25664) );
  XOR U25611 ( .A(n25650), .B(n25648), .Z(n25676) );
  XNOR U25612 ( .A(n25734), .B(n25655), .Z(n25648) );
  XOR U25613 ( .A(p_input[1080]), .B(p_input[2072]), .Z(n25655) );
  XOR U25614 ( .A(n25645), .B(n25654), .Z(n25734) );
  XOR U25615 ( .A(n25735), .B(n25651), .Z(n25654) );
  XOR U25616 ( .A(p_input[1078]), .B(p_input[2070]), .Z(n25651) );
  XOR U25617 ( .A(p_input[1079]), .B(n17295), .Z(n25735) );
  XOR U25618 ( .A(p_input[1074]), .B(p_input[2066]), .Z(n25645) );
  XNOR U25619 ( .A(n25660), .B(n25659), .Z(n25650) );
  XOR U25620 ( .A(n25736), .B(n25656), .Z(n25659) );
  XOR U25621 ( .A(p_input[1075]), .B(p_input[2067]), .Z(n25656) );
  XOR U25622 ( .A(p_input[1076]), .B(n17297), .Z(n25736) );
  XOR U25623 ( .A(p_input[1077]), .B(p_input[2069]), .Z(n25660) );
  XOR U25624 ( .A(n25675), .B(n25737), .Z(n25733) );
  IV U25625 ( .A(n25661), .Z(n25737) );
  XOR U25626 ( .A(p_input[1057]), .B(p_input[2049]), .Z(n25661) );
  XNOR U25627 ( .A(n25738), .B(n25683), .Z(n25675) );
  XNOR U25628 ( .A(n25671), .B(n25670), .Z(n25683) );
  XNOR U25629 ( .A(n25739), .B(n25667), .Z(n25670) );
  XNOR U25630 ( .A(p_input[1082]), .B(p_input[2074]), .Z(n25667) );
  XOR U25631 ( .A(p_input[1083]), .B(n17300), .Z(n25739) );
  XOR U25632 ( .A(p_input[1084]), .B(p_input[2076]), .Z(n25671) );
  XOR U25633 ( .A(n25681), .B(n25740), .Z(n25738) );
  IV U25634 ( .A(n25672), .Z(n25740) );
  XOR U25635 ( .A(p_input[1073]), .B(p_input[2065]), .Z(n25672) );
  XNOR U25636 ( .A(n25741), .B(n25688), .Z(n25681) );
  XNOR U25637 ( .A(p_input[1087]), .B(n17303), .Z(n25688) );
  XOR U25638 ( .A(n25678), .B(n25687), .Z(n25741) );
  XOR U25639 ( .A(n25742), .B(n25684), .Z(n25687) );
  XOR U25640 ( .A(p_input[1085]), .B(p_input[2077]), .Z(n25684) );
  XOR U25641 ( .A(p_input[1086]), .B(n17305), .Z(n25742) );
  XOR U25642 ( .A(p_input[1081]), .B(p_input[2073]), .Z(n25678) );
  XOR U25643 ( .A(n25700), .B(n25699), .Z(n25665) );
  XNOR U25644 ( .A(n25743), .B(n25707), .Z(n25699) );
  XNOR U25645 ( .A(n25695), .B(n25694), .Z(n25707) );
  XNOR U25646 ( .A(n25744), .B(n25691), .Z(n25694) );
  XNOR U25647 ( .A(p_input[1067]), .B(p_input[2059]), .Z(n25691) );
  XOR U25648 ( .A(p_input[1068]), .B(n16451), .Z(n25744) );
  XOR U25649 ( .A(p_input[1069]), .B(p_input[2061]), .Z(n25695) );
  XOR U25650 ( .A(n25705), .B(n25745), .Z(n25743) );
  IV U25651 ( .A(n25696), .Z(n25745) );
  XOR U25652 ( .A(p_input[1058]), .B(p_input[2050]), .Z(n25696) );
  XNOR U25653 ( .A(n25746), .B(n25712), .Z(n25705) );
  XNOR U25654 ( .A(p_input[1072]), .B(n16454), .Z(n25712) );
  XOR U25655 ( .A(n25702), .B(n25711), .Z(n25746) );
  XOR U25656 ( .A(n25747), .B(n25708), .Z(n25711) );
  XOR U25657 ( .A(p_input[1070]), .B(p_input[2062]), .Z(n25708) );
  XOR U25658 ( .A(p_input[1071]), .B(n16456), .Z(n25747) );
  XOR U25659 ( .A(p_input[1066]), .B(p_input[2058]), .Z(n25702) );
  XOR U25660 ( .A(n25719), .B(n25717), .Z(n25700) );
  XNOR U25661 ( .A(n25748), .B(n25724), .Z(n25717) );
  XOR U25662 ( .A(p_input[1065]), .B(p_input[2057]), .Z(n25724) );
  XOR U25663 ( .A(n25714), .B(n25723), .Z(n25748) );
  XOR U25664 ( .A(n25749), .B(n25720), .Z(n25723) );
  XOR U25665 ( .A(p_input[1063]), .B(p_input[2055]), .Z(n25720) );
  XOR U25666 ( .A(p_input[1064]), .B(n17312), .Z(n25749) );
  XOR U25667 ( .A(p_input[1059]), .B(p_input[2051]), .Z(n25714) );
  XNOR U25668 ( .A(n25729), .B(n25728), .Z(n25719) );
  XOR U25669 ( .A(n25750), .B(n25725), .Z(n25728) );
  XOR U25670 ( .A(p_input[1060]), .B(p_input[2052]), .Z(n25725) );
  XOR U25671 ( .A(p_input[1061]), .B(n17314), .Z(n25750) );
  XOR U25672 ( .A(p_input[1062]), .B(p_input[2054]), .Z(n25729) );
  XNOR U25673 ( .A(n25751), .B(n25752), .Z(n25542) );
  AND U25674 ( .A(n430), .B(n25753), .Z(n25752) );
  XNOR U25675 ( .A(n25754), .B(n25755), .Z(n430) );
  AND U25676 ( .A(n25756), .B(n25757), .Z(n25755) );
  XOR U25677 ( .A(n25754), .B(n25552), .Z(n25757) );
  XNOR U25678 ( .A(n25754), .B(n25494), .Z(n25756) );
  XOR U25679 ( .A(n25758), .B(n25759), .Z(n25754) );
  AND U25680 ( .A(n25760), .B(n25761), .Z(n25759) );
  XNOR U25681 ( .A(n25565), .B(n25758), .Z(n25761) );
  XOR U25682 ( .A(n25758), .B(n25506), .Z(n25760) );
  XOR U25683 ( .A(n25762), .B(n25763), .Z(n25758) );
  AND U25684 ( .A(n25764), .B(n25765), .Z(n25763) );
  XNOR U25685 ( .A(n25590), .B(n25762), .Z(n25765) );
  XOR U25686 ( .A(n25762), .B(n25517), .Z(n25764) );
  XOR U25687 ( .A(n25766), .B(n25767), .Z(n25762) );
  AND U25688 ( .A(n25768), .B(n25769), .Z(n25767) );
  XOR U25689 ( .A(n25766), .B(n25527), .Z(n25768) );
  XOR U25690 ( .A(n25770), .B(n25771), .Z(n25483) );
  AND U25691 ( .A(n434), .B(n25753), .Z(n25771) );
  XNOR U25692 ( .A(n25751), .B(n25770), .Z(n25753) );
  XNOR U25693 ( .A(n25772), .B(n25773), .Z(n434) );
  AND U25694 ( .A(n25774), .B(n25775), .Z(n25773) );
  XNOR U25695 ( .A(n25776), .B(n25772), .Z(n25775) );
  IV U25696 ( .A(n25552), .Z(n25776) );
  XNOR U25697 ( .A(n25777), .B(n25778), .Z(n25552) );
  AND U25698 ( .A(n437), .B(n25779), .Z(n25778) );
  XNOR U25699 ( .A(n25777), .B(n25780), .Z(n25779) );
  XNOR U25700 ( .A(n25494), .B(n25772), .Z(n25774) );
  XOR U25701 ( .A(n25781), .B(n25782), .Z(n25494) );
  AND U25702 ( .A(n445), .B(n25783), .Z(n25782) );
  XOR U25703 ( .A(n25784), .B(n25785), .Z(n25772) );
  AND U25704 ( .A(n25786), .B(n25787), .Z(n25785) );
  XNOR U25705 ( .A(n25784), .B(n25565), .Z(n25787) );
  XNOR U25706 ( .A(n25788), .B(n25789), .Z(n25565) );
  AND U25707 ( .A(n437), .B(n25790), .Z(n25789) );
  XOR U25708 ( .A(n25791), .B(n25788), .Z(n25790) );
  XNOR U25709 ( .A(n25792), .B(n25784), .Z(n25786) );
  IV U25710 ( .A(n25506), .Z(n25792) );
  XOR U25711 ( .A(n25793), .B(n25794), .Z(n25506) );
  AND U25712 ( .A(n445), .B(n25795), .Z(n25794) );
  XOR U25713 ( .A(n25796), .B(n25797), .Z(n25784) );
  AND U25714 ( .A(n25798), .B(n25799), .Z(n25797) );
  XNOR U25715 ( .A(n25796), .B(n25590), .Z(n25799) );
  XNOR U25716 ( .A(n25800), .B(n25801), .Z(n25590) );
  AND U25717 ( .A(n437), .B(n25802), .Z(n25801) );
  XNOR U25718 ( .A(n25803), .B(n25800), .Z(n25802) );
  XOR U25719 ( .A(n25517), .B(n25796), .Z(n25798) );
  XOR U25720 ( .A(n25804), .B(n25805), .Z(n25517) );
  AND U25721 ( .A(n445), .B(n25806), .Z(n25805) );
  XOR U25722 ( .A(n25766), .B(n25807), .Z(n25796) );
  AND U25723 ( .A(n25808), .B(n25769), .Z(n25807) );
  XNOR U25724 ( .A(n25636), .B(n25766), .Z(n25769) );
  XNOR U25725 ( .A(n25809), .B(n25810), .Z(n25636) );
  AND U25726 ( .A(n437), .B(n25811), .Z(n25810) );
  XOR U25727 ( .A(n25812), .B(n25809), .Z(n25811) );
  XNOR U25728 ( .A(n25813), .B(n25766), .Z(n25808) );
  IV U25729 ( .A(n25527), .Z(n25813) );
  XOR U25730 ( .A(n25814), .B(n25815), .Z(n25527) );
  AND U25731 ( .A(n445), .B(n25816), .Z(n25815) );
  XOR U25732 ( .A(n25817), .B(n25818), .Z(n25766) );
  AND U25733 ( .A(n25819), .B(n25820), .Z(n25818) );
  XNOR U25734 ( .A(n25817), .B(n25730), .Z(n25820) );
  XNOR U25735 ( .A(n25821), .B(n25822), .Z(n25730) );
  AND U25736 ( .A(n437), .B(n25823), .Z(n25822) );
  XNOR U25737 ( .A(n25824), .B(n25821), .Z(n25823) );
  XNOR U25738 ( .A(n25825), .B(n25817), .Z(n25819) );
  IV U25739 ( .A(n25539), .Z(n25825) );
  XOR U25740 ( .A(n25826), .B(n25827), .Z(n25539) );
  AND U25741 ( .A(n445), .B(n25828), .Z(n25827) );
  AND U25742 ( .A(n25770), .B(n25751), .Z(n25817) );
  XNOR U25743 ( .A(n25829), .B(n25830), .Z(n25751) );
  AND U25744 ( .A(n437), .B(n25831), .Z(n25830) );
  XNOR U25745 ( .A(n25832), .B(n25829), .Z(n25831) );
  XNOR U25746 ( .A(n25833), .B(n25834), .Z(n437) );
  AND U25747 ( .A(n25835), .B(n25836), .Z(n25834) );
  XOR U25748 ( .A(n25780), .B(n25833), .Z(n25836) );
  AND U25749 ( .A(n25837), .B(n25838), .Z(n25780) );
  XOR U25750 ( .A(n25833), .B(n25777), .Z(n25835) );
  XNOR U25751 ( .A(n25839), .B(n25840), .Z(n25777) );
  AND U25752 ( .A(n441), .B(n25783), .Z(n25840) );
  XOR U25753 ( .A(n25781), .B(n25839), .Z(n25783) );
  XOR U25754 ( .A(n25841), .B(n25842), .Z(n25833) );
  AND U25755 ( .A(n25843), .B(n25844), .Z(n25842) );
  XNOR U25756 ( .A(n25841), .B(n25837), .Z(n25844) );
  IV U25757 ( .A(n25791), .Z(n25837) );
  XOR U25758 ( .A(n25845), .B(n25846), .Z(n25791) );
  XOR U25759 ( .A(n25847), .B(n25838), .Z(n25846) );
  AND U25760 ( .A(n25803), .B(n25848), .Z(n25838) );
  AND U25761 ( .A(n25849), .B(n25850), .Z(n25847) );
  XOR U25762 ( .A(n25851), .B(n25845), .Z(n25849) );
  XNOR U25763 ( .A(n25788), .B(n25841), .Z(n25843) );
  XNOR U25764 ( .A(n25852), .B(n25853), .Z(n25788) );
  AND U25765 ( .A(n441), .B(n25795), .Z(n25853) );
  XOR U25766 ( .A(n25852), .B(n25793), .Z(n25795) );
  XOR U25767 ( .A(n25854), .B(n25855), .Z(n25841) );
  AND U25768 ( .A(n25856), .B(n25857), .Z(n25855) );
  XNOR U25769 ( .A(n25854), .B(n25803), .Z(n25857) );
  XOR U25770 ( .A(n25858), .B(n25850), .Z(n25803) );
  XNOR U25771 ( .A(n25859), .B(n25845), .Z(n25850) );
  XOR U25772 ( .A(n25860), .B(n25861), .Z(n25845) );
  AND U25773 ( .A(n25862), .B(n25863), .Z(n25861) );
  XOR U25774 ( .A(n25864), .B(n25860), .Z(n25862) );
  XNOR U25775 ( .A(n25865), .B(n25866), .Z(n25859) );
  AND U25776 ( .A(n25867), .B(n25868), .Z(n25866) );
  XOR U25777 ( .A(n25865), .B(n25869), .Z(n25867) );
  XNOR U25778 ( .A(n25851), .B(n25848), .Z(n25858) );
  AND U25779 ( .A(n25870), .B(n25871), .Z(n25848) );
  XOR U25780 ( .A(n25872), .B(n25873), .Z(n25851) );
  AND U25781 ( .A(n25874), .B(n25875), .Z(n25873) );
  XOR U25782 ( .A(n25872), .B(n25876), .Z(n25874) );
  XNOR U25783 ( .A(n25800), .B(n25854), .Z(n25856) );
  XNOR U25784 ( .A(n25877), .B(n25878), .Z(n25800) );
  AND U25785 ( .A(n441), .B(n25806), .Z(n25878) );
  XOR U25786 ( .A(n25877), .B(n25804), .Z(n25806) );
  XOR U25787 ( .A(n25879), .B(n25880), .Z(n25854) );
  AND U25788 ( .A(n25881), .B(n25882), .Z(n25880) );
  XNOR U25789 ( .A(n25879), .B(n25870), .Z(n25882) );
  IV U25790 ( .A(n25812), .Z(n25870) );
  XNOR U25791 ( .A(n25883), .B(n25863), .Z(n25812) );
  XNOR U25792 ( .A(n25884), .B(n25869), .Z(n25863) );
  XOR U25793 ( .A(n25885), .B(n25886), .Z(n25869) );
  AND U25794 ( .A(n25887), .B(n25888), .Z(n25886) );
  XOR U25795 ( .A(n25885), .B(n25889), .Z(n25887) );
  XNOR U25796 ( .A(n25868), .B(n25860), .Z(n25884) );
  XOR U25797 ( .A(n25890), .B(n25891), .Z(n25860) );
  AND U25798 ( .A(n25892), .B(n25893), .Z(n25891) );
  XNOR U25799 ( .A(n25894), .B(n25890), .Z(n25892) );
  XNOR U25800 ( .A(n25895), .B(n25865), .Z(n25868) );
  XOR U25801 ( .A(n25896), .B(n25897), .Z(n25865) );
  AND U25802 ( .A(n25898), .B(n25899), .Z(n25897) );
  XOR U25803 ( .A(n25896), .B(n25900), .Z(n25898) );
  XNOR U25804 ( .A(n25901), .B(n25902), .Z(n25895) );
  AND U25805 ( .A(n25903), .B(n25904), .Z(n25902) );
  XNOR U25806 ( .A(n25901), .B(n25905), .Z(n25903) );
  XNOR U25807 ( .A(n25864), .B(n25871), .Z(n25883) );
  AND U25808 ( .A(n25824), .B(n25906), .Z(n25871) );
  XOR U25809 ( .A(n25876), .B(n25875), .Z(n25864) );
  XNOR U25810 ( .A(n25907), .B(n25872), .Z(n25875) );
  XOR U25811 ( .A(n25908), .B(n25909), .Z(n25872) );
  AND U25812 ( .A(n25910), .B(n25911), .Z(n25909) );
  XOR U25813 ( .A(n25908), .B(n25912), .Z(n25910) );
  XNOR U25814 ( .A(n25913), .B(n25914), .Z(n25907) );
  AND U25815 ( .A(n25915), .B(n25916), .Z(n25914) );
  XOR U25816 ( .A(n25913), .B(n25917), .Z(n25915) );
  XOR U25817 ( .A(n25918), .B(n25919), .Z(n25876) );
  AND U25818 ( .A(n25920), .B(n25921), .Z(n25919) );
  XOR U25819 ( .A(n25918), .B(n25922), .Z(n25920) );
  XNOR U25820 ( .A(n25809), .B(n25879), .Z(n25881) );
  XNOR U25821 ( .A(n25923), .B(n25924), .Z(n25809) );
  AND U25822 ( .A(n441), .B(n25816), .Z(n25924) );
  XOR U25823 ( .A(n25923), .B(n25814), .Z(n25816) );
  XOR U25824 ( .A(n25925), .B(n25926), .Z(n25879) );
  AND U25825 ( .A(n25927), .B(n25928), .Z(n25926) );
  XNOR U25826 ( .A(n25925), .B(n25824), .Z(n25928) );
  XOR U25827 ( .A(n25929), .B(n25893), .Z(n25824) );
  XNOR U25828 ( .A(n25930), .B(n25900), .Z(n25893) );
  XOR U25829 ( .A(n25889), .B(n25888), .Z(n25900) );
  XNOR U25830 ( .A(n25931), .B(n25885), .Z(n25888) );
  XOR U25831 ( .A(n25932), .B(n25933), .Z(n25885) );
  AND U25832 ( .A(n25934), .B(n25935), .Z(n25933) );
  XNOR U25833 ( .A(n25936), .B(n25937), .Z(n25934) );
  IV U25834 ( .A(n25932), .Z(n25936) );
  XNOR U25835 ( .A(n25938), .B(n25939), .Z(n25931) );
  NOR U25836 ( .A(n25940), .B(n25941), .Z(n25939) );
  XNOR U25837 ( .A(n25938), .B(n25942), .Z(n25940) );
  XOR U25838 ( .A(n25943), .B(n25944), .Z(n25889) );
  NOR U25839 ( .A(n25945), .B(n25946), .Z(n25944) );
  XNOR U25840 ( .A(n25943), .B(n25947), .Z(n25945) );
  XNOR U25841 ( .A(n25899), .B(n25890), .Z(n25930) );
  XOR U25842 ( .A(n25948), .B(n25949), .Z(n25890) );
  AND U25843 ( .A(n25950), .B(n25951), .Z(n25949) );
  XOR U25844 ( .A(n25948), .B(n25952), .Z(n25950) );
  XOR U25845 ( .A(n25953), .B(n25905), .Z(n25899) );
  XOR U25846 ( .A(n25954), .B(n25955), .Z(n25905) );
  NOR U25847 ( .A(n25956), .B(n25957), .Z(n25955) );
  XOR U25848 ( .A(n25954), .B(n25958), .Z(n25956) );
  XNOR U25849 ( .A(n25904), .B(n25896), .Z(n25953) );
  XOR U25850 ( .A(n25959), .B(n25960), .Z(n25896) );
  AND U25851 ( .A(n25961), .B(n25962), .Z(n25960) );
  XOR U25852 ( .A(n25959), .B(n25963), .Z(n25961) );
  XNOR U25853 ( .A(n25964), .B(n25901), .Z(n25904) );
  XOR U25854 ( .A(n25965), .B(n25966), .Z(n25901) );
  AND U25855 ( .A(n25967), .B(n25968), .Z(n25966) );
  XNOR U25856 ( .A(n25969), .B(n25970), .Z(n25967) );
  IV U25857 ( .A(n25965), .Z(n25969) );
  XNOR U25858 ( .A(n25971), .B(n25972), .Z(n25964) );
  NOR U25859 ( .A(n25973), .B(n25974), .Z(n25972) );
  XNOR U25860 ( .A(n25971), .B(n25975), .Z(n25973) );
  XOR U25861 ( .A(n25894), .B(n25906), .Z(n25929) );
  NOR U25862 ( .A(n25832), .B(n25976), .Z(n25906) );
  XNOR U25863 ( .A(n25912), .B(n25911), .Z(n25894) );
  XNOR U25864 ( .A(n25977), .B(n25917), .Z(n25911) );
  XNOR U25865 ( .A(n25978), .B(n25979), .Z(n25917) );
  NOR U25866 ( .A(n25980), .B(n25981), .Z(n25979) );
  XOR U25867 ( .A(n25978), .B(n25982), .Z(n25980) );
  XNOR U25868 ( .A(n25916), .B(n25908), .Z(n25977) );
  XOR U25869 ( .A(n25983), .B(n25984), .Z(n25908) );
  AND U25870 ( .A(n25985), .B(n25986), .Z(n25984) );
  XOR U25871 ( .A(n25983), .B(n25987), .Z(n25985) );
  XNOR U25872 ( .A(n25988), .B(n25913), .Z(n25916) );
  XOR U25873 ( .A(n25989), .B(n25990), .Z(n25913) );
  AND U25874 ( .A(n25991), .B(n25992), .Z(n25990) );
  XNOR U25875 ( .A(n25993), .B(n25994), .Z(n25991) );
  IV U25876 ( .A(n25989), .Z(n25993) );
  XNOR U25877 ( .A(n25995), .B(n25996), .Z(n25988) );
  NOR U25878 ( .A(n25997), .B(n25998), .Z(n25996) );
  XNOR U25879 ( .A(n25995), .B(n25999), .Z(n25997) );
  XOR U25880 ( .A(n25922), .B(n25921), .Z(n25912) );
  XNOR U25881 ( .A(n26000), .B(n25918), .Z(n25921) );
  XOR U25882 ( .A(n26001), .B(n26002), .Z(n25918) );
  AND U25883 ( .A(n26003), .B(n26004), .Z(n26002) );
  XNOR U25884 ( .A(n26005), .B(n26006), .Z(n26003) );
  IV U25885 ( .A(n26001), .Z(n26005) );
  XNOR U25886 ( .A(n26007), .B(n26008), .Z(n26000) );
  NOR U25887 ( .A(n26009), .B(n26010), .Z(n26008) );
  XNOR U25888 ( .A(n26007), .B(n26011), .Z(n26009) );
  XOR U25889 ( .A(n26012), .B(n26013), .Z(n25922) );
  NOR U25890 ( .A(n26014), .B(n26015), .Z(n26013) );
  XNOR U25891 ( .A(n26012), .B(n26016), .Z(n26014) );
  XNOR U25892 ( .A(n25821), .B(n25925), .Z(n25927) );
  XNOR U25893 ( .A(n26017), .B(n26018), .Z(n25821) );
  AND U25894 ( .A(n441), .B(n25828), .Z(n26018) );
  XOR U25895 ( .A(n26017), .B(n25826), .Z(n25828) );
  AND U25896 ( .A(n25829), .B(n25832), .Z(n25925) );
  XOR U25897 ( .A(n26019), .B(n25976), .Z(n25832) );
  XNOR U25898 ( .A(p_input[1088]), .B(p_input[2048]), .Z(n25976) );
  XNOR U25899 ( .A(n25952), .B(n25951), .Z(n26019) );
  XNOR U25900 ( .A(n26020), .B(n25963), .Z(n25951) );
  XOR U25901 ( .A(n25937), .B(n25935), .Z(n25963) );
  XNOR U25902 ( .A(n26021), .B(n25942), .Z(n25935) );
  XOR U25903 ( .A(p_input[1112]), .B(p_input[2072]), .Z(n25942) );
  XOR U25904 ( .A(n25932), .B(n25941), .Z(n26021) );
  XOR U25905 ( .A(n26022), .B(n25938), .Z(n25941) );
  XOR U25906 ( .A(p_input[1110]), .B(p_input[2070]), .Z(n25938) );
  XOR U25907 ( .A(p_input[1111]), .B(n17295), .Z(n26022) );
  XOR U25908 ( .A(p_input[1106]), .B(p_input[2066]), .Z(n25932) );
  XNOR U25909 ( .A(n25947), .B(n25946), .Z(n25937) );
  XOR U25910 ( .A(n26023), .B(n25943), .Z(n25946) );
  XOR U25911 ( .A(p_input[1107]), .B(p_input[2067]), .Z(n25943) );
  XOR U25912 ( .A(p_input[1108]), .B(n17297), .Z(n26023) );
  XOR U25913 ( .A(p_input[1109]), .B(p_input[2069]), .Z(n25947) );
  XOR U25914 ( .A(n25962), .B(n26024), .Z(n26020) );
  IV U25915 ( .A(n25948), .Z(n26024) );
  XOR U25916 ( .A(p_input[1089]), .B(p_input[2049]), .Z(n25948) );
  XNOR U25917 ( .A(n26025), .B(n25970), .Z(n25962) );
  XNOR U25918 ( .A(n25958), .B(n25957), .Z(n25970) );
  XNOR U25919 ( .A(n26026), .B(n25954), .Z(n25957) );
  XNOR U25920 ( .A(p_input[1114]), .B(p_input[2074]), .Z(n25954) );
  XOR U25921 ( .A(p_input[1115]), .B(n17300), .Z(n26026) );
  XOR U25922 ( .A(p_input[1116]), .B(p_input[2076]), .Z(n25958) );
  XOR U25923 ( .A(n25968), .B(n26027), .Z(n26025) );
  IV U25924 ( .A(n25959), .Z(n26027) );
  XOR U25925 ( .A(p_input[1105]), .B(p_input[2065]), .Z(n25959) );
  XNOR U25926 ( .A(n26028), .B(n25975), .Z(n25968) );
  XNOR U25927 ( .A(p_input[1119]), .B(n17303), .Z(n25975) );
  XOR U25928 ( .A(n25965), .B(n25974), .Z(n26028) );
  XOR U25929 ( .A(n26029), .B(n25971), .Z(n25974) );
  XOR U25930 ( .A(p_input[1117]), .B(p_input[2077]), .Z(n25971) );
  XOR U25931 ( .A(p_input[1118]), .B(n17305), .Z(n26029) );
  XOR U25932 ( .A(p_input[1113]), .B(p_input[2073]), .Z(n25965) );
  XOR U25933 ( .A(n25987), .B(n25986), .Z(n25952) );
  XNOR U25934 ( .A(n26030), .B(n25994), .Z(n25986) );
  XNOR U25935 ( .A(n25982), .B(n25981), .Z(n25994) );
  XNOR U25936 ( .A(n26031), .B(n25978), .Z(n25981) );
  XNOR U25937 ( .A(p_input[1099]), .B(p_input[2059]), .Z(n25978) );
  XOR U25938 ( .A(p_input[1100]), .B(n16451), .Z(n26031) );
  XOR U25939 ( .A(p_input[1101]), .B(p_input[2061]), .Z(n25982) );
  XOR U25940 ( .A(n25992), .B(n26032), .Z(n26030) );
  IV U25941 ( .A(n25983), .Z(n26032) );
  XOR U25942 ( .A(p_input[1090]), .B(p_input[2050]), .Z(n25983) );
  XNOR U25943 ( .A(n26033), .B(n25999), .Z(n25992) );
  XNOR U25944 ( .A(p_input[1104]), .B(n16454), .Z(n25999) );
  XOR U25945 ( .A(n25989), .B(n25998), .Z(n26033) );
  XOR U25946 ( .A(n26034), .B(n25995), .Z(n25998) );
  XOR U25947 ( .A(p_input[1102]), .B(p_input[2062]), .Z(n25995) );
  XOR U25948 ( .A(p_input[1103]), .B(n16456), .Z(n26034) );
  XOR U25949 ( .A(p_input[1098]), .B(p_input[2058]), .Z(n25989) );
  XOR U25950 ( .A(n26006), .B(n26004), .Z(n25987) );
  XNOR U25951 ( .A(n26035), .B(n26011), .Z(n26004) );
  XOR U25952 ( .A(p_input[1097]), .B(p_input[2057]), .Z(n26011) );
  XOR U25953 ( .A(n26001), .B(n26010), .Z(n26035) );
  XOR U25954 ( .A(n26036), .B(n26007), .Z(n26010) );
  XOR U25955 ( .A(p_input[1095]), .B(p_input[2055]), .Z(n26007) );
  XOR U25956 ( .A(p_input[1096]), .B(n17312), .Z(n26036) );
  XOR U25957 ( .A(p_input[1091]), .B(p_input[2051]), .Z(n26001) );
  XNOR U25958 ( .A(n26016), .B(n26015), .Z(n26006) );
  XOR U25959 ( .A(n26037), .B(n26012), .Z(n26015) );
  XOR U25960 ( .A(p_input[1092]), .B(p_input[2052]), .Z(n26012) );
  XOR U25961 ( .A(p_input[1093]), .B(n17314), .Z(n26037) );
  XOR U25962 ( .A(p_input[1094]), .B(p_input[2054]), .Z(n26016) );
  XNOR U25963 ( .A(n26038), .B(n26039), .Z(n25829) );
  AND U25964 ( .A(n441), .B(n26040), .Z(n26039) );
  XNOR U25965 ( .A(n26041), .B(n26042), .Z(n441) );
  AND U25966 ( .A(n26043), .B(n26044), .Z(n26042) );
  XOR U25967 ( .A(n26041), .B(n25839), .Z(n26044) );
  XNOR U25968 ( .A(n26041), .B(n25781), .Z(n26043) );
  XOR U25969 ( .A(n26045), .B(n26046), .Z(n26041) );
  AND U25970 ( .A(n26047), .B(n26048), .Z(n26046) );
  XNOR U25971 ( .A(n25852), .B(n26045), .Z(n26048) );
  XOR U25972 ( .A(n26045), .B(n25793), .Z(n26047) );
  XOR U25973 ( .A(n26049), .B(n26050), .Z(n26045) );
  AND U25974 ( .A(n26051), .B(n26052), .Z(n26050) );
  XNOR U25975 ( .A(n25877), .B(n26049), .Z(n26052) );
  XOR U25976 ( .A(n26049), .B(n25804), .Z(n26051) );
  XOR U25977 ( .A(n26053), .B(n26054), .Z(n26049) );
  AND U25978 ( .A(n26055), .B(n26056), .Z(n26054) );
  XOR U25979 ( .A(n26053), .B(n25814), .Z(n26055) );
  XOR U25980 ( .A(n26057), .B(n26058), .Z(n25770) );
  AND U25981 ( .A(n445), .B(n26040), .Z(n26058) );
  XNOR U25982 ( .A(n26038), .B(n26057), .Z(n26040) );
  XNOR U25983 ( .A(n26059), .B(n26060), .Z(n445) );
  AND U25984 ( .A(n26061), .B(n26062), .Z(n26060) );
  XNOR U25985 ( .A(n26063), .B(n26059), .Z(n26062) );
  IV U25986 ( .A(n25839), .Z(n26063) );
  XNOR U25987 ( .A(n26064), .B(n26065), .Z(n25839) );
  AND U25988 ( .A(n448), .B(n26066), .Z(n26065) );
  XNOR U25989 ( .A(n26064), .B(n26067), .Z(n26066) );
  XNOR U25990 ( .A(n25781), .B(n26059), .Z(n26061) );
  XOR U25991 ( .A(n26068), .B(n26069), .Z(n25781) );
  AND U25992 ( .A(n456), .B(n26070), .Z(n26069) );
  XOR U25993 ( .A(n26071), .B(n26072), .Z(n26059) );
  AND U25994 ( .A(n26073), .B(n26074), .Z(n26072) );
  XNOR U25995 ( .A(n26071), .B(n25852), .Z(n26074) );
  XNOR U25996 ( .A(n26075), .B(n26076), .Z(n25852) );
  AND U25997 ( .A(n448), .B(n26077), .Z(n26076) );
  XOR U25998 ( .A(n26078), .B(n26075), .Z(n26077) );
  XNOR U25999 ( .A(n26079), .B(n26071), .Z(n26073) );
  IV U26000 ( .A(n25793), .Z(n26079) );
  XOR U26001 ( .A(n26080), .B(n26081), .Z(n25793) );
  AND U26002 ( .A(n456), .B(n26082), .Z(n26081) );
  XOR U26003 ( .A(n26083), .B(n26084), .Z(n26071) );
  AND U26004 ( .A(n26085), .B(n26086), .Z(n26084) );
  XNOR U26005 ( .A(n26083), .B(n25877), .Z(n26086) );
  XNOR U26006 ( .A(n26087), .B(n26088), .Z(n25877) );
  AND U26007 ( .A(n448), .B(n26089), .Z(n26088) );
  XNOR U26008 ( .A(n26090), .B(n26087), .Z(n26089) );
  XOR U26009 ( .A(n25804), .B(n26083), .Z(n26085) );
  XOR U26010 ( .A(n26091), .B(n26092), .Z(n25804) );
  AND U26011 ( .A(n456), .B(n26093), .Z(n26092) );
  XOR U26012 ( .A(n26053), .B(n26094), .Z(n26083) );
  AND U26013 ( .A(n26095), .B(n26056), .Z(n26094) );
  XNOR U26014 ( .A(n25923), .B(n26053), .Z(n26056) );
  XNOR U26015 ( .A(n26096), .B(n26097), .Z(n25923) );
  AND U26016 ( .A(n448), .B(n26098), .Z(n26097) );
  XOR U26017 ( .A(n26099), .B(n26096), .Z(n26098) );
  XNOR U26018 ( .A(n26100), .B(n26053), .Z(n26095) );
  IV U26019 ( .A(n25814), .Z(n26100) );
  XOR U26020 ( .A(n26101), .B(n26102), .Z(n25814) );
  AND U26021 ( .A(n456), .B(n26103), .Z(n26102) );
  XOR U26022 ( .A(n26104), .B(n26105), .Z(n26053) );
  AND U26023 ( .A(n26106), .B(n26107), .Z(n26105) );
  XNOR U26024 ( .A(n26104), .B(n26017), .Z(n26107) );
  XNOR U26025 ( .A(n26108), .B(n26109), .Z(n26017) );
  AND U26026 ( .A(n448), .B(n26110), .Z(n26109) );
  XNOR U26027 ( .A(n26111), .B(n26108), .Z(n26110) );
  XNOR U26028 ( .A(n26112), .B(n26104), .Z(n26106) );
  IV U26029 ( .A(n25826), .Z(n26112) );
  XOR U26030 ( .A(n26113), .B(n26114), .Z(n25826) );
  AND U26031 ( .A(n456), .B(n26115), .Z(n26114) );
  AND U26032 ( .A(n26057), .B(n26038), .Z(n26104) );
  XNOR U26033 ( .A(n26116), .B(n26117), .Z(n26038) );
  AND U26034 ( .A(n448), .B(n26118), .Z(n26117) );
  XNOR U26035 ( .A(n26119), .B(n26116), .Z(n26118) );
  XNOR U26036 ( .A(n26120), .B(n26121), .Z(n448) );
  AND U26037 ( .A(n26122), .B(n26123), .Z(n26121) );
  XOR U26038 ( .A(n26067), .B(n26120), .Z(n26123) );
  AND U26039 ( .A(n26124), .B(n26125), .Z(n26067) );
  XOR U26040 ( .A(n26120), .B(n26064), .Z(n26122) );
  XNOR U26041 ( .A(n26126), .B(n26127), .Z(n26064) );
  AND U26042 ( .A(n452), .B(n26070), .Z(n26127) );
  XOR U26043 ( .A(n26068), .B(n26126), .Z(n26070) );
  XOR U26044 ( .A(n26128), .B(n26129), .Z(n26120) );
  AND U26045 ( .A(n26130), .B(n26131), .Z(n26129) );
  XNOR U26046 ( .A(n26128), .B(n26124), .Z(n26131) );
  IV U26047 ( .A(n26078), .Z(n26124) );
  XOR U26048 ( .A(n26132), .B(n26133), .Z(n26078) );
  XOR U26049 ( .A(n26134), .B(n26125), .Z(n26133) );
  AND U26050 ( .A(n26090), .B(n26135), .Z(n26125) );
  AND U26051 ( .A(n26136), .B(n26137), .Z(n26134) );
  XOR U26052 ( .A(n26138), .B(n26132), .Z(n26136) );
  XNOR U26053 ( .A(n26075), .B(n26128), .Z(n26130) );
  XNOR U26054 ( .A(n26139), .B(n26140), .Z(n26075) );
  AND U26055 ( .A(n452), .B(n26082), .Z(n26140) );
  XOR U26056 ( .A(n26139), .B(n26080), .Z(n26082) );
  XOR U26057 ( .A(n26141), .B(n26142), .Z(n26128) );
  AND U26058 ( .A(n26143), .B(n26144), .Z(n26142) );
  XNOR U26059 ( .A(n26141), .B(n26090), .Z(n26144) );
  XOR U26060 ( .A(n26145), .B(n26137), .Z(n26090) );
  XNOR U26061 ( .A(n26146), .B(n26132), .Z(n26137) );
  XOR U26062 ( .A(n26147), .B(n26148), .Z(n26132) );
  AND U26063 ( .A(n26149), .B(n26150), .Z(n26148) );
  XOR U26064 ( .A(n26151), .B(n26147), .Z(n26149) );
  XNOR U26065 ( .A(n26152), .B(n26153), .Z(n26146) );
  AND U26066 ( .A(n26154), .B(n26155), .Z(n26153) );
  XOR U26067 ( .A(n26152), .B(n26156), .Z(n26154) );
  XNOR U26068 ( .A(n26138), .B(n26135), .Z(n26145) );
  AND U26069 ( .A(n26157), .B(n26158), .Z(n26135) );
  XOR U26070 ( .A(n26159), .B(n26160), .Z(n26138) );
  AND U26071 ( .A(n26161), .B(n26162), .Z(n26160) );
  XOR U26072 ( .A(n26159), .B(n26163), .Z(n26161) );
  XNOR U26073 ( .A(n26087), .B(n26141), .Z(n26143) );
  XNOR U26074 ( .A(n26164), .B(n26165), .Z(n26087) );
  AND U26075 ( .A(n452), .B(n26093), .Z(n26165) );
  XOR U26076 ( .A(n26164), .B(n26091), .Z(n26093) );
  XOR U26077 ( .A(n26166), .B(n26167), .Z(n26141) );
  AND U26078 ( .A(n26168), .B(n26169), .Z(n26167) );
  XNOR U26079 ( .A(n26166), .B(n26157), .Z(n26169) );
  IV U26080 ( .A(n26099), .Z(n26157) );
  XNOR U26081 ( .A(n26170), .B(n26150), .Z(n26099) );
  XNOR U26082 ( .A(n26171), .B(n26156), .Z(n26150) );
  XOR U26083 ( .A(n26172), .B(n26173), .Z(n26156) );
  AND U26084 ( .A(n26174), .B(n26175), .Z(n26173) );
  XOR U26085 ( .A(n26172), .B(n26176), .Z(n26174) );
  XNOR U26086 ( .A(n26155), .B(n26147), .Z(n26171) );
  XOR U26087 ( .A(n26177), .B(n26178), .Z(n26147) );
  AND U26088 ( .A(n26179), .B(n26180), .Z(n26178) );
  XNOR U26089 ( .A(n26181), .B(n26177), .Z(n26179) );
  XNOR U26090 ( .A(n26182), .B(n26152), .Z(n26155) );
  XOR U26091 ( .A(n26183), .B(n26184), .Z(n26152) );
  AND U26092 ( .A(n26185), .B(n26186), .Z(n26184) );
  XOR U26093 ( .A(n26183), .B(n26187), .Z(n26185) );
  XNOR U26094 ( .A(n26188), .B(n26189), .Z(n26182) );
  AND U26095 ( .A(n26190), .B(n26191), .Z(n26189) );
  XNOR U26096 ( .A(n26188), .B(n26192), .Z(n26190) );
  XNOR U26097 ( .A(n26151), .B(n26158), .Z(n26170) );
  AND U26098 ( .A(n26111), .B(n26193), .Z(n26158) );
  XOR U26099 ( .A(n26163), .B(n26162), .Z(n26151) );
  XNOR U26100 ( .A(n26194), .B(n26159), .Z(n26162) );
  XOR U26101 ( .A(n26195), .B(n26196), .Z(n26159) );
  AND U26102 ( .A(n26197), .B(n26198), .Z(n26196) );
  XOR U26103 ( .A(n26195), .B(n26199), .Z(n26197) );
  XNOR U26104 ( .A(n26200), .B(n26201), .Z(n26194) );
  AND U26105 ( .A(n26202), .B(n26203), .Z(n26201) );
  XOR U26106 ( .A(n26200), .B(n26204), .Z(n26202) );
  XOR U26107 ( .A(n26205), .B(n26206), .Z(n26163) );
  AND U26108 ( .A(n26207), .B(n26208), .Z(n26206) );
  XOR U26109 ( .A(n26205), .B(n26209), .Z(n26207) );
  XNOR U26110 ( .A(n26096), .B(n26166), .Z(n26168) );
  XNOR U26111 ( .A(n26210), .B(n26211), .Z(n26096) );
  AND U26112 ( .A(n452), .B(n26103), .Z(n26211) );
  XOR U26113 ( .A(n26210), .B(n26101), .Z(n26103) );
  XOR U26114 ( .A(n26212), .B(n26213), .Z(n26166) );
  AND U26115 ( .A(n26214), .B(n26215), .Z(n26213) );
  XNOR U26116 ( .A(n26212), .B(n26111), .Z(n26215) );
  XOR U26117 ( .A(n26216), .B(n26180), .Z(n26111) );
  XNOR U26118 ( .A(n26217), .B(n26187), .Z(n26180) );
  XOR U26119 ( .A(n26176), .B(n26175), .Z(n26187) );
  XNOR U26120 ( .A(n26218), .B(n26172), .Z(n26175) );
  XOR U26121 ( .A(n26219), .B(n26220), .Z(n26172) );
  AND U26122 ( .A(n26221), .B(n26222), .Z(n26220) );
  XNOR U26123 ( .A(n26223), .B(n26224), .Z(n26221) );
  IV U26124 ( .A(n26219), .Z(n26223) );
  XNOR U26125 ( .A(n26225), .B(n26226), .Z(n26218) );
  NOR U26126 ( .A(n26227), .B(n26228), .Z(n26226) );
  XNOR U26127 ( .A(n26225), .B(n26229), .Z(n26227) );
  XOR U26128 ( .A(n26230), .B(n26231), .Z(n26176) );
  NOR U26129 ( .A(n26232), .B(n26233), .Z(n26231) );
  XNOR U26130 ( .A(n26230), .B(n26234), .Z(n26232) );
  XNOR U26131 ( .A(n26186), .B(n26177), .Z(n26217) );
  XOR U26132 ( .A(n26235), .B(n26236), .Z(n26177) );
  AND U26133 ( .A(n26237), .B(n26238), .Z(n26236) );
  XOR U26134 ( .A(n26235), .B(n26239), .Z(n26237) );
  XOR U26135 ( .A(n26240), .B(n26192), .Z(n26186) );
  XOR U26136 ( .A(n26241), .B(n26242), .Z(n26192) );
  NOR U26137 ( .A(n26243), .B(n26244), .Z(n26242) );
  XOR U26138 ( .A(n26241), .B(n26245), .Z(n26243) );
  XNOR U26139 ( .A(n26191), .B(n26183), .Z(n26240) );
  XOR U26140 ( .A(n26246), .B(n26247), .Z(n26183) );
  AND U26141 ( .A(n26248), .B(n26249), .Z(n26247) );
  XOR U26142 ( .A(n26246), .B(n26250), .Z(n26248) );
  XNOR U26143 ( .A(n26251), .B(n26188), .Z(n26191) );
  XOR U26144 ( .A(n26252), .B(n26253), .Z(n26188) );
  AND U26145 ( .A(n26254), .B(n26255), .Z(n26253) );
  XNOR U26146 ( .A(n26256), .B(n26257), .Z(n26254) );
  IV U26147 ( .A(n26252), .Z(n26256) );
  XNOR U26148 ( .A(n26258), .B(n26259), .Z(n26251) );
  NOR U26149 ( .A(n26260), .B(n26261), .Z(n26259) );
  XNOR U26150 ( .A(n26258), .B(n26262), .Z(n26260) );
  XOR U26151 ( .A(n26181), .B(n26193), .Z(n26216) );
  NOR U26152 ( .A(n26119), .B(n26263), .Z(n26193) );
  XNOR U26153 ( .A(n26199), .B(n26198), .Z(n26181) );
  XNOR U26154 ( .A(n26264), .B(n26204), .Z(n26198) );
  XNOR U26155 ( .A(n26265), .B(n26266), .Z(n26204) );
  NOR U26156 ( .A(n26267), .B(n26268), .Z(n26266) );
  XOR U26157 ( .A(n26265), .B(n26269), .Z(n26267) );
  XNOR U26158 ( .A(n26203), .B(n26195), .Z(n26264) );
  XOR U26159 ( .A(n26270), .B(n26271), .Z(n26195) );
  AND U26160 ( .A(n26272), .B(n26273), .Z(n26271) );
  XOR U26161 ( .A(n26270), .B(n26274), .Z(n26272) );
  XNOR U26162 ( .A(n26275), .B(n26200), .Z(n26203) );
  XOR U26163 ( .A(n26276), .B(n26277), .Z(n26200) );
  AND U26164 ( .A(n26278), .B(n26279), .Z(n26277) );
  XNOR U26165 ( .A(n26280), .B(n26281), .Z(n26278) );
  IV U26166 ( .A(n26276), .Z(n26280) );
  XNOR U26167 ( .A(n26282), .B(n26283), .Z(n26275) );
  NOR U26168 ( .A(n26284), .B(n26285), .Z(n26283) );
  XNOR U26169 ( .A(n26282), .B(n26286), .Z(n26284) );
  XOR U26170 ( .A(n26209), .B(n26208), .Z(n26199) );
  XNOR U26171 ( .A(n26287), .B(n26205), .Z(n26208) );
  XOR U26172 ( .A(n26288), .B(n26289), .Z(n26205) );
  AND U26173 ( .A(n26290), .B(n26291), .Z(n26289) );
  XNOR U26174 ( .A(n26292), .B(n26293), .Z(n26290) );
  IV U26175 ( .A(n26288), .Z(n26292) );
  XNOR U26176 ( .A(n26294), .B(n26295), .Z(n26287) );
  NOR U26177 ( .A(n26296), .B(n26297), .Z(n26295) );
  XNOR U26178 ( .A(n26294), .B(n26298), .Z(n26296) );
  XOR U26179 ( .A(n26299), .B(n26300), .Z(n26209) );
  NOR U26180 ( .A(n26301), .B(n26302), .Z(n26300) );
  XNOR U26181 ( .A(n26299), .B(n26303), .Z(n26301) );
  XNOR U26182 ( .A(n26108), .B(n26212), .Z(n26214) );
  XNOR U26183 ( .A(n26304), .B(n26305), .Z(n26108) );
  AND U26184 ( .A(n452), .B(n26115), .Z(n26305) );
  XOR U26185 ( .A(n26304), .B(n26113), .Z(n26115) );
  AND U26186 ( .A(n26116), .B(n26119), .Z(n26212) );
  XOR U26187 ( .A(n26306), .B(n26263), .Z(n26119) );
  XNOR U26188 ( .A(p_input[1120]), .B(p_input[2048]), .Z(n26263) );
  XNOR U26189 ( .A(n26239), .B(n26238), .Z(n26306) );
  XNOR U26190 ( .A(n26307), .B(n26250), .Z(n26238) );
  XOR U26191 ( .A(n26224), .B(n26222), .Z(n26250) );
  XNOR U26192 ( .A(n26308), .B(n26229), .Z(n26222) );
  XOR U26193 ( .A(p_input[1144]), .B(p_input[2072]), .Z(n26229) );
  XOR U26194 ( .A(n26219), .B(n26228), .Z(n26308) );
  XOR U26195 ( .A(n26309), .B(n26225), .Z(n26228) );
  XOR U26196 ( .A(p_input[1142]), .B(p_input[2070]), .Z(n26225) );
  XOR U26197 ( .A(p_input[1143]), .B(n17295), .Z(n26309) );
  XOR U26198 ( .A(p_input[1138]), .B(p_input[2066]), .Z(n26219) );
  XNOR U26199 ( .A(n26234), .B(n26233), .Z(n26224) );
  XOR U26200 ( .A(n26310), .B(n26230), .Z(n26233) );
  XOR U26201 ( .A(p_input[1139]), .B(p_input[2067]), .Z(n26230) );
  XOR U26202 ( .A(p_input[1140]), .B(n17297), .Z(n26310) );
  XOR U26203 ( .A(p_input[1141]), .B(p_input[2069]), .Z(n26234) );
  XOR U26204 ( .A(n26249), .B(n26311), .Z(n26307) );
  IV U26205 ( .A(n26235), .Z(n26311) );
  XOR U26206 ( .A(p_input[1121]), .B(p_input[2049]), .Z(n26235) );
  XNOR U26207 ( .A(n26312), .B(n26257), .Z(n26249) );
  XNOR U26208 ( .A(n26245), .B(n26244), .Z(n26257) );
  XNOR U26209 ( .A(n26313), .B(n26241), .Z(n26244) );
  XNOR U26210 ( .A(p_input[1146]), .B(p_input[2074]), .Z(n26241) );
  XOR U26211 ( .A(p_input[1147]), .B(n17300), .Z(n26313) );
  XOR U26212 ( .A(p_input[1148]), .B(p_input[2076]), .Z(n26245) );
  XOR U26213 ( .A(n26255), .B(n26314), .Z(n26312) );
  IV U26214 ( .A(n26246), .Z(n26314) );
  XOR U26215 ( .A(p_input[1137]), .B(p_input[2065]), .Z(n26246) );
  XNOR U26216 ( .A(n26315), .B(n26262), .Z(n26255) );
  XNOR U26217 ( .A(p_input[1151]), .B(n17303), .Z(n26262) );
  XOR U26218 ( .A(n26252), .B(n26261), .Z(n26315) );
  XOR U26219 ( .A(n26316), .B(n26258), .Z(n26261) );
  XOR U26220 ( .A(p_input[1149]), .B(p_input[2077]), .Z(n26258) );
  XOR U26221 ( .A(p_input[1150]), .B(n17305), .Z(n26316) );
  XOR U26222 ( .A(p_input[1145]), .B(p_input[2073]), .Z(n26252) );
  XOR U26223 ( .A(n26274), .B(n26273), .Z(n26239) );
  XNOR U26224 ( .A(n26317), .B(n26281), .Z(n26273) );
  XNOR U26225 ( .A(n26269), .B(n26268), .Z(n26281) );
  XNOR U26226 ( .A(n26318), .B(n26265), .Z(n26268) );
  XNOR U26227 ( .A(p_input[1131]), .B(p_input[2059]), .Z(n26265) );
  XOR U26228 ( .A(p_input[1132]), .B(n16451), .Z(n26318) );
  XOR U26229 ( .A(p_input[1133]), .B(p_input[2061]), .Z(n26269) );
  XOR U26230 ( .A(n26279), .B(n26319), .Z(n26317) );
  IV U26231 ( .A(n26270), .Z(n26319) );
  XOR U26232 ( .A(p_input[1122]), .B(p_input[2050]), .Z(n26270) );
  XNOR U26233 ( .A(n26320), .B(n26286), .Z(n26279) );
  XNOR U26234 ( .A(p_input[1136]), .B(n16454), .Z(n26286) );
  XOR U26235 ( .A(n26276), .B(n26285), .Z(n26320) );
  XOR U26236 ( .A(n26321), .B(n26282), .Z(n26285) );
  XOR U26237 ( .A(p_input[1134]), .B(p_input[2062]), .Z(n26282) );
  XOR U26238 ( .A(p_input[1135]), .B(n16456), .Z(n26321) );
  XOR U26239 ( .A(p_input[1130]), .B(p_input[2058]), .Z(n26276) );
  XOR U26240 ( .A(n26293), .B(n26291), .Z(n26274) );
  XNOR U26241 ( .A(n26322), .B(n26298), .Z(n26291) );
  XOR U26242 ( .A(p_input[1129]), .B(p_input[2057]), .Z(n26298) );
  XOR U26243 ( .A(n26288), .B(n26297), .Z(n26322) );
  XOR U26244 ( .A(n26323), .B(n26294), .Z(n26297) );
  XOR U26245 ( .A(p_input[1127]), .B(p_input[2055]), .Z(n26294) );
  XOR U26246 ( .A(p_input[1128]), .B(n17312), .Z(n26323) );
  XOR U26247 ( .A(p_input[1123]), .B(p_input[2051]), .Z(n26288) );
  XNOR U26248 ( .A(n26303), .B(n26302), .Z(n26293) );
  XOR U26249 ( .A(n26324), .B(n26299), .Z(n26302) );
  XOR U26250 ( .A(p_input[1124]), .B(p_input[2052]), .Z(n26299) );
  XOR U26251 ( .A(p_input[1125]), .B(n17314), .Z(n26324) );
  XOR U26252 ( .A(p_input[1126]), .B(p_input[2054]), .Z(n26303) );
  XNOR U26253 ( .A(n26325), .B(n26326), .Z(n26116) );
  AND U26254 ( .A(n452), .B(n26327), .Z(n26326) );
  XNOR U26255 ( .A(n26328), .B(n26329), .Z(n452) );
  AND U26256 ( .A(n26330), .B(n26331), .Z(n26329) );
  XOR U26257 ( .A(n26328), .B(n26126), .Z(n26331) );
  XNOR U26258 ( .A(n26328), .B(n26068), .Z(n26330) );
  XOR U26259 ( .A(n26332), .B(n26333), .Z(n26328) );
  AND U26260 ( .A(n26334), .B(n26335), .Z(n26333) );
  XNOR U26261 ( .A(n26139), .B(n26332), .Z(n26335) );
  XOR U26262 ( .A(n26332), .B(n26080), .Z(n26334) );
  XOR U26263 ( .A(n26336), .B(n26337), .Z(n26332) );
  AND U26264 ( .A(n26338), .B(n26339), .Z(n26337) );
  XNOR U26265 ( .A(n26164), .B(n26336), .Z(n26339) );
  XOR U26266 ( .A(n26336), .B(n26091), .Z(n26338) );
  XOR U26267 ( .A(n26340), .B(n26341), .Z(n26336) );
  AND U26268 ( .A(n26342), .B(n26343), .Z(n26341) );
  XOR U26269 ( .A(n26340), .B(n26101), .Z(n26342) );
  XOR U26270 ( .A(n26344), .B(n26345), .Z(n26057) );
  AND U26271 ( .A(n456), .B(n26327), .Z(n26345) );
  XNOR U26272 ( .A(n26325), .B(n26344), .Z(n26327) );
  XNOR U26273 ( .A(n26346), .B(n26347), .Z(n456) );
  AND U26274 ( .A(n26348), .B(n26349), .Z(n26347) );
  XNOR U26275 ( .A(n26350), .B(n26346), .Z(n26349) );
  IV U26276 ( .A(n26126), .Z(n26350) );
  XNOR U26277 ( .A(n26351), .B(n26352), .Z(n26126) );
  AND U26278 ( .A(n459), .B(n26353), .Z(n26352) );
  XNOR U26279 ( .A(n26351), .B(n26354), .Z(n26353) );
  XNOR U26280 ( .A(n26068), .B(n26346), .Z(n26348) );
  XOR U26281 ( .A(n26355), .B(n26356), .Z(n26068) );
  AND U26282 ( .A(n467), .B(n26357), .Z(n26356) );
  XOR U26283 ( .A(n26358), .B(n26359), .Z(n26346) );
  AND U26284 ( .A(n26360), .B(n26361), .Z(n26359) );
  XNOR U26285 ( .A(n26358), .B(n26139), .Z(n26361) );
  XNOR U26286 ( .A(n26362), .B(n26363), .Z(n26139) );
  AND U26287 ( .A(n459), .B(n26364), .Z(n26363) );
  XOR U26288 ( .A(n26365), .B(n26362), .Z(n26364) );
  XNOR U26289 ( .A(n26366), .B(n26358), .Z(n26360) );
  IV U26290 ( .A(n26080), .Z(n26366) );
  XOR U26291 ( .A(n26367), .B(n26368), .Z(n26080) );
  AND U26292 ( .A(n467), .B(n26369), .Z(n26368) );
  XOR U26293 ( .A(n26370), .B(n26371), .Z(n26358) );
  AND U26294 ( .A(n26372), .B(n26373), .Z(n26371) );
  XNOR U26295 ( .A(n26370), .B(n26164), .Z(n26373) );
  XNOR U26296 ( .A(n26374), .B(n26375), .Z(n26164) );
  AND U26297 ( .A(n459), .B(n26376), .Z(n26375) );
  XNOR U26298 ( .A(n26377), .B(n26374), .Z(n26376) );
  XOR U26299 ( .A(n26091), .B(n26370), .Z(n26372) );
  XOR U26300 ( .A(n26378), .B(n26379), .Z(n26091) );
  AND U26301 ( .A(n467), .B(n26380), .Z(n26379) );
  XOR U26302 ( .A(n26340), .B(n26381), .Z(n26370) );
  AND U26303 ( .A(n26382), .B(n26343), .Z(n26381) );
  XNOR U26304 ( .A(n26210), .B(n26340), .Z(n26343) );
  XNOR U26305 ( .A(n26383), .B(n26384), .Z(n26210) );
  AND U26306 ( .A(n459), .B(n26385), .Z(n26384) );
  XOR U26307 ( .A(n26386), .B(n26383), .Z(n26385) );
  XNOR U26308 ( .A(n26387), .B(n26340), .Z(n26382) );
  IV U26309 ( .A(n26101), .Z(n26387) );
  XOR U26310 ( .A(n26388), .B(n26389), .Z(n26101) );
  AND U26311 ( .A(n467), .B(n26390), .Z(n26389) );
  XOR U26312 ( .A(n26391), .B(n26392), .Z(n26340) );
  AND U26313 ( .A(n26393), .B(n26394), .Z(n26392) );
  XNOR U26314 ( .A(n26391), .B(n26304), .Z(n26394) );
  XNOR U26315 ( .A(n26395), .B(n26396), .Z(n26304) );
  AND U26316 ( .A(n459), .B(n26397), .Z(n26396) );
  XNOR U26317 ( .A(n26398), .B(n26395), .Z(n26397) );
  XNOR U26318 ( .A(n26399), .B(n26391), .Z(n26393) );
  IV U26319 ( .A(n26113), .Z(n26399) );
  XOR U26320 ( .A(n26400), .B(n26401), .Z(n26113) );
  AND U26321 ( .A(n467), .B(n26402), .Z(n26401) );
  AND U26322 ( .A(n26344), .B(n26325), .Z(n26391) );
  XNOR U26323 ( .A(n26403), .B(n26404), .Z(n26325) );
  AND U26324 ( .A(n459), .B(n26405), .Z(n26404) );
  XNOR U26325 ( .A(n26406), .B(n26403), .Z(n26405) );
  XNOR U26326 ( .A(n26407), .B(n26408), .Z(n459) );
  AND U26327 ( .A(n26409), .B(n26410), .Z(n26408) );
  XOR U26328 ( .A(n26354), .B(n26407), .Z(n26410) );
  AND U26329 ( .A(n26411), .B(n26412), .Z(n26354) );
  XOR U26330 ( .A(n26407), .B(n26351), .Z(n26409) );
  XNOR U26331 ( .A(n26413), .B(n26414), .Z(n26351) );
  AND U26332 ( .A(n463), .B(n26357), .Z(n26414) );
  XOR U26333 ( .A(n26355), .B(n26413), .Z(n26357) );
  XOR U26334 ( .A(n26415), .B(n26416), .Z(n26407) );
  AND U26335 ( .A(n26417), .B(n26418), .Z(n26416) );
  XNOR U26336 ( .A(n26415), .B(n26411), .Z(n26418) );
  IV U26337 ( .A(n26365), .Z(n26411) );
  XOR U26338 ( .A(n26419), .B(n26420), .Z(n26365) );
  XOR U26339 ( .A(n26421), .B(n26412), .Z(n26420) );
  AND U26340 ( .A(n26377), .B(n26422), .Z(n26412) );
  AND U26341 ( .A(n26423), .B(n26424), .Z(n26421) );
  XOR U26342 ( .A(n26425), .B(n26419), .Z(n26423) );
  XNOR U26343 ( .A(n26362), .B(n26415), .Z(n26417) );
  XNOR U26344 ( .A(n26426), .B(n26427), .Z(n26362) );
  AND U26345 ( .A(n463), .B(n26369), .Z(n26427) );
  XOR U26346 ( .A(n26426), .B(n26367), .Z(n26369) );
  XOR U26347 ( .A(n26428), .B(n26429), .Z(n26415) );
  AND U26348 ( .A(n26430), .B(n26431), .Z(n26429) );
  XNOR U26349 ( .A(n26428), .B(n26377), .Z(n26431) );
  XOR U26350 ( .A(n26432), .B(n26424), .Z(n26377) );
  XNOR U26351 ( .A(n26433), .B(n26419), .Z(n26424) );
  XOR U26352 ( .A(n26434), .B(n26435), .Z(n26419) );
  AND U26353 ( .A(n26436), .B(n26437), .Z(n26435) );
  XOR U26354 ( .A(n26438), .B(n26434), .Z(n26436) );
  XNOR U26355 ( .A(n26439), .B(n26440), .Z(n26433) );
  AND U26356 ( .A(n26441), .B(n26442), .Z(n26440) );
  XOR U26357 ( .A(n26439), .B(n26443), .Z(n26441) );
  XNOR U26358 ( .A(n26425), .B(n26422), .Z(n26432) );
  AND U26359 ( .A(n26444), .B(n26445), .Z(n26422) );
  XOR U26360 ( .A(n26446), .B(n26447), .Z(n26425) );
  AND U26361 ( .A(n26448), .B(n26449), .Z(n26447) );
  XOR U26362 ( .A(n26446), .B(n26450), .Z(n26448) );
  XNOR U26363 ( .A(n26374), .B(n26428), .Z(n26430) );
  XNOR U26364 ( .A(n26451), .B(n26452), .Z(n26374) );
  AND U26365 ( .A(n463), .B(n26380), .Z(n26452) );
  XOR U26366 ( .A(n26451), .B(n26378), .Z(n26380) );
  XOR U26367 ( .A(n26453), .B(n26454), .Z(n26428) );
  AND U26368 ( .A(n26455), .B(n26456), .Z(n26454) );
  XNOR U26369 ( .A(n26453), .B(n26444), .Z(n26456) );
  IV U26370 ( .A(n26386), .Z(n26444) );
  XNOR U26371 ( .A(n26457), .B(n26437), .Z(n26386) );
  XNOR U26372 ( .A(n26458), .B(n26443), .Z(n26437) );
  XOR U26373 ( .A(n26459), .B(n26460), .Z(n26443) );
  AND U26374 ( .A(n26461), .B(n26462), .Z(n26460) );
  XOR U26375 ( .A(n26459), .B(n26463), .Z(n26461) );
  XNOR U26376 ( .A(n26442), .B(n26434), .Z(n26458) );
  XOR U26377 ( .A(n26464), .B(n26465), .Z(n26434) );
  AND U26378 ( .A(n26466), .B(n26467), .Z(n26465) );
  XNOR U26379 ( .A(n26468), .B(n26464), .Z(n26466) );
  XNOR U26380 ( .A(n26469), .B(n26439), .Z(n26442) );
  XOR U26381 ( .A(n26470), .B(n26471), .Z(n26439) );
  AND U26382 ( .A(n26472), .B(n26473), .Z(n26471) );
  XOR U26383 ( .A(n26470), .B(n26474), .Z(n26472) );
  XNOR U26384 ( .A(n26475), .B(n26476), .Z(n26469) );
  AND U26385 ( .A(n26477), .B(n26478), .Z(n26476) );
  XNOR U26386 ( .A(n26475), .B(n26479), .Z(n26477) );
  XNOR U26387 ( .A(n26438), .B(n26445), .Z(n26457) );
  AND U26388 ( .A(n26398), .B(n26480), .Z(n26445) );
  XOR U26389 ( .A(n26450), .B(n26449), .Z(n26438) );
  XNOR U26390 ( .A(n26481), .B(n26446), .Z(n26449) );
  XOR U26391 ( .A(n26482), .B(n26483), .Z(n26446) );
  AND U26392 ( .A(n26484), .B(n26485), .Z(n26483) );
  XOR U26393 ( .A(n26482), .B(n26486), .Z(n26484) );
  XNOR U26394 ( .A(n26487), .B(n26488), .Z(n26481) );
  AND U26395 ( .A(n26489), .B(n26490), .Z(n26488) );
  XOR U26396 ( .A(n26487), .B(n26491), .Z(n26489) );
  XOR U26397 ( .A(n26492), .B(n26493), .Z(n26450) );
  AND U26398 ( .A(n26494), .B(n26495), .Z(n26493) );
  XOR U26399 ( .A(n26492), .B(n26496), .Z(n26494) );
  XNOR U26400 ( .A(n26383), .B(n26453), .Z(n26455) );
  XNOR U26401 ( .A(n26497), .B(n26498), .Z(n26383) );
  AND U26402 ( .A(n463), .B(n26390), .Z(n26498) );
  XOR U26403 ( .A(n26497), .B(n26388), .Z(n26390) );
  XOR U26404 ( .A(n26499), .B(n26500), .Z(n26453) );
  AND U26405 ( .A(n26501), .B(n26502), .Z(n26500) );
  XNOR U26406 ( .A(n26499), .B(n26398), .Z(n26502) );
  XOR U26407 ( .A(n26503), .B(n26467), .Z(n26398) );
  XNOR U26408 ( .A(n26504), .B(n26474), .Z(n26467) );
  XOR U26409 ( .A(n26463), .B(n26462), .Z(n26474) );
  XNOR U26410 ( .A(n26505), .B(n26459), .Z(n26462) );
  XOR U26411 ( .A(n26506), .B(n26507), .Z(n26459) );
  AND U26412 ( .A(n26508), .B(n26509), .Z(n26507) );
  XNOR U26413 ( .A(n26510), .B(n26511), .Z(n26508) );
  IV U26414 ( .A(n26506), .Z(n26510) );
  XNOR U26415 ( .A(n26512), .B(n26513), .Z(n26505) );
  NOR U26416 ( .A(n26514), .B(n26515), .Z(n26513) );
  XNOR U26417 ( .A(n26512), .B(n26516), .Z(n26514) );
  XOR U26418 ( .A(n26517), .B(n26518), .Z(n26463) );
  NOR U26419 ( .A(n26519), .B(n26520), .Z(n26518) );
  XNOR U26420 ( .A(n26517), .B(n26521), .Z(n26519) );
  XNOR U26421 ( .A(n26473), .B(n26464), .Z(n26504) );
  XOR U26422 ( .A(n26522), .B(n26523), .Z(n26464) );
  AND U26423 ( .A(n26524), .B(n26525), .Z(n26523) );
  XOR U26424 ( .A(n26522), .B(n26526), .Z(n26524) );
  XOR U26425 ( .A(n26527), .B(n26479), .Z(n26473) );
  XOR U26426 ( .A(n26528), .B(n26529), .Z(n26479) );
  NOR U26427 ( .A(n26530), .B(n26531), .Z(n26529) );
  XOR U26428 ( .A(n26528), .B(n26532), .Z(n26530) );
  XNOR U26429 ( .A(n26478), .B(n26470), .Z(n26527) );
  XOR U26430 ( .A(n26533), .B(n26534), .Z(n26470) );
  AND U26431 ( .A(n26535), .B(n26536), .Z(n26534) );
  XOR U26432 ( .A(n26533), .B(n26537), .Z(n26535) );
  XNOR U26433 ( .A(n26538), .B(n26475), .Z(n26478) );
  XOR U26434 ( .A(n26539), .B(n26540), .Z(n26475) );
  AND U26435 ( .A(n26541), .B(n26542), .Z(n26540) );
  XNOR U26436 ( .A(n26543), .B(n26544), .Z(n26541) );
  IV U26437 ( .A(n26539), .Z(n26543) );
  XNOR U26438 ( .A(n26545), .B(n26546), .Z(n26538) );
  NOR U26439 ( .A(n26547), .B(n26548), .Z(n26546) );
  XNOR U26440 ( .A(n26545), .B(n26549), .Z(n26547) );
  XOR U26441 ( .A(n26468), .B(n26480), .Z(n26503) );
  NOR U26442 ( .A(n26406), .B(n26550), .Z(n26480) );
  XNOR U26443 ( .A(n26486), .B(n26485), .Z(n26468) );
  XNOR U26444 ( .A(n26551), .B(n26491), .Z(n26485) );
  XNOR U26445 ( .A(n26552), .B(n26553), .Z(n26491) );
  NOR U26446 ( .A(n26554), .B(n26555), .Z(n26553) );
  XOR U26447 ( .A(n26552), .B(n26556), .Z(n26554) );
  XNOR U26448 ( .A(n26490), .B(n26482), .Z(n26551) );
  XOR U26449 ( .A(n26557), .B(n26558), .Z(n26482) );
  AND U26450 ( .A(n26559), .B(n26560), .Z(n26558) );
  XOR U26451 ( .A(n26557), .B(n26561), .Z(n26559) );
  XNOR U26452 ( .A(n26562), .B(n26487), .Z(n26490) );
  XOR U26453 ( .A(n26563), .B(n26564), .Z(n26487) );
  AND U26454 ( .A(n26565), .B(n26566), .Z(n26564) );
  XNOR U26455 ( .A(n26567), .B(n26568), .Z(n26565) );
  IV U26456 ( .A(n26563), .Z(n26567) );
  XNOR U26457 ( .A(n26569), .B(n26570), .Z(n26562) );
  NOR U26458 ( .A(n26571), .B(n26572), .Z(n26570) );
  XNOR U26459 ( .A(n26569), .B(n26573), .Z(n26571) );
  XOR U26460 ( .A(n26496), .B(n26495), .Z(n26486) );
  XNOR U26461 ( .A(n26574), .B(n26492), .Z(n26495) );
  XOR U26462 ( .A(n26575), .B(n26576), .Z(n26492) );
  AND U26463 ( .A(n26577), .B(n26578), .Z(n26576) );
  XNOR U26464 ( .A(n26579), .B(n26580), .Z(n26577) );
  IV U26465 ( .A(n26575), .Z(n26579) );
  XNOR U26466 ( .A(n26581), .B(n26582), .Z(n26574) );
  NOR U26467 ( .A(n26583), .B(n26584), .Z(n26582) );
  XNOR U26468 ( .A(n26581), .B(n26585), .Z(n26583) );
  XOR U26469 ( .A(n26586), .B(n26587), .Z(n26496) );
  NOR U26470 ( .A(n26588), .B(n26589), .Z(n26587) );
  XNOR U26471 ( .A(n26586), .B(n26590), .Z(n26588) );
  XNOR U26472 ( .A(n26395), .B(n26499), .Z(n26501) );
  XNOR U26473 ( .A(n26591), .B(n26592), .Z(n26395) );
  AND U26474 ( .A(n463), .B(n26402), .Z(n26592) );
  XOR U26475 ( .A(n26591), .B(n26400), .Z(n26402) );
  AND U26476 ( .A(n26403), .B(n26406), .Z(n26499) );
  XOR U26477 ( .A(n26593), .B(n26550), .Z(n26406) );
  XNOR U26478 ( .A(p_input[1152]), .B(p_input[2048]), .Z(n26550) );
  XNOR U26479 ( .A(n26526), .B(n26525), .Z(n26593) );
  XNOR U26480 ( .A(n26594), .B(n26537), .Z(n26525) );
  XOR U26481 ( .A(n26511), .B(n26509), .Z(n26537) );
  XNOR U26482 ( .A(n26595), .B(n26516), .Z(n26509) );
  XOR U26483 ( .A(p_input[1176]), .B(p_input[2072]), .Z(n26516) );
  XOR U26484 ( .A(n26506), .B(n26515), .Z(n26595) );
  XOR U26485 ( .A(n26596), .B(n26512), .Z(n26515) );
  XOR U26486 ( .A(p_input[1174]), .B(p_input[2070]), .Z(n26512) );
  XOR U26487 ( .A(p_input[1175]), .B(n17295), .Z(n26596) );
  XOR U26488 ( .A(p_input[1170]), .B(p_input[2066]), .Z(n26506) );
  XNOR U26489 ( .A(n26521), .B(n26520), .Z(n26511) );
  XOR U26490 ( .A(n26597), .B(n26517), .Z(n26520) );
  XOR U26491 ( .A(p_input[1171]), .B(p_input[2067]), .Z(n26517) );
  XOR U26492 ( .A(p_input[1172]), .B(n17297), .Z(n26597) );
  XOR U26493 ( .A(p_input[1173]), .B(p_input[2069]), .Z(n26521) );
  XOR U26494 ( .A(n26536), .B(n26598), .Z(n26594) );
  IV U26495 ( .A(n26522), .Z(n26598) );
  XOR U26496 ( .A(p_input[1153]), .B(p_input[2049]), .Z(n26522) );
  XNOR U26497 ( .A(n26599), .B(n26544), .Z(n26536) );
  XNOR U26498 ( .A(n26532), .B(n26531), .Z(n26544) );
  XNOR U26499 ( .A(n26600), .B(n26528), .Z(n26531) );
  XNOR U26500 ( .A(p_input[1178]), .B(p_input[2074]), .Z(n26528) );
  XOR U26501 ( .A(p_input[1179]), .B(n17300), .Z(n26600) );
  XOR U26502 ( .A(p_input[1180]), .B(p_input[2076]), .Z(n26532) );
  XOR U26503 ( .A(n26542), .B(n26601), .Z(n26599) );
  IV U26504 ( .A(n26533), .Z(n26601) );
  XOR U26505 ( .A(p_input[1169]), .B(p_input[2065]), .Z(n26533) );
  XNOR U26506 ( .A(n26602), .B(n26549), .Z(n26542) );
  XNOR U26507 ( .A(p_input[1183]), .B(n17303), .Z(n26549) );
  XOR U26508 ( .A(n26539), .B(n26548), .Z(n26602) );
  XOR U26509 ( .A(n26603), .B(n26545), .Z(n26548) );
  XOR U26510 ( .A(p_input[1181]), .B(p_input[2077]), .Z(n26545) );
  XOR U26511 ( .A(p_input[1182]), .B(n17305), .Z(n26603) );
  XOR U26512 ( .A(p_input[1177]), .B(p_input[2073]), .Z(n26539) );
  XOR U26513 ( .A(n26561), .B(n26560), .Z(n26526) );
  XNOR U26514 ( .A(n26604), .B(n26568), .Z(n26560) );
  XNOR U26515 ( .A(n26556), .B(n26555), .Z(n26568) );
  XNOR U26516 ( .A(n26605), .B(n26552), .Z(n26555) );
  XNOR U26517 ( .A(p_input[1163]), .B(p_input[2059]), .Z(n26552) );
  XOR U26518 ( .A(p_input[1164]), .B(n16451), .Z(n26605) );
  XOR U26519 ( .A(p_input[1165]), .B(p_input[2061]), .Z(n26556) );
  XOR U26520 ( .A(n26566), .B(n26606), .Z(n26604) );
  IV U26521 ( .A(n26557), .Z(n26606) );
  XOR U26522 ( .A(p_input[1154]), .B(p_input[2050]), .Z(n26557) );
  XNOR U26523 ( .A(n26607), .B(n26573), .Z(n26566) );
  XNOR U26524 ( .A(p_input[1168]), .B(n16454), .Z(n26573) );
  XOR U26525 ( .A(n26563), .B(n26572), .Z(n26607) );
  XOR U26526 ( .A(n26608), .B(n26569), .Z(n26572) );
  XOR U26527 ( .A(p_input[1166]), .B(p_input[2062]), .Z(n26569) );
  XOR U26528 ( .A(p_input[1167]), .B(n16456), .Z(n26608) );
  XOR U26529 ( .A(p_input[1162]), .B(p_input[2058]), .Z(n26563) );
  XOR U26530 ( .A(n26580), .B(n26578), .Z(n26561) );
  XNOR U26531 ( .A(n26609), .B(n26585), .Z(n26578) );
  XOR U26532 ( .A(p_input[1161]), .B(p_input[2057]), .Z(n26585) );
  XOR U26533 ( .A(n26575), .B(n26584), .Z(n26609) );
  XOR U26534 ( .A(n26610), .B(n26581), .Z(n26584) );
  XOR U26535 ( .A(p_input[1159]), .B(p_input[2055]), .Z(n26581) );
  XOR U26536 ( .A(p_input[1160]), .B(n17312), .Z(n26610) );
  XOR U26537 ( .A(p_input[1155]), .B(p_input[2051]), .Z(n26575) );
  XNOR U26538 ( .A(n26590), .B(n26589), .Z(n26580) );
  XOR U26539 ( .A(n26611), .B(n26586), .Z(n26589) );
  XOR U26540 ( .A(p_input[1156]), .B(p_input[2052]), .Z(n26586) );
  XOR U26541 ( .A(p_input[1157]), .B(n17314), .Z(n26611) );
  XOR U26542 ( .A(p_input[1158]), .B(p_input[2054]), .Z(n26590) );
  XNOR U26543 ( .A(n26612), .B(n26613), .Z(n26403) );
  AND U26544 ( .A(n463), .B(n26614), .Z(n26613) );
  XNOR U26545 ( .A(n26615), .B(n26616), .Z(n463) );
  AND U26546 ( .A(n26617), .B(n26618), .Z(n26616) );
  XOR U26547 ( .A(n26615), .B(n26413), .Z(n26618) );
  XNOR U26548 ( .A(n26615), .B(n26355), .Z(n26617) );
  XOR U26549 ( .A(n26619), .B(n26620), .Z(n26615) );
  AND U26550 ( .A(n26621), .B(n26622), .Z(n26620) );
  XNOR U26551 ( .A(n26426), .B(n26619), .Z(n26622) );
  XOR U26552 ( .A(n26619), .B(n26367), .Z(n26621) );
  XOR U26553 ( .A(n26623), .B(n26624), .Z(n26619) );
  AND U26554 ( .A(n26625), .B(n26626), .Z(n26624) );
  XNOR U26555 ( .A(n26451), .B(n26623), .Z(n26626) );
  XOR U26556 ( .A(n26623), .B(n26378), .Z(n26625) );
  XOR U26557 ( .A(n26627), .B(n26628), .Z(n26623) );
  AND U26558 ( .A(n26629), .B(n26630), .Z(n26628) );
  XOR U26559 ( .A(n26627), .B(n26388), .Z(n26629) );
  XOR U26560 ( .A(n26631), .B(n26632), .Z(n26344) );
  AND U26561 ( .A(n467), .B(n26614), .Z(n26632) );
  XNOR U26562 ( .A(n26612), .B(n26631), .Z(n26614) );
  XNOR U26563 ( .A(n26633), .B(n26634), .Z(n467) );
  AND U26564 ( .A(n26635), .B(n26636), .Z(n26634) );
  XNOR U26565 ( .A(n26637), .B(n26633), .Z(n26636) );
  IV U26566 ( .A(n26413), .Z(n26637) );
  XNOR U26567 ( .A(n26638), .B(n26639), .Z(n26413) );
  AND U26568 ( .A(n470), .B(n26640), .Z(n26639) );
  XNOR U26569 ( .A(n26638), .B(n26641), .Z(n26640) );
  XNOR U26570 ( .A(n26355), .B(n26633), .Z(n26635) );
  XOR U26571 ( .A(n26642), .B(n26643), .Z(n26355) );
  AND U26572 ( .A(n478), .B(n26644), .Z(n26643) );
  XOR U26573 ( .A(n26645), .B(n26646), .Z(n26633) );
  AND U26574 ( .A(n26647), .B(n26648), .Z(n26646) );
  XNOR U26575 ( .A(n26645), .B(n26426), .Z(n26648) );
  XNOR U26576 ( .A(n26649), .B(n26650), .Z(n26426) );
  AND U26577 ( .A(n470), .B(n26651), .Z(n26650) );
  XOR U26578 ( .A(n26652), .B(n26649), .Z(n26651) );
  XNOR U26579 ( .A(n26653), .B(n26645), .Z(n26647) );
  IV U26580 ( .A(n26367), .Z(n26653) );
  XOR U26581 ( .A(n26654), .B(n26655), .Z(n26367) );
  AND U26582 ( .A(n478), .B(n26656), .Z(n26655) );
  XOR U26583 ( .A(n26657), .B(n26658), .Z(n26645) );
  AND U26584 ( .A(n26659), .B(n26660), .Z(n26658) );
  XNOR U26585 ( .A(n26657), .B(n26451), .Z(n26660) );
  XNOR U26586 ( .A(n26661), .B(n26662), .Z(n26451) );
  AND U26587 ( .A(n470), .B(n26663), .Z(n26662) );
  XNOR U26588 ( .A(n26664), .B(n26661), .Z(n26663) );
  XOR U26589 ( .A(n26378), .B(n26657), .Z(n26659) );
  XOR U26590 ( .A(n26665), .B(n26666), .Z(n26378) );
  AND U26591 ( .A(n478), .B(n26667), .Z(n26666) );
  XOR U26592 ( .A(n26627), .B(n26668), .Z(n26657) );
  AND U26593 ( .A(n26669), .B(n26630), .Z(n26668) );
  XNOR U26594 ( .A(n26497), .B(n26627), .Z(n26630) );
  XNOR U26595 ( .A(n26670), .B(n26671), .Z(n26497) );
  AND U26596 ( .A(n470), .B(n26672), .Z(n26671) );
  XOR U26597 ( .A(n26673), .B(n26670), .Z(n26672) );
  XNOR U26598 ( .A(n26674), .B(n26627), .Z(n26669) );
  IV U26599 ( .A(n26388), .Z(n26674) );
  XOR U26600 ( .A(n26675), .B(n26676), .Z(n26388) );
  AND U26601 ( .A(n478), .B(n26677), .Z(n26676) );
  XOR U26602 ( .A(n26678), .B(n26679), .Z(n26627) );
  AND U26603 ( .A(n26680), .B(n26681), .Z(n26679) );
  XNOR U26604 ( .A(n26678), .B(n26591), .Z(n26681) );
  XNOR U26605 ( .A(n26682), .B(n26683), .Z(n26591) );
  AND U26606 ( .A(n470), .B(n26684), .Z(n26683) );
  XNOR U26607 ( .A(n26685), .B(n26682), .Z(n26684) );
  XNOR U26608 ( .A(n26686), .B(n26678), .Z(n26680) );
  IV U26609 ( .A(n26400), .Z(n26686) );
  XOR U26610 ( .A(n26687), .B(n26688), .Z(n26400) );
  AND U26611 ( .A(n478), .B(n26689), .Z(n26688) );
  AND U26612 ( .A(n26631), .B(n26612), .Z(n26678) );
  XNOR U26613 ( .A(n26690), .B(n26691), .Z(n26612) );
  AND U26614 ( .A(n470), .B(n26692), .Z(n26691) );
  XNOR U26615 ( .A(n26693), .B(n26690), .Z(n26692) );
  XNOR U26616 ( .A(n26694), .B(n26695), .Z(n470) );
  AND U26617 ( .A(n26696), .B(n26697), .Z(n26695) );
  XOR U26618 ( .A(n26641), .B(n26694), .Z(n26697) );
  AND U26619 ( .A(n26698), .B(n26699), .Z(n26641) );
  XOR U26620 ( .A(n26694), .B(n26638), .Z(n26696) );
  XNOR U26621 ( .A(n26700), .B(n26701), .Z(n26638) );
  AND U26622 ( .A(n474), .B(n26644), .Z(n26701) );
  XOR U26623 ( .A(n26642), .B(n26700), .Z(n26644) );
  XOR U26624 ( .A(n26702), .B(n26703), .Z(n26694) );
  AND U26625 ( .A(n26704), .B(n26705), .Z(n26703) );
  XNOR U26626 ( .A(n26702), .B(n26698), .Z(n26705) );
  IV U26627 ( .A(n26652), .Z(n26698) );
  XOR U26628 ( .A(n26706), .B(n26707), .Z(n26652) );
  XOR U26629 ( .A(n26708), .B(n26699), .Z(n26707) );
  AND U26630 ( .A(n26664), .B(n26709), .Z(n26699) );
  AND U26631 ( .A(n26710), .B(n26711), .Z(n26708) );
  XOR U26632 ( .A(n26712), .B(n26706), .Z(n26710) );
  XNOR U26633 ( .A(n26649), .B(n26702), .Z(n26704) );
  XNOR U26634 ( .A(n26713), .B(n26714), .Z(n26649) );
  AND U26635 ( .A(n474), .B(n26656), .Z(n26714) );
  XOR U26636 ( .A(n26713), .B(n26654), .Z(n26656) );
  XOR U26637 ( .A(n26715), .B(n26716), .Z(n26702) );
  AND U26638 ( .A(n26717), .B(n26718), .Z(n26716) );
  XNOR U26639 ( .A(n26715), .B(n26664), .Z(n26718) );
  XOR U26640 ( .A(n26719), .B(n26711), .Z(n26664) );
  XNOR U26641 ( .A(n26720), .B(n26706), .Z(n26711) );
  XOR U26642 ( .A(n26721), .B(n26722), .Z(n26706) );
  AND U26643 ( .A(n26723), .B(n26724), .Z(n26722) );
  XOR U26644 ( .A(n26725), .B(n26721), .Z(n26723) );
  XNOR U26645 ( .A(n26726), .B(n26727), .Z(n26720) );
  AND U26646 ( .A(n26728), .B(n26729), .Z(n26727) );
  XOR U26647 ( .A(n26726), .B(n26730), .Z(n26728) );
  XNOR U26648 ( .A(n26712), .B(n26709), .Z(n26719) );
  AND U26649 ( .A(n26731), .B(n26732), .Z(n26709) );
  XOR U26650 ( .A(n26733), .B(n26734), .Z(n26712) );
  AND U26651 ( .A(n26735), .B(n26736), .Z(n26734) );
  XOR U26652 ( .A(n26733), .B(n26737), .Z(n26735) );
  XNOR U26653 ( .A(n26661), .B(n26715), .Z(n26717) );
  XNOR U26654 ( .A(n26738), .B(n26739), .Z(n26661) );
  AND U26655 ( .A(n474), .B(n26667), .Z(n26739) );
  XOR U26656 ( .A(n26738), .B(n26665), .Z(n26667) );
  XOR U26657 ( .A(n26740), .B(n26741), .Z(n26715) );
  AND U26658 ( .A(n26742), .B(n26743), .Z(n26741) );
  XNOR U26659 ( .A(n26740), .B(n26731), .Z(n26743) );
  IV U26660 ( .A(n26673), .Z(n26731) );
  XNOR U26661 ( .A(n26744), .B(n26724), .Z(n26673) );
  XNOR U26662 ( .A(n26745), .B(n26730), .Z(n26724) );
  XOR U26663 ( .A(n26746), .B(n26747), .Z(n26730) );
  AND U26664 ( .A(n26748), .B(n26749), .Z(n26747) );
  XOR U26665 ( .A(n26746), .B(n26750), .Z(n26748) );
  XNOR U26666 ( .A(n26729), .B(n26721), .Z(n26745) );
  XOR U26667 ( .A(n26751), .B(n26752), .Z(n26721) );
  AND U26668 ( .A(n26753), .B(n26754), .Z(n26752) );
  XNOR U26669 ( .A(n26755), .B(n26751), .Z(n26753) );
  XNOR U26670 ( .A(n26756), .B(n26726), .Z(n26729) );
  XOR U26671 ( .A(n26757), .B(n26758), .Z(n26726) );
  AND U26672 ( .A(n26759), .B(n26760), .Z(n26758) );
  XOR U26673 ( .A(n26757), .B(n26761), .Z(n26759) );
  XNOR U26674 ( .A(n26762), .B(n26763), .Z(n26756) );
  AND U26675 ( .A(n26764), .B(n26765), .Z(n26763) );
  XNOR U26676 ( .A(n26762), .B(n26766), .Z(n26764) );
  XNOR U26677 ( .A(n26725), .B(n26732), .Z(n26744) );
  AND U26678 ( .A(n26685), .B(n26767), .Z(n26732) );
  XOR U26679 ( .A(n26737), .B(n26736), .Z(n26725) );
  XNOR U26680 ( .A(n26768), .B(n26733), .Z(n26736) );
  XOR U26681 ( .A(n26769), .B(n26770), .Z(n26733) );
  AND U26682 ( .A(n26771), .B(n26772), .Z(n26770) );
  XOR U26683 ( .A(n26769), .B(n26773), .Z(n26771) );
  XNOR U26684 ( .A(n26774), .B(n26775), .Z(n26768) );
  AND U26685 ( .A(n26776), .B(n26777), .Z(n26775) );
  XOR U26686 ( .A(n26774), .B(n26778), .Z(n26776) );
  XOR U26687 ( .A(n26779), .B(n26780), .Z(n26737) );
  AND U26688 ( .A(n26781), .B(n26782), .Z(n26780) );
  XOR U26689 ( .A(n26779), .B(n26783), .Z(n26781) );
  XNOR U26690 ( .A(n26670), .B(n26740), .Z(n26742) );
  XNOR U26691 ( .A(n26784), .B(n26785), .Z(n26670) );
  AND U26692 ( .A(n474), .B(n26677), .Z(n26785) );
  XOR U26693 ( .A(n26784), .B(n26675), .Z(n26677) );
  XOR U26694 ( .A(n26786), .B(n26787), .Z(n26740) );
  AND U26695 ( .A(n26788), .B(n26789), .Z(n26787) );
  XNOR U26696 ( .A(n26786), .B(n26685), .Z(n26789) );
  XOR U26697 ( .A(n26790), .B(n26754), .Z(n26685) );
  XNOR U26698 ( .A(n26791), .B(n26761), .Z(n26754) );
  XOR U26699 ( .A(n26750), .B(n26749), .Z(n26761) );
  XNOR U26700 ( .A(n26792), .B(n26746), .Z(n26749) );
  XOR U26701 ( .A(n26793), .B(n26794), .Z(n26746) );
  AND U26702 ( .A(n26795), .B(n26796), .Z(n26794) );
  XNOR U26703 ( .A(n26797), .B(n26798), .Z(n26795) );
  IV U26704 ( .A(n26793), .Z(n26797) );
  XNOR U26705 ( .A(n26799), .B(n26800), .Z(n26792) );
  NOR U26706 ( .A(n26801), .B(n26802), .Z(n26800) );
  XNOR U26707 ( .A(n26799), .B(n26803), .Z(n26801) );
  XOR U26708 ( .A(n26804), .B(n26805), .Z(n26750) );
  NOR U26709 ( .A(n26806), .B(n26807), .Z(n26805) );
  XNOR U26710 ( .A(n26804), .B(n26808), .Z(n26806) );
  XNOR U26711 ( .A(n26760), .B(n26751), .Z(n26791) );
  XOR U26712 ( .A(n26809), .B(n26810), .Z(n26751) );
  AND U26713 ( .A(n26811), .B(n26812), .Z(n26810) );
  XOR U26714 ( .A(n26809), .B(n26813), .Z(n26811) );
  XOR U26715 ( .A(n26814), .B(n26766), .Z(n26760) );
  XOR U26716 ( .A(n26815), .B(n26816), .Z(n26766) );
  NOR U26717 ( .A(n26817), .B(n26818), .Z(n26816) );
  XOR U26718 ( .A(n26815), .B(n26819), .Z(n26817) );
  XNOR U26719 ( .A(n26765), .B(n26757), .Z(n26814) );
  XOR U26720 ( .A(n26820), .B(n26821), .Z(n26757) );
  AND U26721 ( .A(n26822), .B(n26823), .Z(n26821) );
  XOR U26722 ( .A(n26820), .B(n26824), .Z(n26822) );
  XNOR U26723 ( .A(n26825), .B(n26762), .Z(n26765) );
  XOR U26724 ( .A(n26826), .B(n26827), .Z(n26762) );
  AND U26725 ( .A(n26828), .B(n26829), .Z(n26827) );
  XNOR U26726 ( .A(n26830), .B(n26831), .Z(n26828) );
  IV U26727 ( .A(n26826), .Z(n26830) );
  XNOR U26728 ( .A(n26832), .B(n26833), .Z(n26825) );
  NOR U26729 ( .A(n26834), .B(n26835), .Z(n26833) );
  XNOR U26730 ( .A(n26832), .B(n26836), .Z(n26834) );
  XOR U26731 ( .A(n26755), .B(n26767), .Z(n26790) );
  NOR U26732 ( .A(n26693), .B(n26837), .Z(n26767) );
  XNOR U26733 ( .A(n26773), .B(n26772), .Z(n26755) );
  XNOR U26734 ( .A(n26838), .B(n26778), .Z(n26772) );
  XNOR U26735 ( .A(n26839), .B(n26840), .Z(n26778) );
  NOR U26736 ( .A(n26841), .B(n26842), .Z(n26840) );
  XOR U26737 ( .A(n26839), .B(n26843), .Z(n26841) );
  XNOR U26738 ( .A(n26777), .B(n26769), .Z(n26838) );
  XOR U26739 ( .A(n26844), .B(n26845), .Z(n26769) );
  AND U26740 ( .A(n26846), .B(n26847), .Z(n26845) );
  XOR U26741 ( .A(n26844), .B(n26848), .Z(n26846) );
  XNOR U26742 ( .A(n26849), .B(n26774), .Z(n26777) );
  XOR U26743 ( .A(n26850), .B(n26851), .Z(n26774) );
  AND U26744 ( .A(n26852), .B(n26853), .Z(n26851) );
  XNOR U26745 ( .A(n26854), .B(n26855), .Z(n26852) );
  IV U26746 ( .A(n26850), .Z(n26854) );
  XNOR U26747 ( .A(n26856), .B(n26857), .Z(n26849) );
  NOR U26748 ( .A(n26858), .B(n26859), .Z(n26857) );
  XNOR U26749 ( .A(n26856), .B(n26860), .Z(n26858) );
  XOR U26750 ( .A(n26783), .B(n26782), .Z(n26773) );
  XNOR U26751 ( .A(n26861), .B(n26779), .Z(n26782) );
  XOR U26752 ( .A(n26862), .B(n26863), .Z(n26779) );
  AND U26753 ( .A(n26864), .B(n26865), .Z(n26863) );
  XNOR U26754 ( .A(n26866), .B(n26867), .Z(n26864) );
  IV U26755 ( .A(n26862), .Z(n26866) );
  XNOR U26756 ( .A(n26868), .B(n26869), .Z(n26861) );
  NOR U26757 ( .A(n26870), .B(n26871), .Z(n26869) );
  XNOR U26758 ( .A(n26868), .B(n26872), .Z(n26870) );
  XOR U26759 ( .A(n26873), .B(n26874), .Z(n26783) );
  NOR U26760 ( .A(n26875), .B(n26876), .Z(n26874) );
  XNOR U26761 ( .A(n26873), .B(n26877), .Z(n26875) );
  XNOR U26762 ( .A(n26682), .B(n26786), .Z(n26788) );
  XNOR U26763 ( .A(n26878), .B(n26879), .Z(n26682) );
  AND U26764 ( .A(n474), .B(n26689), .Z(n26879) );
  XOR U26765 ( .A(n26878), .B(n26687), .Z(n26689) );
  AND U26766 ( .A(n26690), .B(n26693), .Z(n26786) );
  XOR U26767 ( .A(n26880), .B(n26837), .Z(n26693) );
  XNOR U26768 ( .A(p_input[1184]), .B(p_input[2048]), .Z(n26837) );
  XNOR U26769 ( .A(n26813), .B(n26812), .Z(n26880) );
  XNOR U26770 ( .A(n26881), .B(n26824), .Z(n26812) );
  XOR U26771 ( .A(n26798), .B(n26796), .Z(n26824) );
  XNOR U26772 ( .A(n26882), .B(n26803), .Z(n26796) );
  XOR U26773 ( .A(p_input[1208]), .B(p_input[2072]), .Z(n26803) );
  XOR U26774 ( .A(n26793), .B(n26802), .Z(n26882) );
  XOR U26775 ( .A(n26883), .B(n26799), .Z(n26802) );
  XOR U26776 ( .A(p_input[1206]), .B(p_input[2070]), .Z(n26799) );
  XOR U26777 ( .A(p_input[1207]), .B(n17295), .Z(n26883) );
  XOR U26778 ( .A(p_input[1202]), .B(p_input[2066]), .Z(n26793) );
  XNOR U26779 ( .A(n26808), .B(n26807), .Z(n26798) );
  XOR U26780 ( .A(n26884), .B(n26804), .Z(n26807) );
  XOR U26781 ( .A(p_input[1203]), .B(p_input[2067]), .Z(n26804) );
  XOR U26782 ( .A(p_input[1204]), .B(n17297), .Z(n26884) );
  XOR U26783 ( .A(p_input[1205]), .B(p_input[2069]), .Z(n26808) );
  XOR U26784 ( .A(n26823), .B(n26885), .Z(n26881) );
  IV U26785 ( .A(n26809), .Z(n26885) );
  XOR U26786 ( .A(p_input[1185]), .B(p_input[2049]), .Z(n26809) );
  XNOR U26787 ( .A(n26886), .B(n26831), .Z(n26823) );
  XNOR U26788 ( .A(n26819), .B(n26818), .Z(n26831) );
  XNOR U26789 ( .A(n26887), .B(n26815), .Z(n26818) );
  XNOR U26790 ( .A(p_input[1210]), .B(p_input[2074]), .Z(n26815) );
  XOR U26791 ( .A(p_input[1211]), .B(n17300), .Z(n26887) );
  XOR U26792 ( .A(p_input[1212]), .B(p_input[2076]), .Z(n26819) );
  XOR U26793 ( .A(n26829), .B(n26888), .Z(n26886) );
  IV U26794 ( .A(n26820), .Z(n26888) );
  XOR U26795 ( .A(p_input[1201]), .B(p_input[2065]), .Z(n26820) );
  XNOR U26796 ( .A(n26889), .B(n26836), .Z(n26829) );
  XNOR U26797 ( .A(p_input[1215]), .B(n17303), .Z(n26836) );
  XOR U26798 ( .A(n26826), .B(n26835), .Z(n26889) );
  XOR U26799 ( .A(n26890), .B(n26832), .Z(n26835) );
  XOR U26800 ( .A(p_input[1213]), .B(p_input[2077]), .Z(n26832) );
  XOR U26801 ( .A(p_input[1214]), .B(n17305), .Z(n26890) );
  XOR U26802 ( .A(p_input[1209]), .B(p_input[2073]), .Z(n26826) );
  XOR U26803 ( .A(n26848), .B(n26847), .Z(n26813) );
  XNOR U26804 ( .A(n26891), .B(n26855), .Z(n26847) );
  XNOR U26805 ( .A(n26843), .B(n26842), .Z(n26855) );
  XNOR U26806 ( .A(n26892), .B(n26839), .Z(n26842) );
  XNOR U26807 ( .A(p_input[1195]), .B(p_input[2059]), .Z(n26839) );
  XOR U26808 ( .A(p_input[1196]), .B(n16451), .Z(n26892) );
  XOR U26809 ( .A(p_input[1197]), .B(p_input[2061]), .Z(n26843) );
  XOR U26810 ( .A(n26853), .B(n26893), .Z(n26891) );
  IV U26811 ( .A(n26844), .Z(n26893) );
  XOR U26812 ( .A(p_input[1186]), .B(p_input[2050]), .Z(n26844) );
  XNOR U26813 ( .A(n26894), .B(n26860), .Z(n26853) );
  XNOR U26814 ( .A(p_input[1200]), .B(n16454), .Z(n26860) );
  XOR U26815 ( .A(n26850), .B(n26859), .Z(n26894) );
  XOR U26816 ( .A(n26895), .B(n26856), .Z(n26859) );
  XOR U26817 ( .A(p_input[1198]), .B(p_input[2062]), .Z(n26856) );
  XOR U26818 ( .A(p_input[1199]), .B(n16456), .Z(n26895) );
  XOR U26819 ( .A(p_input[1194]), .B(p_input[2058]), .Z(n26850) );
  XOR U26820 ( .A(n26867), .B(n26865), .Z(n26848) );
  XNOR U26821 ( .A(n26896), .B(n26872), .Z(n26865) );
  XOR U26822 ( .A(p_input[1193]), .B(p_input[2057]), .Z(n26872) );
  XOR U26823 ( .A(n26862), .B(n26871), .Z(n26896) );
  XOR U26824 ( .A(n26897), .B(n26868), .Z(n26871) );
  XOR U26825 ( .A(p_input[1191]), .B(p_input[2055]), .Z(n26868) );
  XOR U26826 ( .A(p_input[1192]), .B(n17312), .Z(n26897) );
  XOR U26827 ( .A(p_input[1187]), .B(p_input[2051]), .Z(n26862) );
  XNOR U26828 ( .A(n26877), .B(n26876), .Z(n26867) );
  XOR U26829 ( .A(n26898), .B(n26873), .Z(n26876) );
  XOR U26830 ( .A(p_input[1188]), .B(p_input[2052]), .Z(n26873) );
  XOR U26831 ( .A(p_input[1189]), .B(n17314), .Z(n26898) );
  XOR U26832 ( .A(p_input[1190]), .B(p_input[2054]), .Z(n26877) );
  XNOR U26833 ( .A(n26899), .B(n26900), .Z(n26690) );
  AND U26834 ( .A(n474), .B(n26901), .Z(n26900) );
  XNOR U26835 ( .A(n26902), .B(n26903), .Z(n474) );
  AND U26836 ( .A(n26904), .B(n26905), .Z(n26903) );
  XOR U26837 ( .A(n26902), .B(n26700), .Z(n26905) );
  XNOR U26838 ( .A(n26902), .B(n26642), .Z(n26904) );
  XOR U26839 ( .A(n26906), .B(n26907), .Z(n26902) );
  AND U26840 ( .A(n26908), .B(n26909), .Z(n26907) );
  XNOR U26841 ( .A(n26713), .B(n26906), .Z(n26909) );
  XOR U26842 ( .A(n26906), .B(n26654), .Z(n26908) );
  XOR U26843 ( .A(n26910), .B(n26911), .Z(n26906) );
  AND U26844 ( .A(n26912), .B(n26913), .Z(n26911) );
  XNOR U26845 ( .A(n26738), .B(n26910), .Z(n26913) );
  XOR U26846 ( .A(n26910), .B(n26665), .Z(n26912) );
  XOR U26847 ( .A(n26914), .B(n26915), .Z(n26910) );
  AND U26848 ( .A(n26916), .B(n26917), .Z(n26915) );
  XOR U26849 ( .A(n26914), .B(n26675), .Z(n26916) );
  XOR U26850 ( .A(n26918), .B(n26919), .Z(n26631) );
  AND U26851 ( .A(n478), .B(n26901), .Z(n26919) );
  XNOR U26852 ( .A(n26899), .B(n26918), .Z(n26901) );
  XNOR U26853 ( .A(n26920), .B(n26921), .Z(n478) );
  AND U26854 ( .A(n26922), .B(n26923), .Z(n26921) );
  XNOR U26855 ( .A(n26924), .B(n26920), .Z(n26923) );
  IV U26856 ( .A(n26700), .Z(n26924) );
  XNOR U26857 ( .A(n26925), .B(n26926), .Z(n26700) );
  AND U26858 ( .A(n481), .B(n26927), .Z(n26926) );
  XNOR U26859 ( .A(n26925), .B(n26928), .Z(n26927) );
  XNOR U26860 ( .A(n26642), .B(n26920), .Z(n26922) );
  XOR U26861 ( .A(n26929), .B(n26930), .Z(n26642) );
  AND U26862 ( .A(n489), .B(n26931), .Z(n26930) );
  XOR U26863 ( .A(n26932), .B(n26933), .Z(n26920) );
  AND U26864 ( .A(n26934), .B(n26935), .Z(n26933) );
  XNOR U26865 ( .A(n26932), .B(n26713), .Z(n26935) );
  XNOR U26866 ( .A(n26936), .B(n26937), .Z(n26713) );
  AND U26867 ( .A(n481), .B(n26938), .Z(n26937) );
  XOR U26868 ( .A(n26939), .B(n26936), .Z(n26938) );
  XNOR U26869 ( .A(n26940), .B(n26932), .Z(n26934) );
  IV U26870 ( .A(n26654), .Z(n26940) );
  XOR U26871 ( .A(n26941), .B(n26942), .Z(n26654) );
  AND U26872 ( .A(n489), .B(n26943), .Z(n26942) );
  XOR U26873 ( .A(n26944), .B(n26945), .Z(n26932) );
  AND U26874 ( .A(n26946), .B(n26947), .Z(n26945) );
  XNOR U26875 ( .A(n26944), .B(n26738), .Z(n26947) );
  XNOR U26876 ( .A(n26948), .B(n26949), .Z(n26738) );
  AND U26877 ( .A(n481), .B(n26950), .Z(n26949) );
  XNOR U26878 ( .A(n26951), .B(n26948), .Z(n26950) );
  XOR U26879 ( .A(n26665), .B(n26944), .Z(n26946) );
  XOR U26880 ( .A(n26952), .B(n26953), .Z(n26665) );
  AND U26881 ( .A(n489), .B(n26954), .Z(n26953) );
  XOR U26882 ( .A(n26914), .B(n26955), .Z(n26944) );
  AND U26883 ( .A(n26956), .B(n26917), .Z(n26955) );
  XNOR U26884 ( .A(n26784), .B(n26914), .Z(n26917) );
  XNOR U26885 ( .A(n26957), .B(n26958), .Z(n26784) );
  AND U26886 ( .A(n481), .B(n26959), .Z(n26958) );
  XOR U26887 ( .A(n26960), .B(n26957), .Z(n26959) );
  XNOR U26888 ( .A(n26961), .B(n26914), .Z(n26956) );
  IV U26889 ( .A(n26675), .Z(n26961) );
  XOR U26890 ( .A(n26962), .B(n26963), .Z(n26675) );
  AND U26891 ( .A(n489), .B(n26964), .Z(n26963) );
  XOR U26892 ( .A(n26965), .B(n26966), .Z(n26914) );
  AND U26893 ( .A(n26967), .B(n26968), .Z(n26966) );
  XNOR U26894 ( .A(n26965), .B(n26878), .Z(n26968) );
  XNOR U26895 ( .A(n26969), .B(n26970), .Z(n26878) );
  AND U26896 ( .A(n481), .B(n26971), .Z(n26970) );
  XNOR U26897 ( .A(n26972), .B(n26969), .Z(n26971) );
  XNOR U26898 ( .A(n26973), .B(n26965), .Z(n26967) );
  IV U26899 ( .A(n26687), .Z(n26973) );
  XOR U26900 ( .A(n26974), .B(n26975), .Z(n26687) );
  AND U26901 ( .A(n489), .B(n26976), .Z(n26975) );
  AND U26902 ( .A(n26918), .B(n26899), .Z(n26965) );
  XNOR U26903 ( .A(n26977), .B(n26978), .Z(n26899) );
  AND U26904 ( .A(n481), .B(n26979), .Z(n26978) );
  XNOR U26905 ( .A(n26980), .B(n26977), .Z(n26979) );
  XNOR U26906 ( .A(n26981), .B(n26982), .Z(n481) );
  AND U26907 ( .A(n26983), .B(n26984), .Z(n26982) );
  XOR U26908 ( .A(n26928), .B(n26981), .Z(n26984) );
  AND U26909 ( .A(n26985), .B(n26986), .Z(n26928) );
  XOR U26910 ( .A(n26981), .B(n26925), .Z(n26983) );
  XNOR U26911 ( .A(n26987), .B(n26988), .Z(n26925) );
  AND U26912 ( .A(n485), .B(n26931), .Z(n26988) );
  XOR U26913 ( .A(n26929), .B(n26987), .Z(n26931) );
  XOR U26914 ( .A(n26989), .B(n26990), .Z(n26981) );
  AND U26915 ( .A(n26991), .B(n26992), .Z(n26990) );
  XNOR U26916 ( .A(n26989), .B(n26985), .Z(n26992) );
  IV U26917 ( .A(n26939), .Z(n26985) );
  XOR U26918 ( .A(n26993), .B(n26994), .Z(n26939) );
  XOR U26919 ( .A(n26995), .B(n26986), .Z(n26994) );
  AND U26920 ( .A(n26951), .B(n26996), .Z(n26986) );
  AND U26921 ( .A(n26997), .B(n26998), .Z(n26995) );
  XOR U26922 ( .A(n26999), .B(n26993), .Z(n26997) );
  XNOR U26923 ( .A(n26936), .B(n26989), .Z(n26991) );
  XNOR U26924 ( .A(n27000), .B(n27001), .Z(n26936) );
  AND U26925 ( .A(n485), .B(n26943), .Z(n27001) );
  XOR U26926 ( .A(n27000), .B(n26941), .Z(n26943) );
  XOR U26927 ( .A(n27002), .B(n27003), .Z(n26989) );
  AND U26928 ( .A(n27004), .B(n27005), .Z(n27003) );
  XNOR U26929 ( .A(n27002), .B(n26951), .Z(n27005) );
  XOR U26930 ( .A(n27006), .B(n26998), .Z(n26951) );
  XNOR U26931 ( .A(n27007), .B(n26993), .Z(n26998) );
  XOR U26932 ( .A(n27008), .B(n27009), .Z(n26993) );
  AND U26933 ( .A(n27010), .B(n27011), .Z(n27009) );
  XOR U26934 ( .A(n27012), .B(n27008), .Z(n27010) );
  XNOR U26935 ( .A(n27013), .B(n27014), .Z(n27007) );
  AND U26936 ( .A(n27015), .B(n27016), .Z(n27014) );
  XOR U26937 ( .A(n27013), .B(n27017), .Z(n27015) );
  XNOR U26938 ( .A(n26999), .B(n26996), .Z(n27006) );
  AND U26939 ( .A(n27018), .B(n27019), .Z(n26996) );
  XOR U26940 ( .A(n27020), .B(n27021), .Z(n26999) );
  AND U26941 ( .A(n27022), .B(n27023), .Z(n27021) );
  XOR U26942 ( .A(n27020), .B(n27024), .Z(n27022) );
  XNOR U26943 ( .A(n26948), .B(n27002), .Z(n27004) );
  XNOR U26944 ( .A(n27025), .B(n27026), .Z(n26948) );
  AND U26945 ( .A(n485), .B(n26954), .Z(n27026) );
  XOR U26946 ( .A(n27025), .B(n26952), .Z(n26954) );
  XOR U26947 ( .A(n27027), .B(n27028), .Z(n27002) );
  AND U26948 ( .A(n27029), .B(n27030), .Z(n27028) );
  XNOR U26949 ( .A(n27027), .B(n27018), .Z(n27030) );
  IV U26950 ( .A(n26960), .Z(n27018) );
  XNOR U26951 ( .A(n27031), .B(n27011), .Z(n26960) );
  XNOR U26952 ( .A(n27032), .B(n27017), .Z(n27011) );
  XOR U26953 ( .A(n27033), .B(n27034), .Z(n27017) );
  AND U26954 ( .A(n27035), .B(n27036), .Z(n27034) );
  XOR U26955 ( .A(n27033), .B(n27037), .Z(n27035) );
  XNOR U26956 ( .A(n27016), .B(n27008), .Z(n27032) );
  XOR U26957 ( .A(n27038), .B(n27039), .Z(n27008) );
  AND U26958 ( .A(n27040), .B(n27041), .Z(n27039) );
  XNOR U26959 ( .A(n27042), .B(n27038), .Z(n27040) );
  XNOR U26960 ( .A(n27043), .B(n27013), .Z(n27016) );
  XOR U26961 ( .A(n27044), .B(n27045), .Z(n27013) );
  AND U26962 ( .A(n27046), .B(n27047), .Z(n27045) );
  XOR U26963 ( .A(n27044), .B(n27048), .Z(n27046) );
  XNOR U26964 ( .A(n27049), .B(n27050), .Z(n27043) );
  AND U26965 ( .A(n27051), .B(n27052), .Z(n27050) );
  XNOR U26966 ( .A(n27049), .B(n27053), .Z(n27051) );
  XNOR U26967 ( .A(n27012), .B(n27019), .Z(n27031) );
  AND U26968 ( .A(n26972), .B(n27054), .Z(n27019) );
  XOR U26969 ( .A(n27024), .B(n27023), .Z(n27012) );
  XNOR U26970 ( .A(n27055), .B(n27020), .Z(n27023) );
  XOR U26971 ( .A(n27056), .B(n27057), .Z(n27020) );
  AND U26972 ( .A(n27058), .B(n27059), .Z(n27057) );
  XOR U26973 ( .A(n27056), .B(n27060), .Z(n27058) );
  XNOR U26974 ( .A(n27061), .B(n27062), .Z(n27055) );
  AND U26975 ( .A(n27063), .B(n27064), .Z(n27062) );
  XOR U26976 ( .A(n27061), .B(n27065), .Z(n27063) );
  XOR U26977 ( .A(n27066), .B(n27067), .Z(n27024) );
  AND U26978 ( .A(n27068), .B(n27069), .Z(n27067) );
  XOR U26979 ( .A(n27066), .B(n27070), .Z(n27068) );
  XNOR U26980 ( .A(n26957), .B(n27027), .Z(n27029) );
  XNOR U26981 ( .A(n27071), .B(n27072), .Z(n26957) );
  AND U26982 ( .A(n485), .B(n26964), .Z(n27072) );
  XOR U26983 ( .A(n27071), .B(n26962), .Z(n26964) );
  XOR U26984 ( .A(n27073), .B(n27074), .Z(n27027) );
  AND U26985 ( .A(n27075), .B(n27076), .Z(n27074) );
  XNOR U26986 ( .A(n27073), .B(n26972), .Z(n27076) );
  XOR U26987 ( .A(n27077), .B(n27041), .Z(n26972) );
  XNOR U26988 ( .A(n27078), .B(n27048), .Z(n27041) );
  XOR U26989 ( .A(n27037), .B(n27036), .Z(n27048) );
  XNOR U26990 ( .A(n27079), .B(n27033), .Z(n27036) );
  XOR U26991 ( .A(n27080), .B(n27081), .Z(n27033) );
  AND U26992 ( .A(n27082), .B(n27083), .Z(n27081) );
  XNOR U26993 ( .A(n27084), .B(n27085), .Z(n27082) );
  IV U26994 ( .A(n27080), .Z(n27084) );
  XNOR U26995 ( .A(n27086), .B(n27087), .Z(n27079) );
  NOR U26996 ( .A(n27088), .B(n27089), .Z(n27087) );
  XNOR U26997 ( .A(n27086), .B(n27090), .Z(n27088) );
  XOR U26998 ( .A(n27091), .B(n27092), .Z(n27037) );
  NOR U26999 ( .A(n27093), .B(n27094), .Z(n27092) );
  XNOR U27000 ( .A(n27091), .B(n27095), .Z(n27093) );
  XNOR U27001 ( .A(n27047), .B(n27038), .Z(n27078) );
  XOR U27002 ( .A(n27096), .B(n27097), .Z(n27038) );
  AND U27003 ( .A(n27098), .B(n27099), .Z(n27097) );
  XOR U27004 ( .A(n27096), .B(n27100), .Z(n27098) );
  XOR U27005 ( .A(n27101), .B(n27053), .Z(n27047) );
  XOR U27006 ( .A(n27102), .B(n27103), .Z(n27053) );
  NOR U27007 ( .A(n27104), .B(n27105), .Z(n27103) );
  XOR U27008 ( .A(n27102), .B(n27106), .Z(n27104) );
  XNOR U27009 ( .A(n27052), .B(n27044), .Z(n27101) );
  XOR U27010 ( .A(n27107), .B(n27108), .Z(n27044) );
  AND U27011 ( .A(n27109), .B(n27110), .Z(n27108) );
  XOR U27012 ( .A(n27107), .B(n27111), .Z(n27109) );
  XNOR U27013 ( .A(n27112), .B(n27049), .Z(n27052) );
  XOR U27014 ( .A(n27113), .B(n27114), .Z(n27049) );
  AND U27015 ( .A(n27115), .B(n27116), .Z(n27114) );
  XNOR U27016 ( .A(n27117), .B(n27118), .Z(n27115) );
  IV U27017 ( .A(n27113), .Z(n27117) );
  XNOR U27018 ( .A(n27119), .B(n27120), .Z(n27112) );
  NOR U27019 ( .A(n27121), .B(n27122), .Z(n27120) );
  XNOR U27020 ( .A(n27119), .B(n27123), .Z(n27121) );
  XOR U27021 ( .A(n27042), .B(n27054), .Z(n27077) );
  NOR U27022 ( .A(n26980), .B(n27124), .Z(n27054) );
  XNOR U27023 ( .A(n27060), .B(n27059), .Z(n27042) );
  XNOR U27024 ( .A(n27125), .B(n27065), .Z(n27059) );
  XNOR U27025 ( .A(n27126), .B(n27127), .Z(n27065) );
  NOR U27026 ( .A(n27128), .B(n27129), .Z(n27127) );
  XOR U27027 ( .A(n27126), .B(n27130), .Z(n27128) );
  XNOR U27028 ( .A(n27064), .B(n27056), .Z(n27125) );
  XOR U27029 ( .A(n27131), .B(n27132), .Z(n27056) );
  AND U27030 ( .A(n27133), .B(n27134), .Z(n27132) );
  XOR U27031 ( .A(n27131), .B(n27135), .Z(n27133) );
  XNOR U27032 ( .A(n27136), .B(n27061), .Z(n27064) );
  XOR U27033 ( .A(n27137), .B(n27138), .Z(n27061) );
  AND U27034 ( .A(n27139), .B(n27140), .Z(n27138) );
  XNOR U27035 ( .A(n27141), .B(n27142), .Z(n27139) );
  IV U27036 ( .A(n27137), .Z(n27141) );
  XNOR U27037 ( .A(n27143), .B(n27144), .Z(n27136) );
  NOR U27038 ( .A(n27145), .B(n27146), .Z(n27144) );
  XNOR U27039 ( .A(n27143), .B(n27147), .Z(n27145) );
  XOR U27040 ( .A(n27070), .B(n27069), .Z(n27060) );
  XNOR U27041 ( .A(n27148), .B(n27066), .Z(n27069) );
  XOR U27042 ( .A(n27149), .B(n27150), .Z(n27066) );
  AND U27043 ( .A(n27151), .B(n27152), .Z(n27150) );
  XNOR U27044 ( .A(n27153), .B(n27154), .Z(n27151) );
  IV U27045 ( .A(n27149), .Z(n27153) );
  XNOR U27046 ( .A(n27155), .B(n27156), .Z(n27148) );
  NOR U27047 ( .A(n27157), .B(n27158), .Z(n27156) );
  XNOR U27048 ( .A(n27155), .B(n27159), .Z(n27157) );
  XOR U27049 ( .A(n27160), .B(n27161), .Z(n27070) );
  NOR U27050 ( .A(n27162), .B(n27163), .Z(n27161) );
  XNOR U27051 ( .A(n27160), .B(n27164), .Z(n27162) );
  XNOR U27052 ( .A(n26969), .B(n27073), .Z(n27075) );
  XNOR U27053 ( .A(n27165), .B(n27166), .Z(n26969) );
  AND U27054 ( .A(n485), .B(n26976), .Z(n27166) );
  XOR U27055 ( .A(n27165), .B(n26974), .Z(n26976) );
  AND U27056 ( .A(n26977), .B(n26980), .Z(n27073) );
  XOR U27057 ( .A(n27167), .B(n27124), .Z(n26980) );
  XNOR U27058 ( .A(p_input[1216]), .B(p_input[2048]), .Z(n27124) );
  XNOR U27059 ( .A(n27100), .B(n27099), .Z(n27167) );
  XNOR U27060 ( .A(n27168), .B(n27111), .Z(n27099) );
  XOR U27061 ( .A(n27085), .B(n27083), .Z(n27111) );
  XNOR U27062 ( .A(n27169), .B(n27090), .Z(n27083) );
  XOR U27063 ( .A(p_input[1240]), .B(p_input[2072]), .Z(n27090) );
  XOR U27064 ( .A(n27080), .B(n27089), .Z(n27169) );
  XOR U27065 ( .A(n27170), .B(n27086), .Z(n27089) );
  XOR U27066 ( .A(p_input[1238]), .B(p_input[2070]), .Z(n27086) );
  XOR U27067 ( .A(p_input[1239]), .B(n17295), .Z(n27170) );
  XOR U27068 ( .A(p_input[1234]), .B(p_input[2066]), .Z(n27080) );
  XNOR U27069 ( .A(n27095), .B(n27094), .Z(n27085) );
  XOR U27070 ( .A(n27171), .B(n27091), .Z(n27094) );
  XOR U27071 ( .A(p_input[1235]), .B(p_input[2067]), .Z(n27091) );
  XOR U27072 ( .A(p_input[1236]), .B(n17297), .Z(n27171) );
  XOR U27073 ( .A(p_input[1237]), .B(p_input[2069]), .Z(n27095) );
  XOR U27074 ( .A(n27110), .B(n27172), .Z(n27168) );
  IV U27075 ( .A(n27096), .Z(n27172) );
  XOR U27076 ( .A(p_input[1217]), .B(p_input[2049]), .Z(n27096) );
  XNOR U27077 ( .A(n27173), .B(n27118), .Z(n27110) );
  XNOR U27078 ( .A(n27106), .B(n27105), .Z(n27118) );
  XNOR U27079 ( .A(n27174), .B(n27102), .Z(n27105) );
  XNOR U27080 ( .A(p_input[1242]), .B(p_input[2074]), .Z(n27102) );
  XOR U27081 ( .A(p_input[1243]), .B(n17300), .Z(n27174) );
  XOR U27082 ( .A(p_input[1244]), .B(p_input[2076]), .Z(n27106) );
  XOR U27083 ( .A(n27116), .B(n27175), .Z(n27173) );
  IV U27084 ( .A(n27107), .Z(n27175) );
  XOR U27085 ( .A(p_input[1233]), .B(p_input[2065]), .Z(n27107) );
  XNOR U27086 ( .A(n27176), .B(n27123), .Z(n27116) );
  XNOR U27087 ( .A(p_input[1247]), .B(n17303), .Z(n27123) );
  XOR U27088 ( .A(n27113), .B(n27122), .Z(n27176) );
  XOR U27089 ( .A(n27177), .B(n27119), .Z(n27122) );
  XOR U27090 ( .A(p_input[1245]), .B(p_input[2077]), .Z(n27119) );
  XOR U27091 ( .A(p_input[1246]), .B(n17305), .Z(n27177) );
  XOR U27092 ( .A(p_input[1241]), .B(p_input[2073]), .Z(n27113) );
  XOR U27093 ( .A(n27135), .B(n27134), .Z(n27100) );
  XNOR U27094 ( .A(n27178), .B(n27142), .Z(n27134) );
  XNOR U27095 ( .A(n27130), .B(n27129), .Z(n27142) );
  XNOR U27096 ( .A(n27179), .B(n27126), .Z(n27129) );
  XNOR U27097 ( .A(p_input[1227]), .B(p_input[2059]), .Z(n27126) );
  XOR U27098 ( .A(p_input[1228]), .B(n16451), .Z(n27179) );
  XOR U27099 ( .A(p_input[1229]), .B(p_input[2061]), .Z(n27130) );
  XOR U27100 ( .A(n27140), .B(n27180), .Z(n27178) );
  IV U27101 ( .A(n27131), .Z(n27180) );
  XOR U27102 ( .A(p_input[1218]), .B(p_input[2050]), .Z(n27131) );
  XNOR U27103 ( .A(n27181), .B(n27147), .Z(n27140) );
  XNOR U27104 ( .A(p_input[1232]), .B(n16454), .Z(n27147) );
  XOR U27105 ( .A(n27137), .B(n27146), .Z(n27181) );
  XOR U27106 ( .A(n27182), .B(n27143), .Z(n27146) );
  XOR U27107 ( .A(p_input[1230]), .B(p_input[2062]), .Z(n27143) );
  XOR U27108 ( .A(p_input[1231]), .B(n16456), .Z(n27182) );
  XOR U27109 ( .A(p_input[1226]), .B(p_input[2058]), .Z(n27137) );
  XOR U27110 ( .A(n27154), .B(n27152), .Z(n27135) );
  XNOR U27111 ( .A(n27183), .B(n27159), .Z(n27152) );
  XOR U27112 ( .A(p_input[1225]), .B(p_input[2057]), .Z(n27159) );
  XOR U27113 ( .A(n27149), .B(n27158), .Z(n27183) );
  XOR U27114 ( .A(n27184), .B(n27155), .Z(n27158) );
  XOR U27115 ( .A(p_input[1223]), .B(p_input[2055]), .Z(n27155) );
  XOR U27116 ( .A(p_input[1224]), .B(n17312), .Z(n27184) );
  XOR U27117 ( .A(p_input[1219]), .B(p_input[2051]), .Z(n27149) );
  XNOR U27118 ( .A(n27164), .B(n27163), .Z(n27154) );
  XOR U27119 ( .A(n27185), .B(n27160), .Z(n27163) );
  XOR U27120 ( .A(p_input[1220]), .B(p_input[2052]), .Z(n27160) );
  XOR U27121 ( .A(p_input[1221]), .B(n17314), .Z(n27185) );
  XOR U27122 ( .A(p_input[1222]), .B(p_input[2054]), .Z(n27164) );
  XNOR U27123 ( .A(n27186), .B(n27187), .Z(n26977) );
  AND U27124 ( .A(n485), .B(n27188), .Z(n27187) );
  XNOR U27125 ( .A(n27189), .B(n27190), .Z(n485) );
  AND U27126 ( .A(n27191), .B(n27192), .Z(n27190) );
  XOR U27127 ( .A(n27189), .B(n26987), .Z(n27192) );
  XNOR U27128 ( .A(n27189), .B(n26929), .Z(n27191) );
  XOR U27129 ( .A(n27193), .B(n27194), .Z(n27189) );
  AND U27130 ( .A(n27195), .B(n27196), .Z(n27194) );
  XNOR U27131 ( .A(n27000), .B(n27193), .Z(n27196) );
  XOR U27132 ( .A(n27193), .B(n26941), .Z(n27195) );
  XOR U27133 ( .A(n27197), .B(n27198), .Z(n27193) );
  AND U27134 ( .A(n27199), .B(n27200), .Z(n27198) );
  XNOR U27135 ( .A(n27025), .B(n27197), .Z(n27200) );
  XOR U27136 ( .A(n27197), .B(n26952), .Z(n27199) );
  XOR U27137 ( .A(n27201), .B(n27202), .Z(n27197) );
  AND U27138 ( .A(n27203), .B(n27204), .Z(n27202) );
  XOR U27139 ( .A(n27201), .B(n26962), .Z(n27203) );
  XOR U27140 ( .A(n27205), .B(n27206), .Z(n26918) );
  AND U27141 ( .A(n489), .B(n27188), .Z(n27206) );
  XNOR U27142 ( .A(n27186), .B(n27205), .Z(n27188) );
  XNOR U27143 ( .A(n27207), .B(n27208), .Z(n489) );
  AND U27144 ( .A(n27209), .B(n27210), .Z(n27208) );
  XNOR U27145 ( .A(n27211), .B(n27207), .Z(n27210) );
  IV U27146 ( .A(n26987), .Z(n27211) );
  XNOR U27147 ( .A(n27212), .B(n27213), .Z(n26987) );
  AND U27148 ( .A(n492), .B(n27214), .Z(n27213) );
  XNOR U27149 ( .A(n27212), .B(n27215), .Z(n27214) );
  XNOR U27150 ( .A(n26929), .B(n27207), .Z(n27209) );
  XOR U27151 ( .A(n27216), .B(n27217), .Z(n26929) );
  AND U27152 ( .A(n500), .B(n27218), .Z(n27217) );
  XOR U27153 ( .A(n27219), .B(n27220), .Z(n27207) );
  AND U27154 ( .A(n27221), .B(n27222), .Z(n27220) );
  XNOR U27155 ( .A(n27219), .B(n27000), .Z(n27222) );
  XNOR U27156 ( .A(n27223), .B(n27224), .Z(n27000) );
  AND U27157 ( .A(n492), .B(n27225), .Z(n27224) );
  XOR U27158 ( .A(n27226), .B(n27223), .Z(n27225) );
  XNOR U27159 ( .A(n27227), .B(n27219), .Z(n27221) );
  IV U27160 ( .A(n26941), .Z(n27227) );
  XOR U27161 ( .A(n27228), .B(n27229), .Z(n26941) );
  AND U27162 ( .A(n500), .B(n27230), .Z(n27229) );
  XOR U27163 ( .A(n27231), .B(n27232), .Z(n27219) );
  AND U27164 ( .A(n27233), .B(n27234), .Z(n27232) );
  XNOR U27165 ( .A(n27231), .B(n27025), .Z(n27234) );
  XNOR U27166 ( .A(n27235), .B(n27236), .Z(n27025) );
  AND U27167 ( .A(n492), .B(n27237), .Z(n27236) );
  XNOR U27168 ( .A(n27238), .B(n27235), .Z(n27237) );
  XOR U27169 ( .A(n26952), .B(n27231), .Z(n27233) );
  XOR U27170 ( .A(n27239), .B(n27240), .Z(n26952) );
  AND U27171 ( .A(n500), .B(n27241), .Z(n27240) );
  XOR U27172 ( .A(n27201), .B(n27242), .Z(n27231) );
  AND U27173 ( .A(n27243), .B(n27204), .Z(n27242) );
  XNOR U27174 ( .A(n27071), .B(n27201), .Z(n27204) );
  XNOR U27175 ( .A(n27244), .B(n27245), .Z(n27071) );
  AND U27176 ( .A(n492), .B(n27246), .Z(n27245) );
  XOR U27177 ( .A(n27247), .B(n27244), .Z(n27246) );
  XNOR U27178 ( .A(n27248), .B(n27201), .Z(n27243) );
  IV U27179 ( .A(n26962), .Z(n27248) );
  XOR U27180 ( .A(n27249), .B(n27250), .Z(n26962) );
  AND U27181 ( .A(n500), .B(n27251), .Z(n27250) );
  XOR U27182 ( .A(n27252), .B(n27253), .Z(n27201) );
  AND U27183 ( .A(n27254), .B(n27255), .Z(n27253) );
  XNOR U27184 ( .A(n27252), .B(n27165), .Z(n27255) );
  XNOR U27185 ( .A(n27256), .B(n27257), .Z(n27165) );
  AND U27186 ( .A(n492), .B(n27258), .Z(n27257) );
  XNOR U27187 ( .A(n27259), .B(n27256), .Z(n27258) );
  XNOR U27188 ( .A(n27260), .B(n27252), .Z(n27254) );
  IV U27189 ( .A(n26974), .Z(n27260) );
  XOR U27190 ( .A(n27261), .B(n27262), .Z(n26974) );
  AND U27191 ( .A(n500), .B(n27263), .Z(n27262) );
  AND U27192 ( .A(n27205), .B(n27186), .Z(n27252) );
  XNOR U27193 ( .A(n27264), .B(n27265), .Z(n27186) );
  AND U27194 ( .A(n492), .B(n27266), .Z(n27265) );
  XNOR U27195 ( .A(n27267), .B(n27264), .Z(n27266) );
  XNOR U27196 ( .A(n27268), .B(n27269), .Z(n492) );
  AND U27197 ( .A(n27270), .B(n27271), .Z(n27269) );
  XOR U27198 ( .A(n27215), .B(n27268), .Z(n27271) );
  AND U27199 ( .A(n27272), .B(n27273), .Z(n27215) );
  XOR U27200 ( .A(n27268), .B(n27212), .Z(n27270) );
  XNOR U27201 ( .A(n27274), .B(n27275), .Z(n27212) );
  AND U27202 ( .A(n496), .B(n27218), .Z(n27275) );
  XOR U27203 ( .A(n27216), .B(n27274), .Z(n27218) );
  XOR U27204 ( .A(n27276), .B(n27277), .Z(n27268) );
  AND U27205 ( .A(n27278), .B(n27279), .Z(n27277) );
  XNOR U27206 ( .A(n27276), .B(n27272), .Z(n27279) );
  IV U27207 ( .A(n27226), .Z(n27272) );
  XOR U27208 ( .A(n27280), .B(n27281), .Z(n27226) );
  XOR U27209 ( .A(n27282), .B(n27273), .Z(n27281) );
  AND U27210 ( .A(n27238), .B(n27283), .Z(n27273) );
  AND U27211 ( .A(n27284), .B(n27285), .Z(n27282) );
  XOR U27212 ( .A(n27286), .B(n27280), .Z(n27284) );
  XNOR U27213 ( .A(n27223), .B(n27276), .Z(n27278) );
  XNOR U27214 ( .A(n27287), .B(n27288), .Z(n27223) );
  AND U27215 ( .A(n496), .B(n27230), .Z(n27288) );
  XOR U27216 ( .A(n27287), .B(n27228), .Z(n27230) );
  XOR U27217 ( .A(n27289), .B(n27290), .Z(n27276) );
  AND U27218 ( .A(n27291), .B(n27292), .Z(n27290) );
  XNOR U27219 ( .A(n27289), .B(n27238), .Z(n27292) );
  XOR U27220 ( .A(n27293), .B(n27285), .Z(n27238) );
  XNOR U27221 ( .A(n27294), .B(n27280), .Z(n27285) );
  XOR U27222 ( .A(n27295), .B(n27296), .Z(n27280) );
  AND U27223 ( .A(n27297), .B(n27298), .Z(n27296) );
  XOR U27224 ( .A(n27299), .B(n27295), .Z(n27297) );
  XNOR U27225 ( .A(n27300), .B(n27301), .Z(n27294) );
  AND U27226 ( .A(n27302), .B(n27303), .Z(n27301) );
  XOR U27227 ( .A(n27300), .B(n27304), .Z(n27302) );
  XNOR U27228 ( .A(n27286), .B(n27283), .Z(n27293) );
  AND U27229 ( .A(n27305), .B(n27306), .Z(n27283) );
  XOR U27230 ( .A(n27307), .B(n27308), .Z(n27286) );
  AND U27231 ( .A(n27309), .B(n27310), .Z(n27308) );
  XOR U27232 ( .A(n27307), .B(n27311), .Z(n27309) );
  XNOR U27233 ( .A(n27235), .B(n27289), .Z(n27291) );
  XNOR U27234 ( .A(n27312), .B(n27313), .Z(n27235) );
  AND U27235 ( .A(n496), .B(n27241), .Z(n27313) );
  XOR U27236 ( .A(n27312), .B(n27239), .Z(n27241) );
  XOR U27237 ( .A(n27314), .B(n27315), .Z(n27289) );
  AND U27238 ( .A(n27316), .B(n27317), .Z(n27315) );
  XNOR U27239 ( .A(n27314), .B(n27305), .Z(n27317) );
  IV U27240 ( .A(n27247), .Z(n27305) );
  XNOR U27241 ( .A(n27318), .B(n27298), .Z(n27247) );
  XNOR U27242 ( .A(n27319), .B(n27304), .Z(n27298) );
  XOR U27243 ( .A(n27320), .B(n27321), .Z(n27304) );
  AND U27244 ( .A(n27322), .B(n27323), .Z(n27321) );
  XOR U27245 ( .A(n27320), .B(n27324), .Z(n27322) );
  XNOR U27246 ( .A(n27303), .B(n27295), .Z(n27319) );
  XOR U27247 ( .A(n27325), .B(n27326), .Z(n27295) );
  AND U27248 ( .A(n27327), .B(n27328), .Z(n27326) );
  XNOR U27249 ( .A(n27329), .B(n27325), .Z(n27327) );
  XNOR U27250 ( .A(n27330), .B(n27300), .Z(n27303) );
  XOR U27251 ( .A(n27331), .B(n27332), .Z(n27300) );
  AND U27252 ( .A(n27333), .B(n27334), .Z(n27332) );
  XOR U27253 ( .A(n27331), .B(n27335), .Z(n27333) );
  XNOR U27254 ( .A(n27336), .B(n27337), .Z(n27330) );
  AND U27255 ( .A(n27338), .B(n27339), .Z(n27337) );
  XNOR U27256 ( .A(n27336), .B(n27340), .Z(n27338) );
  XNOR U27257 ( .A(n27299), .B(n27306), .Z(n27318) );
  AND U27258 ( .A(n27259), .B(n27341), .Z(n27306) );
  XOR U27259 ( .A(n27311), .B(n27310), .Z(n27299) );
  XNOR U27260 ( .A(n27342), .B(n27307), .Z(n27310) );
  XOR U27261 ( .A(n27343), .B(n27344), .Z(n27307) );
  AND U27262 ( .A(n27345), .B(n27346), .Z(n27344) );
  XOR U27263 ( .A(n27343), .B(n27347), .Z(n27345) );
  XNOR U27264 ( .A(n27348), .B(n27349), .Z(n27342) );
  AND U27265 ( .A(n27350), .B(n27351), .Z(n27349) );
  XOR U27266 ( .A(n27348), .B(n27352), .Z(n27350) );
  XOR U27267 ( .A(n27353), .B(n27354), .Z(n27311) );
  AND U27268 ( .A(n27355), .B(n27356), .Z(n27354) );
  XOR U27269 ( .A(n27353), .B(n27357), .Z(n27355) );
  XNOR U27270 ( .A(n27244), .B(n27314), .Z(n27316) );
  XNOR U27271 ( .A(n27358), .B(n27359), .Z(n27244) );
  AND U27272 ( .A(n496), .B(n27251), .Z(n27359) );
  XOR U27273 ( .A(n27358), .B(n27249), .Z(n27251) );
  XOR U27274 ( .A(n27360), .B(n27361), .Z(n27314) );
  AND U27275 ( .A(n27362), .B(n27363), .Z(n27361) );
  XNOR U27276 ( .A(n27360), .B(n27259), .Z(n27363) );
  XOR U27277 ( .A(n27364), .B(n27328), .Z(n27259) );
  XNOR U27278 ( .A(n27365), .B(n27335), .Z(n27328) );
  XOR U27279 ( .A(n27324), .B(n27323), .Z(n27335) );
  XNOR U27280 ( .A(n27366), .B(n27320), .Z(n27323) );
  XOR U27281 ( .A(n27367), .B(n27368), .Z(n27320) );
  AND U27282 ( .A(n27369), .B(n27370), .Z(n27368) );
  XNOR U27283 ( .A(n27371), .B(n27372), .Z(n27369) );
  IV U27284 ( .A(n27367), .Z(n27371) );
  XNOR U27285 ( .A(n27373), .B(n27374), .Z(n27366) );
  NOR U27286 ( .A(n27375), .B(n27376), .Z(n27374) );
  XNOR U27287 ( .A(n27373), .B(n27377), .Z(n27375) );
  XOR U27288 ( .A(n27378), .B(n27379), .Z(n27324) );
  NOR U27289 ( .A(n27380), .B(n27381), .Z(n27379) );
  XNOR U27290 ( .A(n27378), .B(n27382), .Z(n27380) );
  XNOR U27291 ( .A(n27334), .B(n27325), .Z(n27365) );
  XOR U27292 ( .A(n27383), .B(n27384), .Z(n27325) );
  AND U27293 ( .A(n27385), .B(n27386), .Z(n27384) );
  XOR U27294 ( .A(n27383), .B(n27387), .Z(n27385) );
  XOR U27295 ( .A(n27388), .B(n27340), .Z(n27334) );
  XOR U27296 ( .A(n27389), .B(n27390), .Z(n27340) );
  NOR U27297 ( .A(n27391), .B(n27392), .Z(n27390) );
  XOR U27298 ( .A(n27389), .B(n27393), .Z(n27391) );
  XNOR U27299 ( .A(n27339), .B(n27331), .Z(n27388) );
  XOR U27300 ( .A(n27394), .B(n27395), .Z(n27331) );
  AND U27301 ( .A(n27396), .B(n27397), .Z(n27395) );
  XOR U27302 ( .A(n27394), .B(n27398), .Z(n27396) );
  XNOR U27303 ( .A(n27399), .B(n27336), .Z(n27339) );
  XOR U27304 ( .A(n27400), .B(n27401), .Z(n27336) );
  AND U27305 ( .A(n27402), .B(n27403), .Z(n27401) );
  XNOR U27306 ( .A(n27404), .B(n27405), .Z(n27402) );
  IV U27307 ( .A(n27400), .Z(n27404) );
  XNOR U27308 ( .A(n27406), .B(n27407), .Z(n27399) );
  NOR U27309 ( .A(n27408), .B(n27409), .Z(n27407) );
  XNOR U27310 ( .A(n27406), .B(n27410), .Z(n27408) );
  XOR U27311 ( .A(n27329), .B(n27341), .Z(n27364) );
  NOR U27312 ( .A(n27267), .B(n27411), .Z(n27341) );
  XNOR U27313 ( .A(n27347), .B(n27346), .Z(n27329) );
  XNOR U27314 ( .A(n27412), .B(n27352), .Z(n27346) );
  XNOR U27315 ( .A(n27413), .B(n27414), .Z(n27352) );
  NOR U27316 ( .A(n27415), .B(n27416), .Z(n27414) );
  XOR U27317 ( .A(n27413), .B(n27417), .Z(n27415) );
  XNOR U27318 ( .A(n27351), .B(n27343), .Z(n27412) );
  XOR U27319 ( .A(n27418), .B(n27419), .Z(n27343) );
  AND U27320 ( .A(n27420), .B(n27421), .Z(n27419) );
  XOR U27321 ( .A(n27418), .B(n27422), .Z(n27420) );
  XNOR U27322 ( .A(n27423), .B(n27348), .Z(n27351) );
  XOR U27323 ( .A(n27424), .B(n27425), .Z(n27348) );
  AND U27324 ( .A(n27426), .B(n27427), .Z(n27425) );
  XNOR U27325 ( .A(n27428), .B(n27429), .Z(n27426) );
  IV U27326 ( .A(n27424), .Z(n27428) );
  XNOR U27327 ( .A(n27430), .B(n27431), .Z(n27423) );
  NOR U27328 ( .A(n27432), .B(n27433), .Z(n27431) );
  XNOR U27329 ( .A(n27430), .B(n27434), .Z(n27432) );
  XOR U27330 ( .A(n27357), .B(n27356), .Z(n27347) );
  XNOR U27331 ( .A(n27435), .B(n27353), .Z(n27356) );
  XOR U27332 ( .A(n27436), .B(n27437), .Z(n27353) );
  AND U27333 ( .A(n27438), .B(n27439), .Z(n27437) );
  XNOR U27334 ( .A(n27440), .B(n27441), .Z(n27438) );
  IV U27335 ( .A(n27436), .Z(n27440) );
  XNOR U27336 ( .A(n27442), .B(n27443), .Z(n27435) );
  NOR U27337 ( .A(n27444), .B(n27445), .Z(n27443) );
  XNOR U27338 ( .A(n27442), .B(n27446), .Z(n27444) );
  XOR U27339 ( .A(n27447), .B(n27448), .Z(n27357) );
  NOR U27340 ( .A(n27449), .B(n27450), .Z(n27448) );
  XNOR U27341 ( .A(n27447), .B(n27451), .Z(n27449) );
  XNOR U27342 ( .A(n27256), .B(n27360), .Z(n27362) );
  XNOR U27343 ( .A(n27452), .B(n27453), .Z(n27256) );
  AND U27344 ( .A(n496), .B(n27263), .Z(n27453) );
  XOR U27345 ( .A(n27452), .B(n27261), .Z(n27263) );
  AND U27346 ( .A(n27264), .B(n27267), .Z(n27360) );
  XOR U27347 ( .A(n27454), .B(n27411), .Z(n27267) );
  XNOR U27348 ( .A(p_input[1248]), .B(p_input[2048]), .Z(n27411) );
  XNOR U27349 ( .A(n27387), .B(n27386), .Z(n27454) );
  XNOR U27350 ( .A(n27455), .B(n27398), .Z(n27386) );
  XOR U27351 ( .A(n27372), .B(n27370), .Z(n27398) );
  XNOR U27352 ( .A(n27456), .B(n27377), .Z(n27370) );
  XOR U27353 ( .A(p_input[1272]), .B(p_input[2072]), .Z(n27377) );
  XOR U27354 ( .A(n27367), .B(n27376), .Z(n27456) );
  XOR U27355 ( .A(n27457), .B(n27373), .Z(n27376) );
  XOR U27356 ( .A(p_input[1270]), .B(p_input[2070]), .Z(n27373) );
  XOR U27357 ( .A(p_input[1271]), .B(n17295), .Z(n27457) );
  XOR U27358 ( .A(p_input[1266]), .B(p_input[2066]), .Z(n27367) );
  XNOR U27359 ( .A(n27382), .B(n27381), .Z(n27372) );
  XOR U27360 ( .A(n27458), .B(n27378), .Z(n27381) );
  XOR U27361 ( .A(p_input[1267]), .B(p_input[2067]), .Z(n27378) );
  XOR U27362 ( .A(p_input[1268]), .B(n17297), .Z(n27458) );
  XOR U27363 ( .A(p_input[1269]), .B(p_input[2069]), .Z(n27382) );
  XOR U27364 ( .A(n27397), .B(n27459), .Z(n27455) );
  IV U27365 ( .A(n27383), .Z(n27459) );
  XOR U27366 ( .A(p_input[1249]), .B(p_input[2049]), .Z(n27383) );
  XNOR U27367 ( .A(n27460), .B(n27405), .Z(n27397) );
  XNOR U27368 ( .A(n27393), .B(n27392), .Z(n27405) );
  XNOR U27369 ( .A(n27461), .B(n27389), .Z(n27392) );
  XNOR U27370 ( .A(p_input[1274]), .B(p_input[2074]), .Z(n27389) );
  XOR U27371 ( .A(p_input[1275]), .B(n17300), .Z(n27461) );
  XOR U27372 ( .A(p_input[1276]), .B(p_input[2076]), .Z(n27393) );
  XOR U27373 ( .A(n27403), .B(n27462), .Z(n27460) );
  IV U27374 ( .A(n27394), .Z(n27462) );
  XOR U27375 ( .A(p_input[1265]), .B(p_input[2065]), .Z(n27394) );
  XNOR U27376 ( .A(n27463), .B(n27410), .Z(n27403) );
  XNOR U27377 ( .A(p_input[1279]), .B(n17303), .Z(n27410) );
  XOR U27378 ( .A(n27400), .B(n27409), .Z(n27463) );
  XOR U27379 ( .A(n27464), .B(n27406), .Z(n27409) );
  XOR U27380 ( .A(p_input[1277]), .B(p_input[2077]), .Z(n27406) );
  XOR U27381 ( .A(p_input[1278]), .B(n17305), .Z(n27464) );
  XOR U27382 ( .A(p_input[1273]), .B(p_input[2073]), .Z(n27400) );
  XOR U27383 ( .A(n27422), .B(n27421), .Z(n27387) );
  XNOR U27384 ( .A(n27465), .B(n27429), .Z(n27421) );
  XNOR U27385 ( .A(n27417), .B(n27416), .Z(n27429) );
  XNOR U27386 ( .A(n27466), .B(n27413), .Z(n27416) );
  XNOR U27387 ( .A(p_input[1259]), .B(p_input[2059]), .Z(n27413) );
  XOR U27388 ( .A(p_input[1260]), .B(n16451), .Z(n27466) );
  XOR U27389 ( .A(p_input[1261]), .B(p_input[2061]), .Z(n27417) );
  XOR U27390 ( .A(n27427), .B(n27467), .Z(n27465) );
  IV U27391 ( .A(n27418), .Z(n27467) );
  XOR U27392 ( .A(p_input[1250]), .B(p_input[2050]), .Z(n27418) );
  XNOR U27393 ( .A(n27468), .B(n27434), .Z(n27427) );
  XNOR U27394 ( .A(p_input[1264]), .B(n16454), .Z(n27434) );
  XOR U27395 ( .A(n27424), .B(n27433), .Z(n27468) );
  XOR U27396 ( .A(n27469), .B(n27430), .Z(n27433) );
  XOR U27397 ( .A(p_input[1262]), .B(p_input[2062]), .Z(n27430) );
  XOR U27398 ( .A(p_input[1263]), .B(n16456), .Z(n27469) );
  XOR U27399 ( .A(p_input[1258]), .B(p_input[2058]), .Z(n27424) );
  XOR U27400 ( .A(n27441), .B(n27439), .Z(n27422) );
  XNOR U27401 ( .A(n27470), .B(n27446), .Z(n27439) );
  XOR U27402 ( .A(p_input[1257]), .B(p_input[2057]), .Z(n27446) );
  XOR U27403 ( .A(n27436), .B(n27445), .Z(n27470) );
  XOR U27404 ( .A(n27471), .B(n27442), .Z(n27445) );
  XOR U27405 ( .A(p_input[1255]), .B(p_input[2055]), .Z(n27442) );
  XOR U27406 ( .A(p_input[1256]), .B(n17312), .Z(n27471) );
  XOR U27407 ( .A(p_input[1251]), .B(p_input[2051]), .Z(n27436) );
  XNOR U27408 ( .A(n27451), .B(n27450), .Z(n27441) );
  XOR U27409 ( .A(n27472), .B(n27447), .Z(n27450) );
  XOR U27410 ( .A(p_input[1252]), .B(p_input[2052]), .Z(n27447) );
  XOR U27411 ( .A(p_input[1253]), .B(n17314), .Z(n27472) );
  XOR U27412 ( .A(p_input[1254]), .B(p_input[2054]), .Z(n27451) );
  XNOR U27413 ( .A(n27473), .B(n27474), .Z(n27264) );
  AND U27414 ( .A(n496), .B(n27475), .Z(n27474) );
  XNOR U27415 ( .A(n27476), .B(n27477), .Z(n496) );
  AND U27416 ( .A(n27478), .B(n27479), .Z(n27477) );
  XOR U27417 ( .A(n27476), .B(n27274), .Z(n27479) );
  XNOR U27418 ( .A(n27476), .B(n27216), .Z(n27478) );
  XOR U27419 ( .A(n27480), .B(n27481), .Z(n27476) );
  AND U27420 ( .A(n27482), .B(n27483), .Z(n27481) );
  XNOR U27421 ( .A(n27287), .B(n27480), .Z(n27483) );
  XOR U27422 ( .A(n27480), .B(n27228), .Z(n27482) );
  XOR U27423 ( .A(n27484), .B(n27485), .Z(n27480) );
  AND U27424 ( .A(n27486), .B(n27487), .Z(n27485) );
  XNOR U27425 ( .A(n27312), .B(n27484), .Z(n27487) );
  XOR U27426 ( .A(n27484), .B(n27239), .Z(n27486) );
  XOR U27427 ( .A(n27488), .B(n27489), .Z(n27484) );
  AND U27428 ( .A(n27490), .B(n27491), .Z(n27489) );
  XOR U27429 ( .A(n27488), .B(n27249), .Z(n27490) );
  XOR U27430 ( .A(n27492), .B(n27493), .Z(n27205) );
  AND U27431 ( .A(n500), .B(n27475), .Z(n27493) );
  XNOR U27432 ( .A(n27473), .B(n27492), .Z(n27475) );
  XNOR U27433 ( .A(n27494), .B(n27495), .Z(n500) );
  AND U27434 ( .A(n27496), .B(n27497), .Z(n27495) );
  XNOR U27435 ( .A(n27498), .B(n27494), .Z(n27497) );
  IV U27436 ( .A(n27274), .Z(n27498) );
  XNOR U27437 ( .A(n27499), .B(n27500), .Z(n27274) );
  AND U27438 ( .A(n503), .B(n27501), .Z(n27500) );
  XNOR U27439 ( .A(n27499), .B(n27502), .Z(n27501) );
  XNOR U27440 ( .A(n27216), .B(n27494), .Z(n27496) );
  XOR U27441 ( .A(n27503), .B(n27504), .Z(n27216) );
  AND U27442 ( .A(n511), .B(n27505), .Z(n27504) );
  XOR U27443 ( .A(n27506), .B(n27507), .Z(n27494) );
  AND U27444 ( .A(n27508), .B(n27509), .Z(n27507) );
  XNOR U27445 ( .A(n27506), .B(n27287), .Z(n27509) );
  XNOR U27446 ( .A(n27510), .B(n27511), .Z(n27287) );
  AND U27447 ( .A(n503), .B(n27512), .Z(n27511) );
  XOR U27448 ( .A(n27513), .B(n27510), .Z(n27512) );
  XNOR U27449 ( .A(n27514), .B(n27506), .Z(n27508) );
  IV U27450 ( .A(n27228), .Z(n27514) );
  XOR U27451 ( .A(n27515), .B(n27516), .Z(n27228) );
  AND U27452 ( .A(n511), .B(n27517), .Z(n27516) );
  XOR U27453 ( .A(n27518), .B(n27519), .Z(n27506) );
  AND U27454 ( .A(n27520), .B(n27521), .Z(n27519) );
  XNOR U27455 ( .A(n27518), .B(n27312), .Z(n27521) );
  XNOR U27456 ( .A(n27522), .B(n27523), .Z(n27312) );
  AND U27457 ( .A(n503), .B(n27524), .Z(n27523) );
  XNOR U27458 ( .A(n27525), .B(n27522), .Z(n27524) );
  XOR U27459 ( .A(n27239), .B(n27518), .Z(n27520) );
  XOR U27460 ( .A(n27526), .B(n27527), .Z(n27239) );
  AND U27461 ( .A(n511), .B(n27528), .Z(n27527) );
  XOR U27462 ( .A(n27488), .B(n27529), .Z(n27518) );
  AND U27463 ( .A(n27530), .B(n27491), .Z(n27529) );
  XNOR U27464 ( .A(n27358), .B(n27488), .Z(n27491) );
  XNOR U27465 ( .A(n27531), .B(n27532), .Z(n27358) );
  AND U27466 ( .A(n503), .B(n27533), .Z(n27532) );
  XOR U27467 ( .A(n27534), .B(n27531), .Z(n27533) );
  XNOR U27468 ( .A(n27535), .B(n27488), .Z(n27530) );
  IV U27469 ( .A(n27249), .Z(n27535) );
  XOR U27470 ( .A(n27536), .B(n27537), .Z(n27249) );
  AND U27471 ( .A(n511), .B(n27538), .Z(n27537) );
  XOR U27472 ( .A(n27539), .B(n27540), .Z(n27488) );
  AND U27473 ( .A(n27541), .B(n27542), .Z(n27540) );
  XNOR U27474 ( .A(n27539), .B(n27452), .Z(n27542) );
  XNOR U27475 ( .A(n27543), .B(n27544), .Z(n27452) );
  AND U27476 ( .A(n503), .B(n27545), .Z(n27544) );
  XNOR U27477 ( .A(n27546), .B(n27543), .Z(n27545) );
  XNOR U27478 ( .A(n27547), .B(n27539), .Z(n27541) );
  IV U27479 ( .A(n27261), .Z(n27547) );
  XOR U27480 ( .A(n27548), .B(n27549), .Z(n27261) );
  AND U27481 ( .A(n511), .B(n27550), .Z(n27549) );
  AND U27482 ( .A(n27492), .B(n27473), .Z(n27539) );
  XNOR U27483 ( .A(n27551), .B(n27552), .Z(n27473) );
  AND U27484 ( .A(n503), .B(n27553), .Z(n27552) );
  XNOR U27485 ( .A(n27554), .B(n27551), .Z(n27553) );
  XNOR U27486 ( .A(n27555), .B(n27556), .Z(n503) );
  AND U27487 ( .A(n27557), .B(n27558), .Z(n27556) );
  XOR U27488 ( .A(n27502), .B(n27555), .Z(n27558) );
  AND U27489 ( .A(n27559), .B(n27560), .Z(n27502) );
  XOR U27490 ( .A(n27555), .B(n27499), .Z(n27557) );
  XNOR U27491 ( .A(n27561), .B(n27562), .Z(n27499) );
  AND U27492 ( .A(n507), .B(n27505), .Z(n27562) );
  XOR U27493 ( .A(n27503), .B(n27561), .Z(n27505) );
  XOR U27494 ( .A(n27563), .B(n27564), .Z(n27555) );
  AND U27495 ( .A(n27565), .B(n27566), .Z(n27564) );
  XNOR U27496 ( .A(n27563), .B(n27559), .Z(n27566) );
  IV U27497 ( .A(n27513), .Z(n27559) );
  XOR U27498 ( .A(n27567), .B(n27568), .Z(n27513) );
  XOR U27499 ( .A(n27569), .B(n27560), .Z(n27568) );
  AND U27500 ( .A(n27525), .B(n27570), .Z(n27560) );
  AND U27501 ( .A(n27571), .B(n27572), .Z(n27569) );
  XOR U27502 ( .A(n27573), .B(n27567), .Z(n27571) );
  XNOR U27503 ( .A(n27510), .B(n27563), .Z(n27565) );
  XNOR U27504 ( .A(n27574), .B(n27575), .Z(n27510) );
  AND U27505 ( .A(n507), .B(n27517), .Z(n27575) );
  XOR U27506 ( .A(n27574), .B(n27515), .Z(n27517) );
  XOR U27507 ( .A(n27576), .B(n27577), .Z(n27563) );
  AND U27508 ( .A(n27578), .B(n27579), .Z(n27577) );
  XNOR U27509 ( .A(n27576), .B(n27525), .Z(n27579) );
  XOR U27510 ( .A(n27580), .B(n27572), .Z(n27525) );
  XNOR U27511 ( .A(n27581), .B(n27567), .Z(n27572) );
  XOR U27512 ( .A(n27582), .B(n27583), .Z(n27567) );
  AND U27513 ( .A(n27584), .B(n27585), .Z(n27583) );
  XOR U27514 ( .A(n27586), .B(n27582), .Z(n27584) );
  XNOR U27515 ( .A(n27587), .B(n27588), .Z(n27581) );
  AND U27516 ( .A(n27589), .B(n27590), .Z(n27588) );
  XOR U27517 ( .A(n27587), .B(n27591), .Z(n27589) );
  XNOR U27518 ( .A(n27573), .B(n27570), .Z(n27580) );
  AND U27519 ( .A(n27592), .B(n27593), .Z(n27570) );
  XOR U27520 ( .A(n27594), .B(n27595), .Z(n27573) );
  AND U27521 ( .A(n27596), .B(n27597), .Z(n27595) );
  XOR U27522 ( .A(n27594), .B(n27598), .Z(n27596) );
  XNOR U27523 ( .A(n27522), .B(n27576), .Z(n27578) );
  XNOR U27524 ( .A(n27599), .B(n27600), .Z(n27522) );
  AND U27525 ( .A(n507), .B(n27528), .Z(n27600) );
  XOR U27526 ( .A(n27599), .B(n27526), .Z(n27528) );
  XOR U27527 ( .A(n27601), .B(n27602), .Z(n27576) );
  AND U27528 ( .A(n27603), .B(n27604), .Z(n27602) );
  XNOR U27529 ( .A(n27601), .B(n27592), .Z(n27604) );
  IV U27530 ( .A(n27534), .Z(n27592) );
  XNOR U27531 ( .A(n27605), .B(n27585), .Z(n27534) );
  XNOR U27532 ( .A(n27606), .B(n27591), .Z(n27585) );
  XOR U27533 ( .A(n27607), .B(n27608), .Z(n27591) );
  AND U27534 ( .A(n27609), .B(n27610), .Z(n27608) );
  XOR U27535 ( .A(n27607), .B(n27611), .Z(n27609) );
  XNOR U27536 ( .A(n27590), .B(n27582), .Z(n27606) );
  XOR U27537 ( .A(n27612), .B(n27613), .Z(n27582) );
  AND U27538 ( .A(n27614), .B(n27615), .Z(n27613) );
  XNOR U27539 ( .A(n27616), .B(n27612), .Z(n27614) );
  XNOR U27540 ( .A(n27617), .B(n27587), .Z(n27590) );
  XOR U27541 ( .A(n27618), .B(n27619), .Z(n27587) );
  AND U27542 ( .A(n27620), .B(n27621), .Z(n27619) );
  XOR U27543 ( .A(n27618), .B(n27622), .Z(n27620) );
  XNOR U27544 ( .A(n27623), .B(n27624), .Z(n27617) );
  AND U27545 ( .A(n27625), .B(n27626), .Z(n27624) );
  XNOR U27546 ( .A(n27623), .B(n27627), .Z(n27625) );
  XNOR U27547 ( .A(n27586), .B(n27593), .Z(n27605) );
  AND U27548 ( .A(n27546), .B(n27628), .Z(n27593) );
  XOR U27549 ( .A(n27598), .B(n27597), .Z(n27586) );
  XNOR U27550 ( .A(n27629), .B(n27594), .Z(n27597) );
  XOR U27551 ( .A(n27630), .B(n27631), .Z(n27594) );
  AND U27552 ( .A(n27632), .B(n27633), .Z(n27631) );
  XOR U27553 ( .A(n27630), .B(n27634), .Z(n27632) );
  XNOR U27554 ( .A(n27635), .B(n27636), .Z(n27629) );
  AND U27555 ( .A(n27637), .B(n27638), .Z(n27636) );
  XOR U27556 ( .A(n27635), .B(n27639), .Z(n27637) );
  XOR U27557 ( .A(n27640), .B(n27641), .Z(n27598) );
  AND U27558 ( .A(n27642), .B(n27643), .Z(n27641) );
  XOR U27559 ( .A(n27640), .B(n27644), .Z(n27642) );
  XNOR U27560 ( .A(n27531), .B(n27601), .Z(n27603) );
  XNOR U27561 ( .A(n27645), .B(n27646), .Z(n27531) );
  AND U27562 ( .A(n507), .B(n27538), .Z(n27646) );
  XOR U27563 ( .A(n27645), .B(n27536), .Z(n27538) );
  XOR U27564 ( .A(n27647), .B(n27648), .Z(n27601) );
  AND U27565 ( .A(n27649), .B(n27650), .Z(n27648) );
  XNOR U27566 ( .A(n27647), .B(n27546), .Z(n27650) );
  XOR U27567 ( .A(n27651), .B(n27615), .Z(n27546) );
  XNOR U27568 ( .A(n27652), .B(n27622), .Z(n27615) );
  XOR U27569 ( .A(n27611), .B(n27610), .Z(n27622) );
  XNOR U27570 ( .A(n27653), .B(n27607), .Z(n27610) );
  XOR U27571 ( .A(n27654), .B(n27655), .Z(n27607) );
  AND U27572 ( .A(n27656), .B(n27657), .Z(n27655) );
  XNOR U27573 ( .A(n27658), .B(n27659), .Z(n27656) );
  IV U27574 ( .A(n27654), .Z(n27658) );
  XNOR U27575 ( .A(n27660), .B(n27661), .Z(n27653) );
  NOR U27576 ( .A(n27662), .B(n27663), .Z(n27661) );
  XNOR U27577 ( .A(n27660), .B(n27664), .Z(n27662) );
  XOR U27578 ( .A(n27665), .B(n27666), .Z(n27611) );
  NOR U27579 ( .A(n27667), .B(n27668), .Z(n27666) );
  XNOR U27580 ( .A(n27665), .B(n27669), .Z(n27667) );
  XNOR U27581 ( .A(n27621), .B(n27612), .Z(n27652) );
  XOR U27582 ( .A(n27670), .B(n27671), .Z(n27612) );
  AND U27583 ( .A(n27672), .B(n27673), .Z(n27671) );
  XOR U27584 ( .A(n27670), .B(n27674), .Z(n27672) );
  XOR U27585 ( .A(n27675), .B(n27627), .Z(n27621) );
  XOR U27586 ( .A(n27676), .B(n27677), .Z(n27627) );
  NOR U27587 ( .A(n27678), .B(n27679), .Z(n27677) );
  XOR U27588 ( .A(n27676), .B(n27680), .Z(n27678) );
  XNOR U27589 ( .A(n27626), .B(n27618), .Z(n27675) );
  XOR U27590 ( .A(n27681), .B(n27682), .Z(n27618) );
  AND U27591 ( .A(n27683), .B(n27684), .Z(n27682) );
  XOR U27592 ( .A(n27681), .B(n27685), .Z(n27683) );
  XNOR U27593 ( .A(n27686), .B(n27623), .Z(n27626) );
  XOR U27594 ( .A(n27687), .B(n27688), .Z(n27623) );
  AND U27595 ( .A(n27689), .B(n27690), .Z(n27688) );
  XNOR U27596 ( .A(n27691), .B(n27692), .Z(n27689) );
  IV U27597 ( .A(n27687), .Z(n27691) );
  XNOR U27598 ( .A(n27693), .B(n27694), .Z(n27686) );
  NOR U27599 ( .A(n27695), .B(n27696), .Z(n27694) );
  XNOR U27600 ( .A(n27693), .B(n27697), .Z(n27695) );
  XOR U27601 ( .A(n27616), .B(n27628), .Z(n27651) );
  NOR U27602 ( .A(n27554), .B(n27698), .Z(n27628) );
  XNOR U27603 ( .A(n27634), .B(n27633), .Z(n27616) );
  XNOR U27604 ( .A(n27699), .B(n27639), .Z(n27633) );
  XNOR U27605 ( .A(n27700), .B(n27701), .Z(n27639) );
  NOR U27606 ( .A(n27702), .B(n27703), .Z(n27701) );
  XOR U27607 ( .A(n27700), .B(n27704), .Z(n27702) );
  XNOR U27608 ( .A(n27638), .B(n27630), .Z(n27699) );
  XOR U27609 ( .A(n27705), .B(n27706), .Z(n27630) );
  AND U27610 ( .A(n27707), .B(n27708), .Z(n27706) );
  XOR U27611 ( .A(n27705), .B(n27709), .Z(n27707) );
  XNOR U27612 ( .A(n27710), .B(n27635), .Z(n27638) );
  XOR U27613 ( .A(n27711), .B(n27712), .Z(n27635) );
  AND U27614 ( .A(n27713), .B(n27714), .Z(n27712) );
  XNOR U27615 ( .A(n27715), .B(n27716), .Z(n27713) );
  IV U27616 ( .A(n27711), .Z(n27715) );
  XNOR U27617 ( .A(n27717), .B(n27718), .Z(n27710) );
  NOR U27618 ( .A(n27719), .B(n27720), .Z(n27718) );
  XNOR U27619 ( .A(n27717), .B(n27721), .Z(n27719) );
  XOR U27620 ( .A(n27644), .B(n27643), .Z(n27634) );
  XNOR U27621 ( .A(n27722), .B(n27640), .Z(n27643) );
  XOR U27622 ( .A(n27723), .B(n27724), .Z(n27640) );
  AND U27623 ( .A(n27725), .B(n27726), .Z(n27724) );
  XNOR U27624 ( .A(n27727), .B(n27728), .Z(n27725) );
  IV U27625 ( .A(n27723), .Z(n27727) );
  XNOR U27626 ( .A(n27729), .B(n27730), .Z(n27722) );
  NOR U27627 ( .A(n27731), .B(n27732), .Z(n27730) );
  XNOR U27628 ( .A(n27729), .B(n27733), .Z(n27731) );
  XOR U27629 ( .A(n27734), .B(n27735), .Z(n27644) );
  NOR U27630 ( .A(n27736), .B(n27737), .Z(n27735) );
  XNOR U27631 ( .A(n27734), .B(n27738), .Z(n27736) );
  XNOR U27632 ( .A(n27543), .B(n27647), .Z(n27649) );
  XNOR U27633 ( .A(n27739), .B(n27740), .Z(n27543) );
  AND U27634 ( .A(n507), .B(n27550), .Z(n27740) );
  XOR U27635 ( .A(n27739), .B(n27548), .Z(n27550) );
  AND U27636 ( .A(n27551), .B(n27554), .Z(n27647) );
  XOR U27637 ( .A(n27741), .B(n27698), .Z(n27554) );
  XNOR U27638 ( .A(p_input[1280]), .B(p_input[2048]), .Z(n27698) );
  XNOR U27639 ( .A(n27674), .B(n27673), .Z(n27741) );
  XNOR U27640 ( .A(n27742), .B(n27685), .Z(n27673) );
  XOR U27641 ( .A(n27659), .B(n27657), .Z(n27685) );
  XNOR U27642 ( .A(n27743), .B(n27664), .Z(n27657) );
  XOR U27643 ( .A(p_input[1304]), .B(p_input[2072]), .Z(n27664) );
  XOR U27644 ( .A(n27654), .B(n27663), .Z(n27743) );
  XOR U27645 ( .A(n27744), .B(n27660), .Z(n27663) );
  XOR U27646 ( .A(p_input[1302]), .B(p_input[2070]), .Z(n27660) );
  XOR U27647 ( .A(p_input[1303]), .B(n17295), .Z(n27744) );
  XOR U27648 ( .A(p_input[1298]), .B(p_input[2066]), .Z(n27654) );
  XNOR U27649 ( .A(n27669), .B(n27668), .Z(n27659) );
  XOR U27650 ( .A(n27745), .B(n27665), .Z(n27668) );
  XOR U27651 ( .A(p_input[1299]), .B(p_input[2067]), .Z(n27665) );
  XOR U27652 ( .A(p_input[1300]), .B(n17297), .Z(n27745) );
  XOR U27653 ( .A(p_input[1301]), .B(p_input[2069]), .Z(n27669) );
  XOR U27654 ( .A(n27684), .B(n27746), .Z(n27742) );
  IV U27655 ( .A(n27670), .Z(n27746) );
  XOR U27656 ( .A(p_input[1281]), .B(p_input[2049]), .Z(n27670) );
  XNOR U27657 ( .A(n27747), .B(n27692), .Z(n27684) );
  XNOR U27658 ( .A(n27680), .B(n27679), .Z(n27692) );
  XNOR U27659 ( .A(n27748), .B(n27676), .Z(n27679) );
  XNOR U27660 ( .A(p_input[1306]), .B(p_input[2074]), .Z(n27676) );
  XOR U27661 ( .A(p_input[1307]), .B(n17300), .Z(n27748) );
  XOR U27662 ( .A(p_input[1308]), .B(p_input[2076]), .Z(n27680) );
  XOR U27663 ( .A(n27690), .B(n27749), .Z(n27747) );
  IV U27664 ( .A(n27681), .Z(n27749) );
  XOR U27665 ( .A(p_input[1297]), .B(p_input[2065]), .Z(n27681) );
  XNOR U27666 ( .A(n27750), .B(n27697), .Z(n27690) );
  XNOR U27667 ( .A(p_input[1311]), .B(n17303), .Z(n27697) );
  XOR U27668 ( .A(n27687), .B(n27696), .Z(n27750) );
  XOR U27669 ( .A(n27751), .B(n27693), .Z(n27696) );
  XOR U27670 ( .A(p_input[1309]), .B(p_input[2077]), .Z(n27693) );
  XOR U27671 ( .A(p_input[1310]), .B(n17305), .Z(n27751) );
  XOR U27672 ( .A(p_input[1305]), .B(p_input[2073]), .Z(n27687) );
  XOR U27673 ( .A(n27709), .B(n27708), .Z(n27674) );
  XNOR U27674 ( .A(n27752), .B(n27716), .Z(n27708) );
  XNOR U27675 ( .A(n27704), .B(n27703), .Z(n27716) );
  XNOR U27676 ( .A(n27753), .B(n27700), .Z(n27703) );
  XNOR U27677 ( .A(p_input[1291]), .B(p_input[2059]), .Z(n27700) );
  XOR U27678 ( .A(p_input[1292]), .B(n16451), .Z(n27753) );
  XOR U27679 ( .A(p_input[1293]), .B(p_input[2061]), .Z(n27704) );
  XOR U27680 ( .A(n27714), .B(n27754), .Z(n27752) );
  IV U27681 ( .A(n27705), .Z(n27754) );
  XOR U27682 ( .A(p_input[1282]), .B(p_input[2050]), .Z(n27705) );
  XNOR U27683 ( .A(n27755), .B(n27721), .Z(n27714) );
  XNOR U27684 ( .A(p_input[1296]), .B(n16454), .Z(n27721) );
  XOR U27685 ( .A(n27711), .B(n27720), .Z(n27755) );
  XOR U27686 ( .A(n27756), .B(n27717), .Z(n27720) );
  XOR U27687 ( .A(p_input[1294]), .B(p_input[2062]), .Z(n27717) );
  XOR U27688 ( .A(p_input[1295]), .B(n16456), .Z(n27756) );
  XOR U27689 ( .A(p_input[1290]), .B(p_input[2058]), .Z(n27711) );
  XOR U27690 ( .A(n27728), .B(n27726), .Z(n27709) );
  XNOR U27691 ( .A(n27757), .B(n27733), .Z(n27726) );
  XOR U27692 ( .A(p_input[1289]), .B(p_input[2057]), .Z(n27733) );
  XOR U27693 ( .A(n27723), .B(n27732), .Z(n27757) );
  XOR U27694 ( .A(n27758), .B(n27729), .Z(n27732) );
  XOR U27695 ( .A(p_input[1287]), .B(p_input[2055]), .Z(n27729) );
  XOR U27696 ( .A(p_input[1288]), .B(n17312), .Z(n27758) );
  XOR U27697 ( .A(p_input[1283]), .B(p_input[2051]), .Z(n27723) );
  XNOR U27698 ( .A(n27738), .B(n27737), .Z(n27728) );
  XOR U27699 ( .A(n27759), .B(n27734), .Z(n27737) );
  XOR U27700 ( .A(p_input[1284]), .B(p_input[2052]), .Z(n27734) );
  XOR U27701 ( .A(p_input[1285]), .B(n17314), .Z(n27759) );
  XOR U27702 ( .A(p_input[1286]), .B(p_input[2054]), .Z(n27738) );
  XNOR U27703 ( .A(n27760), .B(n27761), .Z(n27551) );
  AND U27704 ( .A(n507), .B(n27762), .Z(n27761) );
  XNOR U27705 ( .A(n27763), .B(n27764), .Z(n507) );
  AND U27706 ( .A(n27765), .B(n27766), .Z(n27764) );
  XOR U27707 ( .A(n27763), .B(n27561), .Z(n27766) );
  XNOR U27708 ( .A(n27763), .B(n27503), .Z(n27765) );
  XOR U27709 ( .A(n27767), .B(n27768), .Z(n27763) );
  AND U27710 ( .A(n27769), .B(n27770), .Z(n27768) );
  XNOR U27711 ( .A(n27574), .B(n27767), .Z(n27770) );
  XOR U27712 ( .A(n27767), .B(n27515), .Z(n27769) );
  XOR U27713 ( .A(n27771), .B(n27772), .Z(n27767) );
  AND U27714 ( .A(n27773), .B(n27774), .Z(n27772) );
  XNOR U27715 ( .A(n27599), .B(n27771), .Z(n27774) );
  XOR U27716 ( .A(n27771), .B(n27526), .Z(n27773) );
  XOR U27717 ( .A(n27775), .B(n27776), .Z(n27771) );
  AND U27718 ( .A(n27777), .B(n27778), .Z(n27776) );
  XOR U27719 ( .A(n27775), .B(n27536), .Z(n27777) );
  XOR U27720 ( .A(n27779), .B(n27780), .Z(n27492) );
  AND U27721 ( .A(n511), .B(n27762), .Z(n27780) );
  XNOR U27722 ( .A(n27760), .B(n27779), .Z(n27762) );
  XNOR U27723 ( .A(n27781), .B(n27782), .Z(n511) );
  AND U27724 ( .A(n27783), .B(n27784), .Z(n27782) );
  XNOR U27725 ( .A(n27785), .B(n27781), .Z(n27784) );
  IV U27726 ( .A(n27561), .Z(n27785) );
  XNOR U27727 ( .A(n27786), .B(n27787), .Z(n27561) );
  AND U27728 ( .A(n514), .B(n27788), .Z(n27787) );
  XNOR U27729 ( .A(n27786), .B(n27789), .Z(n27788) );
  XNOR U27730 ( .A(n27503), .B(n27781), .Z(n27783) );
  XOR U27731 ( .A(n27790), .B(n27791), .Z(n27503) );
  AND U27732 ( .A(n522), .B(n27792), .Z(n27791) );
  XOR U27733 ( .A(n27793), .B(n27794), .Z(n27781) );
  AND U27734 ( .A(n27795), .B(n27796), .Z(n27794) );
  XNOR U27735 ( .A(n27793), .B(n27574), .Z(n27796) );
  XNOR U27736 ( .A(n27797), .B(n27798), .Z(n27574) );
  AND U27737 ( .A(n514), .B(n27799), .Z(n27798) );
  XOR U27738 ( .A(n27800), .B(n27797), .Z(n27799) );
  XNOR U27739 ( .A(n27801), .B(n27793), .Z(n27795) );
  IV U27740 ( .A(n27515), .Z(n27801) );
  XOR U27741 ( .A(n27802), .B(n27803), .Z(n27515) );
  AND U27742 ( .A(n522), .B(n27804), .Z(n27803) );
  XOR U27743 ( .A(n27805), .B(n27806), .Z(n27793) );
  AND U27744 ( .A(n27807), .B(n27808), .Z(n27806) );
  XNOR U27745 ( .A(n27805), .B(n27599), .Z(n27808) );
  XNOR U27746 ( .A(n27809), .B(n27810), .Z(n27599) );
  AND U27747 ( .A(n514), .B(n27811), .Z(n27810) );
  XNOR U27748 ( .A(n27812), .B(n27809), .Z(n27811) );
  XOR U27749 ( .A(n27526), .B(n27805), .Z(n27807) );
  XOR U27750 ( .A(n27813), .B(n27814), .Z(n27526) );
  AND U27751 ( .A(n522), .B(n27815), .Z(n27814) );
  XOR U27752 ( .A(n27775), .B(n27816), .Z(n27805) );
  AND U27753 ( .A(n27817), .B(n27778), .Z(n27816) );
  XNOR U27754 ( .A(n27645), .B(n27775), .Z(n27778) );
  XNOR U27755 ( .A(n27818), .B(n27819), .Z(n27645) );
  AND U27756 ( .A(n514), .B(n27820), .Z(n27819) );
  XOR U27757 ( .A(n27821), .B(n27818), .Z(n27820) );
  XNOR U27758 ( .A(n27822), .B(n27775), .Z(n27817) );
  IV U27759 ( .A(n27536), .Z(n27822) );
  XOR U27760 ( .A(n27823), .B(n27824), .Z(n27536) );
  AND U27761 ( .A(n522), .B(n27825), .Z(n27824) );
  XOR U27762 ( .A(n27826), .B(n27827), .Z(n27775) );
  AND U27763 ( .A(n27828), .B(n27829), .Z(n27827) );
  XNOR U27764 ( .A(n27826), .B(n27739), .Z(n27829) );
  XNOR U27765 ( .A(n27830), .B(n27831), .Z(n27739) );
  AND U27766 ( .A(n514), .B(n27832), .Z(n27831) );
  XNOR U27767 ( .A(n27833), .B(n27830), .Z(n27832) );
  XNOR U27768 ( .A(n27834), .B(n27826), .Z(n27828) );
  IV U27769 ( .A(n27548), .Z(n27834) );
  XOR U27770 ( .A(n27835), .B(n27836), .Z(n27548) );
  AND U27771 ( .A(n522), .B(n27837), .Z(n27836) );
  AND U27772 ( .A(n27779), .B(n27760), .Z(n27826) );
  XNOR U27773 ( .A(n27838), .B(n27839), .Z(n27760) );
  AND U27774 ( .A(n514), .B(n27840), .Z(n27839) );
  XNOR U27775 ( .A(n27841), .B(n27838), .Z(n27840) );
  XNOR U27776 ( .A(n27842), .B(n27843), .Z(n514) );
  AND U27777 ( .A(n27844), .B(n27845), .Z(n27843) );
  XOR U27778 ( .A(n27789), .B(n27842), .Z(n27845) );
  AND U27779 ( .A(n27846), .B(n27847), .Z(n27789) );
  XOR U27780 ( .A(n27842), .B(n27786), .Z(n27844) );
  XNOR U27781 ( .A(n27848), .B(n27849), .Z(n27786) );
  AND U27782 ( .A(n518), .B(n27792), .Z(n27849) );
  XOR U27783 ( .A(n27790), .B(n27848), .Z(n27792) );
  XOR U27784 ( .A(n27850), .B(n27851), .Z(n27842) );
  AND U27785 ( .A(n27852), .B(n27853), .Z(n27851) );
  XNOR U27786 ( .A(n27850), .B(n27846), .Z(n27853) );
  IV U27787 ( .A(n27800), .Z(n27846) );
  XOR U27788 ( .A(n27854), .B(n27855), .Z(n27800) );
  XOR U27789 ( .A(n27856), .B(n27847), .Z(n27855) );
  AND U27790 ( .A(n27812), .B(n27857), .Z(n27847) );
  AND U27791 ( .A(n27858), .B(n27859), .Z(n27856) );
  XOR U27792 ( .A(n27860), .B(n27854), .Z(n27858) );
  XNOR U27793 ( .A(n27797), .B(n27850), .Z(n27852) );
  XNOR U27794 ( .A(n27861), .B(n27862), .Z(n27797) );
  AND U27795 ( .A(n518), .B(n27804), .Z(n27862) );
  XOR U27796 ( .A(n27861), .B(n27802), .Z(n27804) );
  XOR U27797 ( .A(n27863), .B(n27864), .Z(n27850) );
  AND U27798 ( .A(n27865), .B(n27866), .Z(n27864) );
  XNOR U27799 ( .A(n27863), .B(n27812), .Z(n27866) );
  XOR U27800 ( .A(n27867), .B(n27859), .Z(n27812) );
  XNOR U27801 ( .A(n27868), .B(n27854), .Z(n27859) );
  XOR U27802 ( .A(n27869), .B(n27870), .Z(n27854) );
  AND U27803 ( .A(n27871), .B(n27872), .Z(n27870) );
  XOR U27804 ( .A(n27873), .B(n27869), .Z(n27871) );
  XNOR U27805 ( .A(n27874), .B(n27875), .Z(n27868) );
  AND U27806 ( .A(n27876), .B(n27877), .Z(n27875) );
  XOR U27807 ( .A(n27874), .B(n27878), .Z(n27876) );
  XNOR U27808 ( .A(n27860), .B(n27857), .Z(n27867) );
  AND U27809 ( .A(n27879), .B(n27880), .Z(n27857) );
  XOR U27810 ( .A(n27881), .B(n27882), .Z(n27860) );
  AND U27811 ( .A(n27883), .B(n27884), .Z(n27882) );
  XOR U27812 ( .A(n27881), .B(n27885), .Z(n27883) );
  XNOR U27813 ( .A(n27809), .B(n27863), .Z(n27865) );
  XNOR U27814 ( .A(n27886), .B(n27887), .Z(n27809) );
  AND U27815 ( .A(n518), .B(n27815), .Z(n27887) );
  XOR U27816 ( .A(n27886), .B(n27813), .Z(n27815) );
  XOR U27817 ( .A(n27888), .B(n27889), .Z(n27863) );
  AND U27818 ( .A(n27890), .B(n27891), .Z(n27889) );
  XNOR U27819 ( .A(n27888), .B(n27879), .Z(n27891) );
  IV U27820 ( .A(n27821), .Z(n27879) );
  XNOR U27821 ( .A(n27892), .B(n27872), .Z(n27821) );
  XNOR U27822 ( .A(n27893), .B(n27878), .Z(n27872) );
  XOR U27823 ( .A(n27894), .B(n27895), .Z(n27878) );
  AND U27824 ( .A(n27896), .B(n27897), .Z(n27895) );
  XOR U27825 ( .A(n27894), .B(n27898), .Z(n27896) );
  XNOR U27826 ( .A(n27877), .B(n27869), .Z(n27893) );
  XOR U27827 ( .A(n27899), .B(n27900), .Z(n27869) );
  AND U27828 ( .A(n27901), .B(n27902), .Z(n27900) );
  XNOR U27829 ( .A(n27903), .B(n27899), .Z(n27901) );
  XNOR U27830 ( .A(n27904), .B(n27874), .Z(n27877) );
  XOR U27831 ( .A(n27905), .B(n27906), .Z(n27874) );
  AND U27832 ( .A(n27907), .B(n27908), .Z(n27906) );
  XOR U27833 ( .A(n27905), .B(n27909), .Z(n27907) );
  XNOR U27834 ( .A(n27910), .B(n27911), .Z(n27904) );
  AND U27835 ( .A(n27912), .B(n27913), .Z(n27911) );
  XNOR U27836 ( .A(n27910), .B(n27914), .Z(n27912) );
  XNOR U27837 ( .A(n27873), .B(n27880), .Z(n27892) );
  AND U27838 ( .A(n27833), .B(n27915), .Z(n27880) );
  XOR U27839 ( .A(n27885), .B(n27884), .Z(n27873) );
  XNOR U27840 ( .A(n27916), .B(n27881), .Z(n27884) );
  XOR U27841 ( .A(n27917), .B(n27918), .Z(n27881) );
  AND U27842 ( .A(n27919), .B(n27920), .Z(n27918) );
  XOR U27843 ( .A(n27917), .B(n27921), .Z(n27919) );
  XNOR U27844 ( .A(n27922), .B(n27923), .Z(n27916) );
  AND U27845 ( .A(n27924), .B(n27925), .Z(n27923) );
  XOR U27846 ( .A(n27922), .B(n27926), .Z(n27924) );
  XOR U27847 ( .A(n27927), .B(n27928), .Z(n27885) );
  AND U27848 ( .A(n27929), .B(n27930), .Z(n27928) );
  XOR U27849 ( .A(n27927), .B(n27931), .Z(n27929) );
  XNOR U27850 ( .A(n27818), .B(n27888), .Z(n27890) );
  XNOR U27851 ( .A(n27932), .B(n27933), .Z(n27818) );
  AND U27852 ( .A(n518), .B(n27825), .Z(n27933) );
  XOR U27853 ( .A(n27932), .B(n27823), .Z(n27825) );
  XOR U27854 ( .A(n27934), .B(n27935), .Z(n27888) );
  AND U27855 ( .A(n27936), .B(n27937), .Z(n27935) );
  XNOR U27856 ( .A(n27934), .B(n27833), .Z(n27937) );
  XOR U27857 ( .A(n27938), .B(n27902), .Z(n27833) );
  XNOR U27858 ( .A(n27939), .B(n27909), .Z(n27902) );
  XOR U27859 ( .A(n27898), .B(n27897), .Z(n27909) );
  XNOR U27860 ( .A(n27940), .B(n27894), .Z(n27897) );
  XOR U27861 ( .A(n27941), .B(n27942), .Z(n27894) );
  AND U27862 ( .A(n27943), .B(n27944), .Z(n27942) );
  XNOR U27863 ( .A(n27945), .B(n27946), .Z(n27943) );
  IV U27864 ( .A(n27941), .Z(n27945) );
  XNOR U27865 ( .A(n27947), .B(n27948), .Z(n27940) );
  NOR U27866 ( .A(n27949), .B(n27950), .Z(n27948) );
  XNOR U27867 ( .A(n27947), .B(n27951), .Z(n27949) );
  XOR U27868 ( .A(n27952), .B(n27953), .Z(n27898) );
  NOR U27869 ( .A(n27954), .B(n27955), .Z(n27953) );
  XNOR U27870 ( .A(n27952), .B(n27956), .Z(n27954) );
  XNOR U27871 ( .A(n27908), .B(n27899), .Z(n27939) );
  XOR U27872 ( .A(n27957), .B(n27958), .Z(n27899) );
  AND U27873 ( .A(n27959), .B(n27960), .Z(n27958) );
  XOR U27874 ( .A(n27957), .B(n27961), .Z(n27959) );
  XOR U27875 ( .A(n27962), .B(n27914), .Z(n27908) );
  XOR U27876 ( .A(n27963), .B(n27964), .Z(n27914) );
  NOR U27877 ( .A(n27965), .B(n27966), .Z(n27964) );
  XOR U27878 ( .A(n27963), .B(n27967), .Z(n27965) );
  XNOR U27879 ( .A(n27913), .B(n27905), .Z(n27962) );
  XOR U27880 ( .A(n27968), .B(n27969), .Z(n27905) );
  AND U27881 ( .A(n27970), .B(n27971), .Z(n27969) );
  XOR U27882 ( .A(n27968), .B(n27972), .Z(n27970) );
  XNOR U27883 ( .A(n27973), .B(n27910), .Z(n27913) );
  XOR U27884 ( .A(n27974), .B(n27975), .Z(n27910) );
  AND U27885 ( .A(n27976), .B(n27977), .Z(n27975) );
  XNOR U27886 ( .A(n27978), .B(n27979), .Z(n27976) );
  IV U27887 ( .A(n27974), .Z(n27978) );
  XNOR U27888 ( .A(n27980), .B(n27981), .Z(n27973) );
  NOR U27889 ( .A(n27982), .B(n27983), .Z(n27981) );
  XNOR U27890 ( .A(n27980), .B(n27984), .Z(n27982) );
  XOR U27891 ( .A(n27903), .B(n27915), .Z(n27938) );
  NOR U27892 ( .A(n27841), .B(n27985), .Z(n27915) );
  XNOR U27893 ( .A(n27921), .B(n27920), .Z(n27903) );
  XNOR U27894 ( .A(n27986), .B(n27926), .Z(n27920) );
  XNOR U27895 ( .A(n27987), .B(n27988), .Z(n27926) );
  NOR U27896 ( .A(n27989), .B(n27990), .Z(n27988) );
  XOR U27897 ( .A(n27987), .B(n27991), .Z(n27989) );
  XNOR U27898 ( .A(n27925), .B(n27917), .Z(n27986) );
  XOR U27899 ( .A(n27992), .B(n27993), .Z(n27917) );
  AND U27900 ( .A(n27994), .B(n27995), .Z(n27993) );
  XOR U27901 ( .A(n27992), .B(n27996), .Z(n27994) );
  XNOR U27902 ( .A(n27997), .B(n27922), .Z(n27925) );
  XOR U27903 ( .A(n27998), .B(n27999), .Z(n27922) );
  AND U27904 ( .A(n28000), .B(n28001), .Z(n27999) );
  XNOR U27905 ( .A(n28002), .B(n28003), .Z(n28000) );
  IV U27906 ( .A(n27998), .Z(n28002) );
  XNOR U27907 ( .A(n28004), .B(n28005), .Z(n27997) );
  NOR U27908 ( .A(n28006), .B(n28007), .Z(n28005) );
  XNOR U27909 ( .A(n28004), .B(n28008), .Z(n28006) );
  XOR U27910 ( .A(n27931), .B(n27930), .Z(n27921) );
  XNOR U27911 ( .A(n28009), .B(n27927), .Z(n27930) );
  XOR U27912 ( .A(n28010), .B(n28011), .Z(n27927) );
  AND U27913 ( .A(n28012), .B(n28013), .Z(n28011) );
  XNOR U27914 ( .A(n28014), .B(n28015), .Z(n28012) );
  IV U27915 ( .A(n28010), .Z(n28014) );
  XNOR U27916 ( .A(n28016), .B(n28017), .Z(n28009) );
  NOR U27917 ( .A(n28018), .B(n28019), .Z(n28017) );
  XNOR U27918 ( .A(n28016), .B(n28020), .Z(n28018) );
  XOR U27919 ( .A(n28021), .B(n28022), .Z(n27931) );
  NOR U27920 ( .A(n28023), .B(n28024), .Z(n28022) );
  XNOR U27921 ( .A(n28021), .B(n28025), .Z(n28023) );
  XNOR U27922 ( .A(n27830), .B(n27934), .Z(n27936) );
  XNOR U27923 ( .A(n28026), .B(n28027), .Z(n27830) );
  AND U27924 ( .A(n518), .B(n27837), .Z(n28027) );
  XOR U27925 ( .A(n28026), .B(n27835), .Z(n27837) );
  AND U27926 ( .A(n27838), .B(n27841), .Z(n27934) );
  XOR U27927 ( .A(n28028), .B(n27985), .Z(n27841) );
  XNOR U27928 ( .A(p_input[1312]), .B(p_input[2048]), .Z(n27985) );
  XNOR U27929 ( .A(n27961), .B(n27960), .Z(n28028) );
  XNOR U27930 ( .A(n28029), .B(n27972), .Z(n27960) );
  XOR U27931 ( .A(n27946), .B(n27944), .Z(n27972) );
  XNOR U27932 ( .A(n28030), .B(n27951), .Z(n27944) );
  XOR U27933 ( .A(p_input[1336]), .B(p_input[2072]), .Z(n27951) );
  XOR U27934 ( .A(n27941), .B(n27950), .Z(n28030) );
  XOR U27935 ( .A(n28031), .B(n27947), .Z(n27950) );
  XOR U27936 ( .A(p_input[1334]), .B(p_input[2070]), .Z(n27947) );
  XOR U27937 ( .A(p_input[1335]), .B(n17295), .Z(n28031) );
  XOR U27938 ( .A(p_input[1330]), .B(p_input[2066]), .Z(n27941) );
  XNOR U27939 ( .A(n27956), .B(n27955), .Z(n27946) );
  XOR U27940 ( .A(n28032), .B(n27952), .Z(n27955) );
  XOR U27941 ( .A(p_input[1331]), .B(p_input[2067]), .Z(n27952) );
  XOR U27942 ( .A(p_input[1332]), .B(n17297), .Z(n28032) );
  XOR U27943 ( .A(p_input[1333]), .B(p_input[2069]), .Z(n27956) );
  XOR U27944 ( .A(n27971), .B(n28033), .Z(n28029) );
  IV U27945 ( .A(n27957), .Z(n28033) );
  XOR U27946 ( .A(p_input[1313]), .B(p_input[2049]), .Z(n27957) );
  XNOR U27947 ( .A(n28034), .B(n27979), .Z(n27971) );
  XNOR U27948 ( .A(n27967), .B(n27966), .Z(n27979) );
  XNOR U27949 ( .A(n28035), .B(n27963), .Z(n27966) );
  XNOR U27950 ( .A(p_input[1338]), .B(p_input[2074]), .Z(n27963) );
  XOR U27951 ( .A(p_input[1339]), .B(n17300), .Z(n28035) );
  XOR U27952 ( .A(p_input[1340]), .B(p_input[2076]), .Z(n27967) );
  XOR U27953 ( .A(n27977), .B(n28036), .Z(n28034) );
  IV U27954 ( .A(n27968), .Z(n28036) );
  XOR U27955 ( .A(p_input[1329]), .B(p_input[2065]), .Z(n27968) );
  XNOR U27956 ( .A(n28037), .B(n27984), .Z(n27977) );
  XNOR U27957 ( .A(p_input[1343]), .B(n17303), .Z(n27984) );
  XOR U27958 ( .A(n27974), .B(n27983), .Z(n28037) );
  XOR U27959 ( .A(n28038), .B(n27980), .Z(n27983) );
  XOR U27960 ( .A(p_input[1341]), .B(p_input[2077]), .Z(n27980) );
  XOR U27961 ( .A(p_input[1342]), .B(n17305), .Z(n28038) );
  XOR U27962 ( .A(p_input[1337]), .B(p_input[2073]), .Z(n27974) );
  XOR U27963 ( .A(n27996), .B(n27995), .Z(n27961) );
  XNOR U27964 ( .A(n28039), .B(n28003), .Z(n27995) );
  XNOR U27965 ( .A(n27991), .B(n27990), .Z(n28003) );
  XNOR U27966 ( .A(n28040), .B(n27987), .Z(n27990) );
  XNOR U27967 ( .A(p_input[1323]), .B(p_input[2059]), .Z(n27987) );
  XOR U27968 ( .A(p_input[1324]), .B(n16451), .Z(n28040) );
  XOR U27969 ( .A(p_input[1325]), .B(p_input[2061]), .Z(n27991) );
  XOR U27970 ( .A(n28001), .B(n28041), .Z(n28039) );
  IV U27971 ( .A(n27992), .Z(n28041) );
  XOR U27972 ( .A(p_input[1314]), .B(p_input[2050]), .Z(n27992) );
  XNOR U27973 ( .A(n28042), .B(n28008), .Z(n28001) );
  XNOR U27974 ( .A(p_input[1328]), .B(n16454), .Z(n28008) );
  XOR U27975 ( .A(n27998), .B(n28007), .Z(n28042) );
  XOR U27976 ( .A(n28043), .B(n28004), .Z(n28007) );
  XOR U27977 ( .A(p_input[1326]), .B(p_input[2062]), .Z(n28004) );
  XOR U27978 ( .A(p_input[1327]), .B(n16456), .Z(n28043) );
  XOR U27979 ( .A(p_input[1322]), .B(p_input[2058]), .Z(n27998) );
  XOR U27980 ( .A(n28015), .B(n28013), .Z(n27996) );
  XNOR U27981 ( .A(n28044), .B(n28020), .Z(n28013) );
  XOR U27982 ( .A(p_input[1321]), .B(p_input[2057]), .Z(n28020) );
  XOR U27983 ( .A(n28010), .B(n28019), .Z(n28044) );
  XOR U27984 ( .A(n28045), .B(n28016), .Z(n28019) );
  XOR U27985 ( .A(p_input[1319]), .B(p_input[2055]), .Z(n28016) );
  XOR U27986 ( .A(p_input[1320]), .B(n17312), .Z(n28045) );
  XOR U27987 ( .A(p_input[1315]), .B(p_input[2051]), .Z(n28010) );
  XNOR U27988 ( .A(n28025), .B(n28024), .Z(n28015) );
  XOR U27989 ( .A(n28046), .B(n28021), .Z(n28024) );
  XOR U27990 ( .A(p_input[1316]), .B(p_input[2052]), .Z(n28021) );
  XOR U27991 ( .A(p_input[1317]), .B(n17314), .Z(n28046) );
  XOR U27992 ( .A(p_input[1318]), .B(p_input[2054]), .Z(n28025) );
  XNOR U27993 ( .A(n28047), .B(n28048), .Z(n27838) );
  AND U27994 ( .A(n518), .B(n28049), .Z(n28048) );
  XNOR U27995 ( .A(n28050), .B(n28051), .Z(n518) );
  AND U27996 ( .A(n28052), .B(n28053), .Z(n28051) );
  XOR U27997 ( .A(n28050), .B(n27848), .Z(n28053) );
  XNOR U27998 ( .A(n28050), .B(n27790), .Z(n28052) );
  XOR U27999 ( .A(n28054), .B(n28055), .Z(n28050) );
  AND U28000 ( .A(n28056), .B(n28057), .Z(n28055) );
  XNOR U28001 ( .A(n27861), .B(n28054), .Z(n28057) );
  XOR U28002 ( .A(n28054), .B(n27802), .Z(n28056) );
  XOR U28003 ( .A(n28058), .B(n28059), .Z(n28054) );
  AND U28004 ( .A(n28060), .B(n28061), .Z(n28059) );
  XNOR U28005 ( .A(n27886), .B(n28058), .Z(n28061) );
  XOR U28006 ( .A(n28058), .B(n27813), .Z(n28060) );
  XOR U28007 ( .A(n28062), .B(n28063), .Z(n28058) );
  AND U28008 ( .A(n28064), .B(n28065), .Z(n28063) );
  XOR U28009 ( .A(n28062), .B(n27823), .Z(n28064) );
  XOR U28010 ( .A(n28066), .B(n28067), .Z(n27779) );
  AND U28011 ( .A(n522), .B(n28049), .Z(n28067) );
  XNOR U28012 ( .A(n28047), .B(n28066), .Z(n28049) );
  XNOR U28013 ( .A(n28068), .B(n28069), .Z(n522) );
  AND U28014 ( .A(n28070), .B(n28071), .Z(n28069) );
  XNOR U28015 ( .A(n28072), .B(n28068), .Z(n28071) );
  IV U28016 ( .A(n27848), .Z(n28072) );
  XNOR U28017 ( .A(n28073), .B(n28074), .Z(n27848) );
  AND U28018 ( .A(n525), .B(n28075), .Z(n28074) );
  XNOR U28019 ( .A(n28073), .B(n28076), .Z(n28075) );
  XNOR U28020 ( .A(n27790), .B(n28068), .Z(n28070) );
  XOR U28021 ( .A(n28077), .B(n28078), .Z(n27790) );
  AND U28022 ( .A(n533), .B(n28079), .Z(n28078) );
  XOR U28023 ( .A(n28080), .B(n28081), .Z(n28068) );
  AND U28024 ( .A(n28082), .B(n28083), .Z(n28081) );
  XNOR U28025 ( .A(n28080), .B(n27861), .Z(n28083) );
  XNOR U28026 ( .A(n28084), .B(n28085), .Z(n27861) );
  AND U28027 ( .A(n525), .B(n28086), .Z(n28085) );
  XOR U28028 ( .A(n28087), .B(n28084), .Z(n28086) );
  XNOR U28029 ( .A(n28088), .B(n28080), .Z(n28082) );
  IV U28030 ( .A(n27802), .Z(n28088) );
  XOR U28031 ( .A(n28089), .B(n28090), .Z(n27802) );
  AND U28032 ( .A(n533), .B(n28091), .Z(n28090) );
  XOR U28033 ( .A(n28092), .B(n28093), .Z(n28080) );
  AND U28034 ( .A(n28094), .B(n28095), .Z(n28093) );
  XNOR U28035 ( .A(n28092), .B(n27886), .Z(n28095) );
  XNOR U28036 ( .A(n28096), .B(n28097), .Z(n27886) );
  AND U28037 ( .A(n525), .B(n28098), .Z(n28097) );
  XNOR U28038 ( .A(n28099), .B(n28096), .Z(n28098) );
  XOR U28039 ( .A(n27813), .B(n28092), .Z(n28094) );
  XOR U28040 ( .A(n28100), .B(n28101), .Z(n27813) );
  AND U28041 ( .A(n533), .B(n28102), .Z(n28101) );
  XOR U28042 ( .A(n28062), .B(n28103), .Z(n28092) );
  AND U28043 ( .A(n28104), .B(n28065), .Z(n28103) );
  XNOR U28044 ( .A(n27932), .B(n28062), .Z(n28065) );
  XNOR U28045 ( .A(n28105), .B(n28106), .Z(n27932) );
  AND U28046 ( .A(n525), .B(n28107), .Z(n28106) );
  XOR U28047 ( .A(n28108), .B(n28105), .Z(n28107) );
  XNOR U28048 ( .A(n28109), .B(n28062), .Z(n28104) );
  IV U28049 ( .A(n27823), .Z(n28109) );
  XOR U28050 ( .A(n28110), .B(n28111), .Z(n27823) );
  AND U28051 ( .A(n533), .B(n28112), .Z(n28111) );
  XOR U28052 ( .A(n28113), .B(n28114), .Z(n28062) );
  AND U28053 ( .A(n28115), .B(n28116), .Z(n28114) );
  XNOR U28054 ( .A(n28113), .B(n28026), .Z(n28116) );
  XNOR U28055 ( .A(n28117), .B(n28118), .Z(n28026) );
  AND U28056 ( .A(n525), .B(n28119), .Z(n28118) );
  XNOR U28057 ( .A(n28120), .B(n28117), .Z(n28119) );
  XNOR U28058 ( .A(n28121), .B(n28113), .Z(n28115) );
  IV U28059 ( .A(n27835), .Z(n28121) );
  XOR U28060 ( .A(n28122), .B(n28123), .Z(n27835) );
  AND U28061 ( .A(n533), .B(n28124), .Z(n28123) );
  AND U28062 ( .A(n28066), .B(n28047), .Z(n28113) );
  XNOR U28063 ( .A(n28125), .B(n28126), .Z(n28047) );
  AND U28064 ( .A(n525), .B(n28127), .Z(n28126) );
  XNOR U28065 ( .A(n28128), .B(n28125), .Z(n28127) );
  XNOR U28066 ( .A(n28129), .B(n28130), .Z(n525) );
  AND U28067 ( .A(n28131), .B(n28132), .Z(n28130) );
  XOR U28068 ( .A(n28076), .B(n28129), .Z(n28132) );
  AND U28069 ( .A(n28133), .B(n28134), .Z(n28076) );
  XOR U28070 ( .A(n28129), .B(n28073), .Z(n28131) );
  XNOR U28071 ( .A(n28135), .B(n28136), .Z(n28073) );
  AND U28072 ( .A(n529), .B(n28079), .Z(n28136) );
  XOR U28073 ( .A(n28077), .B(n28135), .Z(n28079) );
  XOR U28074 ( .A(n28137), .B(n28138), .Z(n28129) );
  AND U28075 ( .A(n28139), .B(n28140), .Z(n28138) );
  XNOR U28076 ( .A(n28137), .B(n28133), .Z(n28140) );
  IV U28077 ( .A(n28087), .Z(n28133) );
  XOR U28078 ( .A(n28141), .B(n28142), .Z(n28087) );
  XOR U28079 ( .A(n28143), .B(n28134), .Z(n28142) );
  AND U28080 ( .A(n28099), .B(n28144), .Z(n28134) );
  AND U28081 ( .A(n28145), .B(n28146), .Z(n28143) );
  XOR U28082 ( .A(n28147), .B(n28141), .Z(n28145) );
  XNOR U28083 ( .A(n28084), .B(n28137), .Z(n28139) );
  XNOR U28084 ( .A(n28148), .B(n28149), .Z(n28084) );
  AND U28085 ( .A(n529), .B(n28091), .Z(n28149) );
  XOR U28086 ( .A(n28148), .B(n28089), .Z(n28091) );
  XOR U28087 ( .A(n28150), .B(n28151), .Z(n28137) );
  AND U28088 ( .A(n28152), .B(n28153), .Z(n28151) );
  XNOR U28089 ( .A(n28150), .B(n28099), .Z(n28153) );
  XOR U28090 ( .A(n28154), .B(n28146), .Z(n28099) );
  XNOR U28091 ( .A(n28155), .B(n28141), .Z(n28146) );
  XOR U28092 ( .A(n28156), .B(n28157), .Z(n28141) );
  AND U28093 ( .A(n28158), .B(n28159), .Z(n28157) );
  XOR U28094 ( .A(n28160), .B(n28156), .Z(n28158) );
  XNOR U28095 ( .A(n28161), .B(n28162), .Z(n28155) );
  AND U28096 ( .A(n28163), .B(n28164), .Z(n28162) );
  XOR U28097 ( .A(n28161), .B(n28165), .Z(n28163) );
  XNOR U28098 ( .A(n28147), .B(n28144), .Z(n28154) );
  AND U28099 ( .A(n28166), .B(n28167), .Z(n28144) );
  XOR U28100 ( .A(n28168), .B(n28169), .Z(n28147) );
  AND U28101 ( .A(n28170), .B(n28171), .Z(n28169) );
  XOR U28102 ( .A(n28168), .B(n28172), .Z(n28170) );
  XNOR U28103 ( .A(n28096), .B(n28150), .Z(n28152) );
  XNOR U28104 ( .A(n28173), .B(n28174), .Z(n28096) );
  AND U28105 ( .A(n529), .B(n28102), .Z(n28174) );
  XOR U28106 ( .A(n28173), .B(n28100), .Z(n28102) );
  XOR U28107 ( .A(n28175), .B(n28176), .Z(n28150) );
  AND U28108 ( .A(n28177), .B(n28178), .Z(n28176) );
  XNOR U28109 ( .A(n28175), .B(n28166), .Z(n28178) );
  IV U28110 ( .A(n28108), .Z(n28166) );
  XNOR U28111 ( .A(n28179), .B(n28159), .Z(n28108) );
  XNOR U28112 ( .A(n28180), .B(n28165), .Z(n28159) );
  XOR U28113 ( .A(n28181), .B(n28182), .Z(n28165) );
  AND U28114 ( .A(n28183), .B(n28184), .Z(n28182) );
  XOR U28115 ( .A(n28181), .B(n28185), .Z(n28183) );
  XNOR U28116 ( .A(n28164), .B(n28156), .Z(n28180) );
  XOR U28117 ( .A(n28186), .B(n28187), .Z(n28156) );
  AND U28118 ( .A(n28188), .B(n28189), .Z(n28187) );
  XNOR U28119 ( .A(n28190), .B(n28186), .Z(n28188) );
  XNOR U28120 ( .A(n28191), .B(n28161), .Z(n28164) );
  XOR U28121 ( .A(n28192), .B(n28193), .Z(n28161) );
  AND U28122 ( .A(n28194), .B(n28195), .Z(n28193) );
  XOR U28123 ( .A(n28192), .B(n28196), .Z(n28194) );
  XNOR U28124 ( .A(n28197), .B(n28198), .Z(n28191) );
  AND U28125 ( .A(n28199), .B(n28200), .Z(n28198) );
  XNOR U28126 ( .A(n28197), .B(n28201), .Z(n28199) );
  XNOR U28127 ( .A(n28160), .B(n28167), .Z(n28179) );
  AND U28128 ( .A(n28120), .B(n28202), .Z(n28167) );
  XOR U28129 ( .A(n28172), .B(n28171), .Z(n28160) );
  XNOR U28130 ( .A(n28203), .B(n28168), .Z(n28171) );
  XOR U28131 ( .A(n28204), .B(n28205), .Z(n28168) );
  AND U28132 ( .A(n28206), .B(n28207), .Z(n28205) );
  XOR U28133 ( .A(n28204), .B(n28208), .Z(n28206) );
  XNOR U28134 ( .A(n28209), .B(n28210), .Z(n28203) );
  AND U28135 ( .A(n28211), .B(n28212), .Z(n28210) );
  XOR U28136 ( .A(n28209), .B(n28213), .Z(n28211) );
  XOR U28137 ( .A(n28214), .B(n28215), .Z(n28172) );
  AND U28138 ( .A(n28216), .B(n28217), .Z(n28215) );
  XOR U28139 ( .A(n28214), .B(n28218), .Z(n28216) );
  XNOR U28140 ( .A(n28105), .B(n28175), .Z(n28177) );
  XNOR U28141 ( .A(n28219), .B(n28220), .Z(n28105) );
  AND U28142 ( .A(n529), .B(n28112), .Z(n28220) );
  XOR U28143 ( .A(n28219), .B(n28110), .Z(n28112) );
  XOR U28144 ( .A(n28221), .B(n28222), .Z(n28175) );
  AND U28145 ( .A(n28223), .B(n28224), .Z(n28222) );
  XNOR U28146 ( .A(n28221), .B(n28120), .Z(n28224) );
  XOR U28147 ( .A(n28225), .B(n28189), .Z(n28120) );
  XNOR U28148 ( .A(n28226), .B(n28196), .Z(n28189) );
  XOR U28149 ( .A(n28185), .B(n28184), .Z(n28196) );
  XNOR U28150 ( .A(n28227), .B(n28181), .Z(n28184) );
  XOR U28151 ( .A(n28228), .B(n28229), .Z(n28181) );
  AND U28152 ( .A(n28230), .B(n28231), .Z(n28229) );
  XNOR U28153 ( .A(n28232), .B(n28233), .Z(n28230) );
  IV U28154 ( .A(n28228), .Z(n28232) );
  XNOR U28155 ( .A(n28234), .B(n28235), .Z(n28227) );
  NOR U28156 ( .A(n28236), .B(n28237), .Z(n28235) );
  XNOR U28157 ( .A(n28234), .B(n28238), .Z(n28236) );
  XOR U28158 ( .A(n28239), .B(n28240), .Z(n28185) );
  NOR U28159 ( .A(n28241), .B(n28242), .Z(n28240) );
  XNOR U28160 ( .A(n28239), .B(n28243), .Z(n28241) );
  XNOR U28161 ( .A(n28195), .B(n28186), .Z(n28226) );
  XOR U28162 ( .A(n28244), .B(n28245), .Z(n28186) );
  AND U28163 ( .A(n28246), .B(n28247), .Z(n28245) );
  XOR U28164 ( .A(n28244), .B(n28248), .Z(n28246) );
  XOR U28165 ( .A(n28249), .B(n28201), .Z(n28195) );
  XOR U28166 ( .A(n28250), .B(n28251), .Z(n28201) );
  NOR U28167 ( .A(n28252), .B(n28253), .Z(n28251) );
  XOR U28168 ( .A(n28250), .B(n28254), .Z(n28252) );
  XNOR U28169 ( .A(n28200), .B(n28192), .Z(n28249) );
  XOR U28170 ( .A(n28255), .B(n28256), .Z(n28192) );
  AND U28171 ( .A(n28257), .B(n28258), .Z(n28256) );
  XOR U28172 ( .A(n28255), .B(n28259), .Z(n28257) );
  XNOR U28173 ( .A(n28260), .B(n28197), .Z(n28200) );
  XOR U28174 ( .A(n28261), .B(n28262), .Z(n28197) );
  AND U28175 ( .A(n28263), .B(n28264), .Z(n28262) );
  XNOR U28176 ( .A(n28265), .B(n28266), .Z(n28263) );
  IV U28177 ( .A(n28261), .Z(n28265) );
  XNOR U28178 ( .A(n28267), .B(n28268), .Z(n28260) );
  NOR U28179 ( .A(n28269), .B(n28270), .Z(n28268) );
  XNOR U28180 ( .A(n28267), .B(n28271), .Z(n28269) );
  XOR U28181 ( .A(n28190), .B(n28202), .Z(n28225) );
  NOR U28182 ( .A(n28128), .B(n28272), .Z(n28202) );
  XNOR U28183 ( .A(n28208), .B(n28207), .Z(n28190) );
  XNOR U28184 ( .A(n28273), .B(n28213), .Z(n28207) );
  XNOR U28185 ( .A(n28274), .B(n28275), .Z(n28213) );
  NOR U28186 ( .A(n28276), .B(n28277), .Z(n28275) );
  XOR U28187 ( .A(n28274), .B(n28278), .Z(n28276) );
  XNOR U28188 ( .A(n28212), .B(n28204), .Z(n28273) );
  XOR U28189 ( .A(n28279), .B(n28280), .Z(n28204) );
  AND U28190 ( .A(n28281), .B(n28282), .Z(n28280) );
  XOR U28191 ( .A(n28279), .B(n28283), .Z(n28281) );
  XNOR U28192 ( .A(n28284), .B(n28209), .Z(n28212) );
  XOR U28193 ( .A(n28285), .B(n28286), .Z(n28209) );
  AND U28194 ( .A(n28287), .B(n28288), .Z(n28286) );
  XNOR U28195 ( .A(n28289), .B(n28290), .Z(n28287) );
  IV U28196 ( .A(n28285), .Z(n28289) );
  XNOR U28197 ( .A(n28291), .B(n28292), .Z(n28284) );
  NOR U28198 ( .A(n28293), .B(n28294), .Z(n28292) );
  XNOR U28199 ( .A(n28291), .B(n28295), .Z(n28293) );
  XOR U28200 ( .A(n28218), .B(n28217), .Z(n28208) );
  XNOR U28201 ( .A(n28296), .B(n28214), .Z(n28217) );
  XOR U28202 ( .A(n28297), .B(n28298), .Z(n28214) );
  AND U28203 ( .A(n28299), .B(n28300), .Z(n28298) );
  XNOR U28204 ( .A(n28301), .B(n28302), .Z(n28299) );
  IV U28205 ( .A(n28297), .Z(n28301) );
  XNOR U28206 ( .A(n28303), .B(n28304), .Z(n28296) );
  NOR U28207 ( .A(n28305), .B(n28306), .Z(n28304) );
  XNOR U28208 ( .A(n28303), .B(n28307), .Z(n28305) );
  XOR U28209 ( .A(n28308), .B(n28309), .Z(n28218) );
  NOR U28210 ( .A(n28310), .B(n28311), .Z(n28309) );
  XNOR U28211 ( .A(n28308), .B(n28312), .Z(n28310) );
  XNOR U28212 ( .A(n28117), .B(n28221), .Z(n28223) );
  XNOR U28213 ( .A(n28313), .B(n28314), .Z(n28117) );
  AND U28214 ( .A(n529), .B(n28124), .Z(n28314) );
  XOR U28215 ( .A(n28313), .B(n28122), .Z(n28124) );
  AND U28216 ( .A(n28125), .B(n28128), .Z(n28221) );
  XOR U28217 ( .A(n28315), .B(n28272), .Z(n28128) );
  XNOR U28218 ( .A(p_input[1344]), .B(p_input[2048]), .Z(n28272) );
  XNOR U28219 ( .A(n28248), .B(n28247), .Z(n28315) );
  XNOR U28220 ( .A(n28316), .B(n28259), .Z(n28247) );
  XOR U28221 ( .A(n28233), .B(n28231), .Z(n28259) );
  XNOR U28222 ( .A(n28317), .B(n28238), .Z(n28231) );
  XOR U28223 ( .A(p_input[1368]), .B(p_input[2072]), .Z(n28238) );
  XOR U28224 ( .A(n28228), .B(n28237), .Z(n28317) );
  XOR U28225 ( .A(n28318), .B(n28234), .Z(n28237) );
  XOR U28226 ( .A(p_input[1366]), .B(p_input[2070]), .Z(n28234) );
  XOR U28227 ( .A(p_input[1367]), .B(n17295), .Z(n28318) );
  XOR U28228 ( .A(p_input[1362]), .B(p_input[2066]), .Z(n28228) );
  XNOR U28229 ( .A(n28243), .B(n28242), .Z(n28233) );
  XOR U28230 ( .A(n28319), .B(n28239), .Z(n28242) );
  XOR U28231 ( .A(p_input[1363]), .B(p_input[2067]), .Z(n28239) );
  XOR U28232 ( .A(p_input[1364]), .B(n17297), .Z(n28319) );
  XOR U28233 ( .A(p_input[1365]), .B(p_input[2069]), .Z(n28243) );
  XOR U28234 ( .A(n28258), .B(n28320), .Z(n28316) );
  IV U28235 ( .A(n28244), .Z(n28320) );
  XOR U28236 ( .A(p_input[1345]), .B(p_input[2049]), .Z(n28244) );
  XNOR U28237 ( .A(n28321), .B(n28266), .Z(n28258) );
  XNOR U28238 ( .A(n28254), .B(n28253), .Z(n28266) );
  XNOR U28239 ( .A(n28322), .B(n28250), .Z(n28253) );
  XNOR U28240 ( .A(p_input[1370]), .B(p_input[2074]), .Z(n28250) );
  XOR U28241 ( .A(p_input[1371]), .B(n17300), .Z(n28322) );
  XOR U28242 ( .A(p_input[1372]), .B(p_input[2076]), .Z(n28254) );
  XOR U28243 ( .A(n28264), .B(n28323), .Z(n28321) );
  IV U28244 ( .A(n28255), .Z(n28323) );
  XOR U28245 ( .A(p_input[1361]), .B(p_input[2065]), .Z(n28255) );
  XNOR U28246 ( .A(n28324), .B(n28271), .Z(n28264) );
  XNOR U28247 ( .A(p_input[1375]), .B(n17303), .Z(n28271) );
  XOR U28248 ( .A(n28261), .B(n28270), .Z(n28324) );
  XOR U28249 ( .A(n28325), .B(n28267), .Z(n28270) );
  XOR U28250 ( .A(p_input[1373]), .B(p_input[2077]), .Z(n28267) );
  XOR U28251 ( .A(p_input[1374]), .B(n17305), .Z(n28325) );
  XOR U28252 ( .A(p_input[1369]), .B(p_input[2073]), .Z(n28261) );
  XOR U28253 ( .A(n28283), .B(n28282), .Z(n28248) );
  XNOR U28254 ( .A(n28326), .B(n28290), .Z(n28282) );
  XNOR U28255 ( .A(n28278), .B(n28277), .Z(n28290) );
  XNOR U28256 ( .A(n28327), .B(n28274), .Z(n28277) );
  XNOR U28257 ( .A(p_input[1355]), .B(p_input[2059]), .Z(n28274) );
  XOR U28258 ( .A(p_input[1356]), .B(n16451), .Z(n28327) );
  XOR U28259 ( .A(p_input[1357]), .B(p_input[2061]), .Z(n28278) );
  XOR U28260 ( .A(n28288), .B(n28328), .Z(n28326) );
  IV U28261 ( .A(n28279), .Z(n28328) );
  XOR U28262 ( .A(p_input[1346]), .B(p_input[2050]), .Z(n28279) );
  XNOR U28263 ( .A(n28329), .B(n28295), .Z(n28288) );
  XNOR U28264 ( .A(p_input[1360]), .B(n16454), .Z(n28295) );
  XOR U28265 ( .A(n28285), .B(n28294), .Z(n28329) );
  XOR U28266 ( .A(n28330), .B(n28291), .Z(n28294) );
  XOR U28267 ( .A(p_input[1358]), .B(p_input[2062]), .Z(n28291) );
  XOR U28268 ( .A(p_input[1359]), .B(n16456), .Z(n28330) );
  XOR U28269 ( .A(p_input[1354]), .B(p_input[2058]), .Z(n28285) );
  XOR U28270 ( .A(n28302), .B(n28300), .Z(n28283) );
  XNOR U28271 ( .A(n28331), .B(n28307), .Z(n28300) );
  XOR U28272 ( .A(p_input[1353]), .B(p_input[2057]), .Z(n28307) );
  XOR U28273 ( .A(n28297), .B(n28306), .Z(n28331) );
  XOR U28274 ( .A(n28332), .B(n28303), .Z(n28306) );
  XOR U28275 ( .A(p_input[1351]), .B(p_input[2055]), .Z(n28303) );
  XOR U28276 ( .A(p_input[1352]), .B(n17312), .Z(n28332) );
  XOR U28277 ( .A(p_input[1347]), .B(p_input[2051]), .Z(n28297) );
  XNOR U28278 ( .A(n28312), .B(n28311), .Z(n28302) );
  XOR U28279 ( .A(n28333), .B(n28308), .Z(n28311) );
  XOR U28280 ( .A(p_input[1348]), .B(p_input[2052]), .Z(n28308) );
  XOR U28281 ( .A(p_input[1349]), .B(n17314), .Z(n28333) );
  XOR U28282 ( .A(p_input[1350]), .B(p_input[2054]), .Z(n28312) );
  XNOR U28283 ( .A(n28334), .B(n28335), .Z(n28125) );
  AND U28284 ( .A(n529), .B(n28336), .Z(n28335) );
  XNOR U28285 ( .A(n28337), .B(n28338), .Z(n529) );
  AND U28286 ( .A(n28339), .B(n28340), .Z(n28338) );
  XOR U28287 ( .A(n28337), .B(n28135), .Z(n28340) );
  XNOR U28288 ( .A(n28337), .B(n28077), .Z(n28339) );
  XOR U28289 ( .A(n28341), .B(n28342), .Z(n28337) );
  AND U28290 ( .A(n28343), .B(n28344), .Z(n28342) );
  XNOR U28291 ( .A(n28148), .B(n28341), .Z(n28344) );
  XOR U28292 ( .A(n28341), .B(n28089), .Z(n28343) );
  XOR U28293 ( .A(n28345), .B(n28346), .Z(n28341) );
  AND U28294 ( .A(n28347), .B(n28348), .Z(n28346) );
  XNOR U28295 ( .A(n28173), .B(n28345), .Z(n28348) );
  XOR U28296 ( .A(n28345), .B(n28100), .Z(n28347) );
  XOR U28297 ( .A(n28349), .B(n28350), .Z(n28345) );
  AND U28298 ( .A(n28351), .B(n28352), .Z(n28350) );
  XOR U28299 ( .A(n28349), .B(n28110), .Z(n28351) );
  XOR U28300 ( .A(n28353), .B(n28354), .Z(n28066) );
  AND U28301 ( .A(n533), .B(n28336), .Z(n28354) );
  XNOR U28302 ( .A(n28334), .B(n28353), .Z(n28336) );
  XNOR U28303 ( .A(n28355), .B(n28356), .Z(n533) );
  AND U28304 ( .A(n28357), .B(n28358), .Z(n28356) );
  XNOR U28305 ( .A(n28359), .B(n28355), .Z(n28358) );
  IV U28306 ( .A(n28135), .Z(n28359) );
  XNOR U28307 ( .A(n28360), .B(n28361), .Z(n28135) );
  AND U28308 ( .A(n536), .B(n28362), .Z(n28361) );
  XNOR U28309 ( .A(n28360), .B(n28363), .Z(n28362) );
  XNOR U28310 ( .A(n28077), .B(n28355), .Z(n28357) );
  XOR U28311 ( .A(n28364), .B(n28365), .Z(n28077) );
  AND U28312 ( .A(n544), .B(n28366), .Z(n28365) );
  XOR U28313 ( .A(n28367), .B(n28368), .Z(n28355) );
  AND U28314 ( .A(n28369), .B(n28370), .Z(n28368) );
  XNOR U28315 ( .A(n28367), .B(n28148), .Z(n28370) );
  XNOR U28316 ( .A(n28371), .B(n28372), .Z(n28148) );
  AND U28317 ( .A(n536), .B(n28373), .Z(n28372) );
  XOR U28318 ( .A(n28374), .B(n28371), .Z(n28373) );
  XNOR U28319 ( .A(n28375), .B(n28367), .Z(n28369) );
  IV U28320 ( .A(n28089), .Z(n28375) );
  XOR U28321 ( .A(n28376), .B(n28377), .Z(n28089) );
  AND U28322 ( .A(n544), .B(n28378), .Z(n28377) );
  XOR U28323 ( .A(n28379), .B(n28380), .Z(n28367) );
  AND U28324 ( .A(n28381), .B(n28382), .Z(n28380) );
  XNOR U28325 ( .A(n28379), .B(n28173), .Z(n28382) );
  XNOR U28326 ( .A(n28383), .B(n28384), .Z(n28173) );
  AND U28327 ( .A(n536), .B(n28385), .Z(n28384) );
  XNOR U28328 ( .A(n28386), .B(n28383), .Z(n28385) );
  XOR U28329 ( .A(n28100), .B(n28379), .Z(n28381) );
  XOR U28330 ( .A(n28387), .B(n28388), .Z(n28100) );
  AND U28331 ( .A(n544), .B(n28389), .Z(n28388) );
  XOR U28332 ( .A(n28349), .B(n28390), .Z(n28379) );
  AND U28333 ( .A(n28391), .B(n28352), .Z(n28390) );
  XNOR U28334 ( .A(n28219), .B(n28349), .Z(n28352) );
  XNOR U28335 ( .A(n28392), .B(n28393), .Z(n28219) );
  AND U28336 ( .A(n536), .B(n28394), .Z(n28393) );
  XOR U28337 ( .A(n28395), .B(n28392), .Z(n28394) );
  XNOR U28338 ( .A(n28396), .B(n28349), .Z(n28391) );
  IV U28339 ( .A(n28110), .Z(n28396) );
  XOR U28340 ( .A(n28397), .B(n28398), .Z(n28110) );
  AND U28341 ( .A(n544), .B(n28399), .Z(n28398) );
  XOR U28342 ( .A(n28400), .B(n28401), .Z(n28349) );
  AND U28343 ( .A(n28402), .B(n28403), .Z(n28401) );
  XNOR U28344 ( .A(n28400), .B(n28313), .Z(n28403) );
  XNOR U28345 ( .A(n28404), .B(n28405), .Z(n28313) );
  AND U28346 ( .A(n536), .B(n28406), .Z(n28405) );
  XNOR U28347 ( .A(n28407), .B(n28404), .Z(n28406) );
  XNOR U28348 ( .A(n28408), .B(n28400), .Z(n28402) );
  IV U28349 ( .A(n28122), .Z(n28408) );
  XOR U28350 ( .A(n28409), .B(n28410), .Z(n28122) );
  AND U28351 ( .A(n544), .B(n28411), .Z(n28410) );
  AND U28352 ( .A(n28353), .B(n28334), .Z(n28400) );
  XNOR U28353 ( .A(n28412), .B(n28413), .Z(n28334) );
  AND U28354 ( .A(n536), .B(n28414), .Z(n28413) );
  XNOR U28355 ( .A(n28415), .B(n28412), .Z(n28414) );
  XNOR U28356 ( .A(n28416), .B(n28417), .Z(n536) );
  AND U28357 ( .A(n28418), .B(n28419), .Z(n28417) );
  XOR U28358 ( .A(n28363), .B(n28416), .Z(n28419) );
  AND U28359 ( .A(n28420), .B(n28421), .Z(n28363) );
  XOR U28360 ( .A(n28416), .B(n28360), .Z(n28418) );
  XNOR U28361 ( .A(n28422), .B(n28423), .Z(n28360) );
  AND U28362 ( .A(n540), .B(n28366), .Z(n28423) );
  XOR U28363 ( .A(n28364), .B(n28422), .Z(n28366) );
  XOR U28364 ( .A(n28424), .B(n28425), .Z(n28416) );
  AND U28365 ( .A(n28426), .B(n28427), .Z(n28425) );
  XNOR U28366 ( .A(n28424), .B(n28420), .Z(n28427) );
  IV U28367 ( .A(n28374), .Z(n28420) );
  XOR U28368 ( .A(n28428), .B(n28429), .Z(n28374) );
  XOR U28369 ( .A(n28430), .B(n28421), .Z(n28429) );
  AND U28370 ( .A(n28386), .B(n28431), .Z(n28421) );
  AND U28371 ( .A(n28432), .B(n28433), .Z(n28430) );
  XOR U28372 ( .A(n28434), .B(n28428), .Z(n28432) );
  XNOR U28373 ( .A(n28371), .B(n28424), .Z(n28426) );
  XNOR U28374 ( .A(n28435), .B(n28436), .Z(n28371) );
  AND U28375 ( .A(n540), .B(n28378), .Z(n28436) );
  XOR U28376 ( .A(n28435), .B(n28376), .Z(n28378) );
  XOR U28377 ( .A(n28437), .B(n28438), .Z(n28424) );
  AND U28378 ( .A(n28439), .B(n28440), .Z(n28438) );
  XNOR U28379 ( .A(n28437), .B(n28386), .Z(n28440) );
  XOR U28380 ( .A(n28441), .B(n28433), .Z(n28386) );
  XNOR U28381 ( .A(n28442), .B(n28428), .Z(n28433) );
  XOR U28382 ( .A(n28443), .B(n28444), .Z(n28428) );
  AND U28383 ( .A(n28445), .B(n28446), .Z(n28444) );
  XOR U28384 ( .A(n28447), .B(n28443), .Z(n28445) );
  XNOR U28385 ( .A(n28448), .B(n28449), .Z(n28442) );
  AND U28386 ( .A(n28450), .B(n28451), .Z(n28449) );
  XOR U28387 ( .A(n28448), .B(n28452), .Z(n28450) );
  XNOR U28388 ( .A(n28434), .B(n28431), .Z(n28441) );
  AND U28389 ( .A(n28453), .B(n28454), .Z(n28431) );
  XOR U28390 ( .A(n28455), .B(n28456), .Z(n28434) );
  AND U28391 ( .A(n28457), .B(n28458), .Z(n28456) );
  XOR U28392 ( .A(n28455), .B(n28459), .Z(n28457) );
  XNOR U28393 ( .A(n28383), .B(n28437), .Z(n28439) );
  XNOR U28394 ( .A(n28460), .B(n28461), .Z(n28383) );
  AND U28395 ( .A(n540), .B(n28389), .Z(n28461) );
  XOR U28396 ( .A(n28460), .B(n28387), .Z(n28389) );
  XOR U28397 ( .A(n28462), .B(n28463), .Z(n28437) );
  AND U28398 ( .A(n28464), .B(n28465), .Z(n28463) );
  XNOR U28399 ( .A(n28462), .B(n28453), .Z(n28465) );
  IV U28400 ( .A(n28395), .Z(n28453) );
  XNOR U28401 ( .A(n28466), .B(n28446), .Z(n28395) );
  XNOR U28402 ( .A(n28467), .B(n28452), .Z(n28446) );
  XOR U28403 ( .A(n28468), .B(n28469), .Z(n28452) );
  AND U28404 ( .A(n28470), .B(n28471), .Z(n28469) );
  XOR U28405 ( .A(n28468), .B(n28472), .Z(n28470) );
  XNOR U28406 ( .A(n28451), .B(n28443), .Z(n28467) );
  XOR U28407 ( .A(n28473), .B(n28474), .Z(n28443) );
  AND U28408 ( .A(n28475), .B(n28476), .Z(n28474) );
  XNOR U28409 ( .A(n28477), .B(n28473), .Z(n28475) );
  XNOR U28410 ( .A(n28478), .B(n28448), .Z(n28451) );
  XOR U28411 ( .A(n28479), .B(n28480), .Z(n28448) );
  AND U28412 ( .A(n28481), .B(n28482), .Z(n28480) );
  XOR U28413 ( .A(n28479), .B(n28483), .Z(n28481) );
  XNOR U28414 ( .A(n28484), .B(n28485), .Z(n28478) );
  AND U28415 ( .A(n28486), .B(n28487), .Z(n28485) );
  XNOR U28416 ( .A(n28484), .B(n28488), .Z(n28486) );
  XNOR U28417 ( .A(n28447), .B(n28454), .Z(n28466) );
  AND U28418 ( .A(n28407), .B(n28489), .Z(n28454) );
  XOR U28419 ( .A(n28459), .B(n28458), .Z(n28447) );
  XNOR U28420 ( .A(n28490), .B(n28455), .Z(n28458) );
  XOR U28421 ( .A(n28491), .B(n28492), .Z(n28455) );
  AND U28422 ( .A(n28493), .B(n28494), .Z(n28492) );
  XOR U28423 ( .A(n28491), .B(n28495), .Z(n28493) );
  XNOR U28424 ( .A(n28496), .B(n28497), .Z(n28490) );
  AND U28425 ( .A(n28498), .B(n28499), .Z(n28497) );
  XOR U28426 ( .A(n28496), .B(n28500), .Z(n28498) );
  XOR U28427 ( .A(n28501), .B(n28502), .Z(n28459) );
  AND U28428 ( .A(n28503), .B(n28504), .Z(n28502) );
  XOR U28429 ( .A(n28501), .B(n28505), .Z(n28503) );
  XNOR U28430 ( .A(n28392), .B(n28462), .Z(n28464) );
  XNOR U28431 ( .A(n28506), .B(n28507), .Z(n28392) );
  AND U28432 ( .A(n540), .B(n28399), .Z(n28507) );
  XOR U28433 ( .A(n28506), .B(n28397), .Z(n28399) );
  XOR U28434 ( .A(n28508), .B(n28509), .Z(n28462) );
  AND U28435 ( .A(n28510), .B(n28511), .Z(n28509) );
  XNOR U28436 ( .A(n28508), .B(n28407), .Z(n28511) );
  XOR U28437 ( .A(n28512), .B(n28476), .Z(n28407) );
  XNOR U28438 ( .A(n28513), .B(n28483), .Z(n28476) );
  XOR U28439 ( .A(n28472), .B(n28471), .Z(n28483) );
  XNOR U28440 ( .A(n28514), .B(n28468), .Z(n28471) );
  XOR U28441 ( .A(n28515), .B(n28516), .Z(n28468) );
  AND U28442 ( .A(n28517), .B(n28518), .Z(n28516) );
  XNOR U28443 ( .A(n28519), .B(n28520), .Z(n28517) );
  IV U28444 ( .A(n28515), .Z(n28519) );
  XNOR U28445 ( .A(n28521), .B(n28522), .Z(n28514) );
  NOR U28446 ( .A(n28523), .B(n28524), .Z(n28522) );
  XNOR U28447 ( .A(n28521), .B(n28525), .Z(n28523) );
  XOR U28448 ( .A(n28526), .B(n28527), .Z(n28472) );
  NOR U28449 ( .A(n28528), .B(n28529), .Z(n28527) );
  XNOR U28450 ( .A(n28526), .B(n28530), .Z(n28528) );
  XNOR U28451 ( .A(n28482), .B(n28473), .Z(n28513) );
  XOR U28452 ( .A(n28531), .B(n28532), .Z(n28473) );
  AND U28453 ( .A(n28533), .B(n28534), .Z(n28532) );
  XOR U28454 ( .A(n28531), .B(n28535), .Z(n28533) );
  XOR U28455 ( .A(n28536), .B(n28488), .Z(n28482) );
  XOR U28456 ( .A(n28537), .B(n28538), .Z(n28488) );
  NOR U28457 ( .A(n28539), .B(n28540), .Z(n28538) );
  XOR U28458 ( .A(n28537), .B(n28541), .Z(n28539) );
  XNOR U28459 ( .A(n28487), .B(n28479), .Z(n28536) );
  XOR U28460 ( .A(n28542), .B(n28543), .Z(n28479) );
  AND U28461 ( .A(n28544), .B(n28545), .Z(n28543) );
  XOR U28462 ( .A(n28542), .B(n28546), .Z(n28544) );
  XNOR U28463 ( .A(n28547), .B(n28484), .Z(n28487) );
  XOR U28464 ( .A(n28548), .B(n28549), .Z(n28484) );
  AND U28465 ( .A(n28550), .B(n28551), .Z(n28549) );
  XNOR U28466 ( .A(n28552), .B(n28553), .Z(n28550) );
  IV U28467 ( .A(n28548), .Z(n28552) );
  XNOR U28468 ( .A(n28554), .B(n28555), .Z(n28547) );
  NOR U28469 ( .A(n28556), .B(n28557), .Z(n28555) );
  XNOR U28470 ( .A(n28554), .B(n28558), .Z(n28556) );
  XOR U28471 ( .A(n28477), .B(n28489), .Z(n28512) );
  NOR U28472 ( .A(n28415), .B(n28559), .Z(n28489) );
  XNOR U28473 ( .A(n28495), .B(n28494), .Z(n28477) );
  XNOR U28474 ( .A(n28560), .B(n28500), .Z(n28494) );
  XNOR U28475 ( .A(n28561), .B(n28562), .Z(n28500) );
  NOR U28476 ( .A(n28563), .B(n28564), .Z(n28562) );
  XOR U28477 ( .A(n28561), .B(n28565), .Z(n28563) );
  XNOR U28478 ( .A(n28499), .B(n28491), .Z(n28560) );
  XOR U28479 ( .A(n28566), .B(n28567), .Z(n28491) );
  AND U28480 ( .A(n28568), .B(n28569), .Z(n28567) );
  XOR U28481 ( .A(n28566), .B(n28570), .Z(n28568) );
  XNOR U28482 ( .A(n28571), .B(n28496), .Z(n28499) );
  XOR U28483 ( .A(n28572), .B(n28573), .Z(n28496) );
  AND U28484 ( .A(n28574), .B(n28575), .Z(n28573) );
  XNOR U28485 ( .A(n28576), .B(n28577), .Z(n28574) );
  IV U28486 ( .A(n28572), .Z(n28576) );
  XNOR U28487 ( .A(n28578), .B(n28579), .Z(n28571) );
  NOR U28488 ( .A(n28580), .B(n28581), .Z(n28579) );
  XNOR U28489 ( .A(n28578), .B(n28582), .Z(n28580) );
  XOR U28490 ( .A(n28505), .B(n28504), .Z(n28495) );
  XNOR U28491 ( .A(n28583), .B(n28501), .Z(n28504) );
  XOR U28492 ( .A(n28584), .B(n28585), .Z(n28501) );
  AND U28493 ( .A(n28586), .B(n28587), .Z(n28585) );
  XNOR U28494 ( .A(n28588), .B(n28589), .Z(n28586) );
  IV U28495 ( .A(n28584), .Z(n28588) );
  XNOR U28496 ( .A(n28590), .B(n28591), .Z(n28583) );
  NOR U28497 ( .A(n28592), .B(n28593), .Z(n28591) );
  XNOR U28498 ( .A(n28590), .B(n28594), .Z(n28592) );
  XOR U28499 ( .A(n28595), .B(n28596), .Z(n28505) );
  NOR U28500 ( .A(n28597), .B(n28598), .Z(n28596) );
  XNOR U28501 ( .A(n28595), .B(n28599), .Z(n28597) );
  XNOR U28502 ( .A(n28404), .B(n28508), .Z(n28510) );
  XNOR U28503 ( .A(n28600), .B(n28601), .Z(n28404) );
  AND U28504 ( .A(n540), .B(n28411), .Z(n28601) );
  XOR U28505 ( .A(n28600), .B(n28409), .Z(n28411) );
  AND U28506 ( .A(n28412), .B(n28415), .Z(n28508) );
  XOR U28507 ( .A(n28602), .B(n28559), .Z(n28415) );
  XNOR U28508 ( .A(p_input[1376]), .B(p_input[2048]), .Z(n28559) );
  XNOR U28509 ( .A(n28535), .B(n28534), .Z(n28602) );
  XNOR U28510 ( .A(n28603), .B(n28546), .Z(n28534) );
  XOR U28511 ( .A(n28520), .B(n28518), .Z(n28546) );
  XNOR U28512 ( .A(n28604), .B(n28525), .Z(n28518) );
  XOR U28513 ( .A(p_input[1400]), .B(p_input[2072]), .Z(n28525) );
  XOR U28514 ( .A(n28515), .B(n28524), .Z(n28604) );
  XOR U28515 ( .A(n28605), .B(n28521), .Z(n28524) );
  XOR U28516 ( .A(p_input[1398]), .B(p_input[2070]), .Z(n28521) );
  XOR U28517 ( .A(p_input[1399]), .B(n17295), .Z(n28605) );
  XOR U28518 ( .A(p_input[1394]), .B(p_input[2066]), .Z(n28515) );
  XNOR U28519 ( .A(n28530), .B(n28529), .Z(n28520) );
  XOR U28520 ( .A(n28606), .B(n28526), .Z(n28529) );
  XOR U28521 ( .A(p_input[1395]), .B(p_input[2067]), .Z(n28526) );
  XOR U28522 ( .A(p_input[1396]), .B(n17297), .Z(n28606) );
  XOR U28523 ( .A(p_input[1397]), .B(p_input[2069]), .Z(n28530) );
  XOR U28524 ( .A(n28545), .B(n28607), .Z(n28603) );
  IV U28525 ( .A(n28531), .Z(n28607) );
  XOR U28526 ( .A(p_input[1377]), .B(p_input[2049]), .Z(n28531) );
  XNOR U28527 ( .A(n28608), .B(n28553), .Z(n28545) );
  XNOR U28528 ( .A(n28541), .B(n28540), .Z(n28553) );
  XNOR U28529 ( .A(n28609), .B(n28537), .Z(n28540) );
  XNOR U28530 ( .A(p_input[1402]), .B(p_input[2074]), .Z(n28537) );
  XOR U28531 ( .A(p_input[1403]), .B(n17300), .Z(n28609) );
  XOR U28532 ( .A(p_input[1404]), .B(p_input[2076]), .Z(n28541) );
  XOR U28533 ( .A(n28551), .B(n28610), .Z(n28608) );
  IV U28534 ( .A(n28542), .Z(n28610) );
  XOR U28535 ( .A(p_input[1393]), .B(p_input[2065]), .Z(n28542) );
  XNOR U28536 ( .A(n28611), .B(n28558), .Z(n28551) );
  XNOR U28537 ( .A(p_input[1407]), .B(n17303), .Z(n28558) );
  XOR U28538 ( .A(n28548), .B(n28557), .Z(n28611) );
  XOR U28539 ( .A(n28612), .B(n28554), .Z(n28557) );
  XOR U28540 ( .A(p_input[1405]), .B(p_input[2077]), .Z(n28554) );
  XOR U28541 ( .A(p_input[1406]), .B(n17305), .Z(n28612) );
  XOR U28542 ( .A(p_input[1401]), .B(p_input[2073]), .Z(n28548) );
  XOR U28543 ( .A(n28570), .B(n28569), .Z(n28535) );
  XNOR U28544 ( .A(n28613), .B(n28577), .Z(n28569) );
  XNOR U28545 ( .A(n28565), .B(n28564), .Z(n28577) );
  XNOR U28546 ( .A(n28614), .B(n28561), .Z(n28564) );
  XNOR U28547 ( .A(p_input[1387]), .B(p_input[2059]), .Z(n28561) );
  XOR U28548 ( .A(p_input[1388]), .B(n16451), .Z(n28614) );
  XOR U28549 ( .A(p_input[1389]), .B(p_input[2061]), .Z(n28565) );
  XOR U28550 ( .A(n28575), .B(n28615), .Z(n28613) );
  IV U28551 ( .A(n28566), .Z(n28615) );
  XOR U28552 ( .A(p_input[1378]), .B(p_input[2050]), .Z(n28566) );
  XNOR U28553 ( .A(n28616), .B(n28582), .Z(n28575) );
  XNOR U28554 ( .A(p_input[1392]), .B(n16454), .Z(n28582) );
  XOR U28555 ( .A(n28572), .B(n28581), .Z(n28616) );
  XOR U28556 ( .A(n28617), .B(n28578), .Z(n28581) );
  XOR U28557 ( .A(p_input[1390]), .B(p_input[2062]), .Z(n28578) );
  XOR U28558 ( .A(p_input[1391]), .B(n16456), .Z(n28617) );
  XOR U28559 ( .A(p_input[1386]), .B(p_input[2058]), .Z(n28572) );
  XOR U28560 ( .A(n28589), .B(n28587), .Z(n28570) );
  XNOR U28561 ( .A(n28618), .B(n28594), .Z(n28587) );
  XOR U28562 ( .A(p_input[1385]), .B(p_input[2057]), .Z(n28594) );
  XOR U28563 ( .A(n28584), .B(n28593), .Z(n28618) );
  XOR U28564 ( .A(n28619), .B(n28590), .Z(n28593) );
  XOR U28565 ( .A(p_input[1383]), .B(p_input[2055]), .Z(n28590) );
  XOR U28566 ( .A(p_input[1384]), .B(n17312), .Z(n28619) );
  XOR U28567 ( .A(p_input[1379]), .B(p_input[2051]), .Z(n28584) );
  XNOR U28568 ( .A(n28599), .B(n28598), .Z(n28589) );
  XOR U28569 ( .A(n28620), .B(n28595), .Z(n28598) );
  XOR U28570 ( .A(p_input[1380]), .B(p_input[2052]), .Z(n28595) );
  XOR U28571 ( .A(p_input[1381]), .B(n17314), .Z(n28620) );
  XOR U28572 ( .A(p_input[1382]), .B(p_input[2054]), .Z(n28599) );
  XNOR U28573 ( .A(n28621), .B(n28622), .Z(n28412) );
  AND U28574 ( .A(n540), .B(n28623), .Z(n28622) );
  XNOR U28575 ( .A(n28624), .B(n28625), .Z(n540) );
  AND U28576 ( .A(n28626), .B(n28627), .Z(n28625) );
  XOR U28577 ( .A(n28624), .B(n28422), .Z(n28627) );
  XNOR U28578 ( .A(n28624), .B(n28364), .Z(n28626) );
  XOR U28579 ( .A(n28628), .B(n28629), .Z(n28624) );
  AND U28580 ( .A(n28630), .B(n28631), .Z(n28629) );
  XNOR U28581 ( .A(n28435), .B(n28628), .Z(n28631) );
  XOR U28582 ( .A(n28628), .B(n28376), .Z(n28630) );
  XOR U28583 ( .A(n28632), .B(n28633), .Z(n28628) );
  AND U28584 ( .A(n28634), .B(n28635), .Z(n28633) );
  XNOR U28585 ( .A(n28460), .B(n28632), .Z(n28635) );
  XOR U28586 ( .A(n28632), .B(n28387), .Z(n28634) );
  XOR U28587 ( .A(n28636), .B(n28637), .Z(n28632) );
  AND U28588 ( .A(n28638), .B(n28639), .Z(n28637) );
  XOR U28589 ( .A(n28636), .B(n28397), .Z(n28638) );
  XOR U28590 ( .A(n28640), .B(n28641), .Z(n28353) );
  AND U28591 ( .A(n544), .B(n28623), .Z(n28641) );
  XNOR U28592 ( .A(n28621), .B(n28640), .Z(n28623) );
  XNOR U28593 ( .A(n28642), .B(n28643), .Z(n544) );
  AND U28594 ( .A(n28644), .B(n28645), .Z(n28643) );
  XNOR U28595 ( .A(n28646), .B(n28642), .Z(n28645) );
  IV U28596 ( .A(n28422), .Z(n28646) );
  XNOR U28597 ( .A(n28647), .B(n28648), .Z(n28422) );
  AND U28598 ( .A(n547), .B(n28649), .Z(n28648) );
  XNOR U28599 ( .A(n28647), .B(n28650), .Z(n28649) );
  XNOR U28600 ( .A(n28364), .B(n28642), .Z(n28644) );
  XOR U28601 ( .A(n28651), .B(n28652), .Z(n28364) );
  AND U28602 ( .A(n555), .B(n28653), .Z(n28652) );
  XOR U28603 ( .A(n28654), .B(n28655), .Z(n28642) );
  AND U28604 ( .A(n28656), .B(n28657), .Z(n28655) );
  XNOR U28605 ( .A(n28654), .B(n28435), .Z(n28657) );
  XNOR U28606 ( .A(n28658), .B(n28659), .Z(n28435) );
  AND U28607 ( .A(n547), .B(n28660), .Z(n28659) );
  XOR U28608 ( .A(n28661), .B(n28658), .Z(n28660) );
  XNOR U28609 ( .A(n28662), .B(n28654), .Z(n28656) );
  IV U28610 ( .A(n28376), .Z(n28662) );
  XOR U28611 ( .A(n28663), .B(n28664), .Z(n28376) );
  AND U28612 ( .A(n555), .B(n28665), .Z(n28664) );
  XOR U28613 ( .A(n28666), .B(n28667), .Z(n28654) );
  AND U28614 ( .A(n28668), .B(n28669), .Z(n28667) );
  XNOR U28615 ( .A(n28666), .B(n28460), .Z(n28669) );
  XNOR U28616 ( .A(n28670), .B(n28671), .Z(n28460) );
  AND U28617 ( .A(n547), .B(n28672), .Z(n28671) );
  XNOR U28618 ( .A(n28673), .B(n28670), .Z(n28672) );
  XOR U28619 ( .A(n28387), .B(n28666), .Z(n28668) );
  XOR U28620 ( .A(n28674), .B(n28675), .Z(n28387) );
  AND U28621 ( .A(n555), .B(n28676), .Z(n28675) );
  XOR U28622 ( .A(n28636), .B(n28677), .Z(n28666) );
  AND U28623 ( .A(n28678), .B(n28639), .Z(n28677) );
  XNOR U28624 ( .A(n28506), .B(n28636), .Z(n28639) );
  XNOR U28625 ( .A(n28679), .B(n28680), .Z(n28506) );
  AND U28626 ( .A(n547), .B(n28681), .Z(n28680) );
  XOR U28627 ( .A(n28682), .B(n28679), .Z(n28681) );
  XNOR U28628 ( .A(n28683), .B(n28636), .Z(n28678) );
  IV U28629 ( .A(n28397), .Z(n28683) );
  XOR U28630 ( .A(n28684), .B(n28685), .Z(n28397) );
  AND U28631 ( .A(n555), .B(n28686), .Z(n28685) );
  XOR U28632 ( .A(n28687), .B(n28688), .Z(n28636) );
  AND U28633 ( .A(n28689), .B(n28690), .Z(n28688) );
  XNOR U28634 ( .A(n28687), .B(n28600), .Z(n28690) );
  XNOR U28635 ( .A(n28691), .B(n28692), .Z(n28600) );
  AND U28636 ( .A(n547), .B(n28693), .Z(n28692) );
  XNOR U28637 ( .A(n28694), .B(n28691), .Z(n28693) );
  XNOR U28638 ( .A(n28695), .B(n28687), .Z(n28689) );
  IV U28639 ( .A(n28409), .Z(n28695) );
  XOR U28640 ( .A(n28696), .B(n28697), .Z(n28409) );
  AND U28641 ( .A(n555), .B(n28698), .Z(n28697) );
  AND U28642 ( .A(n28640), .B(n28621), .Z(n28687) );
  XNOR U28643 ( .A(n28699), .B(n28700), .Z(n28621) );
  AND U28644 ( .A(n547), .B(n28701), .Z(n28700) );
  XNOR U28645 ( .A(n28702), .B(n28699), .Z(n28701) );
  XNOR U28646 ( .A(n28703), .B(n28704), .Z(n547) );
  AND U28647 ( .A(n28705), .B(n28706), .Z(n28704) );
  XOR U28648 ( .A(n28650), .B(n28703), .Z(n28706) );
  AND U28649 ( .A(n28707), .B(n28708), .Z(n28650) );
  XOR U28650 ( .A(n28703), .B(n28647), .Z(n28705) );
  XNOR U28651 ( .A(n28709), .B(n28710), .Z(n28647) );
  AND U28652 ( .A(n551), .B(n28653), .Z(n28710) );
  XOR U28653 ( .A(n28651), .B(n28709), .Z(n28653) );
  XOR U28654 ( .A(n28711), .B(n28712), .Z(n28703) );
  AND U28655 ( .A(n28713), .B(n28714), .Z(n28712) );
  XNOR U28656 ( .A(n28711), .B(n28707), .Z(n28714) );
  IV U28657 ( .A(n28661), .Z(n28707) );
  XOR U28658 ( .A(n28715), .B(n28716), .Z(n28661) );
  XOR U28659 ( .A(n28717), .B(n28708), .Z(n28716) );
  AND U28660 ( .A(n28673), .B(n28718), .Z(n28708) );
  AND U28661 ( .A(n28719), .B(n28720), .Z(n28717) );
  XOR U28662 ( .A(n28721), .B(n28715), .Z(n28719) );
  XNOR U28663 ( .A(n28658), .B(n28711), .Z(n28713) );
  XNOR U28664 ( .A(n28722), .B(n28723), .Z(n28658) );
  AND U28665 ( .A(n551), .B(n28665), .Z(n28723) );
  XOR U28666 ( .A(n28722), .B(n28663), .Z(n28665) );
  XOR U28667 ( .A(n28724), .B(n28725), .Z(n28711) );
  AND U28668 ( .A(n28726), .B(n28727), .Z(n28725) );
  XNOR U28669 ( .A(n28724), .B(n28673), .Z(n28727) );
  XOR U28670 ( .A(n28728), .B(n28720), .Z(n28673) );
  XNOR U28671 ( .A(n28729), .B(n28715), .Z(n28720) );
  XOR U28672 ( .A(n28730), .B(n28731), .Z(n28715) );
  AND U28673 ( .A(n28732), .B(n28733), .Z(n28731) );
  XOR U28674 ( .A(n28734), .B(n28730), .Z(n28732) );
  XNOR U28675 ( .A(n28735), .B(n28736), .Z(n28729) );
  AND U28676 ( .A(n28737), .B(n28738), .Z(n28736) );
  XOR U28677 ( .A(n28735), .B(n28739), .Z(n28737) );
  XNOR U28678 ( .A(n28721), .B(n28718), .Z(n28728) );
  AND U28679 ( .A(n28740), .B(n28741), .Z(n28718) );
  XOR U28680 ( .A(n28742), .B(n28743), .Z(n28721) );
  AND U28681 ( .A(n28744), .B(n28745), .Z(n28743) );
  XOR U28682 ( .A(n28742), .B(n28746), .Z(n28744) );
  XNOR U28683 ( .A(n28670), .B(n28724), .Z(n28726) );
  XNOR U28684 ( .A(n28747), .B(n28748), .Z(n28670) );
  AND U28685 ( .A(n551), .B(n28676), .Z(n28748) );
  XOR U28686 ( .A(n28747), .B(n28674), .Z(n28676) );
  XOR U28687 ( .A(n28749), .B(n28750), .Z(n28724) );
  AND U28688 ( .A(n28751), .B(n28752), .Z(n28750) );
  XNOR U28689 ( .A(n28749), .B(n28740), .Z(n28752) );
  IV U28690 ( .A(n28682), .Z(n28740) );
  XNOR U28691 ( .A(n28753), .B(n28733), .Z(n28682) );
  XNOR U28692 ( .A(n28754), .B(n28739), .Z(n28733) );
  XOR U28693 ( .A(n28755), .B(n28756), .Z(n28739) );
  AND U28694 ( .A(n28757), .B(n28758), .Z(n28756) );
  XOR U28695 ( .A(n28755), .B(n28759), .Z(n28757) );
  XNOR U28696 ( .A(n28738), .B(n28730), .Z(n28754) );
  XOR U28697 ( .A(n28760), .B(n28761), .Z(n28730) );
  AND U28698 ( .A(n28762), .B(n28763), .Z(n28761) );
  XNOR U28699 ( .A(n28764), .B(n28760), .Z(n28762) );
  XNOR U28700 ( .A(n28765), .B(n28735), .Z(n28738) );
  XOR U28701 ( .A(n28766), .B(n28767), .Z(n28735) );
  AND U28702 ( .A(n28768), .B(n28769), .Z(n28767) );
  XOR U28703 ( .A(n28766), .B(n28770), .Z(n28768) );
  XNOR U28704 ( .A(n28771), .B(n28772), .Z(n28765) );
  AND U28705 ( .A(n28773), .B(n28774), .Z(n28772) );
  XNOR U28706 ( .A(n28771), .B(n28775), .Z(n28773) );
  XNOR U28707 ( .A(n28734), .B(n28741), .Z(n28753) );
  AND U28708 ( .A(n28694), .B(n28776), .Z(n28741) );
  XOR U28709 ( .A(n28746), .B(n28745), .Z(n28734) );
  XNOR U28710 ( .A(n28777), .B(n28742), .Z(n28745) );
  XOR U28711 ( .A(n28778), .B(n28779), .Z(n28742) );
  AND U28712 ( .A(n28780), .B(n28781), .Z(n28779) );
  XOR U28713 ( .A(n28778), .B(n28782), .Z(n28780) );
  XNOR U28714 ( .A(n28783), .B(n28784), .Z(n28777) );
  AND U28715 ( .A(n28785), .B(n28786), .Z(n28784) );
  XOR U28716 ( .A(n28783), .B(n28787), .Z(n28785) );
  XOR U28717 ( .A(n28788), .B(n28789), .Z(n28746) );
  AND U28718 ( .A(n28790), .B(n28791), .Z(n28789) );
  XOR U28719 ( .A(n28788), .B(n28792), .Z(n28790) );
  XNOR U28720 ( .A(n28679), .B(n28749), .Z(n28751) );
  XNOR U28721 ( .A(n28793), .B(n28794), .Z(n28679) );
  AND U28722 ( .A(n551), .B(n28686), .Z(n28794) );
  XOR U28723 ( .A(n28793), .B(n28684), .Z(n28686) );
  XOR U28724 ( .A(n28795), .B(n28796), .Z(n28749) );
  AND U28725 ( .A(n28797), .B(n28798), .Z(n28796) );
  XNOR U28726 ( .A(n28795), .B(n28694), .Z(n28798) );
  XOR U28727 ( .A(n28799), .B(n28763), .Z(n28694) );
  XNOR U28728 ( .A(n28800), .B(n28770), .Z(n28763) );
  XOR U28729 ( .A(n28759), .B(n28758), .Z(n28770) );
  XNOR U28730 ( .A(n28801), .B(n28755), .Z(n28758) );
  XOR U28731 ( .A(n28802), .B(n28803), .Z(n28755) );
  AND U28732 ( .A(n28804), .B(n28805), .Z(n28803) );
  XNOR U28733 ( .A(n28806), .B(n28807), .Z(n28804) );
  IV U28734 ( .A(n28802), .Z(n28806) );
  XNOR U28735 ( .A(n28808), .B(n28809), .Z(n28801) );
  NOR U28736 ( .A(n28810), .B(n28811), .Z(n28809) );
  XNOR U28737 ( .A(n28808), .B(n28812), .Z(n28810) );
  XOR U28738 ( .A(n28813), .B(n28814), .Z(n28759) );
  NOR U28739 ( .A(n28815), .B(n28816), .Z(n28814) );
  XNOR U28740 ( .A(n28813), .B(n28817), .Z(n28815) );
  XNOR U28741 ( .A(n28769), .B(n28760), .Z(n28800) );
  XOR U28742 ( .A(n28818), .B(n28819), .Z(n28760) );
  AND U28743 ( .A(n28820), .B(n28821), .Z(n28819) );
  XOR U28744 ( .A(n28818), .B(n28822), .Z(n28820) );
  XOR U28745 ( .A(n28823), .B(n28775), .Z(n28769) );
  XOR U28746 ( .A(n28824), .B(n28825), .Z(n28775) );
  NOR U28747 ( .A(n28826), .B(n28827), .Z(n28825) );
  XOR U28748 ( .A(n28824), .B(n28828), .Z(n28826) );
  XNOR U28749 ( .A(n28774), .B(n28766), .Z(n28823) );
  XOR U28750 ( .A(n28829), .B(n28830), .Z(n28766) );
  AND U28751 ( .A(n28831), .B(n28832), .Z(n28830) );
  XOR U28752 ( .A(n28829), .B(n28833), .Z(n28831) );
  XNOR U28753 ( .A(n28834), .B(n28771), .Z(n28774) );
  XOR U28754 ( .A(n28835), .B(n28836), .Z(n28771) );
  AND U28755 ( .A(n28837), .B(n28838), .Z(n28836) );
  XNOR U28756 ( .A(n28839), .B(n28840), .Z(n28837) );
  IV U28757 ( .A(n28835), .Z(n28839) );
  XNOR U28758 ( .A(n28841), .B(n28842), .Z(n28834) );
  NOR U28759 ( .A(n28843), .B(n28844), .Z(n28842) );
  XNOR U28760 ( .A(n28841), .B(n28845), .Z(n28843) );
  XOR U28761 ( .A(n28764), .B(n28776), .Z(n28799) );
  NOR U28762 ( .A(n28702), .B(n28846), .Z(n28776) );
  XNOR U28763 ( .A(n28782), .B(n28781), .Z(n28764) );
  XNOR U28764 ( .A(n28847), .B(n28787), .Z(n28781) );
  XNOR U28765 ( .A(n28848), .B(n28849), .Z(n28787) );
  NOR U28766 ( .A(n28850), .B(n28851), .Z(n28849) );
  XOR U28767 ( .A(n28848), .B(n28852), .Z(n28850) );
  XNOR U28768 ( .A(n28786), .B(n28778), .Z(n28847) );
  XOR U28769 ( .A(n28853), .B(n28854), .Z(n28778) );
  AND U28770 ( .A(n28855), .B(n28856), .Z(n28854) );
  XOR U28771 ( .A(n28853), .B(n28857), .Z(n28855) );
  XNOR U28772 ( .A(n28858), .B(n28783), .Z(n28786) );
  XOR U28773 ( .A(n28859), .B(n28860), .Z(n28783) );
  AND U28774 ( .A(n28861), .B(n28862), .Z(n28860) );
  XNOR U28775 ( .A(n28863), .B(n28864), .Z(n28861) );
  IV U28776 ( .A(n28859), .Z(n28863) );
  XNOR U28777 ( .A(n28865), .B(n28866), .Z(n28858) );
  NOR U28778 ( .A(n28867), .B(n28868), .Z(n28866) );
  XNOR U28779 ( .A(n28865), .B(n28869), .Z(n28867) );
  XOR U28780 ( .A(n28792), .B(n28791), .Z(n28782) );
  XNOR U28781 ( .A(n28870), .B(n28788), .Z(n28791) );
  XOR U28782 ( .A(n28871), .B(n28872), .Z(n28788) );
  AND U28783 ( .A(n28873), .B(n28874), .Z(n28872) );
  XNOR U28784 ( .A(n28875), .B(n28876), .Z(n28873) );
  IV U28785 ( .A(n28871), .Z(n28875) );
  XNOR U28786 ( .A(n28877), .B(n28878), .Z(n28870) );
  NOR U28787 ( .A(n28879), .B(n28880), .Z(n28878) );
  XNOR U28788 ( .A(n28877), .B(n28881), .Z(n28879) );
  XOR U28789 ( .A(n28882), .B(n28883), .Z(n28792) );
  NOR U28790 ( .A(n28884), .B(n28885), .Z(n28883) );
  XNOR U28791 ( .A(n28882), .B(n28886), .Z(n28884) );
  XNOR U28792 ( .A(n28691), .B(n28795), .Z(n28797) );
  XNOR U28793 ( .A(n28887), .B(n28888), .Z(n28691) );
  AND U28794 ( .A(n551), .B(n28698), .Z(n28888) );
  XOR U28795 ( .A(n28887), .B(n28696), .Z(n28698) );
  AND U28796 ( .A(n28699), .B(n28702), .Z(n28795) );
  XOR U28797 ( .A(n28889), .B(n28846), .Z(n28702) );
  XNOR U28798 ( .A(p_input[1408]), .B(p_input[2048]), .Z(n28846) );
  XNOR U28799 ( .A(n28822), .B(n28821), .Z(n28889) );
  XNOR U28800 ( .A(n28890), .B(n28833), .Z(n28821) );
  XOR U28801 ( .A(n28807), .B(n28805), .Z(n28833) );
  XNOR U28802 ( .A(n28891), .B(n28812), .Z(n28805) );
  XOR U28803 ( .A(p_input[1432]), .B(p_input[2072]), .Z(n28812) );
  XOR U28804 ( .A(n28802), .B(n28811), .Z(n28891) );
  XOR U28805 ( .A(n28892), .B(n28808), .Z(n28811) );
  XOR U28806 ( .A(p_input[1430]), .B(p_input[2070]), .Z(n28808) );
  XOR U28807 ( .A(p_input[1431]), .B(n17295), .Z(n28892) );
  XOR U28808 ( .A(p_input[1426]), .B(p_input[2066]), .Z(n28802) );
  XNOR U28809 ( .A(n28817), .B(n28816), .Z(n28807) );
  XOR U28810 ( .A(n28893), .B(n28813), .Z(n28816) );
  XOR U28811 ( .A(p_input[1427]), .B(p_input[2067]), .Z(n28813) );
  XOR U28812 ( .A(p_input[1428]), .B(n17297), .Z(n28893) );
  XOR U28813 ( .A(p_input[1429]), .B(p_input[2069]), .Z(n28817) );
  XOR U28814 ( .A(n28832), .B(n28894), .Z(n28890) );
  IV U28815 ( .A(n28818), .Z(n28894) );
  XOR U28816 ( .A(p_input[1409]), .B(p_input[2049]), .Z(n28818) );
  XNOR U28817 ( .A(n28895), .B(n28840), .Z(n28832) );
  XNOR U28818 ( .A(n28828), .B(n28827), .Z(n28840) );
  XNOR U28819 ( .A(n28896), .B(n28824), .Z(n28827) );
  XNOR U28820 ( .A(p_input[1434]), .B(p_input[2074]), .Z(n28824) );
  XOR U28821 ( .A(p_input[1435]), .B(n17300), .Z(n28896) );
  XOR U28822 ( .A(p_input[1436]), .B(p_input[2076]), .Z(n28828) );
  XOR U28823 ( .A(n28838), .B(n28897), .Z(n28895) );
  IV U28824 ( .A(n28829), .Z(n28897) );
  XOR U28825 ( .A(p_input[1425]), .B(p_input[2065]), .Z(n28829) );
  XNOR U28826 ( .A(n28898), .B(n28845), .Z(n28838) );
  XNOR U28827 ( .A(p_input[1439]), .B(n17303), .Z(n28845) );
  XOR U28828 ( .A(n28835), .B(n28844), .Z(n28898) );
  XOR U28829 ( .A(n28899), .B(n28841), .Z(n28844) );
  XOR U28830 ( .A(p_input[1437]), .B(p_input[2077]), .Z(n28841) );
  XOR U28831 ( .A(p_input[1438]), .B(n17305), .Z(n28899) );
  XOR U28832 ( .A(p_input[1433]), .B(p_input[2073]), .Z(n28835) );
  XOR U28833 ( .A(n28857), .B(n28856), .Z(n28822) );
  XNOR U28834 ( .A(n28900), .B(n28864), .Z(n28856) );
  XNOR U28835 ( .A(n28852), .B(n28851), .Z(n28864) );
  XNOR U28836 ( .A(n28901), .B(n28848), .Z(n28851) );
  XNOR U28837 ( .A(p_input[1419]), .B(p_input[2059]), .Z(n28848) );
  XOR U28838 ( .A(p_input[1420]), .B(n16451), .Z(n28901) );
  XOR U28839 ( .A(p_input[1421]), .B(p_input[2061]), .Z(n28852) );
  XOR U28840 ( .A(n28862), .B(n28902), .Z(n28900) );
  IV U28841 ( .A(n28853), .Z(n28902) );
  XOR U28842 ( .A(p_input[1410]), .B(p_input[2050]), .Z(n28853) );
  XNOR U28843 ( .A(n28903), .B(n28869), .Z(n28862) );
  XNOR U28844 ( .A(p_input[1424]), .B(n16454), .Z(n28869) );
  XOR U28845 ( .A(n28859), .B(n28868), .Z(n28903) );
  XOR U28846 ( .A(n28904), .B(n28865), .Z(n28868) );
  XOR U28847 ( .A(p_input[1422]), .B(p_input[2062]), .Z(n28865) );
  XOR U28848 ( .A(p_input[1423]), .B(n16456), .Z(n28904) );
  XOR U28849 ( .A(p_input[1418]), .B(p_input[2058]), .Z(n28859) );
  XOR U28850 ( .A(n28876), .B(n28874), .Z(n28857) );
  XNOR U28851 ( .A(n28905), .B(n28881), .Z(n28874) );
  XOR U28852 ( .A(p_input[1417]), .B(p_input[2057]), .Z(n28881) );
  XOR U28853 ( .A(n28871), .B(n28880), .Z(n28905) );
  XOR U28854 ( .A(n28906), .B(n28877), .Z(n28880) );
  XOR U28855 ( .A(p_input[1415]), .B(p_input[2055]), .Z(n28877) );
  XOR U28856 ( .A(p_input[1416]), .B(n17312), .Z(n28906) );
  XOR U28857 ( .A(p_input[1411]), .B(p_input[2051]), .Z(n28871) );
  XNOR U28858 ( .A(n28886), .B(n28885), .Z(n28876) );
  XOR U28859 ( .A(n28907), .B(n28882), .Z(n28885) );
  XOR U28860 ( .A(p_input[1412]), .B(p_input[2052]), .Z(n28882) );
  XOR U28861 ( .A(p_input[1413]), .B(n17314), .Z(n28907) );
  XOR U28862 ( .A(p_input[1414]), .B(p_input[2054]), .Z(n28886) );
  XNOR U28863 ( .A(n28908), .B(n28909), .Z(n28699) );
  AND U28864 ( .A(n551), .B(n28910), .Z(n28909) );
  XNOR U28865 ( .A(n28911), .B(n28912), .Z(n551) );
  AND U28866 ( .A(n28913), .B(n28914), .Z(n28912) );
  XOR U28867 ( .A(n28911), .B(n28709), .Z(n28914) );
  XNOR U28868 ( .A(n28911), .B(n28651), .Z(n28913) );
  XOR U28869 ( .A(n28915), .B(n28916), .Z(n28911) );
  AND U28870 ( .A(n28917), .B(n28918), .Z(n28916) );
  XNOR U28871 ( .A(n28722), .B(n28915), .Z(n28918) );
  XOR U28872 ( .A(n28915), .B(n28663), .Z(n28917) );
  XOR U28873 ( .A(n28919), .B(n28920), .Z(n28915) );
  AND U28874 ( .A(n28921), .B(n28922), .Z(n28920) );
  XNOR U28875 ( .A(n28747), .B(n28919), .Z(n28922) );
  XOR U28876 ( .A(n28919), .B(n28674), .Z(n28921) );
  XOR U28877 ( .A(n28923), .B(n28924), .Z(n28919) );
  AND U28878 ( .A(n28925), .B(n28926), .Z(n28924) );
  XOR U28879 ( .A(n28923), .B(n28684), .Z(n28925) );
  XOR U28880 ( .A(n28927), .B(n28928), .Z(n28640) );
  AND U28881 ( .A(n555), .B(n28910), .Z(n28928) );
  XNOR U28882 ( .A(n28908), .B(n28927), .Z(n28910) );
  XNOR U28883 ( .A(n28929), .B(n28930), .Z(n555) );
  AND U28884 ( .A(n28931), .B(n28932), .Z(n28930) );
  XNOR U28885 ( .A(n28933), .B(n28929), .Z(n28932) );
  IV U28886 ( .A(n28709), .Z(n28933) );
  XNOR U28887 ( .A(n28934), .B(n28935), .Z(n28709) );
  AND U28888 ( .A(n558), .B(n28936), .Z(n28935) );
  XNOR U28889 ( .A(n28934), .B(n28937), .Z(n28936) );
  XNOR U28890 ( .A(n28651), .B(n28929), .Z(n28931) );
  XOR U28891 ( .A(n28938), .B(n28939), .Z(n28651) );
  AND U28892 ( .A(n566), .B(n28940), .Z(n28939) );
  XOR U28893 ( .A(n28941), .B(n28942), .Z(n28929) );
  AND U28894 ( .A(n28943), .B(n28944), .Z(n28942) );
  XNOR U28895 ( .A(n28941), .B(n28722), .Z(n28944) );
  XNOR U28896 ( .A(n28945), .B(n28946), .Z(n28722) );
  AND U28897 ( .A(n558), .B(n28947), .Z(n28946) );
  XOR U28898 ( .A(n28948), .B(n28945), .Z(n28947) );
  XNOR U28899 ( .A(n28949), .B(n28941), .Z(n28943) );
  IV U28900 ( .A(n28663), .Z(n28949) );
  XOR U28901 ( .A(n28950), .B(n28951), .Z(n28663) );
  AND U28902 ( .A(n566), .B(n28952), .Z(n28951) );
  XOR U28903 ( .A(n28953), .B(n28954), .Z(n28941) );
  AND U28904 ( .A(n28955), .B(n28956), .Z(n28954) );
  XNOR U28905 ( .A(n28953), .B(n28747), .Z(n28956) );
  XNOR U28906 ( .A(n28957), .B(n28958), .Z(n28747) );
  AND U28907 ( .A(n558), .B(n28959), .Z(n28958) );
  XNOR U28908 ( .A(n28960), .B(n28957), .Z(n28959) );
  XOR U28909 ( .A(n28674), .B(n28953), .Z(n28955) );
  XOR U28910 ( .A(n28961), .B(n28962), .Z(n28674) );
  AND U28911 ( .A(n566), .B(n28963), .Z(n28962) );
  XOR U28912 ( .A(n28923), .B(n28964), .Z(n28953) );
  AND U28913 ( .A(n28965), .B(n28926), .Z(n28964) );
  XNOR U28914 ( .A(n28793), .B(n28923), .Z(n28926) );
  XNOR U28915 ( .A(n28966), .B(n28967), .Z(n28793) );
  AND U28916 ( .A(n558), .B(n28968), .Z(n28967) );
  XOR U28917 ( .A(n28969), .B(n28966), .Z(n28968) );
  XNOR U28918 ( .A(n28970), .B(n28923), .Z(n28965) );
  IV U28919 ( .A(n28684), .Z(n28970) );
  XOR U28920 ( .A(n28971), .B(n28972), .Z(n28684) );
  AND U28921 ( .A(n566), .B(n28973), .Z(n28972) );
  XOR U28922 ( .A(n28974), .B(n28975), .Z(n28923) );
  AND U28923 ( .A(n28976), .B(n28977), .Z(n28975) );
  XNOR U28924 ( .A(n28974), .B(n28887), .Z(n28977) );
  XNOR U28925 ( .A(n28978), .B(n28979), .Z(n28887) );
  AND U28926 ( .A(n558), .B(n28980), .Z(n28979) );
  XNOR U28927 ( .A(n28981), .B(n28978), .Z(n28980) );
  XNOR U28928 ( .A(n28982), .B(n28974), .Z(n28976) );
  IV U28929 ( .A(n28696), .Z(n28982) );
  XOR U28930 ( .A(n28983), .B(n28984), .Z(n28696) );
  AND U28931 ( .A(n566), .B(n28985), .Z(n28984) );
  AND U28932 ( .A(n28927), .B(n28908), .Z(n28974) );
  XNOR U28933 ( .A(n28986), .B(n28987), .Z(n28908) );
  AND U28934 ( .A(n558), .B(n28988), .Z(n28987) );
  XNOR U28935 ( .A(n28989), .B(n28986), .Z(n28988) );
  XNOR U28936 ( .A(n28990), .B(n28991), .Z(n558) );
  AND U28937 ( .A(n28992), .B(n28993), .Z(n28991) );
  XOR U28938 ( .A(n28937), .B(n28990), .Z(n28993) );
  AND U28939 ( .A(n28994), .B(n28995), .Z(n28937) );
  XOR U28940 ( .A(n28990), .B(n28934), .Z(n28992) );
  XNOR U28941 ( .A(n28996), .B(n28997), .Z(n28934) );
  AND U28942 ( .A(n562), .B(n28940), .Z(n28997) );
  XOR U28943 ( .A(n28938), .B(n28996), .Z(n28940) );
  XOR U28944 ( .A(n28998), .B(n28999), .Z(n28990) );
  AND U28945 ( .A(n29000), .B(n29001), .Z(n28999) );
  XNOR U28946 ( .A(n28998), .B(n28994), .Z(n29001) );
  IV U28947 ( .A(n28948), .Z(n28994) );
  XOR U28948 ( .A(n29002), .B(n29003), .Z(n28948) );
  XOR U28949 ( .A(n29004), .B(n28995), .Z(n29003) );
  AND U28950 ( .A(n28960), .B(n29005), .Z(n28995) );
  AND U28951 ( .A(n29006), .B(n29007), .Z(n29004) );
  XOR U28952 ( .A(n29008), .B(n29002), .Z(n29006) );
  XNOR U28953 ( .A(n28945), .B(n28998), .Z(n29000) );
  XNOR U28954 ( .A(n29009), .B(n29010), .Z(n28945) );
  AND U28955 ( .A(n562), .B(n28952), .Z(n29010) );
  XOR U28956 ( .A(n29009), .B(n28950), .Z(n28952) );
  XOR U28957 ( .A(n29011), .B(n29012), .Z(n28998) );
  AND U28958 ( .A(n29013), .B(n29014), .Z(n29012) );
  XNOR U28959 ( .A(n29011), .B(n28960), .Z(n29014) );
  XOR U28960 ( .A(n29015), .B(n29007), .Z(n28960) );
  XNOR U28961 ( .A(n29016), .B(n29002), .Z(n29007) );
  XOR U28962 ( .A(n29017), .B(n29018), .Z(n29002) );
  AND U28963 ( .A(n29019), .B(n29020), .Z(n29018) );
  XOR U28964 ( .A(n29021), .B(n29017), .Z(n29019) );
  XNOR U28965 ( .A(n29022), .B(n29023), .Z(n29016) );
  AND U28966 ( .A(n29024), .B(n29025), .Z(n29023) );
  XOR U28967 ( .A(n29022), .B(n29026), .Z(n29024) );
  XNOR U28968 ( .A(n29008), .B(n29005), .Z(n29015) );
  AND U28969 ( .A(n29027), .B(n29028), .Z(n29005) );
  XOR U28970 ( .A(n29029), .B(n29030), .Z(n29008) );
  AND U28971 ( .A(n29031), .B(n29032), .Z(n29030) );
  XOR U28972 ( .A(n29029), .B(n29033), .Z(n29031) );
  XNOR U28973 ( .A(n28957), .B(n29011), .Z(n29013) );
  XNOR U28974 ( .A(n29034), .B(n29035), .Z(n28957) );
  AND U28975 ( .A(n562), .B(n28963), .Z(n29035) );
  XOR U28976 ( .A(n29034), .B(n28961), .Z(n28963) );
  XOR U28977 ( .A(n29036), .B(n29037), .Z(n29011) );
  AND U28978 ( .A(n29038), .B(n29039), .Z(n29037) );
  XNOR U28979 ( .A(n29036), .B(n29027), .Z(n29039) );
  IV U28980 ( .A(n28969), .Z(n29027) );
  XNOR U28981 ( .A(n29040), .B(n29020), .Z(n28969) );
  XNOR U28982 ( .A(n29041), .B(n29026), .Z(n29020) );
  XOR U28983 ( .A(n29042), .B(n29043), .Z(n29026) );
  AND U28984 ( .A(n29044), .B(n29045), .Z(n29043) );
  XOR U28985 ( .A(n29042), .B(n29046), .Z(n29044) );
  XNOR U28986 ( .A(n29025), .B(n29017), .Z(n29041) );
  XOR U28987 ( .A(n29047), .B(n29048), .Z(n29017) );
  AND U28988 ( .A(n29049), .B(n29050), .Z(n29048) );
  XNOR U28989 ( .A(n29051), .B(n29047), .Z(n29049) );
  XNOR U28990 ( .A(n29052), .B(n29022), .Z(n29025) );
  XOR U28991 ( .A(n29053), .B(n29054), .Z(n29022) );
  AND U28992 ( .A(n29055), .B(n29056), .Z(n29054) );
  XOR U28993 ( .A(n29053), .B(n29057), .Z(n29055) );
  XNOR U28994 ( .A(n29058), .B(n29059), .Z(n29052) );
  AND U28995 ( .A(n29060), .B(n29061), .Z(n29059) );
  XNOR U28996 ( .A(n29058), .B(n29062), .Z(n29060) );
  XNOR U28997 ( .A(n29021), .B(n29028), .Z(n29040) );
  AND U28998 ( .A(n28981), .B(n29063), .Z(n29028) );
  XOR U28999 ( .A(n29033), .B(n29032), .Z(n29021) );
  XNOR U29000 ( .A(n29064), .B(n29029), .Z(n29032) );
  XOR U29001 ( .A(n29065), .B(n29066), .Z(n29029) );
  AND U29002 ( .A(n29067), .B(n29068), .Z(n29066) );
  XOR U29003 ( .A(n29065), .B(n29069), .Z(n29067) );
  XNOR U29004 ( .A(n29070), .B(n29071), .Z(n29064) );
  AND U29005 ( .A(n29072), .B(n29073), .Z(n29071) );
  XOR U29006 ( .A(n29070), .B(n29074), .Z(n29072) );
  XOR U29007 ( .A(n29075), .B(n29076), .Z(n29033) );
  AND U29008 ( .A(n29077), .B(n29078), .Z(n29076) );
  XOR U29009 ( .A(n29075), .B(n29079), .Z(n29077) );
  XNOR U29010 ( .A(n28966), .B(n29036), .Z(n29038) );
  XNOR U29011 ( .A(n29080), .B(n29081), .Z(n28966) );
  AND U29012 ( .A(n562), .B(n28973), .Z(n29081) );
  XOR U29013 ( .A(n29080), .B(n28971), .Z(n28973) );
  XOR U29014 ( .A(n29082), .B(n29083), .Z(n29036) );
  AND U29015 ( .A(n29084), .B(n29085), .Z(n29083) );
  XNOR U29016 ( .A(n29082), .B(n28981), .Z(n29085) );
  XOR U29017 ( .A(n29086), .B(n29050), .Z(n28981) );
  XNOR U29018 ( .A(n29087), .B(n29057), .Z(n29050) );
  XOR U29019 ( .A(n29046), .B(n29045), .Z(n29057) );
  XNOR U29020 ( .A(n29088), .B(n29042), .Z(n29045) );
  XOR U29021 ( .A(n29089), .B(n29090), .Z(n29042) );
  AND U29022 ( .A(n29091), .B(n29092), .Z(n29090) );
  XNOR U29023 ( .A(n29093), .B(n29094), .Z(n29091) );
  IV U29024 ( .A(n29089), .Z(n29093) );
  XNOR U29025 ( .A(n29095), .B(n29096), .Z(n29088) );
  NOR U29026 ( .A(n29097), .B(n29098), .Z(n29096) );
  XNOR U29027 ( .A(n29095), .B(n29099), .Z(n29097) );
  XOR U29028 ( .A(n29100), .B(n29101), .Z(n29046) );
  NOR U29029 ( .A(n29102), .B(n29103), .Z(n29101) );
  XNOR U29030 ( .A(n29100), .B(n29104), .Z(n29102) );
  XNOR U29031 ( .A(n29056), .B(n29047), .Z(n29087) );
  XOR U29032 ( .A(n29105), .B(n29106), .Z(n29047) );
  AND U29033 ( .A(n29107), .B(n29108), .Z(n29106) );
  XOR U29034 ( .A(n29105), .B(n29109), .Z(n29107) );
  XOR U29035 ( .A(n29110), .B(n29062), .Z(n29056) );
  XOR U29036 ( .A(n29111), .B(n29112), .Z(n29062) );
  NOR U29037 ( .A(n29113), .B(n29114), .Z(n29112) );
  XOR U29038 ( .A(n29111), .B(n29115), .Z(n29113) );
  XNOR U29039 ( .A(n29061), .B(n29053), .Z(n29110) );
  XOR U29040 ( .A(n29116), .B(n29117), .Z(n29053) );
  AND U29041 ( .A(n29118), .B(n29119), .Z(n29117) );
  XOR U29042 ( .A(n29116), .B(n29120), .Z(n29118) );
  XNOR U29043 ( .A(n29121), .B(n29058), .Z(n29061) );
  XOR U29044 ( .A(n29122), .B(n29123), .Z(n29058) );
  AND U29045 ( .A(n29124), .B(n29125), .Z(n29123) );
  XNOR U29046 ( .A(n29126), .B(n29127), .Z(n29124) );
  IV U29047 ( .A(n29122), .Z(n29126) );
  XNOR U29048 ( .A(n29128), .B(n29129), .Z(n29121) );
  NOR U29049 ( .A(n29130), .B(n29131), .Z(n29129) );
  XNOR U29050 ( .A(n29128), .B(n29132), .Z(n29130) );
  XOR U29051 ( .A(n29051), .B(n29063), .Z(n29086) );
  NOR U29052 ( .A(n28989), .B(n29133), .Z(n29063) );
  XNOR U29053 ( .A(n29069), .B(n29068), .Z(n29051) );
  XNOR U29054 ( .A(n29134), .B(n29074), .Z(n29068) );
  XNOR U29055 ( .A(n29135), .B(n29136), .Z(n29074) );
  NOR U29056 ( .A(n29137), .B(n29138), .Z(n29136) );
  XOR U29057 ( .A(n29135), .B(n29139), .Z(n29137) );
  XNOR U29058 ( .A(n29073), .B(n29065), .Z(n29134) );
  XOR U29059 ( .A(n29140), .B(n29141), .Z(n29065) );
  AND U29060 ( .A(n29142), .B(n29143), .Z(n29141) );
  XOR U29061 ( .A(n29140), .B(n29144), .Z(n29142) );
  XNOR U29062 ( .A(n29145), .B(n29070), .Z(n29073) );
  XOR U29063 ( .A(n29146), .B(n29147), .Z(n29070) );
  AND U29064 ( .A(n29148), .B(n29149), .Z(n29147) );
  XNOR U29065 ( .A(n29150), .B(n29151), .Z(n29148) );
  IV U29066 ( .A(n29146), .Z(n29150) );
  XNOR U29067 ( .A(n29152), .B(n29153), .Z(n29145) );
  NOR U29068 ( .A(n29154), .B(n29155), .Z(n29153) );
  XNOR U29069 ( .A(n29152), .B(n29156), .Z(n29154) );
  XOR U29070 ( .A(n29079), .B(n29078), .Z(n29069) );
  XNOR U29071 ( .A(n29157), .B(n29075), .Z(n29078) );
  XOR U29072 ( .A(n29158), .B(n29159), .Z(n29075) );
  AND U29073 ( .A(n29160), .B(n29161), .Z(n29159) );
  XNOR U29074 ( .A(n29162), .B(n29163), .Z(n29160) );
  IV U29075 ( .A(n29158), .Z(n29162) );
  XNOR U29076 ( .A(n29164), .B(n29165), .Z(n29157) );
  NOR U29077 ( .A(n29166), .B(n29167), .Z(n29165) );
  XNOR U29078 ( .A(n29164), .B(n29168), .Z(n29166) );
  XOR U29079 ( .A(n29169), .B(n29170), .Z(n29079) );
  NOR U29080 ( .A(n29171), .B(n29172), .Z(n29170) );
  XNOR U29081 ( .A(n29169), .B(n29173), .Z(n29171) );
  XNOR U29082 ( .A(n28978), .B(n29082), .Z(n29084) );
  XNOR U29083 ( .A(n29174), .B(n29175), .Z(n28978) );
  AND U29084 ( .A(n562), .B(n28985), .Z(n29175) );
  XOR U29085 ( .A(n29174), .B(n28983), .Z(n28985) );
  AND U29086 ( .A(n28986), .B(n28989), .Z(n29082) );
  XOR U29087 ( .A(n29176), .B(n29133), .Z(n28989) );
  XNOR U29088 ( .A(p_input[1440]), .B(p_input[2048]), .Z(n29133) );
  XNOR U29089 ( .A(n29109), .B(n29108), .Z(n29176) );
  XNOR U29090 ( .A(n29177), .B(n29120), .Z(n29108) );
  XOR U29091 ( .A(n29094), .B(n29092), .Z(n29120) );
  XNOR U29092 ( .A(n29178), .B(n29099), .Z(n29092) );
  XOR U29093 ( .A(p_input[1464]), .B(p_input[2072]), .Z(n29099) );
  XOR U29094 ( .A(n29089), .B(n29098), .Z(n29178) );
  XOR U29095 ( .A(n29179), .B(n29095), .Z(n29098) );
  XOR U29096 ( .A(p_input[1462]), .B(p_input[2070]), .Z(n29095) );
  XOR U29097 ( .A(p_input[1463]), .B(n17295), .Z(n29179) );
  XOR U29098 ( .A(p_input[1458]), .B(p_input[2066]), .Z(n29089) );
  XNOR U29099 ( .A(n29104), .B(n29103), .Z(n29094) );
  XOR U29100 ( .A(n29180), .B(n29100), .Z(n29103) );
  XOR U29101 ( .A(p_input[1459]), .B(p_input[2067]), .Z(n29100) );
  XOR U29102 ( .A(p_input[1460]), .B(n17297), .Z(n29180) );
  XOR U29103 ( .A(p_input[1461]), .B(p_input[2069]), .Z(n29104) );
  XOR U29104 ( .A(n29119), .B(n29181), .Z(n29177) );
  IV U29105 ( .A(n29105), .Z(n29181) );
  XOR U29106 ( .A(p_input[1441]), .B(p_input[2049]), .Z(n29105) );
  XNOR U29107 ( .A(n29182), .B(n29127), .Z(n29119) );
  XNOR U29108 ( .A(n29115), .B(n29114), .Z(n29127) );
  XNOR U29109 ( .A(n29183), .B(n29111), .Z(n29114) );
  XNOR U29110 ( .A(p_input[1466]), .B(p_input[2074]), .Z(n29111) );
  XOR U29111 ( .A(p_input[1467]), .B(n17300), .Z(n29183) );
  XOR U29112 ( .A(p_input[1468]), .B(p_input[2076]), .Z(n29115) );
  XOR U29113 ( .A(n29125), .B(n29184), .Z(n29182) );
  IV U29114 ( .A(n29116), .Z(n29184) );
  XOR U29115 ( .A(p_input[1457]), .B(p_input[2065]), .Z(n29116) );
  XNOR U29116 ( .A(n29185), .B(n29132), .Z(n29125) );
  XNOR U29117 ( .A(p_input[1471]), .B(n17303), .Z(n29132) );
  XOR U29118 ( .A(n29122), .B(n29131), .Z(n29185) );
  XOR U29119 ( .A(n29186), .B(n29128), .Z(n29131) );
  XOR U29120 ( .A(p_input[1469]), .B(p_input[2077]), .Z(n29128) );
  XOR U29121 ( .A(p_input[1470]), .B(n17305), .Z(n29186) );
  XOR U29122 ( .A(p_input[1465]), .B(p_input[2073]), .Z(n29122) );
  XOR U29123 ( .A(n29144), .B(n29143), .Z(n29109) );
  XNOR U29124 ( .A(n29187), .B(n29151), .Z(n29143) );
  XNOR U29125 ( .A(n29139), .B(n29138), .Z(n29151) );
  XNOR U29126 ( .A(n29188), .B(n29135), .Z(n29138) );
  XNOR U29127 ( .A(p_input[1451]), .B(p_input[2059]), .Z(n29135) );
  XOR U29128 ( .A(p_input[1452]), .B(n16451), .Z(n29188) );
  XOR U29129 ( .A(p_input[1453]), .B(p_input[2061]), .Z(n29139) );
  XOR U29130 ( .A(n29149), .B(n29189), .Z(n29187) );
  IV U29131 ( .A(n29140), .Z(n29189) );
  XOR U29132 ( .A(p_input[1442]), .B(p_input[2050]), .Z(n29140) );
  XNOR U29133 ( .A(n29190), .B(n29156), .Z(n29149) );
  XNOR U29134 ( .A(p_input[1456]), .B(n16454), .Z(n29156) );
  XOR U29135 ( .A(n29146), .B(n29155), .Z(n29190) );
  XOR U29136 ( .A(n29191), .B(n29152), .Z(n29155) );
  XOR U29137 ( .A(p_input[1454]), .B(p_input[2062]), .Z(n29152) );
  XOR U29138 ( .A(p_input[1455]), .B(n16456), .Z(n29191) );
  XOR U29139 ( .A(p_input[1450]), .B(p_input[2058]), .Z(n29146) );
  XOR U29140 ( .A(n29163), .B(n29161), .Z(n29144) );
  XNOR U29141 ( .A(n29192), .B(n29168), .Z(n29161) );
  XOR U29142 ( .A(p_input[1449]), .B(p_input[2057]), .Z(n29168) );
  XOR U29143 ( .A(n29158), .B(n29167), .Z(n29192) );
  XOR U29144 ( .A(n29193), .B(n29164), .Z(n29167) );
  XOR U29145 ( .A(p_input[1447]), .B(p_input[2055]), .Z(n29164) );
  XOR U29146 ( .A(p_input[1448]), .B(n17312), .Z(n29193) );
  XOR U29147 ( .A(p_input[1443]), .B(p_input[2051]), .Z(n29158) );
  XNOR U29148 ( .A(n29173), .B(n29172), .Z(n29163) );
  XOR U29149 ( .A(n29194), .B(n29169), .Z(n29172) );
  XOR U29150 ( .A(p_input[1444]), .B(p_input[2052]), .Z(n29169) );
  XOR U29151 ( .A(p_input[1445]), .B(n17314), .Z(n29194) );
  XOR U29152 ( .A(p_input[1446]), .B(p_input[2054]), .Z(n29173) );
  XNOR U29153 ( .A(n29195), .B(n29196), .Z(n28986) );
  AND U29154 ( .A(n562), .B(n29197), .Z(n29196) );
  XNOR U29155 ( .A(n29198), .B(n29199), .Z(n562) );
  AND U29156 ( .A(n29200), .B(n29201), .Z(n29199) );
  XOR U29157 ( .A(n29198), .B(n28996), .Z(n29201) );
  XNOR U29158 ( .A(n29198), .B(n28938), .Z(n29200) );
  XOR U29159 ( .A(n29202), .B(n29203), .Z(n29198) );
  AND U29160 ( .A(n29204), .B(n29205), .Z(n29203) );
  XNOR U29161 ( .A(n29009), .B(n29202), .Z(n29205) );
  XOR U29162 ( .A(n29202), .B(n28950), .Z(n29204) );
  XOR U29163 ( .A(n29206), .B(n29207), .Z(n29202) );
  AND U29164 ( .A(n29208), .B(n29209), .Z(n29207) );
  XNOR U29165 ( .A(n29034), .B(n29206), .Z(n29209) );
  XOR U29166 ( .A(n29206), .B(n28961), .Z(n29208) );
  XOR U29167 ( .A(n29210), .B(n29211), .Z(n29206) );
  AND U29168 ( .A(n29212), .B(n29213), .Z(n29211) );
  XOR U29169 ( .A(n29210), .B(n28971), .Z(n29212) );
  XOR U29170 ( .A(n29214), .B(n29215), .Z(n28927) );
  AND U29171 ( .A(n566), .B(n29197), .Z(n29215) );
  XNOR U29172 ( .A(n29195), .B(n29214), .Z(n29197) );
  XNOR U29173 ( .A(n29216), .B(n29217), .Z(n566) );
  AND U29174 ( .A(n29218), .B(n29219), .Z(n29217) );
  XNOR U29175 ( .A(n29220), .B(n29216), .Z(n29219) );
  IV U29176 ( .A(n28996), .Z(n29220) );
  XNOR U29177 ( .A(n29221), .B(n29222), .Z(n28996) );
  AND U29178 ( .A(n569), .B(n29223), .Z(n29222) );
  XNOR U29179 ( .A(n29221), .B(n29224), .Z(n29223) );
  XNOR U29180 ( .A(n28938), .B(n29216), .Z(n29218) );
  XOR U29181 ( .A(n29225), .B(n29226), .Z(n28938) );
  AND U29182 ( .A(n577), .B(n29227), .Z(n29226) );
  XOR U29183 ( .A(n29228), .B(n29229), .Z(n29216) );
  AND U29184 ( .A(n29230), .B(n29231), .Z(n29229) );
  XNOR U29185 ( .A(n29228), .B(n29009), .Z(n29231) );
  XNOR U29186 ( .A(n29232), .B(n29233), .Z(n29009) );
  AND U29187 ( .A(n569), .B(n29234), .Z(n29233) );
  XOR U29188 ( .A(n29235), .B(n29232), .Z(n29234) );
  XNOR U29189 ( .A(n29236), .B(n29228), .Z(n29230) );
  IV U29190 ( .A(n28950), .Z(n29236) );
  XOR U29191 ( .A(n29237), .B(n29238), .Z(n28950) );
  AND U29192 ( .A(n577), .B(n29239), .Z(n29238) );
  XOR U29193 ( .A(n29240), .B(n29241), .Z(n29228) );
  AND U29194 ( .A(n29242), .B(n29243), .Z(n29241) );
  XNOR U29195 ( .A(n29240), .B(n29034), .Z(n29243) );
  XNOR U29196 ( .A(n29244), .B(n29245), .Z(n29034) );
  AND U29197 ( .A(n569), .B(n29246), .Z(n29245) );
  XNOR U29198 ( .A(n29247), .B(n29244), .Z(n29246) );
  XOR U29199 ( .A(n28961), .B(n29240), .Z(n29242) );
  XOR U29200 ( .A(n29248), .B(n29249), .Z(n28961) );
  AND U29201 ( .A(n577), .B(n29250), .Z(n29249) );
  XOR U29202 ( .A(n29210), .B(n29251), .Z(n29240) );
  AND U29203 ( .A(n29252), .B(n29213), .Z(n29251) );
  XNOR U29204 ( .A(n29080), .B(n29210), .Z(n29213) );
  XNOR U29205 ( .A(n29253), .B(n29254), .Z(n29080) );
  AND U29206 ( .A(n569), .B(n29255), .Z(n29254) );
  XOR U29207 ( .A(n29256), .B(n29253), .Z(n29255) );
  XNOR U29208 ( .A(n29257), .B(n29210), .Z(n29252) );
  IV U29209 ( .A(n28971), .Z(n29257) );
  XOR U29210 ( .A(n29258), .B(n29259), .Z(n28971) );
  AND U29211 ( .A(n577), .B(n29260), .Z(n29259) );
  XOR U29212 ( .A(n29261), .B(n29262), .Z(n29210) );
  AND U29213 ( .A(n29263), .B(n29264), .Z(n29262) );
  XNOR U29214 ( .A(n29261), .B(n29174), .Z(n29264) );
  XNOR U29215 ( .A(n29265), .B(n29266), .Z(n29174) );
  AND U29216 ( .A(n569), .B(n29267), .Z(n29266) );
  XNOR U29217 ( .A(n29268), .B(n29265), .Z(n29267) );
  XNOR U29218 ( .A(n29269), .B(n29261), .Z(n29263) );
  IV U29219 ( .A(n28983), .Z(n29269) );
  XOR U29220 ( .A(n29270), .B(n29271), .Z(n28983) );
  AND U29221 ( .A(n577), .B(n29272), .Z(n29271) );
  AND U29222 ( .A(n29214), .B(n29195), .Z(n29261) );
  XNOR U29223 ( .A(n29273), .B(n29274), .Z(n29195) );
  AND U29224 ( .A(n569), .B(n29275), .Z(n29274) );
  XNOR U29225 ( .A(n29276), .B(n29273), .Z(n29275) );
  XNOR U29226 ( .A(n29277), .B(n29278), .Z(n569) );
  AND U29227 ( .A(n29279), .B(n29280), .Z(n29278) );
  XOR U29228 ( .A(n29224), .B(n29277), .Z(n29280) );
  AND U29229 ( .A(n29281), .B(n29282), .Z(n29224) );
  XOR U29230 ( .A(n29277), .B(n29221), .Z(n29279) );
  XNOR U29231 ( .A(n29283), .B(n29284), .Z(n29221) );
  AND U29232 ( .A(n573), .B(n29227), .Z(n29284) );
  XOR U29233 ( .A(n29225), .B(n29283), .Z(n29227) );
  XOR U29234 ( .A(n29285), .B(n29286), .Z(n29277) );
  AND U29235 ( .A(n29287), .B(n29288), .Z(n29286) );
  XNOR U29236 ( .A(n29285), .B(n29281), .Z(n29288) );
  IV U29237 ( .A(n29235), .Z(n29281) );
  XOR U29238 ( .A(n29289), .B(n29290), .Z(n29235) );
  XOR U29239 ( .A(n29291), .B(n29282), .Z(n29290) );
  AND U29240 ( .A(n29247), .B(n29292), .Z(n29282) );
  AND U29241 ( .A(n29293), .B(n29294), .Z(n29291) );
  XOR U29242 ( .A(n29295), .B(n29289), .Z(n29293) );
  XNOR U29243 ( .A(n29232), .B(n29285), .Z(n29287) );
  XNOR U29244 ( .A(n29296), .B(n29297), .Z(n29232) );
  AND U29245 ( .A(n573), .B(n29239), .Z(n29297) );
  XOR U29246 ( .A(n29296), .B(n29237), .Z(n29239) );
  XOR U29247 ( .A(n29298), .B(n29299), .Z(n29285) );
  AND U29248 ( .A(n29300), .B(n29301), .Z(n29299) );
  XNOR U29249 ( .A(n29298), .B(n29247), .Z(n29301) );
  XOR U29250 ( .A(n29302), .B(n29294), .Z(n29247) );
  XNOR U29251 ( .A(n29303), .B(n29289), .Z(n29294) );
  XOR U29252 ( .A(n29304), .B(n29305), .Z(n29289) );
  AND U29253 ( .A(n29306), .B(n29307), .Z(n29305) );
  XOR U29254 ( .A(n29308), .B(n29304), .Z(n29306) );
  XNOR U29255 ( .A(n29309), .B(n29310), .Z(n29303) );
  AND U29256 ( .A(n29311), .B(n29312), .Z(n29310) );
  XOR U29257 ( .A(n29309), .B(n29313), .Z(n29311) );
  XNOR U29258 ( .A(n29295), .B(n29292), .Z(n29302) );
  AND U29259 ( .A(n29314), .B(n29315), .Z(n29292) );
  XOR U29260 ( .A(n29316), .B(n29317), .Z(n29295) );
  AND U29261 ( .A(n29318), .B(n29319), .Z(n29317) );
  XOR U29262 ( .A(n29316), .B(n29320), .Z(n29318) );
  XNOR U29263 ( .A(n29244), .B(n29298), .Z(n29300) );
  XNOR U29264 ( .A(n29321), .B(n29322), .Z(n29244) );
  AND U29265 ( .A(n573), .B(n29250), .Z(n29322) );
  XOR U29266 ( .A(n29321), .B(n29248), .Z(n29250) );
  XOR U29267 ( .A(n29323), .B(n29324), .Z(n29298) );
  AND U29268 ( .A(n29325), .B(n29326), .Z(n29324) );
  XNOR U29269 ( .A(n29323), .B(n29314), .Z(n29326) );
  IV U29270 ( .A(n29256), .Z(n29314) );
  XNOR U29271 ( .A(n29327), .B(n29307), .Z(n29256) );
  XNOR U29272 ( .A(n29328), .B(n29313), .Z(n29307) );
  XOR U29273 ( .A(n29329), .B(n29330), .Z(n29313) );
  AND U29274 ( .A(n29331), .B(n29332), .Z(n29330) );
  XOR U29275 ( .A(n29329), .B(n29333), .Z(n29331) );
  XNOR U29276 ( .A(n29312), .B(n29304), .Z(n29328) );
  XOR U29277 ( .A(n29334), .B(n29335), .Z(n29304) );
  AND U29278 ( .A(n29336), .B(n29337), .Z(n29335) );
  XNOR U29279 ( .A(n29338), .B(n29334), .Z(n29336) );
  XNOR U29280 ( .A(n29339), .B(n29309), .Z(n29312) );
  XOR U29281 ( .A(n29340), .B(n29341), .Z(n29309) );
  AND U29282 ( .A(n29342), .B(n29343), .Z(n29341) );
  XOR U29283 ( .A(n29340), .B(n29344), .Z(n29342) );
  XNOR U29284 ( .A(n29345), .B(n29346), .Z(n29339) );
  AND U29285 ( .A(n29347), .B(n29348), .Z(n29346) );
  XNOR U29286 ( .A(n29345), .B(n29349), .Z(n29347) );
  XNOR U29287 ( .A(n29308), .B(n29315), .Z(n29327) );
  AND U29288 ( .A(n29268), .B(n29350), .Z(n29315) );
  XOR U29289 ( .A(n29320), .B(n29319), .Z(n29308) );
  XNOR U29290 ( .A(n29351), .B(n29316), .Z(n29319) );
  XOR U29291 ( .A(n29352), .B(n29353), .Z(n29316) );
  AND U29292 ( .A(n29354), .B(n29355), .Z(n29353) );
  XOR U29293 ( .A(n29352), .B(n29356), .Z(n29354) );
  XNOR U29294 ( .A(n29357), .B(n29358), .Z(n29351) );
  AND U29295 ( .A(n29359), .B(n29360), .Z(n29358) );
  XOR U29296 ( .A(n29357), .B(n29361), .Z(n29359) );
  XOR U29297 ( .A(n29362), .B(n29363), .Z(n29320) );
  AND U29298 ( .A(n29364), .B(n29365), .Z(n29363) );
  XOR U29299 ( .A(n29362), .B(n29366), .Z(n29364) );
  XNOR U29300 ( .A(n29253), .B(n29323), .Z(n29325) );
  XNOR U29301 ( .A(n29367), .B(n29368), .Z(n29253) );
  AND U29302 ( .A(n573), .B(n29260), .Z(n29368) );
  XOR U29303 ( .A(n29367), .B(n29258), .Z(n29260) );
  XOR U29304 ( .A(n29369), .B(n29370), .Z(n29323) );
  AND U29305 ( .A(n29371), .B(n29372), .Z(n29370) );
  XNOR U29306 ( .A(n29369), .B(n29268), .Z(n29372) );
  XOR U29307 ( .A(n29373), .B(n29337), .Z(n29268) );
  XNOR U29308 ( .A(n29374), .B(n29344), .Z(n29337) );
  XOR U29309 ( .A(n29333), .B(n29332), .Z(n29344) );
  XNOR U29310 ( .A(n29375), .B(n29329), .Z(n29332) );
  XOR U29311 ( .A(n29376), .B(n29377), .Z(n29329) );
  AND U29312 ( .A(n29378), .B(n29379), .Z(n29377) );
  XNOR U29313 ( .A(n29380), .B(n29381), .Z(n29378) );
  IV U29314 ( .A(n29376), .Z(n29380) );
  XNOR U29315 ( .A(n29382), .B(n29383), .Z(n29375) );
  NOR U29316 ( .A(n29384), .B(n29385), .Z(n29383) );
  XNOR U29317 ( .A(n29382), .B(n29386), .Z(n29384) );
  XOR U29318 ( .A(n29387), .B(n29388), .Z(n29333) );
  NOR U29319 ( .A(n29389), .B(n29390), .Z(n29388) );
  XNOR U29320 ( .A(n29387), .B(n29391), .Z(n29389) );
  XNOR U29321 ( .A(n29343), .B(n29334), .Z(n29374) );
  XOR U29322 ( .A(n29392), .B(n29393), .Z(n29334) );
  AND U29323 ( .A(n29394), .B(n29395), .Z(n29393) );
  XOR U29324 ( .A(n29392), .B(n29396), .Z(n29394) );
  XOR U29325 ( .A(n29397), .B(n29349), .Z(n29343) );
  XOR U29326 ( .A(n29398), .B(n29399), .Z(n29349) );
  NOR U29327 ( .A(n29400), .B(n29401), .Z(n29399) );
  XOR U29328 ( .A(n29398), .B(n29402), .Z(n29400) );
  XNOR U29329 ( .A(n29348), .B(n29340), .Z(n29397) );
  XOR U29330 ( .A(n29403), .B(n29404), .Z(n29340) );
  AND U29331 ( .A(n29405), .B(n29406), .Z(n29404) );
  XOR U29332 ( .A(n29403), .B(n29407), .Z(n29405) );
  XNOR U29333 ( .A(n29408), .B(n29345), .Z(n29348) );
  XOR U29334 ( .A(n29409), .B(n29410), .Z(n29345) );
  AND U29335 ( .A(n29411), .B(n29412), .Z(n29410) );
  XNOR U29336 ( .A(n29413), .B(n29414), .Z(n29411) );
  IV U29337 ( .A(n29409), .Z(n29413) );
  XNOR U29338 ( .A(n29415), .B(n29416), .Z(n29408) );
  NOR U29339 ( .A(n29417), .B(n29418), .Z(n29416) );
  XNOR U29340 ( .A(n29415), .B(n29419), .Z(n29417) );
  XOR U29341 ( .A(n29338), .B(n29350), .Z(n29373) );
  NOR U29342 ( .A(n29276), .B(n29420), .Z(n29350) );
  XNOR U29343 ( .A(n29356), .B(n29355), .Z(n29338) );
  XNOR U29344 ( .A(n29421), .B(n29361), .Z(n29355) );
  XNOR U29345 ( .A(n29422), .B(n29423), .Z(n29361) );
  NOR U29346 ( .A(n29424), .B(n29425), .Z(n29423) );
  XOR U29347 ( .A(n29422), .B(n29426), .Z(n29424) );
  XNOR U29348 ( .A(n29360), .B(n29352), .Z(n29421) );
  XOR U29349 ( .A(n29427), .B(n29428), .Z(n29352) );
  AND U29350 ( .A(n29429), .B(n29430), .Z(n29428) );
  XOR U29351 ( .A(n29427), .B(n29431), .Z(n29429) );
  XNOR U29352 ( .A(n29432), .B(n29357), .Z(n29360) );
  XOR U29353 ( .A(n29433), .B(n29434), .Z(n29357) );
  AND U29354 ( .A(n29435), .B(n29436), .Z(n29434) );
  XNOR U29355 ( .A(n29437), .B(n29438), .Z(n29435) );
  IV U29356 ( .A(n29433), .Z(n29437) );
  XNOR U29357 ( .A(n29439), .B(n29440), .Z(n29432) );
  NOR U29358 ( .A(n29441), .B(n29442), .Z(n29440) );
  XNOR U29359 ( .A(n29439), .B(n29443), .Z(n29441) );
  XOR U29360 ( .A(n29366), .B(n29365), .Z(n29356) );
  XNOR U29361 ( .A(n29444), .B(n29362), .Z(n29365) );
  XOR U29362 ( .A(n29445), .B(n29446), .Z(n29362) );
  AND U29363 ( .A(n29447), .B(n29448), .Z(n29446) );
  XNOR U29364 ( .A(n29449), .B(n29450), .Z(n29447) );
  IV U29365 ( .A(n29445), .Z(n29449) );
  XNOR U29366 ( .A(n29451), .B(n29452), .Z(n29444) );
  NOR U29367 ( .A(n29453), .B(n29454), .Z(n29452) );
  XNOR U29368 ( .A(n29451), .B(n29455), .Z(n29453) );
  XOR U29369 ( .A(n29456), .B(n29457), .Z(n29366) );
  NOR U29370 ( .A(n29458), .B(n29459), .Z(n29457) );
  XNOR U29371 ( .A(n29456), .B(n29460), .Z(n29458) );
  XNOR U29372 ( .A(n29265), .B(n29369), .Z(n29371) );
  XNOR U29373 ( .A(n29461), .B(n29462), .Z(n29265) );
  AND U29374 ( .A(n573), .B(n29272), .Z(n29462) );
  XOR U29375 ( .A(n29461), .B(n29270), .Z(n29272) );
  AND U29376 ( .A(n29273), .B(n29276), .Z(n29369) );
  XOR U29377 ( .A(n29463), .B(n29420), .Z(n29276) );
  XNOR U29378 ( .A(p_input[1472]), .B(p_input[2048]), .Z(n29420) );
  XNOR U29379 ( .A(n29396), .B(n29395), .Z(n29463) );
  XNOR U29380 ( .A(n29464), .B(n29407), .Z(n29395) );
  XOR U29381 ( .A(n29381), .B(n29379), .Z(n29407) );
  XNOR U29382 ( .A(n29465), .B(n29386), .Z(n29379) );
  XOR U29383 ( .A(p_input[1496]), .B(p_input[2072]), .Z(n29386) );
  XOR U29384 ( .A(n29376), .B(n29385), .Z(n29465) );
  XOR U29385 ( .A(n29466), .B(n29382), .Z(n29385) );
  XOR U29386 ( .A(p_input[1494]), .B(p_input[2070]), .Z(n29382) );
  XOR U29387 ( .A(p_input[1495]), .B(n17295), .Z(n29466) );
  XOR U29388 ( .A(p_input[1490]), .B(p_input[2066]), .Z(n29376) );
  XNOR U29389 ( .A(n29391), .B(n29390), .Z(n29381) );
  XOR U29390 ( .A(n29467), .B(n29387), .Z(n29390) );
  XOR U29391 ( .A(p_input[1491]), .B(p_input[2067]), .Z(n29387) );
  XOR U29392 ( .A(p_input[1492]), .B(n17297), .Z(n29467) );
  XOR U29393 ( .A(p_input[1493]), .B(p_input[2069]), .Z(n29391) );
  XOR U29394 ( .A(n29406), .B(n29468), .Z(n29464) );
  IV U29395 ( .A(n29392), .Z(n29468) );
  XOR U29396 ( .A(p_input[1473]), .B(p_input[2049]), .Z(n29392) );
  XNOR U29397 ( .A(n29469), .B(n29414), .Z(n29406) );
  XNOR U29398 ( .A(n29402), .B(n29401), .Z(n29414) );
  XNOR U29399 ( .A(n29470), .B(n29398), .Z(n29401) );
  XNOR U29400 ( .A(p_input[1498]), .B(p_input[2074]), .Z(n29398) );
  XOR U29401 ( .A(p_input[1499]), .B(n17300), .Z(n29470) );
  XOR U29402 ( .A(p_input[1500]), .B(p_input[2076]), .Z(n29402) );
  XOR U29403 ( .A(n29412), .B(n29471), .Z(n29469) );
  IV U29404 ( .A(n29403), .Z(n29471) );
  XOR U29405 ( .A(p_input[1489]), .B(p_input[2065]), .Z(n29403) );
  XNOR U29406 ( .A(n29472), .B(n29419), .Z(n29412) );
  XNOR U29407 ( .A(p_input[1503]), .B(n17303), .Z(n29419) );
  XOR U29408 ( .A(n29409), .B(n29418), .Z(n29472) );
  XOR U29409 ( .A(n29473), .B(n29415), .Z(n29418) );
  XOR U29410 ( .A(p_input[1501]), .B(p_input[2077]), .Z(n29415) );
  XOR U29411 ( .A(p_input[1502]), .B(n17305), .Z(n29473) );
  XOR U29412 ( .A(p_input[1497]), .B(p_input[2073]), .Z(n29409) );
  XOR U29413 ( .A(n29431), .B(n29430), .Z(n29396) );
  XNOR U29414 ( .A(n29474), .B(n29438), .Z(n29430) );
  XNOR U29415 ( .A(n29426), .B(n29425), .Z(n29438) );
  XNOR U29416 ( .A(n29475), .B(n29422), .Z(n29425) );
  XNOR U29417 ( .A(p_input[1483]), .B(p_input[2059]), .Z(n29422) );
  XOR U29418 ( .A(p_input[1484]), .B(n16451), .Z(n29475) );
  XOR U29419 ( .A(p_input[1485]), .B(p_input[2061]), .Z(n29426) );
  XOR U29420 ( .A(n29436), .B(n29476), .Z(n29474) );
  IV U29421 ( .A(n29427), .Z(n29476) );
  XOR U29422 ( .A(p_input[1474]), .B(p_input[2050]), .Z(n29427) );
  XNOR U29423 ( .A(n29477), .B(n29443), .Z(n29436) );
  XNOR U29424 ( .A(p_input[1488]), .B(n16454), .Z(n29443) );
  XOR U29425 ( .A(n29433), .B(n29442), .Z(n29477) );
  XOR U29426 ( .A(n29478), .B(n29439), .Z(n29442) );
  XOR U29427 ( .A(p_input[1486]), .B(p_input[2062]), .Z(n29439) );
  XOR U29428 ( .A(p_input[1487]), .B(n16456), .Z(n29478) );
  XOR U29429 ( .A(p_input[1482]), .B(p_input[2058]), .Z(n29433) );
  XOR U29430 ( .A(n29450), .B(n29448), .Z(n29431) );
  XNOR U29431 ( .A(n29479), .B(n29455), .Z(n29448) );
  XOR U29432 ( .A(p_input[1481]), .B(p_input[2057]), .Z(n29455) );
  XOR U29433 ( .A(n29445), .B(n29454), .Z(n29479) );
  XOR U29434 ( .A(n29480), .B(n29451), .Z(n29454) );
  XOR U29435 ( .A(p_input[1479]), .B(p_input[2055]), .Z(n29451) );
  XOR U29436 ( .A(p_input[1480]), .B(n17312), .Z(n29480) );
  XOR U29437 ( .A(p_input[1475]), .B(p_input[2051]), .Z(n29445) );
  XNOR U29438 ( .A(n29460), .B(n29459), .Z(n29450) );
  XOR U29439 ( .A(n29481), .B(n29456), .Z(n29459) );
  XOR U29440 ( .A(p_input[1476]), .B(p_input[2052]), .Z(n29456) );
  XOR U29441 ( .A(p_input[1477]), .B(n17314), .Z(n29481) );
  XOR U29442 ( .A(p_input[1478]), .B(p_input[2054]), .Z(n29460) );
  XNOR U29443 ( .A(n29482), .B(n29483), .Z(n29273) );
  AND U29444 ( .A(n573), .B(n29484), .Z(n29483) );
  XNOR U29445 ( .A(n29485), .B(n29486), .Z(n573) );
  AND U29446 ( .A(n29487), .B(n29488), .Z(n29486) );
  XOR U29447 ( .A(n29485), .B(n29283), .Z(n29488) );
  XNOR U29448 ( .A(n29485), .B(n29225), .Z(n29487) );
  XOR U29449 ( .A(n29489), .B(n29490), .Z(n29485) );
  AND U29450 ( .A(n29491), .B(n29492), .Z(n29490) );
  XNOR U29451 ( .A(n29296), .B(n29489), .Z(n29492) );
  XOR U29452 ( .A(n29489), .B(n29237), .Z(n29491) );
  XOR U29453 ( .A(n29493), .B(n29494), .Z(n29489) );
  AND U29454 ( .A(n29495), .B(n29496), .Z(n29494) );
  XNOR U29455 ( .A(n29321), .B(n29493), .Z(n29496) );
  XOR U29456 ( .A(n29493), .B(n29248), .Z(n29495) );
  XOR U29457 ( .A(n29497), .B(n29498), .Z(n29493) );
  AND U29458 ( .A(n29499), .B(n29500), .Z(n29498) );
  XOR U29459 ( .A(n29497), .B(n29258), .Z(n29499) );
  XOR U29460 ( .A(n29501), .B(n29502), .Z(n29214) );
  AND U29461 ( .A(n577), .B(n29484), .Z(n29502) );
  XNOR U29462 ( .A(n29482), .B(n29501), .Z(n29484) );
  XNOR U29463 ( .A(n29503), .B(n29504), .Z(n577) );
  AND U29464 ( .A(n29505), .B(n29506), .Z(n29504) );
  XNOR U29465 ( .A(n29507), .B(n29503), .Z(n29506) );
  IV U29466 ( .A(n29283), .Z(n29507) );
  XNOR U29467 ( .A(n29508), .B(n29509), .Z(n29283) );
  AND U29468 ( .A(n580), .B(n29510), .Z(n29509) );
  XNOR U29469 ( .A(n29508), .B(n29511), .Z(n29510) );
  XNOR U29470 ( .A(n29225), .B(n29503), .Z(n29505) );
  XOR U29471 ( .A(n29512), .B(n29513), .Z(n29225) );
  AND U29472 ( .A(n588), .B(n29514), .Z(n29513) );
  XOR U29473 ( .A(n29515), .B(n29516), .Z(n29503) );
  AND U29474 ( .A(n29517), .B(n29518), .Z(n29516) );
  XNOR U29475 ( .A(n29515), .B(n29296), .Z(n29518) );
  XNOR U29476 ( .A(n29519), .B(n29520), .Z(n29296) );
  AND U29477 ( .A(n580), .B(n29521), .Z(n29520) );
  XOR U29478 ( .A(n29522), .B(n29519), .Z(n29521) );
  XNOR U29479 ( .A(n29523), .B(n29515), .Z(n29517) );
  IV U29480 ( .A(n29237), .Z(n29523) );
  XOR U29481 ( .A(n29524), .B(n29525), .Z(n29237) );
  AND U29482 ( .A(n588), .B(n29526), .Z(n29525) );
  XOR U29483 ( .A(n29527), .B(n29528), .Z(n29515) );
  AND U29484 ( .A(n29529), .B(n29530), .Z(n29528) );
  XNOR U29485 ( .A(n29527), .B(n29321), .Z(n29530) );
  XNOR U29486 ( .A(n29531), .B(n29532), .Z(n29321) );
  AND U29487 ( .A(n580), .B(n29533), .Z(n29532) );
  XNOR U29488 ( .A(n29534), .B(n29531), .Z(n29533) );
  XOR U29489 ( .A(n29248), .B(n29527), .Z(n29529) );
  XOR U29490 ( .A(n29535), .B(n29536), .Z(n29248) );
  AND U29491 ( .A(n588), .B(n29537), .Z(n29536) );
  XOR U29492 ( .A(n29497), .B(n29538), .Z(n29527) );
  AND U29493 ( .A(n29539), .B(n29500), .Z(n29538) );
  XNOR U29494 ( .A(n29367), .B(n29497), .Z(n29500) );
  XNOR U29495 ( .A(n29540), .B(n29541), .Z(n29367) );
  AND U29496 ( .A(n580), .B(n29542), .Z(n29541) );
  XOR U29497 ( .A(n29543), .B(n29540), .Z(n29542) );
  XNOR U29498 ( .A(n29544), .B(n29497), .Z(n29539) );
  IV U29499 ( .A(n29258), .Z(n29544) );
  XOR U29500 ( .A(n29545), .B(n29546), .Z(n29258) );
  AND U29501 ( .A(n588), .B(n29547), .Z(n29546) );
  XOR U29502 ( .A(n29548), .B(n29549), .Z(n29497) );
  AND U29503 ( .A(n29550), .B(n29551), .Z(n29549) );
  XNOR U29504 ( .A(n29548), .B(n29461), .Z(n29551) );
  XNOR U29505 ( .A(n29552), .B(n29553), .Z(n29461) );
  AND U29506 ( .A(n580), .B(n29554), .Z(n29553) );
  XNOR U29507 ( .A(n29555), .B(n29552), .Z(n29554) );
  XNOR U29508 ( .A(n29556), .B(n29548), .Z(n29550) );
  IV U29509 ( .A(n29270), .Z(n29556) );
  XOR U29510 ( .A(n29557), .B(n29558), .Z(n29270) );
  AND U29511 ( .A(n588), .B(n29559), .Z(n29558) );
  AND U29512 ( .A(n29501), .B(n29482), .Z(n29548) );
  XNOR U29513 ( .A(n29560), .B(n29561), .Z(n29482) );
  AND U29514 ( .A(n580), .B(n29562), .Z(n29561) );
  XNOR U29515 ( .A(n29563), .B(n29560), .Z(n29562) );
  XNOR U29516 ( .A(n29564), .B(n29565), .Z(n580) );
  AND U29517 ( .A(n29566), .B(n29567), .Z(n29565) );
  XOR U29518 ( .A(n29511), .B(n29564), .Z(n29567) );
  AND U29519 ( .A(n29568), .B(n29569), .Z(n29511) );
  XOR U29520 ( .A(n29564), .B(n29508), .Z(n29566) );
  XNOR U29521 ( .A(n29570), .B(n29571), .Z(n29508) );
  AND U29522 ( .A(n584), .B(n29514), .Z(n29571) );
  XOR U29523 ( .A(n29512), .B(n29570), .Z(n29514) );
  XOR U29524 ( .A(n29572), .B(n29573), .Z(n29564) );
  AND U29525 ( .A(n29574), .B(n29575), .Z(n29573) );
  XNOR U29526 ( .A(n29572), .B(n29568), .Z(n29575) );
  IV U29527 ( .A(n29522), .Z(n29568) );
  XOR U29528 ( .A(n29576), .B(n29577), .Z(n29522) );
  XOR U29529 ( .A(n29578), .B(n29569), .Z(n29577) );
  AND U29530 ( .A(n29534), .B(n29579), .Z(n29569) );
  AND U29531 ( .A(n29580), .B(n29581), .Z(n29578) );
  XOR U29532 ( .A(n29582), .B(n29576), .Z(n29580) );
  XNOR U29533 ( .A(n29519), .B(n29572), .Z(n29574) );
  XNOR U29534 ( .A(n29583), .B(n29584), .Z(n29519) );
  AND U29535 ( .A(n584), .B(n29526), .Z(n29584) );
  XOR U29536 ( .A(n29583), .B(n29524), .Z(n29526) );
  XOR U29537 ( .A(n29585), .B(n29586), .Z(n29572) );
  AND U29538 ( .A(n29587), .B(n29588), .Z(n29586) );
  XNOR U29539 ( .A(n29585), .B(n29534), .Z(n29588) );
  XOR U29540 ( .A(n29589), .B(n29581), .Z(n29534) );
  XNOR U29541 ( .A(n29590), .B(n29576), .Z(n29581) );
  XOR U29542 ( .A(n29591), .B(n29592), .Z(n29576) );
  AND U29543 ( .A(n29593), .B(n29594), .Z(n29592) );
  XOR U29544 ( .A(n29595), .B(n29591), .Z(n29593) );
  XNOR U29545 ( .A(n29596), .B(n29597), .Z(n29590) );
  AND U29546 ( .A(n29598), .B(n29599), .Z(n29597) );
  XOR U29547 ( .A(n29596), .B(n29600), .Z(n29598) );
  XNOR U29548 ( .A(n29582), .B(n29579), .Z(n29589) );
  AND U29549 ( .A(n29601), .B(n29602), .Z(n29579) );
  XOR U29550 ( .A(n29603), .B(n29604), .Z(n29582) );
  AND U29551 ( .A(n29605), .B(n29606), .Z(n29604) );
  XOR U29552 ( .A(n29603), .B(n29607), .Z(n29605) );
  XNOR U29553 ( .A(n29531), .B(n29585), .Z(n29587) );
  XNOR U29554 ( .A(n29608), .B(n29609), .Z(n29531) );
  AND U29555 ( .A(n584), .B(n29537), .Z(n29609) );
  XOR U29556 ( .A(n29608), .B(n29535), .Z(n29537) );
  XOR U29557 ( .A(n29610), .B(n29611), .Z(n29585) );
  AND U29558 ( .A(n29612), .B(n29613), .Z(n29611) );
  XNOR U29559 ( .A(n29610), .B(n29601), .Z(n29613) );
  IV U29560 ( .A(n29543), .Z(n29601) );
  XNOR U29561 ( .A(n29614), .B(n29594), .Z(n29543) );
  XNOR U29562 ( .A(n29615), .B(n29600), .Z(n29594) );
  XOR U29563 ( .A(n29616), .B(n29617), .Z(n29600) );
  AND U29564 ( .A(n29618), .B(n29619), .Z(n29617) );
  XOR U29565 ( .A(n29616), .B(n29620), .Z(n29618) );
  XNOR U29566 ( .A(n29599), .B(n29591), .Z(n29615) );
  XOR U29567 ( .A(n29621), .B(n29622), .Z(n29591) );
  AND U29568 ( .A(n29623), .B(n29624), .Z(n29622) );
  XNOR U29569 ( .A(n29625), .B(n29621), .Z(n29623) );
  XNOR U29570 ( .A(n29626), .B(n29596), .Z(n29599) );
  XOR U29571 ( .A(n29627), .B(n29628), .Z(n29596) );
  AND U29572 ( .A(n29629), .B(n29630), .Z(n29628) );
  XOR U29573 ( .A(n29627), .B(n29631), .Z(n29629) );
  XNOR U29574 ( .A(n29632), .B(n29633), .Z(n29626) );
  AND U29575 ( .A(n29634), .B(n29635), .Z(n29633) );
  XNOR U29576 ( .A(n29632), .B(n29636), .Z(n29634) );
  XNOR U29577 ( .A(n29595), .B(n29602), .Z(n29614) );
  AND U29578 ( .A(n29555), .B(n29637), .Z(n29602) );
  XOR U29579 ( .A(n29607), .B(n29606), .Z(n29595) );
  XNOR U29580 ( .A(n29638), .B(n29603), .Z(n29606) );
  XOR U29581 ( .A(n29639), .B(n29640), .Z(n29603) );
  AND U29582 ( .A(n29641), .B(n29642), .Z(n29640) );
  XOR U29583 ( .A(n29639), .B(n29643), .Z(n29641) );
  XNOR U29584 ( .A(n29644), .B(n29645), .Z(n29638) );
  AND U29585 ( .A(n29646), .B(n29647), .Z(n29645) );
  XOR U29586 ( .A(n29644), .B(n29648), .Z(n29646) );
  XOR U29587 ( .A(n29649), .B(n29650), .Z(n29607) );
  AND U29588 ( .A(n29651), .B(n29652), .Z(n29650) );
  XOR U29589 ( .A(n29649), .B(n29653), .Z(n29651) );
  XNOR U29590 ( .A(n29540), .B(n29610), .Z(n29612) );
  XNOR U29591 ( .A(n29654), .B(n29655), .Z(n29540) );
  AND U29592 ( .A(n584), .B(n29547), .Z(n29655) );
  XOR U29593 ( .A(n29654), .B(n29545), .Z(n29547) );
  XOR U29594 ( .A(n29656), .B(n29657), .Z(n29610) );
  AND U29595 ( .A(n29658), .B(n29659), .Z(n29657) );
  XNOR U29596 ( .A(n29656), .B(n29555), .Z(n29659) );
  XOR U29597 ( .A(n29660), .B(n29624), .Z(n29555) );
  XNOR U29598 ( .A(n29661), .B(n29631), .Z(n29624) );
  XOR U29599 ( .A(n29620), .B(n29619), .Z(n29631) );
  XNOR U29600 ( .A(n29662), .B(n29616), .Z(n29619) );
  XOR U29601 ( .A(n29663), .B(n29664), .Z(n29616) );
  AND U29602 ( .A(n29665), .B(n29666), .Z(n29664) );
  XNOR U29603 ( .A(n29667), .B(n29668), .Z(n29665) );
  IV U29604 ( .A(n29663), .Z(n29667) );
  XNOR U29605 ( .A(n29669), .B(n29670), .Z(n29662) );
  NOR U29606 ( .A(n29671), .B(n29672), .Z(n29670) );
  XNOR U29607 ( .A(n29669), .B(n29673), .Z(n29671) );
  XOR U29608 ( .A(n29674), .B(n29675), .Z(n29620) );
  NOR U29609 ( .A(n29676), .B(n29677), .Z(n29675) );
  XNOR U29610 ( .A(n29674), .B(n29678), .Z(n29676) );
  XNOR U29611 ( .A(n29630), .B(n29621), .Z(n29661) );
  XOR U29612 ( .A(n29679), .B(n29680), .Z(n29621) );
  AND U29613 ( .A(n29681), .B(n29682), .Z(n29680) );
  XOR U29614 ( .A(n29679), .B(n29683), .Z(n29681) );
  XOR U29615 ( .A(n29684), .B(n29636), .Z(n29630) );
  XOR U29616 ( .A(n29685), .B(n29686), .Z(n29636) );
  NOR U29617 ( .A(n29687), .B(n29688), .Z(n29686) );
  XOR U29618 ( .A(n29685), .B(n29689), .Z(n29687) );
  XNOR U29619 ( .A(n29635), .B(n29627), .Z(n29684) );
  XOR U29620 ( .A(n29690), .B(n29691), .Z(n29627) );
  AND U29621 ( .A(n29692), .B(n29693), .Z(n29691) );
  XOR U29622 ( .A(n29690), .B(n29694), .Z(n29692) );
  XNOR U29623 ( .A(n29695), .B(n29632), .Z(n29635) );
  XOR U29624 ( .A(n29696), .B(n29697), .Z(n29632) );
  AND U29625 ( .A(n29698), .B(n29699), .Z(n29697) );
  XNOR U29626 ( .A(n29700), .B(n29701), .Z(n29698) );
  IV U29627 ( .A(n29696), .Z(n29700) );
  XNOR U29628 ( .A(n29702), .B(n29703), .Z(n29695) );
  NOR U29629 ( .A(n29704), .B(n29705), .Z(n29703) );
  XNOR U29630 ( .A(n29702), .B(n29706), .Z(n29704) );
  XOR U29631 ( .A(n29625), .B(n29637), .Z(n29660) );
  NOR U29632 ( .A(n29563), .B(n29707), .Z(n29637) );
  XNOR U29633 ( .A(n29643), .B(n29642), .Z(n29625) );
  XNOR U29634 ( .A(n29708), .B(n29648), .Z(n29642) );
  XNOR U29635 ( .A(n29709), .B(n29710), .Z(n29648) );
  NOR U29636 ( .A(n29711), .B(n29712), .Z(n29710) );
  XOR U29637 ( .A(n29709), .B(n29713), .Z(n29711) );
  XNOR U29638 ( .A(n29647), .B(n29639), .Z(n29708) );
  XOR U29639 ( .A(n29714), .B(n29715), .Z(n29639) );
  AND U29640 ( .A(n29716), .B(n29717), .Z(n29715) );
  XOR U29641 ( .A(n29714), .B(n29718), .Z(n29716) );
  XNOR U29642 ( .A(n29719), .B(n29644), .Z(n29647) );
  XOR U29643 ( .A(n29720), .B(n29721), .Z(n29644) );
  AND U29644 ( .A(n29722), .B(n29723), .Z(n29721) );
  XNOR U29645 ( .A(n29724), .B(n29725), .Z(n29722) );
  IV U29646 ( .A(n29720), .Z(n29724) );
  XNOR U29647 ( .A(n29726), .B(n29727), .Z(n29719) );
  NOR U29648 ( .A(n29728), .B(n29729), .Z(n29727) );
  XNOR U29649 ( .A(n29726), .B(n29730), .Z(n29728) );
  XOR U29650 ( .A(n29653), .B(n29652), .Z(n29643) );
  XNOR U29651 ( .A(n29731), .B(n29649), .Z(n29652) );
  XOR U29652 ( .A(n29732), .B(n29733), .Z(n29649) );
  AND U29653 ( .A(n29734), .B(n29735), .Z(n29733) );
  XNOR U29654 ( .A(n29736), .B(n29737), .Z(n29734) );
  IV U29655 ( .A(n29732), .Z(n29736) );
  XNOR U29656 ( .A(n29738), .B(n29739), .Z(n29731) );
  NOR U29657 ( .A(n29740), .B(n29741), .Z(n29739) );
  XNOR U29658 ( .A(n29738), .B(n29742), .Z(n29740) );
  XOR U29659 ( .A(n29743), .B(n29744), .Z(n29653) );
  NOR U29660 ( .A(n29745), .B(n29746), .Z(n29744) );
  XNOR U29661 ( .A(n29743), .B(n29747), .Z(n29745) );
  XNOR U29662 ( .A(n29552), .B(n29656), .Z(n29658) );
  XNOR U29663 ( .A(n29748), .B(n29749), .Z(n29552) );
  AND U29664 ( .A(n584), .B(n29559), .Z(n29749) );
  XOR U29665 ( .A(n29748), .B(n29557), .Z(n29559) );
  AND U29666 ( .A(n29560), .B(n29563), .Z(n29656) );
  XOR U29667 ( .A(n29750), .B(n29707), .Z(n29563) );
  XNOR U29668 ( .A(p_input[1504]), .B(p_input[2048]), .Z(n29707) );
  XNOR U29669 ( .A(n29683), .B(n29682), .Z(n29750) );
  XNOR U29670 ( .A(n29751), .B(n29694), .Z(n29682) );
  XOR U29671 ( .A(n29668), .B(n29666), .Z(n29694) );
  XNOR U29672 ( .A(n29752), .B(n29673), .Z(n29666) );
  XOR U29673 ( .A(p_input[1528]), .B(p_input[2072]), .Z(n29673) );
  XOR U29674 ( .A(n29663), .B(n29672), .Z(n29752) );
  XOR U29675 ( .A(n29753), .B(n29669), .Z(n29672) );
  XOR U29676 ( .A(p_input[1526]), .B(p_input[2070]), .Z(n29669) );
  XOR U29677 ( .A(p_input[1527]), .B(n17295), .Z(n29753) );
  XOR U29678 ( .A(p_input[1522]), .B(p_input[2066]), .Z(n29663) );
  XNOR U29679 ( .A(n29678), .B(n29677), .Z(n29668) );
  XOR U29680 ( .A(n29754), .B(n29674), .Z(n29677) );
  XOR U29681 ( .A(p_input[1523]), .B(p_input[2067]), .Z(n29674) );
  XOR U29682 ( .A(p_input[1524]), .B(n17297), .Z(n29754) );
  XOR U29683 ( .A(p_input[1525]), .B(p_input[2069]), .Z(n29678) );
  XOR U29684 ( .A(n29693), .B(n29755), .Z(n29751) );
  IV U29685 ( .A(n29679), .Z(n29755) );
  XOR U29686 ( .A(p_input[1505]), .B(p_input[2049]), .Z(n29679) );
  XNOR U29687 ( .A(n29756), .B(n29701), .Z(n29693) );
  XNOR U29688 ( .A(n29689), .B(n29688), .Z(n29701) );
  XNOR U29689 ( .A(n29757), .B(n29685), .Z(n29688) );
  XNOR U29690 ( .A(p_input[1530]), .B(p_input[2074]), .Z(n29685) );
  XOR U29691 ( .A(p_input[1531]), .B(n17300), .Z(n29757) );
  XOR U29692 ( .A(p_input[1532]), .B(p_input[2076]), .Z(n29689) );
  XOR U29693 ( .A(n29699), .B(n29758), .Z(n29756) );
  IV U29694 ( .A(n29690), .Z(n29758) );
  XOR U29695 ( .A(p_input[1521]), .B(p_input[2065]), .Z(n29690) );
  XNOR U29696 ( .A(n29759), .B(n29706), .Z(n29699) );
  XNOR U29697 ( .A(p_input[1535]), .B(n17303), .Z(n29706) );
  XOR U29698 ( .A(n29696), .B(n29705), .Z(n29759) );
  XOR U29699 ( .A(n29760), .B(n29702), .Z(n29705) );
  XOR U29700 ( .A(p_input[1533]), .B(p_input[2077]), .Z(n29702) );
  XOR U29701 ( .A(p_input[1534]), .B(n17305), .Z(n29760) );
  XOR U29702 ( .A(p_input[1529]), .B(p_input[2073]), .Z(n29696) );
  XOR U29703 ( .A(n29718), .B(n29717), .Z(n29683) );
  XNOR U29704 ( .A(n29761), .B(n29725), .Z(n29717) );
  XNOR U29705 ( .A(n29713), .B(n29712), .Z(n29725) );
  XNOR U29706 ( .A(n29762), .B(n29709), .Z(n29712) );
  XNOR U29707 ( .A(p_input[1515]), .B(p_input[2059]), .Z(n29709) );
  XOR U29708 ( .A(p_input[1516]), .B(n16451), .Z(n29762) );
  XOR U29709 ( .A(p_input[1517]), .B(p_input[2061]), .Z(n29713) );
  XOR U29710 ( .A(n29723), .B(n29763), .Z(n29761) );
  IV U29711 ( .A(n29714), .Z(n29763) );
  XOR U29712 ( .A(p_input[1506]), .B(p_input[2050]), .Z(n29714) );
  XNOR U29713 ( .A(n29764), .B(n29730), .Z(n29723) );
  XNOR U29714 ( .A(p_input[1520]), .B(n16454), .Z(n29730) );
  XOR U29715 ( .A(n29720), .B(n29729), .Z(n29764) );
  XOR U29716 ( .A(n29765), .B(n29726), .Z(n29729) );
  XOR U29717 ( .A(p_input[1518]), .B(p_input[2062]), .Z(n29726) );
  XOR U29718 ( .A(p_input[1519]), .B(n16456), .Z(n29765) );
  XOR U29719 ( .A(p_input[1514]), .B(p_input[2058]), .Z(n29720) );
  XOR U29720 ( .A(n29737), .B(n29735), .Z(n29718) );
  XNOR U29721 ( .A(n29766), .B(n29742), .Z(n29735) );
  XOR U29722 ( .A(p_input[1513]), .B(p_input[2057]), .Z(n29742) );
  XOR U29723 ( .A(n29732), .B(n29741), .Z(n29766) );
  XOR U29724 ( .A(n29767), .B(n29738), .Z(n29741) );
  XOR U29725 ( .A(p_input[1511]), .B(p_input[2055]), .Z(n29738) );
  XOR U29726 ( .A(p_input[1512]), .B(n17312), .Z(n29767) );
  XOR U29727 ( .A(p_input[1507]), .B(p_input[2051]), .Z(n29732) );
  XNOR U29728 ( .A(n29747), .B(n29746), .Z(n29737) );
  XOR U29729 ( .A(n29768), .B(n29743), .Z(n29746) );
  XOR U29730 ( .A(p_input[1508]), .B(p_input[2052]), .Z(n29743) );
  XOR U29731 ( .A(p_input[1509]), .B(n17314), .Z(n29768) );
  XOR U29732 ( .A(p_input[1510]), .B(p_input[2054]), .Z(n29747) );
  XNOR U29733 ( .A(n29769), .B(n29770), .Z(n29560) );
  AND U29734 ( .A(n584), .B(n29771), .Z(n29770) );
  XNOR U29735 ( .A(n29772), .B(n29773), .Z(n584) );
  AND U29736 ( .A(n29774), .B(n29775), .Z(n29773) );
  XOR U29737 ( .A(n29772), .B(n29570), .Z(n29775) );
  XNOR U29738 ( .A(n29772), .B(n29512), .Z(n29774) );
  XOR U29739 ( .A(n29776), .B(n29777), .Z(n29772) );
  AND U29740 ( .A(n29778), .B(n29779), .Z(n29777) );
  XNOR U29741 ( .A(n29583), .B(n29776), .Z(n29779) );
  XOR U29742 ( .A(n29776), .B(n29524), .Z(n29778) );
  XOR U29743 ( .A(n29780), .B(n29781), .Z(n29776) );
  AND U29744 ( .A(n29782), .B(n29783), .Z(n29781) );
  XNOR U29745 ( .A(n29608), .B(n29780), .Z(n29783) );
  XOR U29746 ( .A(n29780), .B(n29535), .Z(n29782) );
  XOR U29747 ( .A(n29784), .B(n29785), .Z(n29780) );
  AND U29748 ( .A(n29786), .B(n29787), .Z(n29785) );
  XOR U29749 ( .A(n29784), .B(n29545), .Z(n29786) );
  XOR U29750 ( .A(n29788), .B(n29789), .Z(n29501) );
  AND U29751 ( .A(n588), .B(n29771), .Z(n29789) );
  XNOR U29752 ( .A(n29769), .B(n29788), .Z(n29771) );
  XNOR U29753 ( .A(n29790), .B(n29791), .Z(n588) );
  AND U29754 ( .A(n29792), .B(n29793), .Z(n29791) );
  XNOR U29755 ( .A(n29794), .B(n29790), .Z(n29793) );
  IV U29756 ( .A(n29570), .Z(n29794) );
  XNOR U29757 ( .A(n29795), .B(n29796), .Z(n29570) );
  AND U29758 ( .A(n591), .B(n29797), .Z(n29796) );
  XNOR U29759 ( .A(n29795), .B(n29798), .Z(n29797) );
  XNOR U29760 ( .A(n29512), .B(n29790), .Z(n29792) );
  XOR U29761 ( .A(n29799), .B(n29800), .Z(n29512) );
  AND U29762 ( .A(n599), .B(n29801), .Z(n29800) );
  XOR U29763 ( .A(n29802), .B(n29803), .Z(n29790) );
  AND U29764 ( .A(n29804), .B(n29805), .Z(n29803) );
  XNOR U29765 ( .A(n29802), .B(n29583), .Z(n29805) );
  XNOR U29766 ( .A(n29806), .B(n29807), .Z(n29583) );
  AND U29767 ( .A(n591), .B(n29808), .Z(n29807) );
  XOR U29768 ( .A(n29809), .B(n29806), .Z(n29808) );
  XNOR U29769 ( .A(n29810), .B(n29802), .Z(n29804) );
  IV U29770 ( .A(n29524), .Z(n29810) );
  XOR U29771 ( .A(n29811), .B(n29812), .Z(n29524) );
  AND U29772 ( .A(n599), .B(n29813), .Z(n29812) );
  XOR U29773 ( .A(n29814), .B(n29815), .Z(n29802) );
  AND U29774 ( .A(n29816), .B(n29817), .Z(n29815) );
  XNOR U29775 ( .A(n29814), .B(n29608), .Z(n29817) );
  XNOR U29776 ( .A(n29818), .B(n29819), .Z(n29608) );
  AND U29777 ( .A(n591), .B(n29820), .Z(n29819) );
  XNOR U29778 ( .A(n29821), .B(n29818), .Z(n29820) );
  XOR U29779 ( .A(n29535), .B(n29814), .Z(n29816) );
  XOR U29780 ( .A(n29822), .B(n29823), .Z(n29535) );
  AND U29781 ( .A(n599), .B(n29824), .Z(n29823) );
  XOR U29782 ( .A(n29784), .B(n29825), .Z(n29814) );
  AND U29783 ( .A(n29826), .B(n29787), .Z(n29825) );
  XNOR U29784 ( .A(n29654), .B(n29784), .Z(n29787) );
  XNOR U29785 ( .A(n29827), .B(n29828), .Z(n29654) );
  AND U29786 ( .A(n591), .B(n29829), .Z(n29828) );
  XOR U29787 ( .A(n29830), .B(n29827), .Z(n29829) );
  XNOR U29788 ( .A(n29831), .B(n29784), .Z(n29826) );
  IV U29789 ( .A(n29545), .Z(n29831) );
  XOR U29790 ( .A(n29832), .B(n29833), .Z(n29545) );
  AND U29791 ( .A(n599), .B(n29834), .Z(n29833) );
  XOR U29792 ( .A(n29835), .B(n29836), .Z(n29784) );
  AND U29793 ( .A(n29837), .B(n29838), .Z(n29836) );
  XNOR U29794 ( .A(n29835), .B(n29748), .Z(n29838) );
  XNOR U29795 ( .A(n29839), .B(n29840), .Z(n29748) );
  AND U29796 ( .A(n591), .B(n29841), .Z(n29840) );
  XNOR U29797 ( .A(n29842), .B(n29839), .Z(n29841) );
  XNOR U29798 ( .A(n29843), .B(n29835), .Z(n29837) );
  IV U29799 ( .A(n29557), .Z(n29843) );
  XOR U29800 ( .A(n29844), .B(n29845), .Z(n29557) );
  AND U29801 ( .A(n599), .B(n29846), .Z(n29845) );
  AND U29802 ( .A(n29788), .B(n29769), .Z(n29835) );
  XNOR U29803 ( .A(n29847), .B(n29848), .Z(n29769) );
  AND U29804 ( .A(n591), .B(n29849), .Z(n29848) );
  XNOR U29805 ( .A(n29850), .B(n29847), .Z(n29849) );
  XNOR U29806 ( .A(n29851), .B(n29852), .Z(n591) );
  AND U29807 ( .A(n29853), .B(n29854), .Z(n29852) );
  XOR U29808 ( .A(n29798), .B(n29851), .Z(n29854) );
  AND U29809 ( .A(n29855), .B(n29856), .Z(n29798) );
  XOR U29810 ( .A(n29851), .B(n29795), .Z(n29853) );
  XNOR U29811 ( .A(n29857), .B(n29858), .Z(n29795) );
  AND U29812 ( .A(n595), .B(n29801), .Z(n29858) );
  XOR U29813 ( .A(n29799), .B(n29857), .Z(n29801) );
  XOR U29814 ( .A(n29859), .B(n29860), .Z(n29851) );
  AND U29815 ( .A(n29861), .B(n29862), .Z(n29860) );
  XNOR U29816 ( .A(n29859), .B(n29855), .Z(n29862) );
  IV U29817 ( .A(n29809), .Z(n29855) );
  XOR U29818 ( .A(n29863), .B(n29864), .Z(n29809) );
  XOR U29819 ( .A(n29865), .B(n29856), .Z(n29864) );
  AND U29820 ( .A(n29821), .B(n29866), .Z(n29856) );
  AND U29821 ( .A(n29867), .B(n29868), .Z(n29865) );
  XOR U29822 ( .A(n29869), .B(n29863), .Z(n29867) );
  XNOR U29823 ( .A(n29806), .B(n29859), .Z(n29861) );
  XNOR U29824 ( .A(n29870), .B(n29871), .Z(n29806) );
  AND U29825 ( .A(n595), .B(n29813), .Z(n29871) );
  XOR U29826 ( .A(n29870), .B(n29811), .Z(n29813) );
  XOR U29827 ( .A(n29872), .B(n29873), .Z(n29859) );
  AND U29828 ( .A(n29874), .B(n29875), .Z(n29873) );
  XNOR U29829 ( .A(n29872), .B(n29821), .Z(n29875) );
  XOR U29830 ( .A(n29876), .B(n29868), .Z(n29821) );
  XNOR U29831 ( .A(n29877), .B(n29863), .Z(n29868) );
  XOR U29832 ( .A(n29878), .B(n29879), .Z(n29863) );
  AND U29833 ( .A(n29880), .B(n29881), .Z(n29879) );
  XOR U29834 ( .A(n29882), .B(n29878), .Z(n29880) );
  XNOR U29835 ( .A(n29883), .B(n29884), .Z(n29877) );
  AND U29836 ( .A(n29885), .B(n29886), .Z(n29884) );
  XOR U29837 ( .A(n29883), .B(n29887), .Z(n29885) );
  XNOR U29838 ( .A(n29869), .B(n29866), .Z(n29876) );
  AND U29839 ( .A(n29888), .B(n29889), .Z(n29866) );
  XOR U29840 ( .A(n29890), .B(n29891), .Z(n29869) );
  AND U29841 ( .A(n29892), .B(n29893), .Z(n29891) );
  XOR U29842 ( .A(n29890), .B(n29894), .Z(n29892) );
  XNOR U29843 ( .A(n29818), .B(n29872), .Z(n29874) );
  XNOR U29844 ( .A(n29895), .B(n29896), .Z(n29818) );
  AND U29845 ( .A(n595), .B(n29824), .Z(n29896) );
  XOR U29846 ( .A(n29895), .B(n29822), .Z(n29824) );
  XOR U29847 ( .A(n29897), .B(n29898), .Z(n29872) );
  AND U29848 ( .A(n29899), .B(n29900), .Z(n29898) );
  XNOR U29849 ( .A(n29897), .B(n29888), .Z(n29900) );
  IV U29850 ( .A(n29830), .Z(n29888) );
  XNOR U29851 ( .A(n29901), .B(n29881), .Z(n29830) );
  XNOR U29852 ( .A(n29902), .B(n29887), .Z(n29881) );
  XOR U29853 ( .A(n29903), .B(n29904), .Z(n29887) );
  AND U29854 ( .A(n29905), .B(n29906), .Z(n29904) );
  XOR U29855 ( .A(n29903), .B(n29907), .Z(n29905) );
  XNOR U29856 ( .A(n29886), .B(n29878), .Z(n29902) );
  XOR U29857 ( .A(n29908), .B(n29909), .Z(n29878) );
  AND U29858 ( .A(n29910), .B(n29911), .Z(n29909) );
  XNOR U29859 ( .A(n29912), .B(n29908), .Z(n29910) );
  XNOR U29860 ( .A(n29913), .B(n29883), .Z(n29886) );
  XOR U29861 ( .A(n29914), .B(n29915), .Z(n29883) );
  AND U29862 ( .A(n29916), .B(n29917), .Z(n29915) );
  XOR U29863 ( .A(n29914), .B(n29918), .Z(n29916) );
  XNOR U29864 ( .A(n29919), .B(n29920), .Z(n29913) );
  AND U29865 ( .A(n29921), .B(n29922), .Z(n29920) );
  XNOR U29866 ( .A(n29919), .B(n29923), .Z(n29921) );
  XNOR U29867 ( .A(n29882), .B(n29889), .Z(n29901) );
  AND U29868 ( .A(n29842), .B(n29924), .Z(n29889) );
  XOR U29869 ( .A(n29894), .B(n29893), .Z(n29882) );
  XNOR U29870 ( .A(n29925), .B(n29890), .Z(n29893) );
  XOR U29871 ( .A(n29926), .B(n29927), .Z(n29890) );
  AND U29872 ( .A(n29928), .B(n29929), .Z(n29927) );
  XOR U29873 ( .A(n29926), .B(n29930), .Z(n29928) );
  XNOR U29874 ( .A(n29931), .B(n29932), .Z(n29925) );
  AND U29875 ( .A(n29933), .B(n29934), .Z(n29932) );
  XOR U29876 ( .A(n29931), .B(n29935), .Z(n29933) );
  XOR U29877 ( .A(n29936), .B(n29937), .Z(n29894) );
  AND U29878 ( .A(n29938), .B(n29939), .Z(n29937) );
  XOR U29879 ( .A(n29936), .B(n29940), .Z(n29938) );
  XNOR U29880 ( .A(n29827), .B(n29897), .Z(n29899) );
  XNOR U29881 ( .A(n29941), .B(n29942), .Z(n29827) );
  AND U29882 ( .A(n595), .B(n29834), .Z(n29942) );
  XOR U29883 ( .A(n29941), .B(n29832), .Z(n29834) );
  XOR U29884 ( .A(n29943), .B(n29944), .Z(n29897) );
  AND U29885 ( .A(n29945), .B(n29946), .Z(n29944) );
  XNOR U29886 ( .A(n29943), .B(n29842), .Z(n29946) );
  XOR U29887 ( .A(n29947), .B(n29911), .Z(n29842) );
  XNOR U29888 ( .A(n29948), .B(n29918), .Z(n29911) );
  XOR U29889 ( .A(n29907), .B(n29906), .Z(n29918) );
  XNOR U29890 ( .A(n29949), .B(n29903), .Z(n29906) );
  XOR U29891 ( .A(n29950), .B(n29951), .Z(n29903) );
  AND U29892 ( .A(n29952), .B(n29953), .Z(n29951) );
  XNOR U29893 ( .A(n29954), .B(n29955), .Z(n29952) );
  IV U29894 ( .A(n29950), .Z(n29954) );
  XNOR U29895 ( .A(n29956), .B(n29957), .Z(n29949) );
  NOR U29896 ( .A(n29958), .B(n29959), .Z(n29957) );
  XNOR U29897 ( .A(n29956), .B(n29960), .Z(n29958) );
  XOR U29898 ( .A(n29961), .B(n29962), .Z(n29907) );
  NOR U29899 ( .A(n29963), .B(n29964), .Z(n29962) );
  XNOR U29900 ( .A(n29961), .B(n29965), .Z(n29963) );
  XNOR U29901 ( .A(n29917), .B(n29908), .Z(n29948) );
  XOR U29902 ( .A(n29966), .B(n29967), .Z(n29908) );
  AND U29903 ( .A(n29968), .B(n29969), .Z(n29967) );
  XOR U29904 ( .A(n29966), .B(n29970), .Z(n29968) );
  XOR U29905 ( .A(n29971), .B(n29923), .Z(n29917) );
  XOR U29906 ( .A(n29972), .B(n29973), .Z(n29923) );
  NOR U29907 ( .A(n29974), .B(n29975), .Z(n29973) );
  XOR U29908 ( .A(n29972), .B(n29976), .Z(n29974) );
  XNOR U29909 ( .A(n29922), .B(n29914), .Z(n29971) );
  XOR U29910 ( .A(n29977), .B(n29978), .Z(n29914) );
  AND U29911 ( .A(n29979), .B(n29980), .Z(n29978) );
  XOR U29912 ( .A(n29977), .B(n29981), .Z(n29979) );
  XNOR U29913 ( .A(n29982), .B(n29919), .Z(n29922) );
  XOR U29914 ( .A(n29983), .B(n29984), .Z(n29919) );
  AND U29915 ( .A(n29985), .B(n29986), .Z(n29984) );
  XNOR U29916 ( .A(n29987), .B(n29988), .Z(n29985) );
  IV U29917 ( .A(n29983), .Z(n29987) );
  XNOR U29918 ( .A(n29989), .B(n29990), .Z(n29982) );
  NOR U29919 ( .A(n29991), .B(n29992), .Z(n29990) );
  XNOR U29920 ( .A(n29989), .B(n29993), .Z(n29991) );
  XOR U29921 ( .A(n29912), .B(n29924), .Z(n29947) );
  NOR U29922 ( .A(n29850), .B(n29994), .Z(n29924) );
  XNOR U29923 ( .A(n29930), .B(n29929), .Z(n29912) );
  XNOR U29924 ( .A(n29995), .B(n29935), .Z(n29929) );
  XNOR U29925 ( .A(n29996), .B(n29997), .Z(n29935) );
  NOR U29926 ( .A(n29998), .B(n29999), .Z(n29997) );
  XOR U29927 ( .A(n29996), .B(n30000), .Z(n29998) );
  XNOR U29928 ( .A(n29934), .B(n29926), .Z(n29995) );
  XOR U29929 ( .A(n30001), .B(n30002), .Z(n29926) );
  AND U29930 ( .A(n30003), .B(n30004), .Z(n30002) );
  XOR U29931 ( .A(n30001), .B(n30005), .Z(n30003) );
  XNOR U29932 ( .A(n30006), .B(n29931), .Z(n29934) );
  XOR U29933 ( .A(n30007), .B(n30008), .Z(n29931) );
  AND U29934 ( .A(n30009), .B(n30010), .Z(n30008) );
  XNOR U29935 ( .A(n30011), .B(n30012), .Z(n30009) );
  IV U29936 ( .A(n30007), .Z(n30011) );
  XNOR U29937 ( .A(n30013), .B(n30014), .Z(n30006) );
  NOR U29938 ( .A(n30015), .B(n30016), .Z(n30014) );
  XNOR U29939 ( .A(n30013), .B(n30017), .Z(n30015) );
  XOR U29940 ( .A(n29940), .B(n29939), .Z(n29930) );
  XNOR U29941 ( .A(n30018), .B(n29936), .Z(n29939) );
  XOR U29942 ( .A(n30019), .B(n30020), .Z(n29936) );
  AND U29943 ( .A(n30021), .B(n30022), .Z(n30020) );
  XNOR U29944 ( .A(n30023), .B(n30024), .Z(n30021) );
  IV U29945 ( .A(n30019), .Z(n30023) );
  XNOR U29946 ( .A(n30025), .B(n30026), .Z(n30018) );
  NOR U29947 ( .A(n30027), .B(n30028), .Z(n30026) );
  XNOR U29948 ( .A(n30025), .B(n30029), .Z(n30027) );
  XOR U29949 ( .A(n30030), .B(n30031), .Z(n29940) );
  NOR U29950 ( .A(n30032), .B(n30033), .Z(n30031) );
  XNOR U29951 ( .A(n30030), .B(n30034), .Z(n30032) );
  XNOR U29952 ( .A(n29839), .B(n29943), .Z(n29945) );
  XNOR U29953 ( .A(n30035), .B(n30036), .Z(n29839) );
  AND U29954 ( .A(n595), .B(n29846), .Z(n30036) );
  XOR U29955 ( .A(n30035), .B(n29844), .Z(n29846) );
  AND U29956 ( .A(n29847), .B(n29850), .Z(n29943) );
  XOR U29957 ( .A(n30037), .B(n29994), .Z(n29850) );
  XNOR U29958 ( .A(p_input[1536]), .B(p_input[2048]), .Z(n29994) );
  XNOR U29959 ( .A(n29970), .B(n29969), .Z(n30037) );
  XNOR U29960 ( .A(n30038), .B(n29981), .Z(n29969) );
  XOR U29961 ( .A(n29955), .B(n29953), .Z(n29981) );
  XNOR U29962 ( .A(n30039), .B(n29960), .Z(n29953) );
  XOR U29963 ( .A(p_input[1560]), .B(p_input[2072]), .Z(n29960) );
  XOR U29964 ( .A(n29950), .B(n29959), .Z(n30039) );
  XOR U29965 ( .A(n30040), .B(n29956), .Z(n29959) );
  XOR U29966 ( .A(p_input[1558]), .B(p_input[2070]), .Z(n29956) );
  XOR U29967 ( .A(p_input[1559]), .B(n17295), .Z(n30040) );
  XOR U29968 ( .A(p_input[1554]), .B(p_input[2066]), .Z(n29950) );
  XNOR U29969 ( .A(n29965), .B(n29964), .Z(n29955) );
  XOR U29970 ( .A(n30041), .B(n29961), .Z(n29964) );
  XOR U29971 ( .A(p_input[1555]), .B(p_input[2067]), .Z(n29961) );
  XOR U29972 ( .A(p_input[1556]), .B(n17297), .Z(n30041) );
  XOR U29973 ( .A(p_input[1557]), .B(p_input[2069]), .Z(n29965) );
  XOR U29974 ( .A(n29980), .B(n30042), .Z(n30038) );
  IV U29975 ( .A(n29966), .Z(n30042) );
  XOR U29976 ( .A(p_input[1537]), .B(p_input[2049]), .Z(n29966) );
  XNOR U29977 ( .A(n30043), .B(n29988), .Z(n29980) );
  XNOR U29978 ( .A(n29976), .B(n29975), .Z(n29988) );
  XNOR U29979 ( .A(n30044), .B(n29972), .Z(n29975) );
  XNOR U29980 ( .A(p_input[1562]), .B(p_input[2074]), .Z(n29972) );
  XOR U29981 ( .A(p_input[1563]), .B(n17300), .Z(n30044) );
  XOR U29982 ( .A(p_input[1564]), .B(p_input[2076]), .Z(n29976) );
  XOR U29983 ( .A(n29986), .B(n30045), .Z(n30043) );
  IV U29984 ( .A(n29977), .Z(n30045) );
  XOR U29985 ( .A(p_input[1553]), .B(p_input[2065]), .Z(n29977) );
  XNOR U29986 ( .A(n30046), .B(n29993), .Z(n29986) );
  XNOR U29987 ( .A(p_input[1567]), .B(n17303), .Z(n29993) );
  XOR U29988 ( .A(n29983), .B(n29992), .Z(n30046) );
  XOR U29989 ( .A(n30047), .B(n29989), .Z(n29992) );
  XOR U29990 ( .A(p_input[1565]), .B(p_input[2077]), .Z(n29989) );
  XOR U29991 ( .A(p_input[1566]), .B(n17305), .Z(n30047) );
  XOR U29992 ( .A(p_input[1561]), .B(p_input[2073]), .Z(n29983) );
  XOR U29993 ( .A(n30005), .B(n30004), .Z(n29970) );
  XNOR U29994 ( .A(n30048), .B(n30012), .Z(n30004) );
  XNOR U29995 ( .A(n30000), .B(n29999), .Z(n30012) );
  XNOR U29996 ( .A(n30049), .B(n29996), .Z(n29999) );
  XNOR U29997 ( .A(p_input[1547]), .B(p_input[2059]), .Z(n29996) );
  XOR U29998 ( .A(p_input[1548]), .B(n16451), .Z(n30049) );
  XOR U29999 ( .A(p_input[1549]), .B(p_input[2061]), .Z(n30000) );
  XOR U30000 ( .A(n30010), .B(n30050), .Z(n30048) );
  IV U30001 ( .A(n30001), .Z(n30050) );
  XOR U30002 ( .A(p_input[1538]), .B(p_input[2050]), .Z(n30001) );
  XNOR U30003 ( .A(n30051), .B(n30017), .Z(n30010) );
  XNOR U30004 ( .A(p_input[1552]), .B(n16454), .Z(n30017) );
  XOR U30005 ( .A(n30007), .B(n30016), .Z(n30051) );
  XOR U30006 ( .A(n30052), .B(n30013), .Z(n30016) );
  XOR U30007 ( .A(p_input[1550]), .B(p_input[2062]), .Z(n30013) );
  XOR U30008 ( .A(p_input[1551]), .B(n16456), .Z(n30052) );
  XOR U30009 ( .A(p_input[1546]), .B(p_input[2058]), .Z(n30007) );
  XOR U30010 ( .A(n30024), .B(n30022), .Z(n30005) );
  XNOR U30011 ( .A(n30053), .B(n30029), .Z(n30022) );
  XOR U30012 ( .A(p_input[1545]), .B(p_input[2057]), .Z(n30029) );
  XOR U30013 ( .A(n30019), .B(n30028), .Z(n30053) );
  XOR U30014 ( .A(n30054), .B(n30025), .Z(n30028) );
  XOR U30015 ( .A(p_input[1543]), .B(p_input[2055]), .Z(n30025) );
  XOR U30016 ( .A(p_input[1544]), .B(n17312), .Z(n30054) );
  XOR U30017 ( .A(p_input[1539]), .B(p_input[2051]), .Z(n30019) );
  XNOR U30018 ( .A(n30034), .B(n30033), .Z(n30024) );
  XOR U30019 ( .A(n30055), .B(n30030), .Z(n30033) );
  XOR U30020 ( .A(p_input[1540]), .B(p_input[2052]), .Z(n30030) );
  XOR U30021 ( .A(p_input[1541]), .B(n17314), .Z(n30055) );
  XOR U30022 ( .A(p_input[1542]), .B(p_input[2054]), .Z(n30034) );
  XNOR U30023 ( .A(n30056), .B(n30057), .Z(n29847) );
  AND U30024 ( .A(n595), .B(n30058), .Z(n30057) );
  XNOR U30025 ( .A(n30059), .B(n30060), .Z(n595) );
  AND U30026 ( .A(n30061), .B(n30062), .Z(n30060) );
  XOR U30027 ( .A(n30059), .B(n29857), .Z(n30062) );
  XNOR U30028 ( .A(n30059), .B(n29799), .Z(n30061) );
  XOR U30029 ( .A(n30063), .B(n30064), .Z(n30059) );
  AND U30030 ( .A(n30065), .B(n30066), .Z(n30064) );
  XNOR U30031 ( .A(n29870), .B(n30063), .Z(n30066) );
  XOR U30032 ( .A(n30063), .B(n29811), .Z(n30065) );
  XOR U30033 ( .A(n30067), .B(n30068), .Z(n30063) );
  AND U30034 ( .A(n30069), .B(n30070), .Z(n30068) );
  XNOR U30035 ( .A(n29895), .B(n30067), .Z(n30070) );
  XOR U30036 ( .A(n30067), .B(n29822), .Z(n30069) );
  XOR U30037 ( .A(n30071), .B(n30072), .Z(n30067) );
  AND U30038 ( .A(n30073), .B(n30074), .Z(n30072) );
  XOR U30039 ( .A(n30071), .B(n29832), .Z(n30073) );
  XOR U30040 ( .A(n30075), .B(n30076), .Z(n29788) );
  AND U30041 ( .A(n599), .B(n30058), .Z(n30076) );
  XNOR U30042 ( .A(n30056), .B(n30075), .Z(n30058) );
  XNOR U30043 ( .A(n30077), .B(n30078), .Z(n599) );
  AND U30044 ( .A(n30079), .B(n30080), .Z(n30078) );
  XNOR U30045 ( .A(n30081), .B(n30077), .Z(n30080) );
  IV U30046 ( .A(n29857), .Z(n30081) );
  XNOR U30047 ( .A(n30082), .B(n30083), .Z(n29857) );
  AND U30048 ( .A(n602), .B(n30084), .Z(n30083) );
  XNOR U30049 ( .A(n30082), .B(n30085), .Z(n30084) );
  XNOR U30050 ( .A(n29799), .B(n30077), .Z(n30079) );
  XOR U30051 ( .A(n30086), .B(n30087), .Z(n29799) );
  AND U30052 ( .A(n610), .B(n30088), .Z(n30087) );
  XOR U30053 ( .A(n30089), .B(n30090), .Z(n30077) );
  AND U30054 ( .A(n30091), .B(n30092), .Z(n30090) );
  XNOR U30055 ( .A(n30089), .B(n29870), .Z(n30092) );
  XNOR U30056 ( .A(n30093), .B(n30094), .Z(n29870) );
  AND U30057 ( .A(n602), .B(n30095), .Z(n30094) );
  XOR U30058 ( .A(n30096), .B(n30093), .Z(n30095) );
  XNOR U30059 ( .A(n30097), .B(n30089), .Z(n30091) );
  IV U30060 ( .A(n29811), .Z(n30097) );
  XOR U30061 ( .A(n30098), .B(n30099), .Z(n29811) );
  AND U30062 ( .A(n610), .B(n30100), .Z(n30099) );
  XOR U30063 ( .A(n30101), .B(n30102), .Z(n30089) );
  AND U30064 ( .A(n30103), .B(n30104), .Z(n30102) );
  XNOR U30065 ( .A(n30101), .B(n29895), .Z(n30104) );
  XNOR U30066 ( .A(n30105), .B(n30106), .Z(n29895) );
  AND U30067 ( .A(n602), .B(n30107), .Z(n30106) );
  XNOR U30068 ( .A(n30108), .B(n30105), .Z(n30107) );
  XOR U30069 ( .A(n29822), .B(n30101), .Z(n30103) );
  XOR U30070 ( .A(n30109), .B(n30110), .Z(n29822) );
  AND U30071 ( .A(n610), .B(n30111), .Z(n30110) );
  XOR U30072 ( .A(n30071), .B(n30112), .Z(n30101) );
  AND U30073 ( .A(n30113), .B(n30074), .Z(n30112) );
  XNOR U30074 ( .A(n29941), .B(n30071), .Z(n30074) );
  XNOR U30075 ( .A(n30114), .B(n30115), .Z(n29941) );
  AND U30076 ( .A(n602), .B(n30116), .Z(n30115) );
  XOR U30077 ( .A(n30117), .B(n30114), .Z(n30116) );
  XNOR U30078 ( .A(n30118), .B(n30071), .Z(n30113) );
  IV U30079 ( .A(n29832), .Z(n30118) );
  XOR U30080 ( .A(n30119), .B(n30120), .Z(n29832) );
  AND U30081 ( .A(n610), .B(n30121), .Z(n30120) );
  XOR U30082 ( .A(n30122), .B(n30123), .Z(n30071) );
  AND U30083 ( .A(n30124), .B(n30125), .Z(n30123) );
  XNOR U30084 ( .A(n30122), .B(n30035), .Z(n30125) );
  XNOR U30085 ( .A(n30126), .B(n30127), .Z(n30035) );
  AND U30086 ( .A(n602), .B(n30128), .Z(n30127) );
  XNOR U30087 ( .A(n30129), .B(n30126), .Z(n30128) );
  XNOR U30088 ( .A(n30130), .B(n30122), .Z(n30124) );
  IV U30089 ( .A(n29844), .Z(n30130) );
  XOR U30090 ( .A(n30131), .B(n30132), .Z(n29844) );
  AND U30091 ( .A(n610), .B(n30133), .Z(n30132) );
  AND U30092 ( .A(n30075), .B(n30056), .Z(n30122) );
  XNOR U30093 ( .A(n30134), .B(n30135), .Z(n30056) );
  AND U30094 ( .A(n602), .B(n30136), .Z(n30135) );
  XNOR U30095 ( .A(n30137), .B(n30134), .Z(n30136) );
  XNOR U30096 ( .A(n30138), .B(n30139), .Z(n602) );
  AND U30097 ( .A(n30140), .B(n30141), .Z(n30139) );
  XOR U30098 ( .A(n30085), .B(n30138), .Z(n30141) );
  AND U30099 ( .A(n30142), .B(n30143), .Z(n30085) );
  XOR U30100 ( .A(n30138), .B(n30082), .Z(n30140) );
  XNOR U30101 ( .A(n30144), .B(n30145), .Z(n30082) );
  AND U30102 ( .A(n606), .B(n30088), .Z(n30145) );
  XOR U30103 ( .A(n30086), .B(n30144), .Z(n30088) );
  XOR U30104 ( .A(n30146), .B(n30147), .Z(n30138) );
  AND U30105 ( .A(n30148), .B(n30149), .Z(n30147) );
  XNOR U30106 ( .A(n30146), .B(n30142), .Z(n30149) );
  IV U30107 ( .A(n30096), .Z(n30142) );
  XOR U30108 ( .A(n30150), .B(n30151), .Z(n30096) );
  XOR U30109 ( .A(n30152), .B(n30143), .Z(n30151) );
  AND U30110 ( .A(n30108), .B(n30153), .Z(n30143) );
  AND U30111 ( .A(n30154), .B(n30155), .Z(n30152) );
  XOR U30112 ( .A(n30156), .B(n30150), .Z(n30154) );
  XNOR U30113 ( .A(n30093), .B(n30146), .Z(n30148) );
  XNOR U30114 ( .A(n30157), .B(n30158), .Z(n30093) );
  AND U30115 ( .A(n606), .B(n30100), .Z(n30158) );
  XOR U30116 ( .A(n30157), .B(n30098), .Z(n30100) );
  XOR U30117 ( .A(n30159), .B(n30160), .Z(n30146) );
  AND U30118 ( .A(n30161), .B(n30162), .Z(n30160) );
  XNOR U30119 ( .A(n30159), .B(n30108), .Z(n30162) );
  XOR U30120 ( .A(n30163), .B(n30155), .Z(n30108) );
  XNOR U30121 ( .A(n30164), .B(n30150), .Z(n30155) );
  XOR U30122 ( .A(n30165), .B(n30166), .Z(n30150) );
  AND U30123 ( .A(n30167), .B(n30168), .Z(n30166) );
  XOR U30124 ( .A(n30169), .B(n30165), .Z(n30167) );
  XNOR U30125 ( .A(n30170), .B(n30171), .Z(n30164) );
  AND U30126 ( .A(n30172), .B(n30173), .Z(n30171) );
  XOR U30127 ( .A(n30170), .B(n30174), .Z(n30172) );
  XNOR U30128 ( .A(n30156), .B(n30153), .Z(n30163) );
  AND U30129 ( .A(n30175), .B(n30176), .Z(n30153) );
  XOR U30130 ( .A(n30177), .B(n30178), .Z(n30156) );
  AND U30131 ( .A(n30179), .B(n30180), .Z(n30178) );
  XOR U30132 ( .A(n30177), .B(n30181), .Z(n30179) );
  XNOR U30133 ( .A(n30105), .B(n30159), .Z(n30161) );
  XNOR U30134 ( .A(n30182), .B(n30183), .Z(n30105) );
  AND U30135 ( .A(n606), .B(n30111), .Z(n30183) );
  XOR U30136 ( .A(n30182), .B(n30109), .Z(n30111) );
  XOR U30137 ( .A(n30184), .B(n30185), .Z(n30159) );
  AND U30138 ( .A(n30186), .B(n30187), .Z(n30185) );
  XNOR U30139 ( .A(n30184), .B(n30175), .Z(n30187) );
  IV U30140 ( .A(n30117), .Z(n30175) );
  XNOR U30141 ( .A(n30188), .B(n30168), .Z(n30117) );
  XNOR U30142 ( .A(n30189), .B(n30174), .Z(n30168) );
  XOR U30143 ( .A(n30190), .B(n30191), .Z(n30174) );
  AND U30144 ( .A(n30192), .B(n30193), .Z(n30191) );
  XOR U30145 ( .A(n30190), .B(n30194), .Z(n30192) );
  XNOR U30146 ( .A(n30173), .B(n30165), .Z(n30189) );
  XOR U30147 ( .A(n30195), .B(n30196), .Z(n30165) );
  AND U30148 ( .A(n30197), .B(n30198), .Z(n30196) );
  XNOR U30149 ( .A(n30199), .B(n30195), .Z(n30197) );
  XNOR U30150 ( .A(n30200), .B(n30170), .Z(n30173) );
  XOR U30151 ( .A(n30201), .B(n30202), .Z(n30170) );
  AND U30152 ( .A(n30203), .B(n30204), .Z(n30202) );
  XOR U30153 ( .A(n30201), .B(n30205), .Z(n30203) );
  XNOR U30154 ( .A(n30206), .B(n30207), .Z(n30200) );
  AND U30155 ( .A(n30208), .B(n30209), .Z(n30207) );
  XNOR U30156 ( .A(n30206), .B(n30210), .Z(n30208) );
  XNOR U30157 ( .A(n30169), .B(n30176), .Z(n30188) );
  AND U30158 ( .A(n30129), .B(n30211), .Z(n30176) );
  XOR U30159 ( .A(n30181), .B(n30180), .Z(n30169) );
  XNOR U30160 ( .A(n30212), .B(n30177), .Z(n30180) );
  XOR U30161 ( .A(n30213), .B(n30214), .Z(n30177) );
  AND U30162 ( .A(n30215), .B(n30216), .Z(n30214) );
  XOR U30163 ( .A(n30213), .B(n30217), .Z(n30215) );
  XNOR U30164 ( .A(n30218), .B(n30219), .Z(n30212) );
  AND U30165 ( .A(n30220), .B(n30221), .Z(n30219) );
  XOR U30166 ( .A(n30218), .B(n30222), .Z(n30220) );
  XOR U30167 ( .A(n30223), .B(n30224), .Z(n30181) );
  AND U30168 ( .A(n30225), .B(n30226), .Z(n30224) );
  XOR U30169 ( .A(n30223), .B(n30227), .Z(n30225) );
  XNOR U30170 ( .A(n30114), .B(n30184), .Z(n30186) );
  XNOR U30171 ( .A(n30228), .B(n30229), .Z(n30114) );
  AND U30172 ( .A(n606), .B(n30121), .Z(n30229) );
  XOR U30173 ( .A(n30228), .B(n30119), .Z(n30121) );
  XOR U30174 ( .A(n30230), .B(n30231), .Z(n30184) );
  AND U30175 ( .A(n30232), .B(n30233), .Z(n30231) );
  XNOR U30176 ( .A(n30230), .B(n30129), .Z(n30233) );
  XOR U30177 ( .A(n30234), .B(n30198), .Z(n30129) );
  XNOR U30178 ( .A(n30235), .B(n30205), .Z(n30198) );
  XOR U30179 ( .A(n30194), .B(n30193), .Z(n30205) );
  XNOR U30180 ( .A(n30236), .B(n30190), .Z(n30193) );
  XOR U30181 ( .A(n30237), .B(n30238), .Z(n30190) );
  AND U30182 ( .A(n30239), .B(n30240), .Z(n30238) );
  XNOR U30183 ( .A(n30241), .B(n30242), .Z(n30239) );
  IV U30184 ( .A(n30237), .Z(n30241) );
  XNOR U30185 ( .A(n30243), .B(n30244), .Z(n30236) );
  NOR U30186 ( .A(n30245), .B(n30246), .Z(n30244) );
  XNOR U30187 ( .A(n30243), .B(n30247), .Z(n30245) );
  XOR U30188 ( .A(n30248), .B(n30249), .Z(n30194) );
  NOR U30189 ( .A(n30250), .B(n30251), .Z(n30249) );
  XNOR U30190 ( .A(n30248), .B(n30252), .Z(n30250) );
  XNOR U30191 ( .A(n30204), .B(n30195), .Z(n30235) );
  XOR U30192 ( .A(n30253), .B(n30254), .Z(n30195) );
  AND U30193 ( .A(n30255), .B(n30256), .Z(n30254) );
  XOR U30194 ( .A(n30253), .B(n30257), .Z(n30255) );
  XOR U30195 ( .A(n30258), .B(n30210), .Z(n30204) );
  XOR U30196 ( .A(n30259), .B(n30260), .Z(n30210) );
  NOR U30197 ( .A(n30261), .B(n30262), .Z(n30260) );
  XOR U30198 ( .A(n30259), .B(n30263), .Z(n30261) );
  XNOR U30199 ( .A(n30209), .B(n30201), .Z(n30258) );
  XOR U30200 ( .A(n30264), .B(n30265), .Z(n30201) );
  AND U30201 ( .A(n30266), .B(n30267), .Z(n30265) );
  XOR U30202 ( .A(n30264), .B(n30268), .Z(n30266) );
  XNOR U30203 ( .A(n30269), .B(n30206), .Z(n30209) );
  XOR U30204 ( .A(n30270), .B(n30271), .Z(n30206) );
  AND U30205 ( .A(n30272), .B(n30273), .Z(n30271) );
  XNOR U30206 ( .A(n30274), .B(n30275), .Z(n30272) );
  IV U30207 ( .A(n30270), .Z(n30274) );
  XNOR U30208 ( .A(n30276), .B(n30277), .Z(n30269) );
  NOR U30209 ( .A(n30278), .B(n30279), .Z(n30277) );
  XNOR U30210 ( .A(n30276), .B(n30280), .Z(n30278) );
  XOR U30211 ( .A(n30199), .B(n30211), .Z(n30234) );
  NOR U30212 ( .A(n30137), .B(n30281), .Z(n30211) );
  XNOR U30213 ( .A(n30217), .B(n30216), .Z(n30199) );
  XNOR U30214 ( .A(n30282), .B(n30222), .Z(n30216) );
  XNOR U30215 ( .A(n30283), .B(n30284), .Z(n30222) );
  NOR U30216 ( .A(n30285), .B(n30286), .Z(n30284) );
  XOR U30217 ( .A(n30283), .B(n30287), .Z(n30285) );
  XNOR U30218 ( .A(n30221), .B(n30213), .Z(n30282) );
  XOR U30219 ( .A(n30288), .B(n30289), .Z(n30213) );
  AND U30220 ( .A(n30290), .B(n30291), .Z(n30289) );
  XOR U30221 ( .A(n30288), .B(n30292), .Z(n30290) );
  XNOR U30222 ( .A(n30293), .B(n30218), .Z(n30221) );
  XOR U30223 ( .A(n30294), .B(n30295), .Z(n30218) );
  AND U30224 ( .A(n30296), .B(n30297), .Z(n30295) );
  XNOR U30225 ( .A(n30298), .B(n30299), .Z(n30296) );
  IV U30226 ( .A(n30294), .Z(n30298) );
  XNOR U30227 ( .A(n30300), .B(n30301), .Z(n30293) );
  NOR U30228 ( .A(n30302), .B(n30303), .Z(n30301) );
  XNOR U30229 ( .A(n30300), .B(n30304), .Z(n30302) );
  XOR U30230 ( .A(n30227), .B(n30226), .Z(n30217) );
  XNOR U30231 ( .A(n30305), .B(n30223), .Z(n30226) );
  XOR U30232 ( .A(n30306), .B(n30307), .Z(n30223) );
  AND U30233 ( .A(n30308), .B(n30309), .Z(n30307) );
  XNOR U30234 ( .A(n30310), .B(n30311), .Z(n30308) );
  IV U30235 ( .A(n30306), .Z(n30310) );
  XNOR U30236 ( .A(n30312), .B(n30313), .Z(n30305) );
  NOR U30237 ( .A(n30314), .B(n30315), .Z(n30313) );
  XNOR U30238 ( .A(n30312), .B(n30316), .Z(n30314) );
  XOR U30239 ( .A(n30317), .B(n30318), .Z(n30227) );
  NOR U30240 ( .A(n30319), .B(n30320), .Z(n30318) );
  XNOR U30241 ( .A(n30317), .B(n30321), .Z(n30319) );
  XNOR U30242 ( .A(n30126), .B(n30230), .Z(n30232) );
  XNOR U30243 ( .A(n30322), .B(n30323), .Z(n30126) );
  AND U30244 ( .A(n606), .B(n30133), .Z(n30323) );
  XOR U30245 ( .A(n30322), .B(n30131), .Z(n30133) );
  AND U30246 ( .A(n30134), .B(n30137), .Z(n30230) );
  XOR U30247 ( .A(n30324), .B(n30281), .Z(n30137) );
  XNOR U30248 ( .A(p_input[1568]), .B(p_input[2048]), .Z(n30281) );
  XNOR U30249 ( .A(n30257), .B(n30256), .Z(n30324) );
  XNOR U30250 ( .A(n30325), .B(n30268), .Z(n30256) );
  XOR U30251 ( .A(n30242), .B(n30240), .Z(n30268) );
  XNOR U30252 ( .A(n30326), .B(n30247), .Z(n30240) );
  XOR U30253 ( .A(p_input[1592]), .B(p_input[2072]), .Z(n30247) );
  XOR U30254 ( .A(n30237), .B(n30246), .Z(n30326) );
  XOR U30255 ( .A(n30327), .B(n30243), .Z(n30246) );
  XOR U30256 ( .A(p_input[1590]), .B(p_input[2070]), .Z(n30243) );
  XOR U30257 ( .A(p_input[1591]), .B(n17295), .Z(n30327) );
  XOR U30258 ( .A(p_input[1586]), .B(p_input[2066]), .Z(n30237) );
  XNOR U30259 ( .A(n30252), .B(n30251), .Z(n30242) );
  XOR U30260 ( .A(n30328), .B(n30248), .Z(n30251) );
  XOR U30261 ( .A(p_input[1587]), .B(p_input[2067]), .Z(n30248) );
  XOR U30262 ( .A(p_input[1588]), .B(n17297), .Z(n30328) );
  XOR U30263 ( .A(p_input[1589]), .B(p_input[2069]), .Z(n30252) );
  XOR U30264 ( .A(n30267), .B(n30329), .Z(n30325) );
  IV U30265 ( .A(n30253), .Z(n30329) );
  XOR U30266 ( .A(p_input[1569]), .B(p_input[2049]), .Z(n30253) );
  XNOR U30267 ( .A(n30330), .B(n30275), .Z(n30267) );
  XNOR U30268 ( .A(n30263), .B(n30262), .Z(n30275) );
  XNOR U30269 ( .A(n30331), .B(n30259), .Z(n30262) );
  XNOR U30270 ( .A(p_input[1594]), .B(p_input[2074]), .Z(n30259) );
  XOR U30271 ( .A(p_input[1595]), .B(n17300), .Z(n30331) );
  XOR U30272 ( .A(p_input[1596]), .B(p_input[2076]), .Z(n30263) );
  XOR U30273 ( .A(n30273), .B(n30332), .Z(n30330) );
  IV U30274 ( .A(n30264), .Z(n30332) );
  XOR U30275 ( .A(p_input[1585]), .B(p_input[2065]), .Z(n30264) );
  XNOR U30276 ( .A(n30333), .B(n30280), .Z(n30273) );
  XNOR U30277 ( .A(p_input[1599]), .B(n17303), .Z(n30280) );
  XOR U30278 ( .A(n30270), .B(n30279), .Z(n30333) );
  XOR U30279 ( .A(n30334), .B(n30276), .Z(n30279) );
  XOR U30280 ( .A(p_input[1597]), .B(p_input[2077]), .Z(n30276) );
  XOR U30281 ( .A(p_input[1598]), .B(n17305), .Z(n30334) );
  XOR U30282 ( .A(p_input[1593]), .B(p_input[2073]), .Z(n30270) );
  XOR U30283 ( .A(n30292), .B(n30291), .Z(n30257) );
  XNOR U30284 ( .A(n30335), .B(n30299), .Z(n30291) );
  XNOR U30285 ( .A(n30287), .B(n30286), .Z(n30299) );
  XNOR U30286 ( .A(n30336), .B(n30283), .Z(n30286) );
  XNOR U30287 ( .A(p_input[1579]), .B(p_input[2059]), .Z(n30283) );
  XOR U30288 ( .A(p_input[1580]), .B(n16451), .Z(n30336) );
  XOR U30289 ( .A(p_input[1581]), .B(p_input[2061]), .Z(n30287) );
  XOR U30290 ( .A(n30297), .B(n30337), .Z(n30335) );
  IV U30291 ( .A(n30288), .Z(n30337) );
  XOR U30292 ( .A(p_input[1570]), .B(p_input[2050]), .Z(n30288) );
  XNOR U30293 ( .A(n30338), .B(n30304), .Z(n30297) );
  XNOR U30294 ( .A(p_input[1584]), .B(n16454), .Z(n30304) );
  XOR U30295 ( .A(n30294), .B(n30303), .Z(n30338) );
  XOR U30296 ( .A(n30339), .B(n30300), .Z(n30303) );
  XOR U30297 ( .A(p_input[1582]), .B(p_input[2062]), .Z(n30300) );
  XOR U30298 ( .A(p_input[1583]), .B(n16456), .Z(n30339) );
  XOR U30299 ( .A(p_input[1578]), .B(p_input[2058]), .Z(n30294) );
  XOR U30300 ( .A(n30311), .B(n30309), .Z(n30292) );
  XNOR U30301 ( .A(n30340), .B(n30316), .Z(n30309) );
  XOR U30302 ( .A(p_input[1577]), .B(p_input[2057]), .Z(n30316) );
  XOR U30303 ( .A(n30306), .B(n30315), .Z(n30340) );
  XOR U30304 ( .A(n30341), .B(n30312), .Z(n30315) );
  XOR U30305 ( .A(p_input[1575]), .B(p_input[2055]), .Z(n30312) );
  XOR U30306 ( .A(p_input[1576]), .B(n17312), .Z(n30341) );
  XOR U30307 ( .A(p_input[1571]), .B(p_input[2051]), .Z(n30306) );
  XNOR U30308 ( .A(n30321), .B(n30320), .Z(n30311) );
  XOR U30309 ( .A(n30342), .B(n30317), .Z(n30320) );
  XOR U30310 ( .A(p_input[1572]), .B(p_input[2052]), .Z(n30317) );
  XOR U30311 ( .A(p_input[1573]), .B(n17314), .Z(n30342) );
  XOR U30312 ( .A(p_input[1574]), .B(p_input[2054]), .Z(n30321) );
  XNOR U30313 ( .A(n30343), .B(n30344), .Z(n30134) );
  AND U30314 ( .A(n606), .B(n30345), .Z(n30344) );
  XNOR U30315 ( .A(n30346), .B(n30347), .Z(n606) );
  AND U30316 ( .A(n30348), .B(n30349), .Z(n30347) );
  XOR U30317 ( .A(n30346), .B(n30144), .Z(n30349) );
  XNOR U30318 ( .A(n30346), .B(n30086), .Z(n30348) );
  XOR U30319 ( .A(n30350), .B(n30351), .Z(n30346) );
  AND U30320 ( .A(n30352), .B(n30353), .Z(n30351) );
  XNOR U30321 ( .A(n30157), .B(n30350), .Z(n30353) );
  XOR U30322 ( .A(n30350), .B(n30098), .Z(n30352) );
  XOR U30323 ( .A(n30354), .B(n30355), .Z(n30350) );
  AND U30324 ( .A(n30356), .B(n30357), .Z(n30355) );
  XNOR U30325 ( .A(n30182), .B(n30354), .Z(n30357) );
  XOR U30326 ( .A(n30354), .B(n30109), .Z(n30356) );
  XOR U30327 ( .A(n30358), .B(n30359), .Z(n30354) );
  AND U30328 ( .A(n30360), .B(n30361), .Z(n30359) );
  XOR U30329 ( .A(n30358), .B(n30119), .Z(n30360) );
  XOR U30330 ( .A(n30362), .B(n30363), .Z(n30075) );
  AND U30331 ( .A(n610), .B(n30345), .Z(n30363) );
  XNOR U30332 ( .A(n30343), .B(n30362), .Z(n30345) );
  XNOR U30333 ( .A(n30364), .B(n30365), .Z(n610) );
  AND U30334 ( .A(n30366), .B(n30367), .Z(n30365) );
  XNOR U30335 ( .A(n30368), .B(n30364), .Z(n30367) );
  IV U30336 ( .A(n30144), .Z(n30368) );
  XNOR U30337 ( .A(n30369), .B(n30370), .Z(n30144) );
  AND U30338 ( .A(n613), .B(n30371), .Z(n30370) );
  XNOR U30339 ( .A(n30369), .B(n30372), .Z(n30371) );
  XNOR U30340 ( .A(n30086), .B(n30364), .Z(n30366) );
  XOR U30341 ( .A(n30373), .B(n30374), .Z(n30086) );
  AND U30342 ( .A(n621), .B(n30375), .Z(n30374) );
  XOR U30343 ( .A(n30376), .B(n30377), .Z(n30364) );
  AND U30344 ( .A(n30378), .B(n30379), .Z(n30377) );
  XNOR U30345 ( .A(n30376), .B(n30157), .Z(n30379) );
  XNOR U30346 ( .A(n30380), .B(n30381), .Z(n30157) );
  AND U30347 ( .A(n613), .B(n30382), .Z(n30381) );
  XOR U30348 ( .A(n30383), .B(n30380), .Z(n30382) );
  XNOR U30349 ( .A(n30384), .B(n30376), .Z(n30378) );
  IV U30350 ( .A(n30098), .Z(n30384) );
  XOR U30351 ( .A(n30385), .B(n30386), .Z(n30098) );
  AND U30352 ( .A(n621), .B(n30387), .Z(n30386) );
  XOR U30353 ( .A(n30388), .B(n30389), .Z(n30376) );
  AND U30354 ( .A(n30390), .B(n30391), .Z(n30389) );
  XNOR U30355 ( .A(n30388), .B(n30182), .Z(n30391) );
  XNOR U30356 ( .A(n30392), .B(n30393), .Z(n30182) );
  AND U30357 ( .A(n613), .B(n30394), .Z(n30393) );
  XNOR U30358 ( .A(n30395), .B(n30392), .Z(n30394) );
  XOR U30359 ( .A(n30109), .B(n30388), .Z(n30390) );
  XOR U30360 ( .A(n30396), .B(n30397), .Z(n30109) );
  AND U30361 ( .A(n621), .B(n30398), .Z(n30397) );
  XOR U30362 ( .A(n30358), .B(n30399), .Z(n30388) );
  AND U30363 ( .A(n30400), .B(n30361), .Z(n30399) );
  XNOR U30364 ( .A(n30228), .B(n30358), .Z(n30361) );
  XNOR U30365 ( .A(n30401), .B(n30402), .Z(n30228) );
  AND U30366 ( .A(n613), .B(n30403), .Z(n30402) );
  XOR U30367 ( .A(n30404), .B(n30401), .Z(n30403) );
  XNOR U30368 ( .A(n30405), .B(n30358), .Z(n30400) );
  IV U30369 ( .A(n30119), .Z(n30405) );
  XOR U30370 ( .A(n30406), .B(n30407), .Z(n30119) );
  AND U30371 ( .A(n621), .B(n30408), .Z(n30407) );
  XOR U30372 ( .A(n30409), .B(n30410), .Z(n30358) );
  AND U30373 ( .A(n30411), .B(n30412), .Z(n30410) );
  XNOR U30374 ( .A(n30409), .B(n30322), .Z(n30412) );
  XNOR U30375 ( .A(n30413), .B(n30414), .Z(n30322) );
  AND U30376 ( .A(n613), .B(n30415), .Z(n30414) );
  XNOR U30377 ( .A(n30416), .B(n30413), .Z(n30415) );
  XNOR U30378 ( .A(n30417), .B(n30409), .Z(n30411) );
  IV U30379 ( .A(n30131), .Z(n30417) );
  XOR U30380 ( .A(n30418), .B(n30419), .Z(n30131) );
  AND U30381 ( .A(n621), .B(n30420), .Z(n30419) );
  AND U30382 ( .A(n30362), .B(n30343), .Z(n30409) );
  XNOR U30383 ( .A(n30421), .B(n30422), .Z(n30343) );
  AND U30384 ( .A(n613), .B(n30423), .Z(n30422) );
  XNOR U30385 ( .A(n30424), .B(n30421), .Z(n30423) );
  XNOR U30386 ( .A(n30425), .B(n30426), .Z(n613) );
  AND U30387 ( .A(n30427), .B(n30428), .Z(n30426) );
  XOR U30388 ( .A(n30372), .B(n30425), .Z(n30428) );
  AND U30389 ( .A(n30429), .B(n30430), .Z(n30372) );
  XOR U30390 ( .A(n30425), .B(n30369), .Z(n30427) );
  XNOR U30391 ( .A(n30431), .B(n30432), .Z(n30369) );
  AND U30392 ( .A(n617), .B(n30375), .Z(n30432) );
  XOR U30393 ( .A(n30373), .B(n30431), .Z(n30375) );
  XOR U30394 ( .A(n30433), .B(n30434), .Z(n30425) );
  AND U30395 ( .A(n30435), .B(n30436), .Z(n30434) );
  XNOR U30396 ( .A(n30433), .B(n30429), .Z(n30436) );
  IV U30397 ( .A(n30383), .Z(n30429) );
  XOR U30398 ( .A(n30437), .B(n30438), .Z(n30383) );
  XOR U30399 ( .A(n30439), .B(n30430), .Z(n30438) );
  AND U30400 ( .A(n30395), .B(n30440), .Z(n30430) );
  AND U30401 ( .A(n30441), .B(n30442), .Z(n30439) );
  XOR U30402 ( .A(n30443), .B(n30437), .Z(n30441) );
  XNOR U30403 ( .A(n30380), .B(n30433), .Z(n30435) );
  XNOR U30404 ( .A(n30444), .B(n30445), .Z(n30380) );
  AND U30405 ( .A(n617), .B(n30387), .Z(n30445) );
  XOR U30406 ( .A(n30444), .B(n30385), .Z(n30387) );
  XOR U30407 ( .A(n30446), .B(n30447), .Z(n30433) );
  AND U30408 ( .A(n30448), .B(n30449), .Z(n30447) );
  XNOR U30409 ( .A(n30446), .B(n30395), .Z(n30449) );
  XOR U30410 ( .A(n30450), .B(n30442), .Z(n30395) );
  XNOR U30411 ( .A(n30451), .B(n30437), .Z(n30442) );
  XOR U30412 ( .A(n30452), .B(n30453), .Z(n30437) );
  AND U30413 ( .A(n30454), .B(n30455), .Z(n30453) );
  XOR U30414 ( .A(n30456), .B(n30452), .Z(n30454) );
  XNOR U30415 ( .A(n30457), .B(n30458), .Z(n30451) );
  AND U30416 ( .A(n30459), .B(n30460), .Z(n30458) );
  XOR U30417 ( .A(n30457), .B(n30461), .Z(n30459) );
  XNOR U30418 ( .A(n30443), .B(n30440), .Z(n30450) );
  AND U30419 ( .A(n30462), .B(n30463), .Z(n30440) );
  XOR U30420 ( .A(n30464), .B(n30465), .Z(n30443) );
  AND U30421 ( .A(n30466), .B(n30467), .Z(n30465) );
  XOR U30422 ( .A(n30464), .B(n30468), .Z(n30466) );
  XNOR U30423 ( .A(n30392), .B(n30446), .Z(n30448) );
  XNOR U30424 ( .A(n30469), .B(n30470), .Z(n30392) );
  AND U30425 ( .A(n617), .B(n30398), .Z(n30470) );
  XOR U30426 ( .A(n30469), .B(n30396), .Z(n30398) );
  XOR U30427 ( .A(n30471), .B(n30472), .Z(n30446) );
  AND U30428 ( .A(n30473), .B(n30474), .Z(n30472) );
  XNOR U30429 ( .A(n30471), .B(n30462), .Z(n30474) );
  IV U30430 ( .A(n30404), .Z(n30462) );
  XNOR U30431 ( .A(n30475), .B(n30455), .Z(n30404) );
  XNOR U30432 ( .A(n30476), .B(n30461), .Z(n30455) );
  XOR U30433 ( .A(n30477), .B(n30478), .Z(n30461) );
  AND U30434 ( .A(n30479), .B(n30480), .Z(n30478) );
  XOR U30435 ( .A(n30477), .B(n30481), .Z(n30479) );
  XNOR U30436 ( .A(n30460), .B(n30452), .Z(n30476) );
  XOR U30437 ( .A(n30482), .B(n30483), .Z(n30452) );
  AND U30438 ( .A(n30484), .B(n30485), .Z(n30483) );
  XNOR U30439 ( .A(n30486), .B(n30482), .Z(n30484) );
  XNOR U30440 ( .A(n30487), .B(n30457), .Z(n30460) );
  XOR U30441 ( .A(n30488), .B(n30489), .Z(n30457) );
  AND U30442 ( .A(n30490), .B(n30491), .Z(n30489) );
  XOR U30443 ( .A(n30488), .B(n30492), .Z(n30490) );
  XNOR U30444 ( .A(n30493), .B(n30494), .Z(n30487) );
  AND U30445 ( .A(n30495), .B(n30496), .Z(n30494) );
  XNOR U30446 ( .A(n30493), .B(n30497), .Z(n30495) );
  XNOR U30447 ( .A(n30456), .B(n30463), .Z(n30475) );
  AND U30448 ( .A(n30416), .B(n30498), .Z(n30463) );
  XOR U30449 ( .A(n30468), .B(n30467), .Z(n30456) );
  XNOR U30450 ( .A(n30499), .B(n30464), .Z(n30467) );
  XOR U30451 ( .A(n30500), .B(n30501), .Z(n30464) );
  AND U30452 ( .A(n30502), .B(n30503), .Z(n30501) );
  XOR U30453 ( .A(n30500), .B(n30504), .Z(n30502) );
  XNOR U30454 ( .A(n30505), .B(n30506), .Z(n30499) );
  AND U30455 ( .A(n30507), .B(n30508), .Z(n30506) );
  XOR U30456 ( .A(n30505), .B(n30509), .Z(n30507) );
  XOR U30457 ( .A(n30510), .B(n30511), .Z(n30468) );
  AND U30458 ( .A(n30512), .B(n30513), .Z(n30511) );
  XOR U30459 ( .A(n30510), .B(n30514), .Z(n30512) );
  XNOR U30460 ( .A(n30401), .B(n30471), .Z(n30473) );
  XNOR U30461 ( .A(n30515), .B(n30516), .Z(n30401) );
  AND U30462 ( .A(n617), .B(n30408), .Z(n30516) );
  XOR U30463 ( .A(n30515), .B(n30406), .Z(n30408) );
  XOR U30464 ( .A(n30517), .B(n30518), .Z(n30471) );
  AND U30465 ( .A(n30519), .B(n30520), .Z(n30518) );
  XNOR U30466 ( .A(n30517), .B(n30416), .Z(n30520) );
  XOR U30467 ( .A(n30521), .B(n30485), .Z(n30416) );
  XNOR U30468 ( .A(n30522), .B(n30492), .Z(n30485) );
  XOR U30469 ( .A(n30481), .B(n30480), .Z(n30492) );
  XNOR U30470 ( .A(n30523), .B(n30477), .Z(n30480) );
  XOR U30471 ( .A(n30524), .B(n30525), .Z(n30477) );
  AND U30472 ( .A(n30526), .B(n30527), .Z(n30525) );
  XNOR U30473 ( .A(n30528), .B(n30529), .Z(n30526) );
  IV U30474 ( .A(n30524), .Z(n30528) );
  XNOR U30475 ( .A(n30530), .B(n30531), .Z(n30523) );
  NOR U30476 ( .A(n30532), .B(n30533), .Z(n30531) );
  XNOR U30477 ( .A(n30530), .B(n30534), .Z(n30532) );
  XOR U30478 ( .A(n30535), .B(n30536), .Z(n30481) );
  NOR U30479 ( .A(n30537), .B(n30538), .Z(n30536) );
  XNOR U30480 ( .A(n30535), .B(n30539), .Z(n30537) );
  XNOR U30481 ( .A(n30491), .B(n30482), .Z(n30522) );
  XOR U30482 ( .A(n30540), .B(n30541), .Z(n30482) );
  AND U30483 ( .A(n30542), .B(n30543), .Z(n30541) );
  XOR U30484 ( .A(n30540), .B(n30544), .Z(n30542) );
  XOR U30485 ( .A(n30545), .B(n30497), .Z(n30491) );
  XOR U30486 ( .A(n30546), .B(n30547), .Z(n30497) );
  NOR U30487 ( .A(n30548), .B(n30549), .Z(n30547) );
  XOR U30488 ( .A(n30546), .B(n30550), .Z(n30548) );
  XNOR U30489 ( .A(n30496), .B(n30488), .Z(n30545) );
  XOR U30490 ( .A(n30551), .B(n30552), .Z(n30488) );
  AND U30491 ( .A(n30553), .B(n30554), .Z(n30552) );
  XOR U30492 ( .A(n30551), .B(n30555), .Z(n30553) );
  XNOR U30493 ( .A(n30556), .B(n30493), .Z(n30496) );
  XOR U30494 ( .A(n30557), .B(n30558), .Z(n30493) );
  AND U30495 ( .A(n30559), .B(n30560), .Z(n30558) );
  XNOR U30496 ( .A(n30561), .B(n30562), .Z(n30559) );
  IV U30497 ( .A(n30557), .Z(n30561) );
  XNOR U30498 ( .A(n30563), .B(n30564), .Z(n30556) );
  NOR U30499 ( .A(n30565), .B(n30566), .Z(n30564) );
  XNOR U30500 ( .A(n30563), .B(n30567), .Z(n30565) );
  XOR U30501 ( .A(n30486), .B(n30498), .Z(n30521) );
  NOR U30502 ( .A(n30424), .B(n30568), .Z(n30498) );
  XNOR U30503 ( .A(n30504), .B(n30503), .Z(n30486) );
  XNOR U30504 ( .A(n30569), .B(n30509), .Z(n30503) );
  XNOR U30505 ( .A(n30570), .B(n30571), .Z(n30509) );
  NOR U30506 ( .A(n30572), .B(n30573), .Z(n30571) );
  XOR U30507 ( .A(n30570), .B(n30574), .Z(n30572) );
  XNOR U30508 ( .A(n30508), .B(n30500), .Z(n30569) );
  XOR U30509 ( .A(n30575), .B(n30576), .Z(n30500) );
  AND U30510 ( .A(n30577), .B(n30578), .Z(n30576) );
  XOR U30511 ( .A(n30575), .B(n30579), .Z(n30577) );
  XNOR U30512 ( .A(n30580), .B(n30505), .Z(n30508) );
  XOR U30513 ( .A(n30581), .B(n30582), .Z(n30505) );
  AND U30514 ( .A(n30583), .B(n30584), .Z(n30582) );
  XNOR U30515 ( .A(n30585), .B(n30586), .Z(n30583) );
  IV U30516 ( .A(n30581), .Z(n30585) );
  XNOR U30517 ( .A(n30587), .B(n30588), .Z(n30580) );
  NOR U30518 ( .A(n30589), .B(n30590), .Z(n30588) );
  XNOR U30519 ( .A(n30587), .B(n30591), .Z(n30589) );
  XOR U30520 ( .A(n30514), .B(n30513), .Z(n30504) );
  XNOR U30521 ( .A(n30592), .B(n30510), .Z(n30513) );
  XOR U30522 ( .A(n30593), .B(n30594), .Z(n30510) );
  AND U30523 ( .A(n30595), .B(n30596), .Z(n30594) );
  XNOR U30524 ( .A(n30597), .B(n30598), .Z(n30595) );
  IV U30525 ( .A(n30593), .Z(n30597) );
  XNOR U30526 ( .A(n30599), .B(n30600), .Z(n30592) );
  NOR U30527 ( .A(n30601), .B(n30602), .Z(n30600) );
  XNOR U30528 ( .A(n30599), .B(n30603), .Z(n30601) );
  XOR U30529 ( .A(n30604), .B(n30605), .Z(n30514) );
  NOR U30530 ( .A(n30606), .B(n30607), .Z(n30605) );
  XNOR U30531 ( .A(n30604), .B(n30608), .Z(n30606) );
  XNOR U30532 ( .A(n30413), .B(n30517), .Z(n30519) );
  XNOR U30533 ( .A(n30609), .B(n30610), .Z(n30413) );
  AND U30534 ( .A(n617), .B(n30420), .Z(n30610) );
  XOR U30535 ( .A(n30609), .B(n30418), .Z(n30420) );
  AND U30536 ( .A(n30421), .B(n30424), .Z(n30517) );
  XOR U30537 ( .A(n30611), .B(n30568), .Z(n30424) );
  XNOR U30538 ( .A(p_input[1600]), .B(p_input[2048]), .Z(n30568) );
  XNOR U30539 ( .A(n30544), .B(n30543), .Z(n30611) );
  XNOR U30540 ( .A(n30612), .B(n30555), .Z(n30543) );
  XOR U30541 ( .A(n30529), .B(n30527), .Z(n30555) );
  XNOR U30542 ( .A(n30613), .B(n30534), .Z(n30527) );
  XOR U30543 ( .A(p_input[1624]), .B(p_input[2072]), .Z(n30534) );
  XOR U30544 ( .A(n30524), .B(n30533), .Z(n30613) );
  XOR U30545 ( .A(n30614), .B(n30530), .Z(n30533) );
  XOR U30546 ( .A(p_input[1622]), .B(p_input[2070]), .Z(n30530) );
  XOR U30547 ( .A(p_input[1623]), .B(n17295), .Z(n30614) );
  XOR U30548 ( .A(p_input[1618]), .B(p_input[2066]), .Z(n30524) );
  XNOR U30549 ( .A(n30539), .B(n30538), .Z(n30529) );
  XOR U30550 ( .A(n30615), .B(n30535), .Z(n30538) );
  XOR U30551 ( .A(p_input[1619]), .B(p_input[2067]), .Z(n30535) );
  XOR U30552 ( .A(p_input[1620]), .B(n17297), .Z(n30615) );
  XOR U30553 ( .A(p_input[1621]), .B(p_input[2069]), .Z(n30539) );
  XOR U30554 ( .A(n30554), .B(n30616), .Z(n30612) );
  IV U30555 ( .A(n30540), .Z(n30616) );
  XOR U30556 ( .A(p_input[1601]), .B(p_input[2049]), .Z(n30540) );
  XNOR U30557 ( .A(n30617), .B(n30562), .Z(n30554) );
  XNOR U30558 ( .A(n30550), .B(n30549), .Z(n30562) );
  XNOR U30559 ( .A(n30618), .B(n30546), .Z(n30549) );
  XNOR U30560 ( .A(p_input[1626]), .B(p_input[2074]), .Z(n30546) );
  XOR U30561 ( .A(p_input[1627]), .B(n17300), .Z(n30618) );
  XOR U30562 ( .A(p_input[1628]), .B(p_input[2076]), .Z(n30550) );
  XOR U30563 ( .A(n30560), .B(n30619), .Z(n30617) );
  IV U30564 ( .A(n30551), .Z(n30619) );
  XOR U30565 ( .A(p_input[1617]), .B(p_input[2065]), .Z(n30551) );
  XNOR U30566 ( .A(n30620), .B(n30567), .Z(n30560) );
  XNOR U30567 ( .A(p_input[1631]), .B(n17303), .Z(n30567) );
  XOR U30568 ( .A(n30557), .B(n30566), .Z(n30620) );
  XOR U30569 ( .A(n30621), .B(n30563), .Z(n30566) );
  XOR U30570 ( .A(p_input[1629]), .B(p_input[2077]), .Z(n30563) );
  XOR U30571 ( .A(p_input[1630]), .B(n17305), .Z(n30621) );
  XOR U30572 ( .A(p_input[1625]), .B(p_input[2073]), .Z(n30557) );
  XOR U30573 ( .A(n30579), .B(n30578), .Z(n30544) );
  XNOR U30574 ( .A(n30622), .B(n30586), .Z(n30578) );
  XNOR U30575 ( .A(n30574), .B(n30573), .Z(n30586) );
  XNOR U30576 ( .A(n30623), .B(n30570), .Z(n30573) );
  XNOR U30577 ( .A(p_input[1611]), .B(p_input[2059]), .Z(n30570) );
  XOR U30578 ( .A(p_input[1612]), .B(n16451), .Z(n30623) );
  XOR U30579 ( .A(p_input[1613]), .B(p_input[2061]), .Z(n30574) );
  XOR U30580 ( .A(n30584), .B(n30624), .Z(n30622) );
  IV U30581 ( .A(n30575), .Z(n30624) );
  XOR U30582 ( .A(p_input[1602]), .B(p_input[2050]), .Z(n30575) );
  XNOR U30583 ( .A(n30625), .B(n30591), .Z(n30584) );
  XNOR U30584 ( .A(p_input[1616]), .B(n16454), .Z(n30591) );
  XOR U30585 ( .A(n30581), .B(n30590), .Z(n30625) );
  XOR U30586 ( .A(n30626), .B(n30587), .Z(n30590) );
  XOR U30587 ( .A(p_input[1614]), .B(p_input[2062]), .Z(n30587) );
  XOR U30588 ( .A(p_input[1615]), .B(n16456), .Z(n30626) );
  XOR U30589 ( .A(p_input[1610]), .B(p_input[2058]), .Z(n30581) );
  XOR U30590 ( .A(n30598), .B(n30596), .Z(n30579) );
  XNOR U30591 ( .A(n30627), .B(n30603), .Z(n30596) );
  XOR U30592 ( .A(p_input[1609]), .B(p_input[2057]), .Z(n30603) );
  XOR U30593 ( .A(n30593), .B(n30602), .Z(n30627) );
  XOR U30594 ( .A(n30628), .B(n30599), .Z(n30602) );
  XOR U30595 ( .A(p_input[1607]), .B(p_input[2055]), .Z(n30599) );
  XOR U30596 ( .A(p_input[1608]), .B(n17312), .Z(n30628) );
  XOR U30597 ( .A(p_input[1603]), .B(p_input[2051]), .Z(n30593) );
  XNOR U30598 ( .A(n30608), .B(n30607), .Z(n30598) );
  XOR U30599 ( .A(n30629), .B(n30604), .Z(n30607) );
  XOR U30600 ( .A(p_input[1604]), .B(p_input[2052]), .Z(n30604) );
  XOR U30601 ( .A(p_input[1605]), .B(n17314), .Z(n30629) );
  XOR U30602 ( .A(p_input[1606]), .B(p_input[2054]), .Z(n30608) );
  XNOR U30603 ( .A(n30630), .B(n30631), .Z(n30421) );
  AND U30604 ( .A(n617), .B(n30632), .Z(n30631) );
  XNOR U30605 ( .A(n30633), .B(n30634), .Z(n617) );
  AND U30606 ( .A(n30635), .B(n30636), .Z(n30634) );
  XOR U30607 ( .A(n30633), .B(n30431), .Z(n30636) );
  XNOR U30608 ( .A(n30633), .B(n30373), .Z(n30635) );
  XOR U30609 ( .A(n30637), .B(n30638), .Z(n30633) );
  AND U30610 ( .A(n30639), .B(n30640), .Z(n30638) );
  XNOR U30611 ( .A(n30444), .B(n30637), .Z(n30640) );
  XOR U30612 ( .A(n30637), .B(n30385), .Z(n30639) );
  XOR U30613 ( .A(n30641), .B(n30642), .Z(n30637) );
  AND U30614 ( .A(n30643), .B(n30644), .Z(n30642) );
  XNOR U30615 ( .A(n30469), .B(n30641), .Z(n30644) );
  XOR U30616 ( .A(n30641), .B(n30396), .Z(n30643) );
  XOR U30617 ( .A(n30645), .B(n30646), .Z(n30641) );
  AND U30618 ( .A(n30647), .B(n30648), .Z(n30646) );
  XOR U30619 ( .A(n30645), .B(n30406), .Z(n30647) );
  XOR U30620 ( .A(n30649), .B(n30650), .Z(n30362) );
  AND U30621 ( .A(n621), .B(n30632), .Z(n30650) );
  XNOR U30622 ( .A(n30630), .B(n30649), .Z(n30632) );
  XNOR U30623 ( .A(n30651), .B(n30652), .Z(n621) );
  AND U30624 ( .A(n30653), .B(n30654), .Z(n30652) );
  XNOR U30625 ( .A(n30655), .B(n30651), .Z(n30654) );
  IV U30626 ( .A(n30431), .Z(n30655) );
  XNOR U30627 ( .A(n30656), .B(n30657), .Z(n30431) );
  AND U30628 ( .A(n624), .B(n30658), .Z(n30657) );
  XNOR U30629 ( .A(n30656), .B(n30659), .Z(n30658) );
  XNOR U30630 ( .A(n30373), .B(n30651), .Z(n30653) );
  XOR U30631 ( .A(n30660), .B(n30661), .Z(n30373) );
  AND U30632 ( .A(n632), .B(n30662), .Z(n30661) );
  XOR U30633 ( .A(n30663), .B(n30664), .Z(n30651) );
  AND U30634 ( .A(n30665), .B(n30666), .Z(n30664) );
  XNOR U30635 ( .A(n30663), .B(n30444), .Z(n30666) );
  XNOR U30636 ( .A(n30667), .B(n30668), .Z(n30444) );
  AND U30637 ( .A(n624), .B(n30669), .Z(n30668) );
  XOR U30638 ( .A(n30670), .B(n30667), .Z(n30669) );
  XNOR U30639 ( .A(n30671), .B(n30663), .Z(n30665) );
  IV U30640 ( .A(n30385), .Z(n30671) );
  XOR U30641 ( .A(n30672), .B(n30673), .Z(n30385) );
  AND U30642 ( .A(n632), .B(n30674), .Z(n30673) );
  XOR U30643 ( .A(n30675), .B(n30676), .Z(n30663) );
  AND U30644 ( .A(n30677), .B(n30678), .Z(n30676) );
  XNOR U30645 ( .A(n30675), .B(n30469), .Z(n30678) );
  XNOR U30646 ( .A(n30679), .B(n30680), .Z(n30469) );
  AND U30647 ( .A(n624), .B(n30681), .Z(n30680) );
  XNOR U30648 ( .A(n30682), .B(n30679), .Z(n30681) );
  XOR U30649 ( .A(n30396), .B(n30675), .Z(n30677) );
  XOR U30650 ( .A(n30683), .B(n30684), .Z(n30396) );
  AND U30651 ( .A(n632), .B(n30685), .Z(n30684) );
  XOR U30652 ( .A(n30645), .B(n30686), .Z(n30675) );
  AND U30653 ( .A(n30687), .B(n30648), .Z(n30686) );
  XNOR U30654 ( .A(n30515), .B(n30645), .Z(n30648) );
  XNOR U30655 ( .A(n30688), .B(n30689), .Z(n30515) );
  AND U30656 ( .A(n624), .B(n30690), .Z(n30689) );
  XOR U30657 ( .A(n30691), .B(n30688), .Z(n30690) );
  XNOR U30658 ( .A(n30692), .B(n30645), .Z(n30687) );
  IV U30659 ( .A(n30406), .Z(n30692) );
  XOR U30660 ( .A(n30693), .B(n30694), .Z(n30406) );
  AND U30661 ( .A(n632), .B(n30695), .Z(n30694) );
  XOR U30662 ( .A(n30696), .B(n30697), .Z(n30645) );
  AND U30663 ( .A(n30698), .B(n30699), .Z(n30697) );
  XNOR U30664 ( .A(n30696), .B(n30609), .Z(n30699) );
  XNOR U30665 ( .A(n30700), .B(n30701), .Z(n30609) );
  AND U30666 ( .A(n624), .B(n30702), .Z(n30701) );
  XNOR U30667 ( .A(n30703), .B(n30700), .Z(n30702) );
  XNOR U30668 ( .A(n30704), .B(n30696), .Z(n30698) );
  IV U30669 ( .A(n30418), .Z(n30704) );
  XOR U30670 ( .A(n30705), .B(n30706), .Z(n30418) );
  AND U30671 ( .A(n632), .B(n30707), .Z(n30706) );
  AND U30672 ( .A(n30649), .B(n30630), .Z(n30696) );
  XNOR U30673 ( .A(n30708), .B(n30709), .Z(n30630) );
  AND U30674 ( .A(n624), .B(n30710), .Z(n30709) );
  XNOR U30675 ( .A(n30711), .B(n30708), .Z(n30710) );
  XNOR U30676 ( .A(n30712), .B(n30713), .Z(n624) );
  AND U30677 ( .A(n30714), .B(n30715), .Z(n30713) );
  XOR U30678 ( .A(n30659), .B(n30712), .Z(n30715) );
  AND U30679 ( .A(n30716), .B(n30717), .Z(n30659) );
  XOR U30680 ( .A(n30712), .B(n30656), .Z(n30714) );
  XNOR U30681 ( .A(n30718), .B(n30719), .Z(n30656) );
  AND U30682 ( .A(n628), .B(n30662), .Z(n30719) );
  XOR U30683 ( .A(n30660), .B(n30718), .Z(n30662) );
  XOR U30684 ( .A(n30720), .B(n30721), .Z(n30712) );
  AND U30685 ( .A(n30722), .B(n30723), .Z(n30721) );
  XNOR U30686 ( .A(n30720), .B(n30716), .Z(n30723) );
  IV U30687 ( .A(n30670), .Z(n30716) );
  XOR U30688 ( .A(n30724), .B(n30725), .Z(n30670) );
  XOR U30689 ( .A(n30726), .B(n30717), .Z(n30725) );
  AND U30690 ( .A(n30682), .B(n30727), .Z(n30717) );
  AND U30691 ( .A(n30728), .B(n30729), .Z(n30726) );
  XOR U30692 ( .A(n30730), .B(n30724), .Z(n30728) );
  XNOR U30693 ( .A(n30667), .B(n30720), .Z(n30722) );
  XNOR U30694 ( .A(n30731), .B(n30732), .Z(n30667) );
  AND U30695 ( .A(n628), .B(n30674), .Z(n30732) );
  XOR U30696 ( .A(n30731), .B(n30672), .Z(n30674) );
  XOR U30697 ( .A(n30733), .B(n30734), .Z(n30720) );
  AND U30698 ( .A(n30735), .B(n30736), .Z(n30734) );
  XNOR U30699 ( .A(n30733), .B(n30682), .Z(n30736) );
  XOR U30700 ( .A(n30737), .B(n30729), .Z(n30682) );
  XNOR U30701 ( .A(n30738), .B(n30724), .Z(n30729) );
  XOR U30702 ( .A(n30739), .B(n30740), .Z(n30724) );
  AND U30703 ( .A(n30741), .B(n30742), .Z(n30740) );
  XOR U30704 ( .A(n30743), .B(n30739), .Z(n30741) );
  XNOR U30705 ( .A(n30744), .B(n30745), .Z(n30738) );
  AND U30706 ( .A(n30746), .B(n30747), .Z(n30745) );
  XOR U30707 ( .A(n30744), .B(n30748), .Z(n30746) );
  XNOR U30708 ( .A(n30730), .B(n30727), .Z(n30737) );
  AND U30709 ( .A(n30749), .B(n30750), .Z(n30727) );
  XOR U30710 ( .A(n30751), .B(n30752), .Z(n30730) );
  AND U30711 ( .A(n30753), .B(n30754), .Z(n30752) );
  XOR U30712 ( .A(n30751), .B(n30755), .Z(n30753) );
  XNOR U30713 ( .A(n30679), .B(n30733), .Z(n30735) );
  XNOR U30714 ( .A(n30756), .B(n30757), .Z(n30679) );
  AND U30715 ( .A(n628), .B(n30685), .Z(n30757) );
  XOR U30716 ( .A(n30756), .B(n30683), .Z(n30685) );
  XOR U30717 ( .A(n30758), .B(n30759), .Z(n30733) );
  AND U30718 ( .A(n30760), .B(n30761), .Z(n30759) );
  XNOR U30719 ( .A(n30758), .B(n30749), .Z(n30761) );
  IV U30720 ( .A(n30691), .Z(n30749) );
  XNOR U30721 ( .A(n30762), .B(n30742), .Z(n30691) );
  XNOR U30722 ( .A(n30763), .B(n30748), .Z(n30742) );
  XOR U30723 ( .A(n30764), .B(n30765), .Z(n30748) );
  AND U30724 ( .A(n30766), .B(n30767), .Z(n30765) );
  XOR U30725 ( .A(n30764), .B(n30768), .Z(n30766) );
  XNOR U30726 ( .A(n30747), .B(n30739), .Z(n30763) );
  XOR U30727 ( .A(n30769), .B(n30770), .Z(n30739) );
  AND U30728 ( .A(n30771), .B(n30772), .Z(n30770) );
  XNOR U30729 ( .A(n30773), .B(n30769), .Z(n30771) );
  XNOR U30730 ( .A(n30774), .B(n30744), .Z(n30747) );
  XOR U30731 ( .A(n30775), .B(n30776), .Z(n30744) );
  AND U30732 ( .A(n30777), .B(n30778), .Z(n30776) );
  XOR U30733 ( .A(n30775), .B(n30779), .Z(n30777) );
  XNOR U30734 ( .A(n30780), .B(n30781), .Z(n30774) );
  AND U30735 ( .A(n30782), .B(n30783), .Z(n30781) );
  XNOR U30736 ( .A(n30780), .B(n30784), .Z(n30782) );
  XNOR U30737 ( .A(n30743), .B(n30750), .Z(n30762) );
  AND U30738 ( .A(n30703), .B(n30785), .Z(n30750) );
  XOR U30739 ( .A(n30755), .B(n30754), .Z(n30743) );
  XNOR U30740 ( .A(n30786), .B(n30751), .Z(n30754) );
  XOR U30741 ( .A(n30787), .B(n30788), .Z(n30751) );
  AND U30742 ( .A(n30789), .B(n30790), .Z(n30788) );
  XOR U30743 ( .A(n30787), .B(n30791), .Z(n30789) );
  XNOR U30744 ( .A(n30792), .B(n30793), .Z(n30786) );
  AND U30745 ( .A(n30794), .B(n30795), .Z(n30793) );
  XOR U30746 ( .A(n30792), .B(n30796), .Z(n30794) );
  XOR U30747 ( .A(n30797), .B(n30798), .Z(n30755) );
  AND U30748 ( .A(n30799), .B(n30800), .Z(n30798) );
  XOR U30749 ( .A(n30797), .B(n30801), .Z(n30799) );
  XNOR U30750 ( .A(n30688), .B(n30758), .Z(n30760) );
  XNOR U30751 ( .A(n30802), .B(n30803), .Z(n30688) );
  AND U30752 ( .A(n628), .B(n30695), .Z(n30803) );
  XOR U30753 ( .A(n30802), .B(n30693), .Z(n30695) );
  XOR U30754 ( .A(n30804), .B(n30805), .Z(n30758) );
  AND U30755 ( .A(n30806), .B(n30807), .Z(n30805) );
  XNOR U30756 ( .A(n30804), .B(n30703), .Z(n30807) );
  XOR U30757 ( .A(n30808), .B(n30772), .Z(n30703) );
  XNOR U30758 ( .A(n30809), .B(n30779), .Z(n30772) );
  XOR U30759 ( .A(n30768), .B(n30767), .Z(n30779) );
  XNOR U30760 ( .A(n30810), .B(n30764), .Z(n30767) );
  XOR U30761 ( .A(n30811), .B(n30812), .Z(n30764) );
  AND U30762 ( .A(n30813), .B(n30814), .Z(n30812) );
  XNOR U30763 ( .A(n30815), .B(n30816), .Z(n30813) );
  IV U30764 ( .A(n30811), .Z(n30815) );
  XNOR U30765 ( .A(n30817), .B(n30818), .Z(n30810) );
  NOR U30766 ( .A(n30819), .B(n30820), .Z(n30818) );
  XNOR U30767 ( .A(n30817), .B(n30821), .Z(n30819) );
  XOR U30768 ( .A(n30822), .B(n30823), .Z(n30768) );
  NOR U30769 ( .A(n30824), .B(n30825), .Z(n30823) );
  XNOR U30770 ( .A(n30822), .B(n30826), .Z(n30824) );
  XNOR U30771 ( .A(n30778), .B(n30769), .Z(n30809) );
  XOR U30772 ( .A(n30827), .B(n30828), .Z(n30769) );
  AND U30773 ( .A(n30829), .B(n30830), .Z(n30828) );
  XOR U30774 ( .A(n30827), .B(n30831), .Z(n30829) );
  XOR U30775 ( .A(n30832), .B(n30784), .Z(n30778) );
  XOR U30776 ( .A(n30833), .B(n30834), .Z(n30784) );
  NOR U30777 ( .A(n30835), .B(n30836), .Z(n30834) );
  XOR U30778 ( .A(n30833), .B(n30837), .Z(n30835) );
  XNOR U30779 ( .A(n30783), .B(n30775), .Z(n30832) );
  XOR U30780 ( .A(n30838), .B(n30839), .Z(n30775) );
  AND U30781 ( .A(n30840), .B(n30841), .Z(n30839) );
  XOR U30782 ( .A(n30838), .B(n30842), .Z(n30840) );
  XNOR U30783 ( .A(n30843), .B(n30780), .Z(n30783) );
  XOR U30784 ( .A(n30844), .B(n30845), .Z(n30780) );
  AND U30785 ( .A(n30846), .B(n30847), .Z(n30845) );
  XNOR U30786 ( .A(n30848), .B(n30849), .Z(n30846) );
  IV U30787 ( .A(n30844), .Z(n30848) );
  XNOR U30788 ( .A(n30850), .B(n30851), .Z(n30843) );
  NOR U30789 ( .A(n30852), .B(n30853), .Z(n30851) );
  XNOR U30790 ( .A(n30850), .B(n30854), .Z(n30852) );
  XOR U30791 ( .A(n30773), .B(n30785), .Z(n30808) );
  NOR U30792 ( .A(n30711), .B(n30855), .Z(n30785) );
  XNOR U30793 ( .A(n30791), .B(n30790), .Z(n30773) );
  XNOR U30794 ( .A(n30856), .B(n30796), .Z(n30790) );
  XNOR U30795 ( .A(n30857), .B(n30858), .Z(n30796) );
  NOR U30796 ( .A(n30859), .B(n30860), .Z(n30858) );
  XOR U30797 ( .A(n30857), .B(n30861), .Z(n30859) );
  XNOR U30798 ( .A(n30795), .B(n30787), .Z(n30856) );
  XOR U30799 ( .A(n30862), .B(n30863), .Z(n30787) );
  AND U30800 ( .A(n30864), .B(n30865), .Z(n30863) );
  XOR U30801 ( .A(n30862), .B(n30866), .Z(n30864) );
  XNOR U30802 ( .A(n30867), .B(n30792), .Z(n30795) );
  XOR U30803 ( .A(n30868), .B(n30869), .Z(n30792) );
  AND U30804 ( .A(n30870), .B(n30871), .Z(n30869) );
  XNOR U30805 ( .A(n30872), .B(n30873), .Z(n30870) );
  IV U30806 ( .A(n30868), .Z(n30872) );
  XNOR U30807 ( .A(n30874), .B(n30875), .Z(n30867) );
  NOR U30808 ( .A(n30876), .B(n30877), .Z(n30875) );
  XNOR U30809 ( .A(n30874), .B(n30878), .Z(n30876) );
  XOR U30810 ( .A(n30801), .B(n30800), .Z(n30791) );
  XNOR U30811 ( .A(n30879), .B(n30797), .Z(n30800) );
  XOR U30812 ( .A(n30880), .B(n30881), .Z(n30797) );
  AND U30813 ( .A(n30882), .B(n30883), .Z(n30881) );
  XNOR U30814 ( .A(n30884), .B(n30885), .Z(n30882) );
  IV U30815 ( .A(n30880), .Z(n30884) );
  XNOR U30816 ( .A(n30886), .B(n30887), .Z(n30879) );
  NOR U30817 ( .A(n30888), .B(n30889), .Z(n30887) );
  XNOR U30818 ( .A(n30886), .B(n30890), .Z(n30888) );
  XOR U30819 ( .A(n30891), .B(n30892), .Z(n30801) );
  NOR U30820 ( .A(n30893), .B(n30894), .Z(n30892) );
  XNOR U30821 ( .A(n30891), .B(n30895), .Z(n30893) );
  XNOR U30822 ( .A(n30700), .B(n30804), .Z(n30806) );
  XNOR U30823 ( .A(n30896), .B(n30897), .Z(n30700) );
  AND U30824 ( .A(n628), .B(n30707), .Z(n30897) );
  XOR U30825 ( .A(n30896), .B(n30705), .Z(n30707) );
  AND U30826 ( .A(n30708), .B(n30711), .Z(n30804) );
  XOR U30827 ( .A(n30898), .B(n30855), .Z(n30711) );
  XNOR U30828 ( .A(p_input[1632]), .B(p_input[2048]), .Z(n30855) );
  XNOR U30829 ( .A(n30831), .B(n30830), .Z(n30898) );
  XNOR U30830 ( .A(n30899), .B(n30842), .Z(n30830) );
  XOR U30831 ( .A(n30816), .B(n30814), .Z(n30842) );
  XNOR U30832 ( .A(n30900), .B(n30821), .Z(n30814) );
  XOR U30833 ( .A(p_input[1656]), .B(p_input[2072]), .Z(n30821) );
  XOR U30834 ( .A(n30811), .B(n30820), .Z(n30900) );
  XOR U30835 ( .A(n30901), .B(n30817), .Z(n30820) );
  XOR U30836 ( .A(p_input[1654]), .B(p_input[2070]), .Z(n30817) );
  XOR U30837 ( .A(p_input[1655]), .B(n17295), .Z(n30901) );
  XOR U30838 ( .A(p_input[1650]), .B(p_input[2066]), .Z(n30811) );
  XNOR U30839 ( .A(n30826), .B(n30825), .Z(n30816) );
  XOR U30840 ( .A(n30902), .B(n30822), .Z(n30825) );
  XOR U30841 ( .A(p_input[1651]), .B(p_input[2067]), .Z(n30822) );
  XOR U30842 ( .A(p_input[1652]), .B(n17297), .Z(n30902) );
  XOR U30843 ( .A(p_input[1653]), .B(p_input[2069]), .Z(n30826) );
  XOR U30844 ( .A(n30841), .B(n30903), .Z(n30899) );
  IV U30845 ( .A(n30827), .Z(n30903) );
  XOR U30846 ( .A(p_input[1633]), .B(p_input[2049]), .Z(n30827) );
  XNOR U30847 ( .A(n30904), .B(n30849), .Z(n30841) );
  XNOR U30848 ( .A(n30837), .B(n30836), .Z(n30849) );
  XNOR U30849 ( .A(n30905), .B(n30833), .Z(n30836) );
  XNOR U30850 ( .A(p_input[1658]), .B(p_input[2074]), .Z(n30833) );
  XOR U30851 ( .A(p_input[1659]), .B(n17300), .Z(n30905) );
  XOR U30852 ( .A(p_input[1660]), .B(p_input[2076]), .Z(n30837) );
  XOR U30853 ( .A(n30847), .B(n30906), .Z(n30904) );
  IV U30854 ( .A(n30838), .Z(n30906) );
  XOR U30855 ( .A(p_input[1649]), .B(p_input[2065]), .Z(n30838) );
  XNOR U30856 ( .A(n30907), .B(n30854), .Z(n30847) );
  XNOR U30857 ( .A(p_input[1663]), .B(n17303), .Z(n30854) );
  XOR U30858 ( .A(n30844), .B(n30853), .Z(n30907) );
  XOR U30859 ( .A(n30908), .B(n30850), .Z(n30853) );
  XOR U30860 ( .A(p_input[1661]), .B(p_input[2077]), .Z(n30850) );
  XOR U30861 ( .A(p_input[1662]), .B(n17305), .Z(n30908) );
  XOR U30862 ( .A(p_input[1657]), .B(p_input[2073]), .Z(n30844) );
  XOR U30863 ( .A(n30866), .B(n30865), .Z(n30831) );
  XNOR U30864 ( .A(n30909), .B(n30873), .Z(n30865) );
  XNOR U30865 ( .A(n30861), .B(n30860), .Z(n30873) );
  XNOR U30866 ( .A(n30910), .B(n30857), .Z(n30860) );
  XNOR U30867 ( .A(p_input[1643]), .B(p_input[2059]), .Z(n30857) );
  XOR U30868 ( .A(p_input[1644]), .B(n16451), .Z(n30910) );
  XOR U30869 ( .A(p_input[1645]), .B(p_input[2061]), .Z(n30861) );
  XOR U30870 ( .A(n30871), .B(n30911), .Z(n30909) );
  IV U30871 ( .A(n30862), .Z(n30911) );
  XOR U30872 ( .A(p_input[1634]), .B(p_input[2050]), .Z(n30862) );
  XNOR U30873 ( .A(n30912), .B(n30878), .Z(n30871) );
  XNOR U30874 ( .A(p_input[1648]), .B(n16454), .Z(n30878) );
  XOR U30875 ( .A(n30868), .B(n30877), .Z(n30912) );
  XOR U30876 ( .A(n30913), .B(n30874), .Z(n30877) );
  XOR U30877 ( .A(p_input[1646]), .B(p_input[2062]), .Z(n30874) );
  XOR U30878 ( .A(p_input[1647]), .B(n16456), .Z(n30913) );
  XOR U30879 ( .A(p_input[1642]), .B(p_input[2058]), .Z(n30868) );
  XOR U30880 ( .A(n30885), .B(n30883), .Z(n30866) );
  XNOR U30881 ( .A(n30914), .B(n30890), .Z(n30883) );
  XOR U30882 ( .A(p_input[1641]), .B(p_input[2057]), .Z(n30890) );
  XOR U30883 ( .A(n30880), .B(n30889), .Z(n30914) );
  XOR U30884 ( .A(n30915), .B(n30886), .Z(n30889) );
  XOR U30885 ( .A(p_input[1639]), .B(p_input[2055]), .Z(n30886) );
  XOR U30886 ( .A(p_input[1640]), .B(n17312), .Z(n30915) );
  XOR U30887 ( .A(p_input[1635]), .B(p_input[2051]), .Z(n30880) );
  XNOR U30888 ( .A(n30895), .B(n30894), .Z(n30885) );
  XOR U30889 ( .A(n30916), .B(n30891), .Z(n30894) );
  XOR U30890 ( .A(p_input[1636]), .B(p_input[2052]), .Z(n30891) );
  XOR U30891 ( .A(p_input[1637]), .B(n17314), .Z(n30916) );
  XOR U30892 ( .A(p_input[1638]), .B(p_input[2054]), .Z(n30895) );
  XNOR U30893 ( .A(n30917), .B(n30918), .Z(n30708) );
  AND U30894 ( .A(n628), .B(n30919), .Z(n30918) );
  XNOR U30895 ( .A(n30920), .B(n30921), .Z(n628) );
  AND U30896 ( .A(n30922), .B(n30923), .Z(n30921) );
  XOR U30897 ( .A(n30920), .B(n30718), .Z(n30923) );
  XNOR U30898 ( .A(n30920), .B(n30660), .Z(n30922) );
  XOR U30899 ( .A(n30924), .B(n30925), .Z(n30920) );
  AND U30900 ( .A(n30926), .B(n30927), .Z(n30925) );
  XNOR U30901 ( .A(n30731), .B(n30924), .Z(n30927) );
  XOR U30902 ( .A(n30924), .B(n30672), .Z(n30926) );
  XOR U30903 ( .A(n30928), .B(n30929), .Z(n30924) );
  AND U30904 ( .A(n30930), .B(n30931), .Z(n30929) );
  XNOR U30905 ( .A(n30756), .B(n30928), .Z(n30931) );
  XOR U30906 ( .A(n30928), .B(n30683), .Z(n30930) );
  XOR U30907 ( .A(n30932), .B(n30933), .Z(n30928) );
  AND U30908 ( .A(n30934), .B(n30935), .Z(n30933) );
  XOR U30909 ( .A(n30932), .B(n30693), .Z(n30934) );
  XOR U30910 ( .A(n30936), .B(n30937), .Z(n30649) );
  AND U30911 ( .A(n632), .B(n30919), .Z(n30937) );
  XNOR U30912 ( .A(n30917), .B(n30936), .Z(n30919) );
  XNOR U30913 ( .A(n30938), .B(n30939), .Z(n632) );
  AND U30914 ( .A(n30940), .B(n30941), .Z(n30939) );
  XNOR U30915 ( .A(n30942), .B(n30938), .Z(n30941) );
  IV U30916 ( .A(n30718), .Z(n30942) );
  XNOR U30917 ( .A(n30943), .B(n30944), .Z(n30718) );
  AND U30918 ( .A(n635), .B(n30945), .Z(n30944) );
  XNOR U30919 ( .A(n30943), .B(n30946), .Z(n30945) );
  XNOR U30920 ( .A(n30660), .B(n30938), .Z(n30940) );
  XOR U30921 ( .A(n30947), .B(n30948), .Z(n30660) );
  AND U30922 ( .A(n643), .B(n30949), .Z(n30948) );
  XOR U30923 ( .A(n30950), .B(n30951), .Z(n30938) );
  AND U30924 ( .A(n30952), .B(n30953), .Z(n30951) );
  XNOR U30925 ( .A(n30950), .B(n30731), .Z(n30953) );
  XNOR U30926 ( .A(n30954), .B(n30955), .Z(n30731) );
  AND U30927 ( .A(n635), .B(n30956), .Z(n30955) );
  XOR U30928 ( .A(n30957), .B(n30954), .Z(n30956) );
  XNOR U30929 ( .A(n30958), .B(n30950), .Z(n30952) );
  IV U30930 ( .A(n30672), .Z(n30958) );
  XOR U30931 ( .A(n30959), .B(n30960), .Z(n30672) );
  AND U30932 ( .A(n643), .B(n30961), .Z(n30960) );
  XOR U30933 ( .A(n30962), .B(n30963), .Z(n30950) );
  AND U30934 ( .A(n30964), .B(n30965), .Z(n30963) );
  XNOR U30935 ( .A(n30962), .B(n30756), .Z(n30965) );
  XNOR U30936 ( .A(n30966), .B(n30967), .Z(n30756) );
  AND U30937 ( .A(n635), .B(n30968), .Z(n30967) );
  XNOR U30938 ( .A(n30969), .B(n30966), .Z(n30968) );
  XOR U30939 ( .A(n30683), .B(n30962), .Z(n30964) );
  XOR U30940 ( .A(n30970), .B(n30971), .Z(n30683) );
  AND U30941 ( .A(n643), .B(n30972), .Z(n30971) );
  XOR U30942 ( .A(n30932), .B(n30973), .Z(n30962) );
  AND U30943 ( .A(n30974), .B(n30935), .Z(n30973) );
  XNOR U30944 ( .A(n30802), .B(n30932), .Z(n30935) );
  XNOR U30945 ( .A(n30975), .B(n30976), .Z(n30802) );
  AND U30946 ( .A(n635), .B(n30977), .Z(n30976) );
  XOR U30947 ( .A(n30978), .B(n30975), .Z(n30977) );
  XNOR U30948 ( .A(n30979), .B(n30932), .Z(n30974) );
  IV U30949 ( .A(n30693), .Z(n30979) );
  XOR U30950 ( .A(n30980), .B(n30981), .Z(n30693) );
  AND U30951 ( .A(n643), .B(n30982), .Z(n30981) );
  XOR U30952 ( .A(n30983), .B(n30984), .Z(n30932) );
  AND U30953 ( .A(n30985), .B(n30986), .Z(n30984) );
  XNOR U30954 ( .A(n30983), .B(n30896), .Z(n30986) );
  XNOR U30955 ( .A(n30987), .B(n30988), .Z(n30896) );
  AND U30956 ( .A(n635), .B(n30989), .Z(n30988) );
  XNOR U30957 ( .A(n30990), .B(n30987), .Z(n30989) );
  XNOR U30958 ( .A(n30991), .B(n30983), .Z(n30985) );
  IV U30959 ( .A(n30705), .Z(n30991) );
  XOR U30960 ( .A(n30992), .B(n30993), .Z(n30705) );
  AND U30961 ( .A(n643), .B(n30994), .Z(n30993) );
  AND U30962 ( .A(n30936), .B(n30917), .Z(n30983) );
  XNOR U30963 ( .A(n30995), .B(n30996), .Z(n30917) );
  AND U30964 ( .A(n635), .B(n30997), .Z(n30996) );
  XNOR U30965 ( .A(n30998), .B(n30995), .Z(n30997) );
  XNOR U30966 ( .A(n30999), .B(n31000), .Z(n635) );
  AND U30967 ( .A(n31001), .B(n31002), .Z(n31000) );
  XOR U30968 ( .A(n30946), .B(n30999), .Z(n31002) );
  AND U30969 ( .A(n31003), .B(n31004), .Z(n30946) );
  XOR U30970 ( .A(n30999), .B(n30943), .Z(n31001) );
  XNOR U30971 ( .A(n31005), .B(n31006), .Z(n30943) );
  AND U30972 ( .A(n639), .B(n30949), .Z(n31006) );
  XOR U30973 ( .A(n30947), .B(n31005), .Z(n30949) );
  XOR U30974 ( .A(n31007), .B(n31008), .Z(n30999) );
  AND U30975 ( .A(n31009), .B(n31010), .Z(n31008) );
  XNOR U30976 ( .A(n31007), .B(n31003), .Z(n31010) );
  IV U30977 ( .A(n30957), .Z(n31003) );
  XOR U30978 ( .A(n31011), .B(n31012), .Z(n30957) );
  XOR U30979 ( .A(n31013), .B(n31004), .Z(n31012) );
  AND U30980 ( .A(n30969), .B(n31014), .Z(n31004) );
  AND U30981 ( .A(n31015), .B(n31016), .Z(n31013) );
  XOR U30982 ( .A(n31017), .B(n31011), .Z(n31015) );
  XNOR U30983 ( .A(n30954), .B(n31007), .Z(n31009) );
  XNOR U30984 ( .A(n31018), .B(n31019), .Z(n30954) );
  AND U30985 ( .A(n639), .B(n30961), .Z(n31019) );
  XOR U30986 ( .A(n31018), .B(n30959), .Z(n30961) );
  XOR U30987 ( .A(n31020), .B(n31021), .Z(n31007) );
  AND U30988 ( .A(n31022), .B(n31023), .Z(n31021) );
  XNOR U30989 ( .A(n31020), .B(n30969), .Z(n31023) );
  XOR U30990 ( .A(n31024), .B(n31016), .Z(n30969) );
  XNOR U30991 ( .A(n31025), .B(n31011), .Z(n31016) );
  XOR U30992 ( .A(n31026), .B(n31027), .Z(n31011) );
  AND U30993 ( .A(n31028), .B(n31029), .Z(n31027) );
  XOR U30994 ( .A(n31030), .B(n31026), .Z(n31028) );
  XNOR U30995 ( .A(n31031), .B(n31032), .Z(n31025) );
  AND U30996 ( .A(n31033), .B(n31034), .Z(n31032) );
  XOR U30997 ( .A(n31031), .B(n31035), .Z(n31033) );
  XNOR U30998 ( .A(n31017), .B(n31014), .Z(n31024) );
  AND U30999 ( .A(n31036), .B(n31037), .Z(n31014) );
  XOR U31000 ( .A(n31038), .B(n31039), .Z(n31017) );
  AND U31001 ( .A(n31040), .B(n31041), .Z(n31039) );
  XOR U31002 ( .A(n31038), .B(n31042), .Z(n31040) );
  XNOR U31003 ( .A(n30966), .B(n31020), .Z(n31022) );
  XNOR U31004 ( .A(n31043), .B(n31044), .Z(n30966) );
  AND U31005 ( .A(n639), .B(n30972), .Z(n31044) );
  XOR U31006 ( .A(n31043), .B(n30970), .Z(n30972) );
  XOR U31007 ( .A(n31045), .B(n31046), .Z(n31020) );
  AND U31008 ( .A(n31047), .B(n31048), .Z(n31046) );
  XNOR U31009 ( .A(n31045), .B(n31036), .Z(n31048) );
  IV U31010 ( .A(n30978), .Z(n31036) );
  XNOR U31011 ( .A(n31049), .B(n31029), .Z(n30978) );
  XNOR U31012 ( .A(n31050), .B(n31035), .Z(n31029) );
  XOR U31013 ( .A(n31051), .B(n31052), .Z(n31035) );
  AND U31014 ( .A(n31053), .B(n31054), .Z(n31052) );
  XOR U31015 ( .A(n31051), .B(n31055), .Z(n31053) );
  XNOR U31016 ( .A(n31034), .B(n31026), .Z(n31050) );
  XOR U31017 ( .A(n31056), .B(n31057), .Z(n31026) );
  AND U31018 ( .A(n31058), .B(n31059), .Z(n31057) );
  XNOR U31019 ( .A(n31060), .B(n31056), .Z(n31058) );
  XNOR U31020 ( .A(n31061), .B(n31031), .Z(n31034) );
  XOR U31021 ( .A(n31062), .B(n31063), .Z(n31031) );
  AND U31022 ( .A(n31064), .B(n31065), .Z(n31063) );
  XOR U31023 ( .A(n31062), .B(n31066), .Z(n31064) );
  XNOR U31024 ( .A(n31067), .B(n31068), .Z(n31061) );
  AND U31025 ( .A(n31069), .B(n31070), .Z(n31068) );
  XNOR U31026 ( .A(n31067), .B(n31071), .Z(n31069) );
  XNOR U31027 ( .A(n31030), .B(n31037), .Z(n31049) );
  AND U31028 ( .A(n30990), .B(n31072), .Z(n31037) );
  XOR U31029 ( .A(n31042), .B(n31041), .Z(n31030) );
  XNOR U31030 ( .A(n31073), .B(n31038), .Z(n31041) );
  XOR U31031 ( .A(n31074), .B(n31075), .Z(n31038) );
  AND U31032 ( .A(n31076), .B(n31077), .Z(n31075) );
  XOR U31033 ( .A(n31074), .B(n31078), .Z(n31076) );
  XNOR U31034 ( .A(n31079), .B(n31080), .Z(n31073) );
  AND U31035 ( .A(n31081), .B(n31082), .Z(n31080) );
  XOR U31036 ( .A(n31079), .B(n31083), .Z(n31081) );
  XOR U31037 ( .A(n31084), .B(n31085), .Z(n31042) );
  AND U31038 ( .A(n31086), .B(n31087), .Z(n31085) );
  XOR U31039 ( .A(n31084), .B(n31088), .Z(n31086) );
  XNOR U31040 ( .A(n30975), .B(n31045), .Z(n31047) );
  XNOR U31041 ( .A(n31089), .B(n31090), .Z(n30975) );
  AND U31042 ( .A(n639), .B(n30982), .Z(n31090) );
  XOR U31043 ( .A(n31089), .B(n30980), .Z(n30982) );
  XOR U31044 ( .A(n31091), .B(n31092), .Z(n31045) );
  AND U31045 ( .A(n31093), .B(n31094), .Z(n31092) );
  XNOR U31046 ( .A(n31091), .B(n30990), .Z(n31094) );
  XOR U31047 ( .A(n31095), .B(n31059), .Z(n30990) );
  XNOR U31048 ( .A(n31096), .B(n31066), .Z(n31059) );
  XOR U31049 ( .A(n31055), .B(n31054), .Z(n31066) );
  XNOR U31050 ( .A(n31097), .B(n31051), .Z(n31054) );
  XOR U31051 ( .A(n31098), .B(n31099), .Z(n31051) );
  AND U31052 ( .A(n31100), .B(n31101), .Z(n31099) );
  XNOR U31053 ( .A(n31102), .B(n31103), .Z(n31100) );
  IV U31054 ( .A(n31098), .Z(n31102) );
  XNOR U31055 ( .A(n31104), .B(n31105), .Z(n31097) );
  NOR U31056 ( .A(n31106), .B(n31107), .Z(n31105) );
  XNOR U31057 ( .A(n31104), .B(n31108), .Z(n31106) );
  XOR U31058 ( .A(n31109), .B(n31110), .Z(n31055) );
  NOR U31059 ( .A(n31111), .B(n31112), .Z(n31110) );
  XNOR U31060 ( .A(n31109), .B(n31113), .Z(n31111) );
  XNOR U31061 ( .A(n31065), .B(n31056), .Z(n31096) );
  XOR U31062 ( .A(n31114), .B(n31115), .Z(n31056) );
  AND U31063 ( .A(n31116), .B(n31117), .Z(n31115) );
  XOR U31064 ( .A(n31114), .B(n31118), .Z(n31116) );
  XOR U31065 ( .A(n31119), .B(n31071), .Z(n31065) );
  XOR U31066 ( .A(n31120), .B(n31121), .Z(n31071) );
  NOR U31067 ( .A(n31122), .B(n31123), .Z(n31121) );
  XOR U31068 ( .A(n31120), .B(n31124), .Z(n31122) );
  XNOR U31069 ( .A(n31070), .B(n31062), .Z(n31119) );
  XOR U31070 ( .A(n31125), .B(n31126), .Z(n31062) );
  AND U31071 ( .A(n31127), .B(n31128), .Z(n31126) );
  XOR U31072 ( .A(n31125), .B(n31129), .Z(n31127) );
  XNOR U31073 ( .A(n31130), .B(n31067), .Z(n31070) );
  XOR U31074 ( .A(n31131), .B(n31132), .Z(n31067) );
  AND U31075 ( .A(n31133), .B(n31134), .Z(n31132) );
  XNOR U31076 ( .A(n31135), .B(n31136), .Z(n31133) );
  IV U31077 ( .A(n31131), .Z(n31135) );
  XNOR U31078 ( .A(n31137), .B(n31138), .Z(n31130) );
  NOR U31079 ( .A(n31139), .B(n31140), .Z(n31138) );
  XNOR U31080 ( .A(n31137), .B(n31141), .Z(n31139) );
  XOR U31081 ( .A(n31060), .B(n31072), .Z(n31095) );
  NOR U31082 ( .A(n30998), .B(n31142), .Z(n31072) );
  XNOR U31083 ( .A(n31078), .B(n31077), .Z(n31060) );
  XNOR U31084 ( .A(n31143), .B(n31083), .Z(n31077) );
  XNOR U31085 ( .A(n31144), .B(n31145), .Z(n31083) );
  NOR U31086 ( .A(n31146), .B(n31147), .Z(n31145) );
  XOR U31087 ( .A(n31144), .B(n31148), .Z(n31146) );
  XNOR U31088 ( .A(n31082), .B(n31074), .Z(n31143) );
  XOR U31089 ( .A(n31149), .B(n31150), .Z(n31074) );
  AND U31090 ( .A(n31151), .B(n31152), .Z(n31150) );
  XOR U31091 ( .A(n31149), .B(n31153), .Z(n31151) );
  XNOR U31092 ( .A(n31154), .B(n31079), .Z(n31082) );
  XOR U31093 ( .A(n31155), .B(n31156), .Z(n31079) );
  AND U31094 ( .A(n31157), .B(n31158), .Z(n31156) );
  XNOR U31095 ( .A(n31159), .B(n31160), .Z(n31157) );
  IV U31096 ( .A(n31155), .Z(n31159) );
  XNOR U31097 ( .A(n31161), .B(n31162), .Z(n31154) );
  NOR U31098 ( .A(n31163), .B(n31164), .Z(n31162) );
  XNOR U31099 ( .A(n31161), .B(n31165), .Z(n31163) );
  XOR U31100 ( .A(n31088), .B(n31087), .Z(n31078) );
  XNOR U31101 ( .A(n31166), .B(n31084), .Z(n31087) );
  XOR U31102 ( .A(n31167), .B(n31168), .Z(n31084) );
  AND U31103 ( .A(n31169), .B(n31170), .Z(n31168) );
  XNOR U31104 ( .A(n31171), .B(n31172), .Z(n31169) );
  IV U31105 ( .A(n31167), .Z(n31171) );
  XNOR U31106 ( .A(n31173), .B(n31174), .Z(n31166) );
  NOR U31107 ( .A(n31175), .B(n31176), .Z(n31174) );
  XNOR U31108 ( .A(n31173), .B(n31177), .Z(n31175) );
  XOR U31109 ( .A(n31178), .B(n31179), .Z(n31088) );
  NOR U31110 ( .A(n31180), .B(n31181), .Z(n31179) );
  XNOR U31111 ( .A(n31178), .B(n31182), .Z(n31180) );
  XNOR U31112 ( .A(n30987), .B(n31091), .Z(n31093) );
  XNOR U31113 ( .A(n31183), .B(n31184), .Z(n30987) );
  AND U31114 ( .A(n639), .B(n30994), .Z(n31184) );
  XOR U31115 ( .A(n31183), .B(n30992), .Z(n30994) );
  AND U31116 ( .A(n30995), .B(n30998), .Z(n31091) );
  XOR U31117 ( .A(n31185), .B(n31142), .Z(n30998) );
  XNOR U31118 ( .A(p_input[1664]), .B(p_input[2048]), .Z(n31142) );
  XNOR U31119 ( .A(n31118), .B(n31117), .Z(n31185) );
  XNOR U31120 ( .A(n31186), .B(n31129), .Z(n31117) );
  XOR U31121 ( .A(n31103), .B(n31101), .Z(n31129) );
  XNOR U31122 ( .A(n31187), .B(n31108), .Z(n31101) );
  XOR U31123 ( .A(p_input[1688]), .B(p_input[2072]), .Z(n31108) );
  XOR U31124 ( .A(n31098), .B(n31107), .Z(n31187) );
  XOR U31125 ( .A(n31188), .B(n31104), .Z(n31107) );
  XOR U31126 ( .A(p_input[1686]), .B(p_input[2070]), .Z(n31104) );
  XOR U31127 ( .A(p_input[1687]), .B(n17295), .Z(n31188) );
  XOR U31128 ( .A(p_input[1682]), .B(p_input[2066]), .Z(n31098) );
  XNOR U31129 ( .A(n31113), .B(n31112), .Z(n31103) );
  XOR U31130 ( .A(n31189), .B(n31109), .Z(n31112) );
  XOR U31131 ( .A(p_input[1683]), .B(p_input[2067]), .Z(n31109) );
  XOR U31132 ( .A(p_input[1684]), .B(n17297), .Z(n31189) );
  XOR U31133 ( .A(p_input[1685]), .B(p_input[2069]), .Z(n31113) );
  XOR U31134 ( .A(n31128), .B(n31190), .Z(n31186) );
  IV U31135 ( .A(n31114), .Z(n31190) );
  XOR U31136 ( .A(p_input[1665]), .B(p_input[2049]), .Z(n31114) );
  XNOR U31137 ( .A(n31191), .B(n31136), .Z(n31128) );
  XNOR U31138 ( .A(n31124), .B(n31123), .Z(n31136) );
  XNOR U31139 ( .A(n31192), .B(n31120), .Z(n31123) );
  XNOR U31140 ( .A(p_input[1690]), .B(p_input[2074]), .Z(n31120) );
  XOR U31141 ( .A(p_input[1691]), .B(n17300), .Z(n31192) );
  XOR U31142 ( .A(p_input[1692]), .B(p_input[2076]), .Z(n31124) );
  XOR U31143 ( .A(n31134), .B(n31193), .Z(n31191) );
  IV U31144 ( .A(n31125), .Z(n31193) );
  XOR U31145 ( .A(p_input[1681]), .B(p_input[2065]), .Z(n31125) );
  XNOR U31146 ( .A(n31194), .B(n31141), .Z(n31134) );
  XNOR U31147 ( .A(p_input[1695]), .B(n17303), .Z(n31141) );
  XOR U31148 ( .A(n31131), .B(n31140), .Z(n31194) );
  XOR U31149 ( .A(n31195), .B(n31137), .Z(n31140) );
  XOR U31150 ( .A(p_input[1693]), .B(p_input[2077]), .Z(n31137) );
  XOR U31151 ( .A(p_input[1694]), .B(n17305), .Z(n31195) );
  XOR U31152 ( .A(p_input[1689]), .B(p_input[2073]), .Z(n31131) );
  XOR U31153 ( .A(n31153), .B(n31152), .Z(n31118) );
  XNOR U31154 ( .A(n31196), .B(n31160), .Z(n31152) );
  XNOR U31155 ( .A(n31148), .B(n31147), .Z(n31160) );
  XNOR U31156 ( .A(n31197), .B(n31144), .Z(n31147) );
  XNOR U31157 ( .A(p_input[1675]), .B(p_input[2059]), .Z(n31144) );
  XOR U31158 ( .A(p_input[1676]), .B(n16451), .Z(n31197) );
  XOR U31159 ( .A(p_input[1677]), .B(p_input[2061]), .Z(n31148) );
  XOR U31160 ( .A(n31158), .B(n31198), .Z(n31196) );
  IV U31161 ( .A(n31149), .Z(n31198) );
  XOR U31162 ( .A(p_input[1666]), .B(p_input[2050]), .Z(n31149) );
  XNOR U31163 ( .A(n31199), .B(n31165), .Z(n31158) );
  XNOR U31164 ( .A(p_input[1680]), .B(n16454), .Z(n31165) );
  XOR U31165 ( .A(n31155), .B(n31164), .Z(n31199) );
  XOR U31166 ( .A(n31200), .B(n31161), .Z(n31164) );
  XOR U31167 ( .A(p_input[1678]), .B(p_input[2062]), .Z(n31161) );
  XOR U31168 ( .A(p_input[1679]), .B(n16456), .Z(n31200) );
  XOR U31169 ( .A(p_input[1674]), .B(p_input[2058]), .Z(n31155) );
  XOR U31170 ( .A(n31172), .B(n31170), .Z(n31153) );
  XNOR U31171 ( .A(n31201), .B(n31177), .Z(n31170) );
  XOR U31172 ( .A(p_input[1673]), .B(p_input[2057]), .Z(n31177) );
  XOR U31173 ( .A(n31167), .B(n31176), .Z(n31201) );
  XOR U31174 ( .A(n31202), .B(n31173), .Z(n31176) );
  XOR U31175 ( .A(p_input[1671]), .B(p_input[2055]), .Z(n31173) );
  XOR U31176 ( .A(p_input[1672]), .B(n17312), .Z(n31202) );
  XOR U31177 ( .A(p_input[1667]), .B(p_input[2051]), .Z(n31167) );
  XNOR U31178 ( .A(n31182), .B(n31181), .Z(n31172) );
  XOR U31179 ( .A(n31203), .B(n31178), .Z(n31181) );
  XOR U31180 ( .A(p_input[1668]), .B(p_input[2052]), .Z(n31178) );
  XOR U31181 ( .A(p_input[1669]), .B(n17314), .Z(n31203) );
  XOR U31182 ( .A(p_input[1670]), .B(p_input[2054]), .Z(n31182) );
  XNOR U31183 ( .A(n31204), .B(n31205), .Z(n30995) );
  AND U31184 ( .A(n639), .B(n31206), .Z(n31205) );
  XNOR U31185 ( .A(n31207), .B(n31208), .Z(n639) );
  AND U31186 ( .A(n31209), .B(n31210), .Z(n31208) );
  XOR U31187 ( .A(n31207), .B(n31005), .Z(n31210) );
  XNOR U31188 ( .A(n31207), .B(n30947), .Z(n31209) );
  XOR U31189 ( .A(n31211), .B(n31212), .Z(n31207) );
  AND U31190 ( .A(n31213), .B(n31214), .Z(n31212) );
  XNOR U31191 ( .A(n31018), .B(n31211), .Z(n31214) );
  XOR U31192 ( .A(n31211), .B(n30959), .Z(n31213) );
  XOR U31193 ( .A(n31215), .B(n31216), .Z(n31211) );
  AND U31194 ( .A(n31217), .B(n31218), .Z(n31216) );
  XNOR U31195 ( .A(n31043), .B(n31215), .Z(n31218) );
  XOR U31196 ( .A(n31215), .B(n30970), .Z(n31217) );
  XOR U31197 ( .A(n31219), .B(n31220), .Z(n31215) );
  AND U31198 ( .A(n31221), .B(n31222), .Z(n31220) );
  XOR U31199 ( .A(n31219), .B(n30980), .Z(n31221) );
  XOR U31200 ( .A(n31223), .B(n31224), .Z(n30936) );
  AND U31201 ( .A(n643), .B(n31206), .Z(n31224) );
  XNOR U31202 ( .A(n31204), .B(n31223), .Z(n31206) );
  XNOR U31203 ( .A(n31225), .B(n31226), .Z(n643) );
  AND U31204 ( .A(n31227), .B(n31228), .Z(n31226) );
  XNOR U31205 ( .A(n31229), .B(n31225), .Z(n31228) );
  IV U31206 ( .A(n31005), .Z(n31229) );
  XNOR U31207 ( .A(n31230), .B(n31231), .Z(n31005) );
  AND U31208 ( .A(n646), .B(n31232), .Z(n31231) );
  XNOR U31209 ( .A(n31230), .B(n31233), .Z(n31232) );
  XNOR U31210 ( .A(n30947), .B(n31225), .Z(n31227) );
  XOR U31211 ( .A(n31234), .B(n31235), .Z(n30947) );
  AND U31212 ( .A(n654), .B(n31236), .Z(n31235) );
  XOR U31213 ( .A(n31237), .B(n31238), .Z(n31225) );
  AND U31214 ( .A(n31239), .B(n31240), .Z(n31238) );
  XNOR U31215 ( .A(n31237), .B(n31018), .Z(n31240) );
  XNOR U31216 ( .A(n31241), .B(n31242), .Z(n31018) );
  AND U31217 ( .A(n646), .B(n31243), .Z(n31242) );
  XOR U31218 ( .A(n31244), .B(n31241), .Z(n31243) );
  XNOR U31219 ( .A(n31245), .B(n31237), .Z(n31239) );
  IV U31220 ( .A(n30959), .Z(n31245) );
  XOR U31221 ( .A(n31246), .B(n31247), .Z(n30959) );
  AND U31222 ( .A(n654), .B(n31248), .Z(n31247) );
  XOR U31223 ( .A(n31249), .B(n31250), .Z(n31237) );
  AND U31224 ( .A(n31251), .B(n31252), .Z(n31250) );
  XNOR U31225 ( .A(n31249), .B(n31043), .Z(n31252) );
  XNOR U31226 ( .A(n31253), .B(n31254), .Z(n31043) );
  AND U31227 ( .A(n646), .B(n31255), .Z(n31254) );
  XNOR U31228 ( .A(n31256), .B(n31253), .Z(n31255) );
  XOR U31229 ( .A(n30970), .B(n31249), .Z(n31251) );
  XOR U31230 ( .A(n31257), .B(n31258), .Z(n30970) );
  AND U31231 ( .A(n654), .B(n31259), .Z(n31258) );
  XOR U31232 ( .A(n31219), .B(n31260), .Z(n31249) );
  AND U31233 ( .A(n31261), .B(n31222), .Z(n31260) );
  XNOR U31234 ( .A(n31089), .B(n31219), .Z(n31222) );
  XNOR U31235 ( .A(n31262), .B(n31263), .Z(n31089) );
  AND U31236 ( .A(n646), .B(n31264), .Z(n31263) );
  XOR U31237 ( .A(n31265), .B(n31262), .Z(n31264) );
  XNOR U31238 ( .A(n31266), .B(n31219), .Z(n31261) );
  IV U31239 ( .A(n30980), .Z(n31266) );
  XOR U31240 ( .A(n31267), .B(n31268), .Z(n30980) );
  AND U31241 ( .A(n654), .B(n31269), .Z(n31268) );
  XOR U31242 ( .A(n31270), .B(n31271), .Z(n31219) );
  AND U31243 ( .A(n31272), .B(n31273), .Z(n31271) );
  XNOR U31244 ( .A(n31270), .B(n31183), .Z(n31273) );
  XNOR U31245 ( .A(n31274), .B(n31275), .Z(n31183) );
  AND U31246 ( .A(n646), .B(n31276), .Z(n31275) );
  XNOR U31247 ( .A(n31277), .B(n31274), .Z(n31276) );
  XNOR U31248 ( .A(n31278), .B(n31270), .Z(n31272) );
  IV U31249 ( .A(n30992), .Z(n31278) );
  XOR U31250 ( .A(n31279), .B(n31280), .Z(n30992) );
  AND U31251 ( .A(n654), .B(n31281), .Z(n31280) );
  AND U31252 ( .A(n31223), .B(n31204), .Z(n31270) );
  XNOR U31253 ( .A(n31282), .B(n31283), .Z(n31204) );
  AND U31254 ( .A(n646), .B(n31284), .Z(n31283) );
  XNOR U31255 ( .A(n31285), .B(n31282), .Z(n31284) );
  XNOR U31256 ( .A(n31286), .B(n31287), .Z(n646) );
  AND U31257 ( .A(n31288), .B(n31289), .Z(n31287) );
  XOR U31258 ( .A(n31233), .B(n31286), .Z(n31289) );
  AND U31259 ( .A(n31290), .B(n31291), .Z(n31233) );
  XOR U31260 ( .A(n31286), .B(n31230), .Z(n31288) );
  XNOR U31261 ( .A(n31292), .B(n31293), .Z(n31230) );
  AND U31262 ( .A(n650), .B(n31236), .Z(n31293) );
  XOR U31263 ( .A(n31234), .B(n31292), .Z(n31236) );
  XOR U31264 ( .A(n31294), .B(n31295), .Z(n31286) );
  AND U31265 ( .A(n31296), .B(n31297), .Z(n31295) );
  XNOR U31266 ( .A(n31294), .B(n31290), .Z(n31297) );
  IV U31267 ( .A(n31244), .Z(n31290) );
  XOR U31268 ( .A(n31298), .B(n31299), .Z(n31244) );
  XOR U31269 ( .A(n31300), .B(n31291), .Z(n31299) );
  AND U31270 ( .A(n31256), .B(n31301), .Z(n31291) );
  AND U31271 ( .A(n31302), .B(n31303), .Z(n31300) );
  XOR U31272 ( .A(n31304), .B(n31298), .Z(n31302) );
  XNOR U31273 ( .A(n31241), .B(n31294), .Z(n31296) );
  XNOR U31274 ( .A(n31305), .B(n31306), .Z(n31241) );
  AND U31275 ( .A(n650), .B(n31248), .Z(n31306) );
  XOR U31276 ( .A(n31305), .B(n31246), .Z(n31248) );
  XOR U31277 ( .A(n31307), .B(n31308), .Z(n31294) );
  AND U31278 ( .A(n31309), .B(n31310), .Z(n31308) );
  XNOR U31279 ( .A(n31307), .B(n31256), .Z(n31310) );
  XOR U31280 ( .A(n31311), .B(n31303), .Z(n31256) );
  XNOR U31281 ( .A(n31312), .B(n31298), .Z(n31303) );
  XOR U31282 ( .A(n31313), .B(n31314), .Z(n31298) );
  AND U31283 ( .A(n31315), .B(n31316), .Z(n31314) );
  XOR U31284 ( .A(n31317), .B(n31313), .Z(n31315) );
  XNOR U31285 ( .A(n31318), .B(n31319), .Z(n31312) );
  AND U31286 ( .A(n31320), .B(n31321), .Z(n31319) );
  XOR U31287 ( .A(n31318), .B(n31322), .Z(n31320) );
  XNOR U31288 ( .A(n31304), .B(n31301), .Z(n31311) );
  AND U31289 ( .A(n31323), .B(n31324), .Z(n31301) );
  XOR U31290 ( .A(n31325), .B(n31326), .Z(n31304) );
  AND U31291 ( .A(n31327), .B(n31328), .Z(n31326) );
  XOR U31292 ( .A(n31325), .B(n31329), .Z(n31327) );
  XNOR U31293 ( .A(n31253), .B(n31307), .Z(n31309) );
  XNOR U31294 ( .A(n31330), .B(n31331), .Z(n31253) );
  AND U31295 ( .A(n650), .B(n31259), .Z(n31331) );
  XOR U31296 ( .A(n31330), .B(n31257), .Z(n31259) );
  XOR U31297 ( .A(n31332), .B(n31333), .Z(n31307) );
  AND U31298 ( .A(n31334), .B(n31335), .Z(n31333) );
  XNOR U31299 ( .A(n31332), .B(n31323), .Z(n31335) );
  IV U31300 ( .A(n31265), .Z(n31323) );
  XNOR U31301 ( .A(n31336), .B(n31316), .Z(n31265) );
  XNOR U31302 ( .A(n31337), .B(n31322), .Z(n31316) );
  XOR U31303 ( .A(n31338), .B(n31339), .Z(n31322) );
  AND U31304 ( .A(n31340), .B(n31341), .Z(n31339) );
  XOR U31305 ( .A(n31338), .B(n31342), .Z(n31340) );
  XNOR U31306 ( .A(n31321), .B(n31313), .Z(n31337) );
  XOR U31307 ( .A(n31343), .B(n31344), .Z(n31313) );
  AND U31308 ( .A(n31345), .B(n31346), .Z(n31344) );
  XNOR U31309 ( .A(n31347), .B(n31343), .Z(n31345) );
  XNOR U31310 ( .A(n31348), .B(n31318), .Z(n31321) );
  XOR U31311 ( .A(n31349), .B(n31350), .Z(n31318) );
  AND U31312 ( .A(n31351), .B(n31352), .Z(n31350) );
  XOR U31313 ( .A(n31349), .B(n31353), .Z(n31351) );
  XNOR U31314 ( .A(n31354), .B(n31355), .Z(n31348) );
  AND U31315 ( .A(n31356), .B(n31357), .Z(n31355) );
  XNOR U31316 ( .A(n31354), .B(n31358), .Z(n31356) );
  XNOR U31317 ( .A(n31317), .B(n31324), .Z(n31336) );
  AND U31318 ( .A(n31277), .B(n31359), .Z(n31324) );
  XOR U31319 ( .A(n31329), .B(n31328), .Z(n31317) );
  XNOR U31320 ( .A(n31360), .B(n31325), .Z(n31328) );
  XOR U31321 ( .A(n31361), .B(n31362), .Z(n31325) );
  AND U31322 ( .A(n31363), .B(n31364), .Z(n31362) );
  XOR U31323 ( .A(n31361), .B(n31365), .Z(n31363) );
  XNOR U31324 ( .A(n31366), .B(n31367), .Z(n31360) );
  AND U31325 ( .A(n31368), .B(n31369), .Z(n31367) );
  XOR U31326 ( .A(n31366), .B(n31370), .Z(n31368) );
  XOR U31327 ( .A(n31371), .B(n31372), .Z(n31329) );
  AND U31328 ( .A(n31373), .B(n31374), .Z(n31372) );
  XOR U31329 ( .A(n31371), .B(n31375), .Z(n31373) );
  XNOR U31330 ( .A(n31262), .B(n31332), .Z(n31334) );
  XNOR U31331 ( .A(n31376), .B(n31377), .Z(n31262) );
  AND U31332 ( .A(n650), .B(n31269), .Z(n31377) );
  XOR U31333 ( .A(n31376), .B(n31267), .Z(n31269) );
  XOR U31334 ( .A(n31378), .B(n31379), .Z(n31332) );
  AND U31335 ( .A(n31380), .B(n31381), .Z(n31379) );
  XNOR U31336 ( .A(n31378), .B(n31277), .Z(n31381) );
  XOR U31337 ( .A(n31382), .B(n31346), .Z(n31277) );
  XNOR U31338 ( .A(n31383), .B(n31353), .Z(n31346) );
  XOR U31339 ( .A(n31342), .B(n31341), .Z(n31353) );
  XNOR U31340 ( .A(n31384), .B(n31338), .Z(n31341) );
  XOR U31341 ( .A(n31385), .B(n31386), .Z(n31338) );
  AND U31342 ( .A(n31387), .B(n31388), .Z(n31386) );
  XNOR U31343 ( .A(n31389), .B(n31390), .Z(n31387) );
  IV U31344 ( .A(n31385), .Z(n31389) );
  XNOR U31345 ( .A(n31391), .B(n31392), .Z(n31384) );
  NOR U31346 ( .A(n31393), .B(n31394), .Z(n31392) );
  XNOR U31347 ( .A(n31391), .B(n31395), .Z(n31393) );
  XOR U31348 ( .A(n31396), .B(n31397), .Z(n31342) );
  NOR U31349 ( .A(n31398), .B(n31399), .Z(n31397) );
  XNOR U31350 ( .A(n31396), .B(n31400), .Z(n31398) );
  XNOR U31351 ( .A(n31352), .B(n31343), .Z(n31383) );
  XOR U31352 ( .A(n31401), .B(n31402), .Z(n31343) );
  AND U31353 ( .A(n31403), .B(n31404), .Z(n31402) );
  XOR U31354 ( .A(n31401), .B(n31405), .Z(n31403) );
  XOR U31355 ( .A(n31406), .B(n31358), .Z(n31352) );
  XOR U31356 ( .A(n31407), .B(n31408), .Z(n31358) );
  NOR U31357 ( .A(n31409), .B(n31410), .Z(n31408) );
  XOR U31358 ( .A(n31407), .B(n31411), .Z(n31409) );
  XNOR U31359 ( .A(n31357), .B(n31349), .Z(n31406) );
  XOR U31360 ( .A(n31412), .B(n31413), .Z(n31349) );
  AND U31361 ( .A(n31414), .B(n31415), .Z(n31413) );
  XOR U31362 ( .A(n31412), .B(n31416), .Z(n31414) );
  XNOR U31363 ( .A(n31417), .B(n31354), .Z(n31357) );
  XOR U31364 ( .A(n31418), .B(n31419), .Z(n31354) );
  AND U31365 ( .A(n31420), .B(n31421), .Z(n31419) );
  XNOR U31366 ( .A(n31422), .B(n31423), .Z(n31420) );
  IV U31367 ( .A(n31418), .Z(n31422) );
  XNOR U31368 ( .A(n31424), .B(n31425), .Z(n31417) );
  NOR U31369 ( .A(n31426), .B(n31427), .Z(n31425) );
  XNOR U31370 ( .A(n31424), .B(n31428), .Z(n31426) );
  XOR U31371 ( .A(n31347), .B(n31359), .Z(n31382) );
  NOR U31372 ( .A(n31285), .B(n31429), .Z(n31359) );
  XNOR U31373 ( .A(n31365), .B(n31364), .Z(n31347) );
  XNOR U31374 ( .A(n31430), .B(n31370), .Z(n31364) );
  XNOR U31375 ( .A(n31431), .B(n31432), .Z(n31370) );
  NOR U31376 ( .A(n31433), .B(n31434), .Z(n31432) );
  XOR U31377 ( .A(n31431), .B(n31435), .Z(n31433) );
  XNOR U31378 ( .A(n31369), .B(n31361), .Z(n31430) );
  XOR U31379 ( .A(n31436), .B(n31437), .Z(n31361) );
  AND U31380 ( .A(n31438), .B(n31439), .Z(n31437) );
  XOR U31381 ( .A(n31436), .B(n31440), .Z(n31438) );
  XNOR U31382 ( .A(n31441), .B(n31366), .Z(n31369) );
  XOR U31383 ( .A(n31442), .B(n31443), .Z(n31366) );
  AND U31384 ( .A(n31444), .B(n31445), .Z(n31443) );
  XNOR U31385 ( .A(n31446), .B(n31447), .Z(n31444) );
  IV U31386 ( .A(n31442), .Z(n31446) );
  XNOR U31387 ( .A(n31448), .B(n31449), .Z(n31441) );
  NOR U31388 ( .A(n31450), .B(n31451), .Z(n31449) );
  XNOR U31389 ( .A(n31448), .B(n31452), .Z(n31450) );
  XOR U31390 ( .A(n31375), .B(n31374), .Z(n31365) );
  XNOR U31391 ( .A(n31453), .B(n31371), .Z(n31374) );
  XOR U31392 ( .A(n31454), .B(n31455), .Z(n31371) );
  AND U31393 ( .A(n31456), .B(n31457), .Z(n31455) );
  XNOR U31394 ( .A(n31458), .B(n31459), .Z(n31456) );
  IV U31395 ( .A(n31454), .Z(n31458) );
  XNOR U31396 ( .A(n31460), .B(n31461), .Z(n31453) );
  NOR U31397 ( .A(n31462), .B(n31463), .Z(n31461) );
  XNOR U31398 ( .A(n31460), .B(n31464), .Z(n31462) );
  XOR U31399 ( .A(n31465), .B(n31466), .Z(n31375) );
  NOR U31400 ( .A(n31467), .B(n31468), .Z(n31466) );
  XNOR U31401 ( .A(n31465), .B(n31469), .Z(n31467) );
  XNOR U31402 ( .A(n31274), .B(n31378), .Z(n31380) );
  XNOR U31403 ( .A(n31470), .B(n31471), .Z(n31274) );
  AND U31404 ( .A(n650), .B(n31281), .Z(n31471) );
  XOR U31405 ( .A(n31470), .B(n31279), .Z(n31281) );
  AND U31406 ( .A(n31282), .B(n31285), .Z(n31378) );
  XOR U31407 ( .A(n31472), .B(n31429), .Z(n31285) );
  XNOR U31408 ( .A(p_input[1696]), .B(p_input[2048]), .Z(n31429) );
  XNOR U31409 ( .A(n31405), .B(n31404), .Z(n31472) );
  XNOR U31410 ( .A(n31473), .B(n31416), .Z(n31404) );
  XOR U31411 ( .A(n31390), .B(n31388), .Z(n31416) );
  XNOR U31412 ( .A(n31474), .B(n31395), .Z(n31388) );
  XOR U31413 ( .A(p_input[1720]), .B(p_input[2072]), .Z(n31395) );
  XOR U31414 ( .A(n31385), .B(n31394), .Z(n31474) );
  XOR U31415 ( .A(n31475), .B(n31391), .Z(n31394) );
  XOR U31416 ( .A(p_input[1718]), .B(p_input[2070]), .Z(n31391) );
  XOR U31417 ( .A(p_input[1719]), .B(n17295), .Z(n31475) );
  XOR U31418 ( .A(p_input[1714]), .B(p_input[2066]), .Z(n31385) );
  XNOR U31419 ( .A(n31400), .B(n31399), .Z(n31390) );
  XOR U31420 ( .A(n31476), .B(n31396), .Z(n31399) );
  XOR U31421 ( .A(p_input[1715]), .B(p_input[2067]), .Z(n31396) );
  XOR U31422 ( .A(p_input[1716]), .B(n17297), .Z(n31476) );
  XOR U31423 ( .A(p_input[1717]), .B(p_input[2069]), .Z(n31400) );
  XOR U31424 ( .A(n31415), .B(n31477), .Z(n31473) );
  IV U31425 ( .A(n31401), .Z(n31477) );
  XOR U31426 ( .A(p_input[1697]), .B(p_input[2049]), .Z(n31401) );
  XNOR U31427 ( .A(n31478), .B(n31423), .Z(n31415) );
  XNOR U31428 ( .A(n31411), .B(n31410), .Z(n31423) );
  XNOR U31429 ( .A(n31479), .B(n31407), .Z(n31410) );
  XNOR U31430 ( .A(p_input[1722]), .B(p_input[2074]), .Z(n31407) );
  XOR U31431 ( .A(p_input[1723]), .B(n17300), .Z(n31479) );
  XOR U31432 ( .A(p_input[1724]), .B(p_input[2076]), .Z(n31411) );
  XOR U31433 ( .A(n31421), .B(n31480), .Z(n31478) );
  IV U31434 ( .A(n31412), .Z(n31480) );
  XOR U31435 ( .A(p_input[1713]), .B(p_input[2065]), .Z(n31412) );
  XNOR U31436 ( .A(n31481), .B(n31428), .Z(n31421) );
  XNOR U31437 ( .A(p_input[1727]), .B(n17303), .Z(n31428) );
  XOR U31438 ( .A(n31418), .B(n31427), .Z(n31481) );
  XOR U31439 ( .A(n31482), .B(n31424), .Z(n31427) );
  XOR U31440 ( .A(p_input[1725]), .B(p_input[2077]), .Z(n31424) );
  XOR U31441 ( .A(p_input[1726]), .B(n17305), .Z(n31482) );
  XOR U31442 ( .A(p_input[1721]), .B(p_input[2073]), .Z(n31418) );
  XOR U31443 ( .A(n31440), .B(n31439), .Z(n31405) );
  XNOR U31444 ( .A(n31483), .B(n31447), .Z(n31439) );
  XNOR U31445 ( .A(n31435), .B(n31434), .Z(n31447) );
  XNOR U31446 ( .A(n31484), .B(n31431), .Z(n31434) );
  XNOR U31447 ( .A(p_input[1707]), .B(p_input[2059]), .Z(n31431) );
  XOR U31448 ( .A(p_input[1708]), .B(n16451), .Z(n31484) );
  XOR U31449 ( .A(p_input[1709]), .B(p_input[2061]), .Z(n31435) );
  XOR U31450 ( .A(n31445), .B(n31485), .Z(n31483) );
  IV U31451 ( .A(n31436), .Z(n31485) );
  XOR U31452 ( .A(p_input[1698]), .B(p_input[2050]), .Z(n31436) );
  XNOR U31453 ( .A(n31486), .B(n31452), .Z(n31445) );
  XNOR U31454 ( .A(p_input[1712]), .B(n16454), .Z(n31452) );
  XOR U31455 ( .A(n31442), .B(n31451), .Z(n31486) );
  XOR U31456 ( .A(n31487), .B(n31448), .Z(n31451) );
  XOR U31457 ( .A(p_input[1710]), .B(p_input[2062]), .Z(n31448) );
  XOR U31458 ( .A(p_input[1711]), .B(n16456), .Z(n31487) );
  XOR U31459 ( .A(p_input[1706]), .B(p_input[2058]), .Z(n31442) );
  XOR U31460 ( .A(n31459), .B(n31457), .Z(n31440) );
  XNOR U31461 ( .A(n31488), .B(n31464), .Z(n31457) );
  XOR U31462 ( .A(p_input[1705]), .B(p_input[2057]), .Z(n31464) );
  XOR U31463 ( .A(n31454), .B(n31463), .Z(n31488) );
  XOR U31464 ( .A(n31489), .B(n31460), .Z(n31463) );
  XOR U31465 ( .A(p_input[1703]), .B(p_input[2055]), .Z(n31460) );
  XOR U31466 ( .A(p_input[1704]), .B(n17312), .Z(n31489) );
  XOR U31467 ( .A(p_input[1699]), .B(p_input[2051]), .Z(n31454) );
  XNOR U31468 ( .A(n31469), .B(n31468), .Z(n31459) );
  XOR U31469 ( .A(n31490), .B(n31465), .Z(n31468) );
  XOR U31470 ( .A(p_input[1700]), .B(p_input[2052]), .Z(n31465) );
  XOR U31471 ( .A(p_input[1701]), .B(n17314), .Z(n31490) );
  XOR U31472 ( .A(p_input[1702]), .B(p_input[2054]), .Z(n31469) );
  XNOR U31473 ( .A(n31491), .B(n31492), .Z(n31282) );
  AND U31474 ( .A(n650), .B(n31493), .Z(n31492) );
  XNOR U31475 ( .A(n31494), .B(n31495), .Z(n650) );
  AND U31476 ( .A(n31496), .B(n31497), .Z(n31495) );
  XOR U31477 ( .A(n31494), .B(n31292), .Z(n31497) );
  XNOR U31478 ( .A(n31494), .B(n31234), .Z(n31496) );
  XOR U31479 ( .A(n31498), .B(n31499), .Z(n31494) );
  AND U31480 ( .A(n31500), .B(n31501), .Z(n31499) );
  XNOR U31481 ( .A(n31305), .B(n31498), .Z(n31501) );
  XOR U31482 ( .A(n31498), .B(n31246), .Z(n31500) );
  XOR U31483 ( .A(n31502), .B(n31503), .Z(n31498) );
  AND U31484 ( .A(n31504), .B(n31505), .Z(n31503) );
  XNOR U31485 ( .A(n31330), .B(n31502), .Z(n31505) );
  XOR U31486 ( .A(n31502), .B(n31257), .Z(n31504) );
  XOR U31487 ( .A(n31506), .B(n31507), .Z(n31502) );
  AND U31488 ( .A(n31508), .B(n31509), .Z(n31507) );
  XOR U31489 ( .A(n31506), .B(n31267), .Z(n31508) );
  XOR U31490 ( .A(n31510), .B(n31511), .Z(n31223) );
  AND U31491 ( .A(n654), .B(n31493), .Z(n31511) );
  XNOR U31492 ( .A(n31491), .B(n31510), .Z(n31493) );
  XNOR U31493 ( .A(n31512), .B(n31513), .Z(n654) );
  AND U31494 ( .A(n31514), .B(n31515), .Z(n31513) );
  XNOR U31495 ( .A(n31516), .B(n31512), .Z(n31515) );
  IV U31496 ( .A(n31292), .Z(n31516) );
  XNOR U31497 ( .A(n31517), .B(n31518), .Z(n31292) );
  AND U31498 ( .A(n657), .B(n31519), .Z(n31518) );
  XNOR U31499 ( .A(n31517), .B(n31520), .Z(n31519) );
  XNOR U31500 ( .A(n31234), .B(n31512), .Z(n31514) );
  XOR U31501 ( .A(n31521), .B(n31522), .Z(n31234) );
  AND U31502 ( .A(n665), .B(n31523), .Z(n31522) );
  XOR U31503 ( .A(n31524), .B(n31525), .Z(n31512) );
  AND U31504 ( .A(n31526), .B(n31527), .Z(n31525) );
  XNOR U31505 ( .A(n31524), .B(n31305), .Z(n31527) );
  XNOR U31506 ( .A(n31528), .B(n31529), .Z(n31305) );
  AND U31507 ( .A(n657), .B(n31530), .Z(n31529) );
  XOR U31508 ( .A(n31531), .B(n31528), .Z(n31530) );
  XNOR U31509 ( .A(n31532), .B(n31524), .Z(n31526) );
  IV U31510 ( .A(n31246), .Z(n31532) );
  XOR U31511 ( .A(n31533), .B(n31534), .Z(n31246) );
  AND U31512 ( .A(n665), .B(n31535), .Z(n31534) );
  XOR U31513 ( .A(n31536), .B(n31537), .Z(n31524) );
  AND U31514 ( .A(n31538), .B(n31539), .Z(n31537) );
  XNOR U31515 ( .A(n31536), .B(n31330), .Z(n31539) );
  XNOR U31516 ( .A(n31540), .B(n31541), .Z(n31330) );
  AND U31517 ( .A(n657), .B(n31542), .Z(n31541) );
  XNOR U31518 ( .A(n31543), .B(n31540), .Z(n31542) );
  XOR U31519 ( .A(n31257), .B(n31536), .Z(n31538) );
  XOR U31520 ( .A(n31544), .B(n31545), .Z(n31257) );
  AND U31521 ( .A(n665), .B(n31546), .Z(n31545) );
  XOR U31522 ( .A(n31506), .B(n31547), .Z(n31536) );
  AND U31523 ( .A(n31548), .B(n31509), .Z(n31547) );
  XNOR U31524 ( .A(n31376), .B(n31506), .Z(n31509) );
  XNOR U31525 ( .A(n31549), .B(n31550), .Z(n31376) );
  AND U31526 ( .A(n657), .B(n31551), .Z(n31550) );
  XOR U31527 ( .A(n31552), .B(n31549), .Z(n31551) );
  XNOR U31528 ( .A(n31553), .B(n31506), .Z(n31548) );
  IV U31529 ( .A(n31267), .Z(n31553) );
  XOR U31530 ( .A(n31554), .B(n31555), .Z(n31267) );
  AND U31531 ( .A(n665), .B(n31556), .Z(n31555) );
  XOR U31532 ( .A(n31557), .B(n31558), .Z(n31506) );
  AND U31533 ( .A(n31559), .B(n31560), .Z(n31558) );
  XNOR U31534 ( .A(n31557), .B(n31470), .Z(n31560) );
  XNOR U31535 ( .A(n31561), .B(n31562), .Z(n31470) );
  AND U31536 ( .A(n657), .B(n31563), .Z(n31562) );
  XNOR U31537 ( .A(n31564), .B(n31561), .Z(n31563) );
  XNOR U31538 ( .A(n31565), .B(n31557), .Z(n31559) );
  IV U31539 ( .A(n31279), .Z(n31565) );
  XOR U31540 ( .A(n31566), .B(n31567), .Z(n31279) );
  AND U31541 ( .A(n665), .B(n31568), .Z(n31567) );
  AND U31542 ( .A(n31510), .B(n31491), .Z(n31557) );
  XNOR U31543 ( .A(n31569), .B(n31570), .Z(n31491) );
  AND U31544 ( .A(n657), .B(n31571), .Z(n31570) );
  XNOR U31545 ( .A(n31572), .B(n31569), .Z(n31571) );
  XNOR U31546 ( .A(n31573), .B(n31574), .Z(n657) );
  AND U31547 ( .A(n31575), .B(n31576), .Z(n31574) );
  XOR U31548 ( .A(n31520), .B(n31573), .Z(n31576) );
  AND U31549 ( .A(n31577), .B(n31578), .Z(n31520) );
  XOR U31550 ( .A(n31573), .B(n31517), .Z(n31575) );
  XNOR U31551 ( .A(n31579), .B(n31580), .Z(n31517) );
  AND U31552 ( .A(n661), .B(n31523), .Z(n31580) );
  XOR U31553 ( .A(n31521), .B(n31579), .Z(n31523) );
  XOR U31554 ( .A(n31581), .B(n31582), .Z(n31573) );
  AND U31555 ( .A(n31583), .B(n31584), .Z(n31582) );
  XNOR U31556 ( .A(n31581), .B(n31577), .Z(n31584) );
  IV U31557 ( .A(n31531), .Z(n31577) );
  XOR U31558 ( .A(n31585), .B(n31586), .Z(n31531) );
  XOR U31559 ( .A(n31587), .B(n31578), .Z(n31586) );
  AND U31560 ( .A(n31543), .B(n31588), .Z(n31578) );
  AND U31561 ( .A(n31589), .B(n31590), .Z(n31587) );
  XOR U31562 ( .A(n31591), .B(n31585), .Z(n31589) );
  XNOR U31563 ( .A(n31528), .B(n31581), .Z(n31583) );
  XNOR U31564 ( .A(n31592), .B(n31593), .Z(n31528) );
  AND U31565 ( .A(n661), .B(n31535), .Z(n31593) );
  XOR U31566 ( .A(n31592), .B(n31533), .Z(n31535) );
  XOR U31567 ( .A(n31594), .B(n31595), .Z(n31581) );
  AND U31568 ( .A(n31596), .B(n31597), .Z(n31595) );
  XNOR U31569 ( .A(n31594), .B(n31543), .Z(n31597) );
  XOR U31570 ( .A(n31598), .B(n31590), .Z(n31543) );
  XNOR U31571 ( .A(n31599), .B(n31585), .Z(n31590) );
  XOR U31572 ( .A(n31600), .B(n31601), .Z(n31585) );
  AND U31573 ( .A(n31602), .B(n31603), .Z(n31601) );
  XOR U31574 ( .A(n31604), .B(n31600), .Z(n31602) );
  XNOR U31575 ( .A(n31605), .B(n31606), .Z(n31599) );
  AND U31576 ( .A(n31607), .B(n31608), .Z(n31606) );
  XOR U31577 ( .A(n31605), .B(n31609), .Z(n31607) );
  XNOR U31578 ( .A(n31591), .B(n31588), .Z(n31598) );
  AND U31579 ( .A(n31610), .B(n31611), .Z(n31588) );
  XOR U31580 ( .A(n31612), .B(n31613), .Z(n31591) );
  AND U31581 ( .A(n31614), .B(n31615), .Z(n31613) );
  XOR U31582 ( .A(n31612), .B(n31616), .Z(n31614) );
  XNOR U31583 ( .A(n31540), .B(n31594), .Z(n31596) );
  XNOR U31584 ( .A(n31617), .B(n31618), .Z(n31540) );
  AND U31585 ( .A(n661), .B(n31546), .Z(n31618) );
  XOR U31586 ( .A(n31617), .B(n31544), .Z(n31546) );
  XOR U31587 ( .A(n31619), .B(n31620), .Z(n31594) );
  AND U31588 ( .A(n31621), .B(n31622), .Z(n31620) );
  XNOR U31589 ( .A(n31619), .B(n31610), .Z(n31622) );
  IV U31590 ( .A(n31552), .Z(n31610) );
  XNOR U31591 ( .A(n31623), .B(n31603), .Z(n31552) );
  XNOR U31592 ( .A(n31624), .B(n31609), .Z(n31603) );
  XOR U31593 ( .A(n31625), .B(n31626), .Z(n31609) );
  AND U31594 ( .A(n31627), .B(n31628), .Z(n31626) );
  XOR U31595 ( .A(n31625), .B(n31629), .Z(n31627) );
  XNOR U31596 ( .A(n31608), .B(n31600), .Z(n31624) );
  XOR U31597 ( .A(n31630), .B(n31631), .Z(n31600) );
  AND U31598 ( .A(n31632), .B(n31633), .Z(n31631) );
  XNOR U31599 ( .A(n31634), .B(n31630), .Z(n31632) );
  XNOR U31600 ( .A(n31635), .B(n31605), .Z(n31608) );
  XOR U31601 ( .A(n31636), .B(n31637), .Z(n31605) );
  AND U31602 ( .A(n31638), .B(n31639), .Z(n31637) );
  XOR U31603 ( .A(n31636), .B(n31640), .Z(n31638) );
  XNOR U31604 ( .A(n31641), .B(n31642), .Z(n31635) );
  AND U31605 ( .A(n31643), .B(n31644), .Z(n31642) );
  XNOR U31606 ( .A(n31641), .B(n31645), .Z(n31643) );
  XNOR U31607 ( .A(n31604), .B(n31611), .Z(n31623) );
  AND U31608 ( .A(n31564), .B(n31646), .Z(n31611) );
  XOR U31609 ( .A(n31616), .B(n31615), .Z(n31604) );
  XNOR U31610 ( .A(n31647), .B(n31612), .Z(n31615) );
  XOR U31611 ( .A(n31648), .B(n31649), .Z(n31612) );
  AND U31612 ( .A(n31650), .B(n31651), .Z(n31649) );
  XOR U31613 ( .A(n31648), .B(n31652), .Z(n31650) );
  XNOR U31614 ( .A(n31653), .B(n31654), .Z(n31647) );
  AND U31615 ( .A(n31655), .B(n31656), .Z(n31654) );
  XOR U31616 ( .A(n31653), .B(n31657), .Z(n31655) );
  XOR U31617 ( .A(n31658), .B(n31659), .Z(n31616) );
  AND U31618 ( .A(n31660), .B(n31661), .Z(n31659) );
  XOR U31619 ( .A(n31658), .B(n31662), .Z(n31660) );
  XNOR U31620 ( .A(n31549), .B(n31619), .Z(n31621) );
  XNOR U31621 ( .A(n31663), .B(n31664), .Z(n31549) );
  AND U31622 ( .A(n661), .B(n31556), .Z(n31664) );
  XOR U31623 ( .A(n31663), .B(n31554), .Z(n31556) );
  XOR U31624 ( .A(n31665), .B(n31666), .Z(n31619) );
  AND U31625 ( .A(n31667), .B(n31668), .Z(n31666) );
  XNOR U31626 ( .A(n31665), .B(n31564), .Z(n31668) );
  XOR U31627 ( .A(n31669), .B(n31633), .Z(n31564) );
  XNOR U31628 ( .A(n31670), .B(n31640), .Z(n31633) );
  XOR U31629 ( .A(n31629), .B(n31628), .Z(n31640) );
  XNOR U31630 ( .A(n31671), .B(n31625), .Z(n31628) );
  XOR U31631 ( .A(n31672), .B(n31673), .Z(n31625) );
  AND U31632 ( .A(n31674), .B(n31675), .Z(n31673) );
  XNOR U31633 ( .A(n31676), .B(n31677), .Z(n31674) );
  IV U31634 ( .A(n31672), .Z(n31676) );
  XNOR U31635 ( .A(n31678), .B(n31679), .Z(n31671) );
  NOR U31636 ( .A(n31680), .B(n31681), .Z(n31679) );
  XNOR U31637 ( .A(n31678), .B(n31682), .Z(n31680) );
  XOR U31638 ( .A(n31683), .B(n31684), .Z(n31629) );
  NOR U31639 ( .A(n31685), .B(n31686), .Z(n31684) );
  XNOR U31640 ( .A(n31683), .B(n31687), .Z(n31685) );
  XNOR U31641 ( .A(n31639), .B(n31630), .Z(n31670) );
  XOR U31642 ( .A(n31688), .B(n31689), .Z(n31630) );
  AND U31643 ( .A(n31690), .B(n31691), .Z(n31689) );
  XOR U31644 ( .A(n31688), .B(n31692), .Z(n31690) );
  XOR U31645 ( .A(n31693), .B(n31645), .Z(n31639) );
  XOR U31646 ( .A(n31694), .B(n31695), .Z(n31645) );
  NOR U31647 ( .A(n31696), .B(n31697), .Z(n31695) );
  XOR U31648 ( .A(n31694), .B(n31698), .Z(n31696) );
  XNOR U31649 ( .A(n31644), .B(n31636), .Z(n31693) );
  XOR U31650 ( .A(n31699), .B(n31700), .Z(n31636) );
  AND U31651 ( .A(n31701), .B(n31702), .Z(n31700) );
  XOR U31652 ( .A(n31699), .B(n31703), .Z(n31701) );
  XNOR U31653 ( .A(n31704), .B(n31641), .Z(n31644) );
  XOR U31654 ( .A(n31705), .B(n31706), .Z(n31641) );
  AND U31655 ( .A(n31707), .B(n31708), .Z(n31706) );
  XNOR U31656 ( .A(n31709), .B(n31710), .Z(n31707) );
  IV U31657 ( .A(n31705), .Z(n31709) );
  XNOR U31658 ( .A(n31711), .B(n31712), .Z(n31704) );
  NOR U31659 ( .A(n31713), .B(n31714), .Z(n31712) );
  XNOR U31660 ( .A(n31711), .B(n31715), .Z(n31713) );
  XOR U31661 ( .A(n31634), .B(n31646), .Z(n31669) );
  NOR U31662 ( .A(n31572), .B(n31716), .Z(n31646) );
  XNOR U31663 ( .A(n31652), .B(n31651), .Z(n31634) );
  XNOR U31664 ( .A(n31717), .B(n31657), .Z(n31651) );
  XNOR U31665 ( .A(n31718), .B(n31719), .Z(n31657) );
  NOR U31666 ( .A(n31720), .B(n31721), .Z(n31719) );
  XOR U31667 ( .A(n31718), .B(n31722), .Z(n31720) );
  XNOR U31668 ( .A(n31656), .B(n31648), .Z(n31717) );
  XOR U31669 ( .A(n31723), .B(n31724), .Z(n31648) );
  AND U31670 ( .A(n31725), .B(n31726), .Z(n31724) );
  XOR U31671 ( .A(n31723), .B(n31727), .Z(n31725) );
  XNOR U31672 ( .A(n31728), .B(n31653), .Z(n31656) );
  XOR U31673 ( .A(n31729), .B(n31730), .Z(n31653) );
  AND U31674 ( .A(n31731), .B(n31732), .Z(n31730) );
  XNOR U31675 ( .A(n31733), .B(n31734), .Z(n31731) );
  IV U31676 ( .A(n31729), .Z(n31733) );
  XNOR U31677 ( .A(n31735), .B(n31736), .Z(n31728) );
  NOR U31678 ( .A(n31737), .B(n31738), .Z(n31736) );
  XNOR U31679 ( .A(n31735), .B(n31739), .Z(n31737) );
  XOR U31680 ( .A(n31662), .B(n31661), .Z(n31652) );
  XNOR U31681 ( .A(n31740), .B(n31658), .Z(n31661) );
  XOR U31682 ( .A(n31741), .B(n31742), .Z(n31658) );
  AND U31683 ( .A(n31743), .B(n31744), .Z(n31742) );
  XNOR U31684 ( .A(n31745), .B(n31746), .Z(n31743) );
  IV U31685 ( .A(n31741), .Z(n31745) );
  XNOR U31686 ( .A(n31747), .B(n31748), .Z(n31740) );
  NOR U31687 ( .A(n31749), .B(n31750), .Z(n31748) );
  XNOR U31688 ( .A(n31747), .B(n31751), .Z(n31749) );
  XOR U31689 ( .A(n31752), .B(n31753), .Z(n31662) );
  NOR U31690 ( .A(n31754), .B(n31755), .Z(n31753) );
  XNOR U31691 ( .A(n31752), .B(n31756), .Z(n31754) );
  XNOR U31692 ( .A(n31561), .B(n31665), .Z(n31667) );
  XNOR U31693 ( .A(n31757), .B(n31758), .Z(n31561) );
  AND U31694 ( .A(n661), .B(n31568), .Z(n31758) );
  XOR U31695 ( .A(n31757), .B(n31566), .Z(n31568) );
  AND U31696 ( .A(n31569), .B(n31572), .Z(n31665) );
  XOR U31697 ( .A(n31759), .B(n31716), .Z(n31572) );
  XNOR U31698 ( .A(p_input[1728]), .B(p_input[2048]), .Z(n31716) );
  XNOR U31699 ( .A(n31692), .B(n31691), .Z(n31759) );
  XNOR U31700 ( .A(n31760), .B(n31703), .Z(n31691) );
  XOR U31701 ( .A(n31677), .B(n31675), .Z(n31703) );
  XNOR U31702 ( .A(n31761), .B(n31682), .Z(n31675) );
  XOR U31703 ( .A(p_input[1752]), .B(p_input[2072]), .Z(n31682) );
  XOR U31704 ( .A(n31672), .B(n31681), .Z(n31761) );
  XOR U31705 ( .A(n31762), .B(n31678), .Z(n31681) );
  XOR U31706 ( .A(p_input[1750]), .B(p_input[2070]), .Z(n31678) );
  XOR U31707 ( .A(p_input[1751]), .B(n17295), .Z(n31762) );
  XOR U31708 ( .A(p_input[1746]), .B(p_input[2066]), .Z(n31672) );
  XNOR U31709 ( .A(n31687), .B(n31686), .Z(n31677) );
  XOR U31710 ( .A(n31763), .B(n31683), .Z(n31686) );
  XOR U31711 ( .A(p_input[1747]), .B(p_input[2067]), .Z(n31683) );
  XOR U31712 ( .A(p_input[1748]), .B(n17297), .Z(n31763) );
  XOR U31713 ( .A(p_input[1749]), .B(p_input[2069]), .Z(n31687) );
  XOR U31714 ( .A(n31702), .B(n31764), .Z(n31760) );
  IV U31715 ( .A(n31688), .Z(n31764) );
  XOR U31716 ( .A(p_input[1729]), .B(p_input[2049]), .Z(n31688) );
  XNOR U31717 ( .A(n31765), .B(n31710), .Z(n31702) );
  XNOR U31718 ( .A(n31698), .B(n31697), .Z(n31710) );
  XNOR U31719 ( .A(n31766), .B(n31694), .Z(n31697) );
  XNOR U31720 ( .A(p_input[1754]), .B(p_input[2074]), .Z(n31694) );
  XOR U31721 ( .A(p_input[1755]), .B(n17300), .Z(n31766) );
  XOR U31722 ( .A(p_input[1756]), .B(p_input[2076]), .Z(n31698) );
  XOR U31723 ( .A(n31708), .B(n31767), .Z(n31765) );
  IV U31724 ( .A(n31699), .Z(n31767) );
  XOR U31725 ( .A(p_input[1745]), .B(p_input[2065]), .Z(n31699) );
  XNOR U31726 ( .A(n31768), .B(n31715), .Z(n31708) );
  XNOR U31727 ( .A(p_input[1759]), .B(n17303), .Z(n31715) );
  XOR U31728 ( .A(n31705), .B(n31714), .Z(n31768) );
  XOR U31729 ( .A(n31769), .B(n31711), .Z(n31714) );
  XOR U31730 ( .A(p_input[1757]), .B(p_input[2077]), .Z(n31711) );
  XOR U31731 ( .A(p_input[1758]), .B(n17305), .Z(n31769) );
  XOR U31732 ( .A(p_input[1753]), .B(p_input[2073]), .Z(n31705) );
  XOR U31733 ( .A(n31727), .B(n31726), .Z(n31692) );
  XNOR U31734 ( .A(n31770), .B(n31734), .Z(n31726) );
  XNOR U31735 ( .A(n31722), .B(n31721), .Z(n31734) );
  XNOR U31736 ( .A(n31771), .B(n31718), .Z(n31721) );
  XNOR U31737 ( .A(p_input[1739]), .B(p_input[2059]), .Z(n31718) );
  XOR U31738 ( .A(p_input[1740]), .B(n16451), .Z(n31771) );
  XOR U31739 ( .A(p_input[1741]), .B(p_input[2061]), .Z(n31722) );
  XOR U31740 ( .A(n31732), .B(n31772), .Z(n31770) );
  IV U31741 ( .A(n31723), .Z(n31772) );
  XOR U31742 ( .A(p_input[1730]), .B(p_input[2050]), .Z(n31723) );
  XNOR U31743 ( .A(n31773), .B(n31739), .Z(n31732) );
  XNOR U31744 ( .A(p_input[1744]), .B(n16454), .Z(n31739) );
  XOR U31745 ( .A(n31729), .B(n31738), .Z(n31773) );
  XOR U31746 ( .A(n31774), .B(n31735), .Z(n31738) );
  XOR U31747 ( .A(p_input[1742]), .B(p_input[2062]), .Z(n31735) );
  XOR U31748 ( .A(p_input[1743]), .B(n16456), .Z(n31774) );
  XOR U31749 ( .A(p_input[1738]), .B(p_input[2058]), .Z(n31729) );
  XOR U31750 ( .A(n31746), .B(n31744), .Z(n31727) );
  XNOR U31751 ( .A(n31775), .B(n31751), .Z(n31744) );
  XOR U31752 ( .A(p_input[1737]), .B(p_input[2057]), .Z(n31751) );
  XOR U31753 ( .A(n31741), .B(n31750), .Z(n31775) );
  XOR U31754 ( .A(n31776), .B(n31747), .Z(n31750) );
  XOR U31755 ( .A(p_input[1735]), .B(p_input[2055]), .Z(n31747) );
  XOR U31756 ( .A(p_input[1736]), .B(n17312), .Z(n31776) );
  XOR U31757 ( .A(p_input[1731]), .B(p_input[2051]), .Z(n31741) );
  XNOR U31758 ( .A(n31756), .B(n31755), .Z(n31746) );
  XOR U31759 ( .A(n31777), .B(n31752), .Z(n31755) );
  XOR U31760 ( .A(p_input[1732]), .B(p_input[2052]), .Z(n31752) );
  XOR U31761 ( .A(p_input[1733]), .B(n17314), .Z(n31777) );
  XOR U31762 ( .A(p_input[1734]), .B(p_input[2054]), .Z(n31756) );
  XNOR U31763 ( .A(n31778), .B(n31779), .Z(n31569) );
  AND U31764 ( .A(n661), .B(n31780), .Z(n31779) );
  XNOR U31765 ( .A(n31781), .B(n31782), .Z(n661) );
  AND U31766 ( .A(n31783), .B(n31784), .Z(n31782) );
  XOR U31767 ( .A(n31781), .B(n31579), .Z(n31784) );
  XNOR U31768 ( .A(n31781), .B(n31521), .Z(n31783) );
  XOR U31769 ( .A(n31785), .B(n31786), .Z(n31781) );
  AND U31770 ( .A(n31787), .B(n31788), .Z(n31786) );
  XNOR U31771 ( .A(n31592), .B(n31785), .Z(n31788) );
  XOR U31772 ( .A(n31785), .B(n31533), .Z(n31787) );
  XOR U31773 ( .A(n31789), .B(n31790), .Z(n31785) );
  AND U31774 ( .A(n31791), .B(n31792), .Z(n31790) );
  XNOR U31775 ( .A(n31617), .B(n31789), .Z(n31792) );
  XOR U31776 ( .A(n31789), .B(n31544), .Z(n31791) );
  XOR U31777 ( .A(n31793), .B(n31794), .Z(n31789) );
  AND U31778 ( .A(n31795), .B(n31796), .Z(n31794) );
  XOR U31779 ( .A(n31793), .B(n31554), .Z(n31795) );
  XOR U31780 ( .A(n31797), .B(n31798), .Z(n31510) );
  AND U31781 ( .A(n665), .B(n31780), .Z(n31798) );
  XNOR U31782 ( .A(n31778), .B(n31797), .Z(n31780) );
  XNOR U31783 ( .A(n31799), .B(n31800), .Z(n665) );
  AND U31784 ( .A(n31801), .B(n31802), .Z(n31800) );
  XNOR U31785 ( .A(n31803), .B(n31799), .Z(n31802) );
  IV U31786 ( .A(n31579), .Z(n31803) );
  XNOR U31787 ( .A(n31804), .B(n31805), .Z(n31579) );
  AND U31788 ( .A(n668), .B(n31806), .Z(n31805) );
  XNOR U31789 ( .A(n31804), .B(n31807), .Z(n31806) );
  XNOR U31790 ( .A(n31521), .B(n31799), .Z(n31801) );
  XOR U31791 ( .A(n31808), .B(n31809), .Z(n31521) );
  AND U31792 ( .A(n676), .B(n31810), .Z(n31809) );
  XOR U31793 ( .A(n31811), .B(n31812), .Z(n31799) );
  AND U31794 ( .A(n31813), .B(n31814), .Z(n31812) );
  XNOR U31795 ( .A(n31811), .B(n31592), .Z(n31814) );
  XNOR U31796 ( .A(n31815), .B(n31816), .Z(n31592) );
  AND U31797 ( .A(n668), .B(n31817), .Z(n31816) );
  XOR U31798 ( .A(n31818), .B(n31815), .Z(n31817) );
  XNOR U31799 ( .A(n31819), .B(n31811), .Z(n31813) );
  IV U31800 ( .A(n31533), .Z(n31819) );
  XOR U31801 ( .A(n31820), .B(n31821), .Z(n31533) );
  AND U31802 ( .A(n676), .B(n31822), .Z(n31821) );
  XOR U31803 ( .A(n31823), .B(n31824), .Z(n31811) );
  AND U31804 ( .A(n31825), .B(n31826), .Z(n31824) );
  XNOR U31805 ( .A(n31823), .B(n31617), .Z(n31826) );
  XNOR U31806 ( .A(n31827), .B(n31828), .Z(n31617) );
  AND U31807 ( .A(n668), .B(n31829), .Z(n31828) );
  XNOR U31808 ( .A(n31830), .B(n31827), .Z(n31829) );
  XOR U31809 ( .A(n31544), .B(n31823), .Z(n31825) );
  XOR U31810 ( .A(n31831), .B(n31832), .Z(n31544) );
  AND U31811 ( .A(n676), .B(n31833), .Z(n31832) );
  XOR U31812 ( .A(n31793), .B(n31834), .Z(n31823) );
  AND U31813 ( .A(n31835), .B(n31796), .Z(n31834) );
  XNOR U31814 ( .A(n31663), .B(n31793), .Z(n31796) );
  XNOR U31815 ( .A(n31836), .B(n31837), .Z(n31663) );
  AND U31816 ( .A(n668), .B(n31838), .Z(n31837) );
  XOR U31817 ( .A(n31839), .B(n31836), .Z(n31838) );
  XNOR U31818 ( .A(n31840), .B(n31793), .Z(n31835) );
  IV U31819 ( .A(n31554), .Z(n31840) );
  XOR U31820 ( .A(n31841), .B(n31842), .Z(n31554) );
  AND U31821 ( .A(n676), .B(n31843), .Z(n31842) );
  XOR U31822 ( .A(n31844), .B(n31845), .Z(n31793) );
  AND U31823 ( .A(n31846), .B(n31847), .Z(n31845) );
  XNOR U31824 ( .A(n31844), .B(n31757), .Z(n31847) );
  XNOR U31825 ( .A(n31848), .B(n31849), .Z(n31757) );
  AND U31826 ( .A(n668), .B(n31850), .Z(n31849) );
  XNOR U31827 ( .A(n31851), .B(n31848), .Z(n31850) );
  XNOR U31828 ( .A(n31852), .B(n31844), .Z(n31846) );
  IV U31829 ( .A(n31566), .Z(n31852) );
  XOR U31830 ( .A(n31853), .B(n31854), .Z(n31566) );
  AND U31831 ( .A(n676), .B(n31855), .Z(n31854) );
  AND U31832 ( .A(n31797), .B(n31778), .Z(n31844) );
  XNOR U31833 ( .A(n31856), .B(n31857), .Z(n31778) );
  AND U31834 ( .A(n668), .B(n31858), .Z(n31857) );
  XNOR U31835 ( .A(n31859), .B(n31856), .Z(n31858) );
  XNOR U31836 ( .A(n31860), .B(n31861), .Z(n668) );
  AND U31837 ( .A(n31862), .B(n31863), .Z(n31861) );
  XOR U31838 ( .A(n31807), .B(n31860), .Z(n31863) );
  AND U31839 ( .A(n31864), .B(n31865), .Z(n31807) );
  XOR U31840 ( .A(n31860), .B(n31804), .Z(n31862) );
  XNOR U31841 ( .A(n31866), .B(n31867), .Z(n31804) );
  AND U31842 ( .A(n672), .B(n31810), .Z(n31867) );
  XOR U31843 ( .A(n31808), .B(n31866), .Z(n31810) );
  XOR U31844 ( .A(n31868), .B(n31869), .Z(n31860) );
  AND U31845 ( .A(n31870), .B(n31871), .Z(n31869) );
  XNOR U31846 ( .A(n31868), .B(n31864), .Z(n31871) );
  IV U31847 ( .A(n31818), .Z(n31864) );
  XOR U31848 ( .A(n31872), .B(n31873), .Z(n31818) );
  XOR U31849 ( .A(n31874), .B(n31865), .Z(n31873) );
  AND U31850 ( .A(n31830), .B(n31875), .Z(n31865) );
  AND U31851 ( .A(n31876), .B(n31877), .Z(n31874) );
  XOR U31852 ( .A(n31878), .B(n31872), .Z(n31876) );
  XNOR U31853 ( .A(n31815), .B(n31868), .Z(n31870) );
  XNOR U31854 ( .A(n31879), .B(n31880), .Z(n31815) );
  AND U31855 ( .A(n672), .B(n31822), .Z(n31880) );
  XOR U31856 ( .A(n31879), .B(n31820), .Z(n31822) );
  XOR U31857 ( .A(n31881), .B(n31882), .Z(n31868) );
  AND U31858 ( .A(n31883), .B(n31884), .Z(n31882) );
  XNOR U31859 ( .A(n31881), .B(n31830), .Z(n31884) );
  XOR U31860 ( .A(n31885), .B(n31877), .Z(n31830) );
  XNOR U31861 ( .A(n31886), .B(n31872), .Z(n31877) );
  XOR U31862 ( .A(n31887), .B(n31888), .Z(n31872) );
  AND U31863 ( .A(n31889), .B(n31890), .Z(n31888) );
  XOR U31864 ( .A(n31891), .B(n31887), .Z(n31889) );
  XNOR U31865 ( .A(n31892), .B(n31893), .Z(n31886) );
  AND U31866 ( .A(n31894), .B(n31895), .Z(n31893) );
  XOR U31867 ( .A(n31892), .B(n31896), .Z(n31894) );
  XNOR U31868 ( .A(n31878), .B(n31875), .Z(n31885) );
  AND U31869 ( .A(n31897), .B(n31898), .Z(n31875) );
  XOR U31870 ( .A(n31899), .B(n31900), .Z(n31878) );
  AND U31871 ( .A(n31901), .B(n31902), .Z(n31900) );
  XOR U31872 ( .A(n31899), .B(n31903), .Z(n31901) );
  XNOR U31873 ( .A(n31827), .B(n31881), .Z(n31883) );
  XNOR U31874 ( .A(n31904), .B(n31905), .Z(n31827) );
  AND U31875 ( .A(n672), .B(n31833), .Z(n31905) );
  XOR U31876 ( .A(n31904), .B(n31831), .Z(n31833) );
  XOR U31877 ( .A(n31906), .B(n31907), .Z(n31881) );
  AND U31878 ( .A(n31908), .B(n31909), .Z(n31907) );
  XNOR U31879 ( .A(n31906), .B(n31897), .Z(n31909) );
  IV U31880 ( .A(n31839), .Z(n31897) );
  XNOR U31881 ( .A(n31910), .B(n31890), .Z(n31839) );
  XNOR U31882 ( .A(n31911), .B(n31896), .Z(n31890) );
  XOR U31883 ( .A(n31912), .B(n31913), .Z(n31896) );
  AND U31884 ( .A(n31914), .B(n31915), .Z(n31913) );
  XOR U31885 ( .A(n31912), .B(n31916), .Z(n31914) );
  XNOR U31886 ( .A(n31895), .B(n31887), .Z(n31911) );
  XOR U31887 ( .A(n31917), .B(n31918), .Z(n31887) );
  AND U31888 ( .A(n31919), .B(n31920), .Z(n31918) );
  XNOR U31889 ( .A(n31921), .B(n31917), .Z(n31919) );
  XNOR U31890 ( .A(n31922), .B(n31892), .Z(n31895) );
  XOR U31891 ( .A(n31923), .B(n31924), .Z(n31892) );
  AND U31892 ( .A(n31925), .B(n31926), .Z(n31924) );
  XOR U31893 ( .A(n31923), .B(n31927), .Z(n31925) );
  XNOR U31894 ( .A(n31928), .B(n31929), .Z(n31922) );
  AND U31895 ( .A(n31930), .B(n31931), .Z(n31929) );
  XNOR U31896 ( .A(n31928), .B(n31932), .Z(n31930) );
  XNOR U31897 ( .A(n31891), .B(n31898), .Z(n31910) );
  AND U31898 ( .A(n31851), .B(n31933), .Z(n31898) );
  XOR U31899 ( .A(n31903), .B(n31902), .Z(n31891) );
  XNOR U31900 ( .A(n31934), .B(n31899), .Z(n31902) );
  XOR U31901 ( .A(n31935), .B(n31936), .Z(n31899) );
  AND U31902 ( .A(n31937), .B(n31938), .Z(n31936) );
  XOR U31903 ( .A(n31935), .B(n31939), .Z(n31937) );
  XNOR U31904 ( .A(n31940), .B(n31941), .Z(n31934) );
  AND U31905 ( .A(n31942), .B(n31943), .Z(n31941) );
  XOR U31906 ( .A(n31940), .B(n31944), .Z(n31942) );
  XOR U31907 ( .A(n31945), .B(n31946), .Z(n31903) );
  AND U31908 ( .A(n31947), .B(n31948), .Z(n31946) );
  XOR U31909 ( .A(n31945), .B(n31949), .Z(n31947) );
  XNOR U31910 ( .A(n31836), .B(n31906), .Z(n31908) );
  XNOR U31911 ( .A(n31950), .B(n31951), .Z(n31836) );
  AND U31912 ( .A(n672), .B(n31843), .Z(n31951) );
  XOR U31913 ( .A(n31950), .B(n31841), .Z(n31843) );
  XOR U31914 ( .A(n31952), .B(n31953), .Z(n31906) );
  AND U31915 ( .A(n31954), .B(n31955), .Z(n31953) );
  XNOR U31916 ( .A(n31952), .B(n31851), .Z(n31955) );
  XOR U31917 ( .A(n31956), .B(n31920), .Z(n31851) );
  XNOR U31918 ( .A(n31957), .B(n31927), .Z(n31920) );
  XOR U31919 ( .A(n31916), .B(n31915), .Z(n31927) );
  XNOR U31920 ( .A(n31958), .B(n31912), .Z(n31915) );
  XOR U31921 ( .A(n31959), .B(n31960), .Z(n31912) );
  AND U31922 ( .A(n31961), .B(n31962), .Z(n31960) );
  XNOR U31923 ( .A(n31963), .B(n31964), .Z(n31961) );
  IV U31924 ( .A(n31959), .Z(n31963) );
  XNOR U31925 ( .A(n31965), .B(n31966), .Z(n31958) );
  NOR U31926 ( .A(n31967), .B(n31968), .Z(n31966) );
  XNOR U31927 ( .A(n31965), .B(n31969), .Z(n31967) );
  XOR U31928 ( .A(n31970), .B(n31971), .Z(n31916) );
  NOR U31929 ( .A(n31972), .B(n31973), .Z(n31971) );
  XNOR U31930 ( .A(n31970), .B(n31974), .Z(n31972) );
  XNOR U31931 ( .A(n31926), .B(n31917), .Z(n31957) );
  XOR U31932 ( .A(n31975), .B(n31976), .Z(n31917) );
  AND U31933 ( .A(n31977), .B(n31978), .Z(n31976) );
  XOR U31934 ( .A(n31975), .B(n31979), .Z(n31977) );
  XOR U31935 ( .A(n31980), .B(n31932), .Z(n31926) );
  XOR U31936 ( .A(n31981), .B(n31982), .Z(n31932) );
  NOR U31937 ( .A(n31983), .B(n31984), .Z(n31982) );
  XOR U31938 ( .A(n31981), .B(n31985), .Z(n31983) );
  XNOR U31939 ( .A(n31931), .B(n31923), .Z(n31980) );
  XOR U31940 ( .A(n31986), .B(n31987), .Z(n31923) );
  AND U31941 ( .A(n31988), .B(n31989), .Z(n31987) );
  XOR U31942 ( .A(n31986), .B(n31990), .Z(n31988) );
  XNOR U31943 ( .A(n31991), .B(n31928), .Z(n31931) );
  XOR U31944 ( .A(n31992), .B(n31993), .Z(n31928) );
  AND U31945 ( .A(n31994), .B(n31995), .Z(n31993) );
  XNOR U31946 ( .A(n31996), .B(n31997), .Z(n31994) );
  IV U31947 ( .A(n31992), .Z(n31996) );
  XNOR U31948 ( .A(n31998), .B(n31999), .Z(n31991) );
  NOR U31949 ( .A(n32000), .B(n32001), .Z(n31999) );
  XNOR U31950 ( .A(n31998), .B(n32002), .Z(n32000) );
  XOR U31951 ( .A(n31921), .B(n31933), .Z(n31956) );
  NOR U31952 ( .A(n31859), .B(n32003), .Z(n31933) );
  XNOR U31953 ( .A(n31939), .B(n31938), .Z(n31921) );
  XNOR U31954 ( .A(n32004), .B(n31944), .Z(n31938) );
  XNOR U31955 ( .A(n32005), .B(n32006), .Z(n31944) );
  NOR U31956 ( .A(n32007), .B(n32008), .Z(n32006) );
  XOR U31957 ( .A(n32005), .B(n32009), .Z(n32007) );
  XNOR U31958 ( .A(n31943), .B(n31935), .Z(n32004) );
  XOR U31959 ( .A(n32010), .B(n32011), .Z(n31935) );
  AND U31960 ( .A(n32012), .B(n32013), .Z(n32011) );
  XOR U31961 ( .A(n32010), .B(n32014), .Z(n32012) );
  XNOR U31962 ( .A(n32015), .B(n31940), .Z(n31943) );
  XOR U31963 ( .A(n32016), .B(n32017), .Z(n31940) );
  AND U31964 ( .A(n32018), .B(n32019), .Z(n32017) );
  XNOR U31965 ( .A(n32020), .B(n32021), .Z(n32018) );
  IV U31966 ( .A(n32016), .Z(n32020) );
  XNOR U31967 ( .A(n32022), .B(n32023), .Z(n32015) );
  NOR U31968 ( .A(n32024), .B(n32025), .Z(n32023) );
  XNOR U31969 ( .A(n32022), .B(n32026), .Z(n32024) );
  XOR U31970 ( .A(n31949), .B(n31948), .Z(n31939) );
  XNOR U31971 ( .A(n32027), .B(n31945), .Z(n31948) );
  XOR U31972 ( .A(n32028), .B(n32029), .Z(n31945) );
  AND U31973 ( .A(n32030), .B(n32031), .Z(n32029) );
  XNOR U31974 ( .A(n32032), .B(n32033), .Z(n32030) );
  IV U31975 ( .A(n32028), .Z(n32032) );
  XNOR U31976 ( .A(n32034), .B(n32035), .Z(n32027) );
  NOR U31977 ( .A(n32036), .B(n32037), .Z(n32035) );
  XNOR U31978 ( .A(n32034), .B(n32038), .Z(n32036) );
  XOR U31979 ( .A(n32039), .B(n32040), .Z(n31949) );
  NOR U31980 ( .A(n32041), .B(n32042), .Z(n32040) );
  XNOR U31981 ( .A(n32039), .B(n32043), .Z(n32041) );
  XNOR U31982 ( .A(n31848), .B(n31952), .Z(n31954) );
  XNOR U31983 ( .A(n32044), .B(n32045), .Z(n31848) );
  AND U31984 ( .A(n672), .B(n31855), .Z(n32045) );
  XOR U31985 ( .A(n32044), .B(n31853), .Z(n31855) );
  AND U31986 ( .A(n31856), .B(n31859), .Z(n31952) );
  XOR U31987 ( .A(n32046), .B(n32003), .Z(n31859) );
  XNOR U31988 ( .A(p_input[1760]), .B(p_input[2048]), .Z(n32003) );
  XNOR U31989 ( .A(n31979), .B(n31978), .Z(n32046) );
  XNOR U31990 ( .A(n32047), .B(n31990), .Z(n31978) );
  XOR U31991 ( .A(n31964), .B(n31962), .Z(n31990) );
  XNOR U31992 ( .A(n32048), .B(n31969), .Z(n31962) );
  XOR U31993 ( .A(p_input[1784]), .B(p_input[2072]), .Z(n31969) );
  XOR U31994 ( .A(n31959), .B(n31968), .Z(n32048) );
  XOR U31995 ( .A(n32049), .B(n31965), .Z(n31968) );
  XOR U31996 ( .A(p_input[1782]), .B(p_input[2070]), .Z(n31965) );
  XOR U31997 ( .A(p_input[1783]), .B(n17295), .Z(n32049) );
  XOR U31998 ( .A(p_input[1778]), .B(p_input[2066]), .Z(n31959) );
  XNOR U31999 ( .A(n31974), .B(n31973), .Z(n31964) );
  XOR U32000 ( .A(n32050), .B(n31970), .Z(n31973) );
  XOR U32001 ( .A(p_input[1779]), .B(p_input[2067]), .Z(n31970) );
  XOR U32002 ( .A(p_input[1780]), .B(n17297), .Z(n32050) );
  XOR U32003 ( .A(p_input[1781]), .B(p_input[2069]), .Z(n31974) );
  XOR U32004 ( .A(n31989), .B(n32051), .Z(n32047) );
  IV U32005 ( .A(n31975), .Z(n32051) );
  XOR U32006 ( .A(p_input[1761]), .B(p_input[2049]), .Z(n31975) );
  XNOR U32007 ( .A(n32052), .B(n31997), .Z(n31989) );
  XNOR U32008 ( .A(n31985), .B(n31984), .Z(n31997) );
  XNOR U32009 ( .A(n32053), .B(n31981), .Z(n31984) );
  XNOR U32010 ( .A(p_input[1786]), .B(p_input[2074]), .Z(n31981) );
  XOR U32011 ( .A(p_input[1787]), .B(n17300), .Z(n32053) );
  XOR U32012 ( .A(p_input[1788]), .B(p_input[2076]), .Z(n31985) );
  XOR U32013 ( .A(n31995), .B(n32054), .Z(n32052) );
  IV U32014 ( .A(n31986), .Z(n32054) );
  XOR U32015 ( .A(p_input[1777]), .B(p_input[2065]), .Z(n31986) );
  XNOR U32016 ( .A(n32055), .B(n32002), .Z(n31995) );
  XNOR U32017 ( .A(p_input[1791]), .B(n17303), .Z(n32002) );
  XOR U32018 ( .A(n31992), .B(n32001), .Z(n32055) );
  XOR U32019 ( .A(n32056), .B(n31998), .Z(n32001) );
  XOR U32020 ( .A(p_input[1789]), .B(p_input[2077]), .Z(n31998) );
  XOR U32021 ( .A(p_input[1790]), .B(n17305), .Z(n32056) );
  XOR U32022 ( .A(p_input[1785]), .B(p_input[2073]), .Z(n31992) );
  XOR U32023 ( .A(n32014), .B(n32013), .Z(n31979) );
  XNOR U32024 ( .A(n32057), .B(n32021), .Z(n32013) );
  XNOR U32025 ( .A(n32009), .B(n32008), .Z(n32021) );
  XNOR U32026 ( .A(n32058), .B(n32005), .Z(n32008) );
  XNOR U32027 ( .A(p_input[1771]), .B(p_input[2059]), .Z(n32005) );
  XOR U32028 ( .A(p_input[1772]), .B(n16451), .Z(n32058) );
  XOR U32029 ( .A(p_input[1773]), .B(p_input[2061]), .Z(n32009) );
  XOR U32030 ( .A(n32019), .B(n32059), .Z(n32057) );
  IV U32031 ( .A(n32010), .Z(n32059) );
  XOR U32032 ( .A(p_input[1762]), .B(p_input[2050]), .Z(n32010) );
  XNOR U32033 ( .A(n32060), .B(n32026), .Z(n32019) );
  XNOR U32034 ( .A(p_input[1776]), .B(n16454), .Z(n32026) );
  XOR U32035 ( .A(n32016), .B(n32025), .Z(n32060) );
  XOR U32036 ( .A(n32061), .B(n32022), .Z(n32025) );
  XOR U32037 ( .A(p_input[1774]), .B(p_input[2062]), .Z(n32022) );
  XOR U32038 ( .A(p_input[1775]), .B(n16456), .Z(n32061) );
  XOR U32039 ( .A(p_input[1770]), .B(p_input[2058]), .Z(n32016) );
  XOR U32040 ( .A(n32033), .B(n32031), .Z(n32014) );
  XNOR U32041 ( .A(n32062), .B(n32038), .Z(n32031) );
  XOR U32042 ( .A(p_input[1769]), .B(p_input[2057]), .Z(n32038) );
  XOR U32043 ( .A(n32028), .B(n32037), .Z(n32062) );
  XOR U32044 ( .A(n32063), .B(n32034), .Z(n32037) );
  XOR U32045 ( .A(p_input[1767]), .B(p_input[2055]), .Z(n32034) );
  XOR U32046 ( .A(p_input[1768]), .B(n17312), .Z(n32063) );
  XOR U32047 ( .A(p_input[1763]), .B(p_input[2051]), .Z(n32028) );
  XNOR U32048 ( .A(n32043), .B(n32042), .Z(n32033) );
  XOR U32049 ( .A(n32064), .B(n32039), .Z(n32042) );
  XOR U32050 ( .A(p_input[1764]), .B(p_input[2052]), .Z(n32039) );
  XOR U32051 ( .A(p_input[1765]), .B(n17314), .Z(n32064) );
  XOR U32052 ( .A(p_input[1766]), .B(p_input[2054]), .Z(n32043) );
  XNOR U32053 ( .A(n32065), .B(n32066), .Z(n31856) );
  AND U32054 ( .A(n672), .B(n32067), .Z(n32066) );
  XNOR U32055 ( .A(n32068), .B(n32069), .Z(n672) );
  AND U32056 ( .A(n32070), .B(n32071), .Z(n32069) );
  XOR U32057 ( .A(n32068), .B(n31866), .Z(n32071) );
  XNOR U32058 ( .A(n32068), .B(n31808), .Z(n32070) );
  XOR U32059 ( .A(n32072), .B(n32073), .Z(n32068) );
  AND U32060 ( .A(n32074), .B(n32075), .Z(n32073) );
  XNOR U32061 ( .A(n31879), .B(n32072), .Z(n32075) );
  XOR U32062 ( .A(n32072), .B(n31820), .Z(n32074) );
  XOR U32063 ( .A(n32076), .B(n32077), .Z(n32072) );
  AND U32064 ( .A(n32078), .B(n32079), .Z(n32077) );
  XNOR U32065 ( .A(n31904), .B(n32076), .Z(n32079) );
  XOR U32066 ( .A(n32076), .B(n31831), .Z(n32078) );
  XOR U32067 ( .A(n32080), .B(n32081), .Z(n32076) );
  AND U32068 ( .A(n32082), .B(n32083), .Z(n32081) );
  XOR U32069 ( .A(n32080), .B(n31841), .Z(n32082) );
  XOR U32070 ( .A(n32084), .B(n32085), .Z(n31797) );
  AND U32071 ( .A(n676), .B(n32067), .Z(n32085) );
  XNOR U32072 ( .A(n32065), .B(n32084), .Z(n32067) );
  XNOR U32073 ( .A(n32086), .B(n32087), .Z(n676) );
  AND U32074 ( .A(n32088), .B(n32089), .Z(n32087) );
  XNOR U32075 ( .A(n32090), .B(n32086), .Z(n32089) );
  IV U32076 ( .A(n31866), .Z(n32090) );
  XNOR U32077 ( .A(n32091), .B(n32092), .Z(n31866) );
  AND U32078 ( .A(n679), .B(n32093), .Z(n32092) );
  XNOR U32079 ( .A(n32091), .B(n32094), .Z(n32093) );
  XNOR U32080 ( .A(n31808), .B(n32086), .Z(n32088) );
  XOR U32081 ( .A(n32095), .B(n32096), .Z(n31808) );
  AND U32082 ( .A(n687), .B(n32097), .Z(n32096) );
  XOR U32083 ( .A(n32098), .B(n32099), .Z(n32086) );
  AND U32084 ( .A(n32100), .B(n32101), .Z(n32099) );
  XNOR U32085 ( .A(n32098), .B(n31879), .Z(n32101) );
  XNOR U32086 ( .A(n32102), .B(n32103), .Z(n31879) );
  AND U32087 ( .A(n679), .B(n32104), .Z(n32103) );
  XOR U32088 ( .A(n32105), .B(n32102), .Z(n32104) );
  XNOR U32089 ( .A(n32106), .B(n32098), .Z(n32100) );
  IV U32090 ( .A(n31820), .Z(n32106) );
  XOR U32091 ( .A(n32107), .B(n32108), .Z(n31820) );
  AND U32092 ( .A(n687), .B(n32109), .Z(n32108) );
  XOR U32093 ( .A(n32110), .B(n32111), .Z(n32098) );
  AND U32094 ( .A(n32112), .B(n32113), .Z(n32111) );
  XNOR U32095 ( .A(n32110), .B(n31904), .Z(n32113) );
  XNOR U32096 ( .A(n32114), .B(n32115), .Z(n31904) );
  AND U32097 ( .A(n679), .B(n32116), .Z(n32115) );
  XNOR U32098 ( .A(n32117), .B(n32114), .Z(n32116) );
  XOR U32099 ( .A(n31831), .B(n32110), .Z(n32112) );
  XOR U32100 ( .A(n32118), .B(n32119), .Z(n31831) );
  AND U32101 ( .A(n687), .B(n32120), .Z(n32119) );
  XOR U32102 ( .A(n32080), .B(n32121), .Z(n32110) );
  AND U32103 ( .A(n32122), .B(n32083), .Z(n32121) );
  XNOR U32104 ( .A(n31950), .B(n32080), .Z(n32083) );
  XNOR U32105 ( .A(n32123), .B(n32124), .Z(n31950) );
  AND U32106 ( .A(n679), .B(n32125), .Z(n32124) );
  XOR U32107 ( .A(n32126), .B(n32123), .Z(n32125) );
  XNOR U32108 ( .A(n32127), .B(n32080), .Z(n32122) );
  IV U32109 ( .A(n31841), .Z(n32127) );
  XOR U32110 ( .A(n32128), .B(n32129), .Z(n31841) );
  AND U32111 ( .A(n687), .B(n32130), .Z(n32129) );
  XOR U32112 ( .A(n32131), .B(n32132), .Z(n32080) );
  AND U32113 ( .A(n32133), .B(n32134), .Z(n32132) );
  XNOR U32114 ( .A(n32131), .B(n32044), .Z(n32134) );
  XNOR U32115 ( .A(n32135), .B(n32136), .Z(n32044) );
  AND U32116 ( .A(n679), .B(n32137), .Z(n32136) );
  XNOR U32117 ( .A(n32138), .B(n32135), .Z(n32137) );
  XNOR U32118 ( .A(n32139), .B(n32131), .Z(n32133) );
  IV U32119 ( .A(n31853), .Z(n32139) );
  XOR U32120 ( .A(n32140), .B(n32141), .Z(n31853) );
  AND U32121 ( .A(n687), .B(n32142), .Z(n32141) );
  AND U32122 ( .A(n32084), .B(n32065), .Z(n32131) );
  XNOR U32123 ( .A(n32143), .B(n32144), .Z(n32065) );
  AND U32124 ( .A(n679), .B(n32145), .Z(n32144) );
  XNOR U32125 ( .A(n32146), .B(n32143), .Z(n32145) );
  XNOR U32126 ( .A(n32147), .B(n32148), .Z(n679) );
  AND U32127 ( .A(n32149), .B(n32150), .Z(n32148) );
  XOR U32128 ( .A(n32094), .B(n32147), .Z(n32150) );
  AND U32129 ( .A(n32151), .B(n32152), .Z(n32094) );
  XOR U32130 ( .A(n32147), .B(n32091), .Z(n32149) );
  XNOR U32131 ( .A(n32153), .B(n32154), .Z(n32091) );
  AND U32132 ( .A(n683), .B(n32097), .Z(n32154) );
  XOR U32133 ( .A(n32095), .B(n32153), .Z(n32097) );
  XOR U32134 ( .A(n32155), .B(n32156), .Z(n32147) );
  AND U32135 ( .A(n32157), .B(n32158), .Z(n32156) );
  XNOR U32136 ( .A(n32155), .B(n32151), .Z(n32158) );
  IV U32137 ( .A(n32105), .Z(n32151) );
  XOR U32138 ( .A(n32159), .B(n32160), .Z(n32105) );
  XOR U32139 ( .A(n32161), .B(n32152), .Z(n32160) );
  AND U32140 ( .A(n32117), .B(n32162), .Z(n32152) );
  AND U32141 ( .A(n32163), .B(n32164), .Z(n32161) );
  XOR U32142 ( .A(n32165), .B(n32159), .Z(n32163) );
  XNOR U32143 ( .A(n32102), .B(n32155), .Z(n32157) );
  XNOR U32144 ( .A(n32166), .B(n32167), .Z(n32102) );
  AND U32145 ( .A(n683), .B(n32109), .Z(n32167) );
  XOR U32146 ( .A(n32166), .B(n32107), .Z(n32109) );
  XOR U32147 ( .A(n32168), .B(n32169), .Z(n32155) );
  AND U32148 ( .A(n32170), .B(n32171), .Z(n32169) );
  XNOR U32149 ( .A(n32168), .B(n32117), .Z(n32171) );
  XOR U32150 ( .A(n32172), .B(n32164), .Z(n32117) );
  XNOR U32151 ( .A(n32173), .B(n32159), .Z(n32164) );
  XOR U32152 ( .A(n32174), .B(n32175), .Z(n32159) );
  AND U32153 ( .A(n32176), .B(n32177), .Z(n32175) );
  XOR U32154 ( .A(n32178), .B(n32174), .Z(n32176) );
  XNOR U32155 ( .A(n32179), .B(n32180), .Z(n32173) );
  AND U32156 ( .A(n32181), .B(n32182), .Z(n32180) );
  XOR U32157 ( .A(n32179), .B(n32183), .Z(n32181) );
  XNOR U32158 ( .A(n32165), .B(n32162), .Z(n32172) );
  AND U32159 ( .A(n32184), .B(n32185), .Z(n32162) );
  XOR U32160 ( .A(n32186), .B(n32187), .Z(n32165) );
  AND U32161 ( .A(n32188), .B(n32189), .Z(n32187) );
  XOR U32162 ( .A(n32186), .B(n32190), .Z(n32188) );
  XNOR U32163 ( .A(n32114), .B(n32168), .Z(n32170) );
  XNOR U32164 ( .A(n32191), .B(n32192), .Z(n32114) );
  AND U32165 ( .A(n683), .B(n32120), .Z(n32192) );
  XOR U32166 ( .A(n32191), .B(n32118), .Z(n32120) );
  XOR U32167 ( .A(n32193), .B(n32194), .Z(n32168) );
  AND U32168 ( .A(n32195), .B(n32196), .Z(n32194) );
  XNOR U32169 ( .A(n32193), .B(n32184), .Z(n32196) );
  IV U32170 ( .A(n32126), .Z(n32184) );
  XNOR U32171 ( .A(n32197), .B(n32177), .Z(n32126) );
  XNOR U32172 ( .A(n32198), .B(n32183), .Z(n32177) );
  XOR U32173 ( .A(n32199), .B(n32200), .Z(n32183) );
  AND U32174 ( .A(n32201), .B(n32202), .Z(n32200) );
  XOR U32175 ( .A(n32199), .B(n32203), .Z(n32201) );
  XNOR U32176 ( .A(n32182), .B(n32174), .Z(n32198) );
  XOR U32177 ( .A(n32204), .B(n32205), .Z(n32174) );
  AND U32178 ( .A(n32206), .B(n32207), .Z(n32205) );
  XNOR U32179 ( .A(n32208), .B(n32204), .Z(n32206) );
  XNOR U32180 ( .A(n32209), .B(n32179), .Z(n32182) );
  XOR U32181 ( .A(n32210), .B(n32211), .Z(n32179) );
  AND U32182 ( .A(n32212), .B(n32213), .Z(n32211) );
  XOR U32183 ( .A(n32210), .B(n32214), .Z(n32212) );
  XNOR U32184 ( .A(n32215), .B(n32216), .Z(n32209) );
  AND U32185 ( .A(n32217), .B(n32218), .Z(n32216) );
  XNOR U32186 ( .A(n32215), .B(n32219), .Z(n32217) );
  XNOR U32187 ( .A(n32178), .B(n32185), .Z(n32197) );
  AND U32188 ( .A(n32138), .B(n32220), .Z(n32185) );
  XOR U32189 ( .A(n32190), .B(n32189), .Z(n32178) );
  XNOR U32190 ( .A(n32221), .B(n32186), .Z(n32189) );
  XOR U32191 ( .A(n32222), .B(n32223), .Z(n32186) );
  AND U32192 ( .A(n32224), .B(n32225), .Z(n32223) );
  XOR U32193 ( .A(n32222), .B(n32226), .Z(n32224) );
  XNOR U32194 ( .A(n32227), .B(n32228), .Z(n32221) );
  AND U32195 ( .A(n32229), .B(n32230), .Z(n32228) );
  XOR U32196 ( .A(n32227), .B(n32231), .Z(n32229) );
  XOR U32197 ( .A(n32232), .B(n32233), .Z(n32190) );
  AND U32198 ( .A(n32234), .B(n32235), .Z(n32233) );
  XOR U32199 ( .A(n32232), .B(n32236), .Z(n32234) );
  XNOR U32200 ( .A(n32123), .B(n32193), .Z(n32195) );
  XNOR U32201 ( .A(n32237), .B(n32238), .Z(n32123) );
  AND U32202 ( .A(n683), .B(n32130), .Z(n32238) );
  XOR U32203 ( .A(n32237), .B(n32128), .Z(n32130) );
  XOR U32204 ( .A(n32239), .B(n32240), .Z(n32193) );
  AND U32205 ( .A(n32241), .B(n32242), .Z(n32240) );
  XNOR U32206 ( .A(n32239), .B(n32138), .Z(n32242) );
  XOR U32207 ( .A(n32243), .B(n32207), .Z(n32138) );
  XNOR U32208 ( .A(n32244), .B(n32214), .Z(n32207) );
  XOR U32209 ( .A(n32203), .B(n32202), .Z(n32214) );
  XNOR U32210 ( .A(n32245), .B(n32199), .Z(n32202) );
  XOR U32211 ( .A(n32246), .B(n32247), .Z(n32199) );
  AND U32212 ( .A(n32248), .B(n32249), .Z(n32247) );
  XNOR U32213 ( .A(n32250), .B(n32251), .Z(n32248) );
  IV U32214 ( .A(n32246), .Z(n32250) );
  XNOR U32215 ( .A(n32252), .B(n32253), .Z(n32245) );
  NOR U32216 ( .A(n32254), .B(n32255), .Z(n32253) );
  XNOR U32217 ( .A(n32252), .B(n32256), .Z(n32254) );
  XOR U32218 ( .A(n32257), .B(n32258), .Z(n32203) );
  NOR U32219 ( .A(n32259), .B(n32260), .Z(n32258) );
  XNOR U32220 ( .A(n32257), .B(n32261), .Z(n32259) );
  XNOR U32221 ( .A(n32213), .B(n32204), .Z(n32244) );
  XOR U32222 ( .A(n32262), .B(n32263), .Z(n32204) );
  AND U32223 ( .A(n32264), .B(n32265), .Z(n32263) );
  XOR U32224 ( .A(n32262), .B(n32266), .Z(n32264) );
  XOR U32225 ( .A(n32267), .B(n32219), .Z(n32213) );
  XOR U32226 ( .A(n32268), .B(n32269), .Z(n32219) );
  NOR U32227 ( .A(n32270), .B(n32271), .Z(n32269) );
  XOR U32228 ( .A(n32268), .B(n32272), .Z(n32270) );
  XNOR U32229 ( .A(n32218), .B(n32210), .Z(n32267) );
  XOR U32230 ( .A(n32273), .B(n32274), .Z(n32210) );
  AND U32231 ( .A(n32275), .B(n32276), .Z(n32274) );
  XOR U32232 ( .A(n32273), .B(n32277), .Z(n32275) );
  XNOR U32233 ( .A(n32278), .B(n32215), .Z(n32218) );
  XOR U32234 ( .A(n32279), .B(n32280), .Z(n32215) );
  AND U32235 ( .A(n32281), .B(n32282), .Z(n32280) );
  XNOR U32236 ( .A(n32283), .B(n32284), .Z(n32281) );
  IV U32237 ( .A(n32279), .Z(n32283) );
  XNOR U32238 ( .A(n32285), .B(n32286), .Z(n32278) );
  NOR U32239 ( .A(n32287), .B(n32288), .Z(n32286) );
  XNOR U32240 ( .A(n32285), .B(n32289), .Z(n32287) );
  XOR U32241 ( .A(n32208), .B(n32220), .Z(n32243) );
  NOR U32242 ( .A(n32146), .B(n32290), .Z(n32220) );
  XNOR U32243 ( .A(n32226), .B(n32225), .Z(n32208) );
  XNOR U32244 ( .A(n32291), .B(n32231), .Z(n32225) );
  XNOR U32245 ( .A(n32292), .B(n32293), .Z(n32231) );
  NOR U32246 ( .A(n32294), .B(n32295), .Z(n32293) );
  XOR U32247 ( .A(n32292), .B(n32296), .Z(n32294) );
  XNOR U32248 ( .A(n32230), .B(n32222), .Z(n32291) );
  XOR U32249 ( .A(n32297), .B(n32298), .Z(n32222) );
  AND U32250 ( .A(n32299), .B(n32300), .Z(n32298) );
  XOR U32251 ( .A(n32297), .B(n32301), .Z(n32299) );
  XNOR U32252 ( .A(n32302), .B(n32227), .Z(n32230) );
  XOR U32253 ( .A(n32303), .B(n32304), .Z(n32227) );
  AND U32254 ( .A(n32305), .B(n32306), .Z(n32304) );
  XNOR U32255 ( .A(n32307), .B(n32308), .Z(n32305) );
  IV U32256 ( .A(n32303), .Z(n32307) );
  XNOR U32257 ( .A(n32309), .B(n32310), .Z(n32302) );
  NOR U32258 ( .A(n32311), .B(n32312), .Z(n32310) );
  XNOR U32259 ( .A(n32309), .B(n32313), .Z(n32311) );
  XOR U32260 ( .A(n32236), .B(n32235), .Z(n32226) );
  XNOR U32261 ( .A(n32314), .B(n32232), .Z(n32235) );
  XOR U32262 ( .A(n32315), .B(n32316), .Z(n32232) );
  AND U32263 ( .A(n32317), .B(n32318), .Z(n32316) );
  XNOR U32264 ( .A(n32319), .B(n32320), .Z(n32317) );
  IV U32265 ( .A(n32315), .Z(n32319) );
  XNOR U32266 ( .A(n32321), .B(n32322), .Z(n32314) );
  NOR U32267 ( .A(n32323), .B(n32324), .Z(n32322) );
  XNOR U32268 ( .A(n32321), .B(n32325), .Z(n32323) );
  XOR U32269 ( .A(n32326), .B(n32327), .Z(n32236) );
  NOR U32270 ( .A(n32328), .B(n32329), .Z(n32327) );
  XNOR U32271 ( .A(n32326), .B(n32330), .Z(n32328) );
  XNOR U32272 ( .A(n32135), .B(n32239), .Z(n32241) );
  XNOR U32273 ( .A(n32331), .B(n32332), .Z(n32135) );
  AND U32274 ( .A(n683), .B(n32142), .Z(n32332) );
  XOR U32275 ( .A(n32331), .B(n32140), .Z(n32142) );
  AND U32276 ( .A(n32143), .B(n32146), .Z(n32239) );
  XOR U32277 ( .A(n32333), .B(n32290), .Z(n32146) );
  XNOR U32278 ( .A(p_input[1792]), .B(p_input[2048]), .Z(n32290) );
  XNOR U32279 ( .A(n32266), .B(n32265), .Z(n32333) );
  XNOR U32280 ( .A(n32334), .B(n32277), .Z(n32265) );
  XOR U32281 ( .A(n32251), .B(n32249), .Z(n32277) );
  XNOR U32282 ( .A(n32335), .B(n32256), .Z(n32249) );
  XOR U32283 ( .A(p_input[1816]), .B(p_input[2072]), .Z(n32256) );
  XOR U32284 ( .A(n32246), .B(n32255), .Z(n32335) );
  XOR U32285 ( .A(n32336), .B(n32252), .Z(n32255) );
  XOR U32286 ( .A(p_input[1814]), .B(p_input[2070]), .Z(n32252) );
  XOR U32287 ( .A(p_input[1815]), .B(n17295), .Z(n32336) );
  XOR U32288 ( .A(p_input[1810]), .B(p_input[2066]), .Z(n32246) );
  XNOR U32289 ( .A(n32261), .B(n32260), .Z(n32251) );
  XOR U32290 ( .A(n32337), .B(n32257), .Z(n32260) );
  XOR U32291 ( .A(p_input[1811]), .B(p_input[2067]), .Z(n32257) );
  XOR U32292 ( .A(p_input[1812]), .B(n17297), .Z(n32337) );
  XOR U32293 ( .A(p_input[1813]), .B(p_input[2069]), .Z(n32261) );
  XOR U32294 ( .A(n32276), .B(n32338), .Z(n32334) );
  IV U32295 ( .A(n32262), .Z(n32338) );
  XOR U32296 ( .A(p_input[1793]), .B(p_input[2049]), .Z(n32262) );
  XNOR U32297 ( .A(n32339), .B(n32284), .Z(n32276) );
  XNOR U32298 ( .A(n32272), .B(n32271), .Z(n32284) );
  XNOR U32299 ( .A(n32340), .B(n32268), .Z(n32271) );
  XNOR U32300 ( .A(p_input[1818]), .B(p_input[2074]), .Z(n32268) );
  XOR U32301 ( .A(p_input[1819]), .B(n17300), .Z(n32340) );
  XOR U32302 ( .A(p_input[1820]), .B(p_input[2076]), .Z(n32272) );
  XOR U32303 ( .A(n32282), .B(n32341), .Z(n32339) );
  IV U32304 ( .A(n32273), .Z(n32341) );
  XOR U32305 ( .A(p_input[1809]), .B(p_input[2065]), .Z(n32273) );
  XNOR U32306 ( .A(n32342), .B(n32289), .Z(n32282) );
  XNOR U32307 ( .A(p_input[1823]), .B(n17303), .Z(n32289) );
  XOR U32308 ( .A(n32279), .B(n32288), .Z(n32342) );
  XOR U32309 ( .A(n32343), .B(n32285), .Z(n32288) );
  XOR U32310 ( .A(p_input[1821]), .B(p_input[2077]), .Z(n32285) );
  XOR U32311 ( .A(p_input[1822]), .B(n17305), .Z(n32343) );
  XOR U32312 ( .A(p_input[1817]), .B(p_input[2073]), .Z(n32279) );
  XOR U32313 ( .A(n32301), .B(n32300), .Z(n32266) );
  XNOR U32314 ( .A(n32344), .B(n32308), .Z(n32300) );
  XNOR U32315 ( .A(n32296), .B(n32295), .Z(n32308) );
  XNOR U32316 ( .A(n32345), .B(n32292), .Z(n32295) );
  XNOR U32317 ( .A(p_input[1803]), .B(p_input[2059]), .Z(n32292) );
  XOR U32318 ( .A(p_input[1804]), .B(n16451), .Z(n32345) );
  XOR U32319 ( .A(p_input[1805]), .B(p_input[2061]), .Z(n32296) );
  XOR U32320 ( .A(n32306), .B(n32346), .Z(n32344) );
  IV U32321 ( .A(n32297), .Z(n32346) );
  XOR U32322 ( .A(p_input[1794]), .B(p_input[2050]), .Z(n32297) );
  XNOR U32323 ( .A(n32347), .B(n32313), .Z(n32306) );
  XNOR U32324 ( .A(p_input[1808]), .B(n16454), .Z(n32313) );
  XOR U32325 ( .A(n32303), .B(n32312), .Z(n32347) );
  XOR U32326 ( .A(n32348), .B(n32309), .Z(n32312) );
  XOR U32327 ( .A(p_input[1806]), .B(p_input[2062]), .Z(n32309) );
  XOR U32328 ( .A(p_input[1807]), .B(n16456), .Z(n32348) );
  XOR U32329 ( .A(p_input[1802]), .B(p_input[2058]), .Z(n32303) );
  XOR U32330 ( .A(n32320), .B(n32318), .Z(n32301) );
  XNOR U32331 ( .A(n32349), .B(n32325), .Z(n32318) );
  XOR U32332 ( .A(p_input[1801]), .B(p_input[2057]), .Z(n32325) );
  XOR U32333 ( .A(n32315), .B(n32324), .Z(n32349) );
  XOR U32334 ( .A(n32350), .B(n32321), .Z(n32324) );
  XOR U32335 ( .A(p_input[1799]), .B(p_input[2055]), .Z(n32321) );
  XOR U32336 ( .A(p_input[1800]), .B(n17312), .Z(n32350) );
  XOR U32337 ( .A(p_input[1795]), .B(p_input[2051]), .Z(n32315) );
  XNOR U32338 ( .A(n32330), .B(n32329), .Z(n32320) );
  XOR U32339 ( .A(n32351), .B(n32326), .Z(n32329) );
  XOR U32340 ( .A(p_input[1796]), .B(p_input[2052]), .Z(n32326) );
  XOR U32341 ( .A(p_input[1797]), .B(n17314), .Z(n32351) );
  XOR U32342 ( .A(p_input[1798]), .B(p_input[2054]), .Z(n32330) );
  XNOR U32343 ( .A(n32352), .B(n32353), .Z(n32143) );
  AND U32344 ( .A(n683), .B(n32354), .Z(n32353) );
  XNOR U32345 ( .A(n32355), .B(n32356), .Z(n683) );
  AND U32346 ( .A(n32357), .B(n32358), .Z(n32356) );
  XOR U32347 ( .A(n32355), .B(n32153), .Z(n32358) );
  XNOR U32348 ( .A(n32355), .B(n32095), .Z(n32357) );
  XOR U32349 ( .A(n32359), .B(n32360), .Z(n32355) );
  AND U32350 ( .A(n32361), .B(n32362), .Z(n32360) );
  XNOR U32351 ( .A(n32166), .B(n32359), .Z(n32362) );
  XOR U32352 ( .A(n32359), .B(n32107), .Z(n32361) );
  XOR U32353 ( .A(n32363), .B(n32364), .Z(n32359) );
  AND U32354 ( .A(n32365), .B(n32366), .Z(n32364) );
  XNOR U32355 ( .A(n32191), .B(n32363), .Z(n32366) );
  XOR U32356 ( .A(n32363), .B(n32118), .Z(n32365) );
  XOR U32357 ( .A(n32367), .B(n32368), .Z(n32363) );
  AND U32358 ( .A(n32369), .B(n32370), .Z(n32368) );
  XOR U32359 ( .A(n32367), .B(n32128), .Z(n32369) );
  XOR U32360 ( .A(n32371), .B(n32372), .Z(n32084) );
  AND U32361 ( .A(n687), .B(n32354), .Z(n32372) );
  XNOR U32362 ( .A(n32352), .B(n32371), .Z(n32354) );
  XNOR U32363 ( .A(n32373), .B(n32374), .Z(n687) );
  AND U32364 ( .A(n32375), .B(n32376), .Z(n32374) );
  XNOR U32365 ( .A(n32377), .B(n32373), .Z(n32376) );
  IV U32366 ( .A(n32153), .Z(n32377) );
  XNOR U32367 ( .A(n32378), .B(n32379), .Z(n32153) );
  AND U32368 ( .A(n690), .B(n32380), .Z(n32379) );
  XNOR U32369 ( .A(n32378), .B(n32381), .Z(n32380) );
  XNOR U32370 ( .A(n32095), .B(n32373), .Z(n32375) );
  XNOR U32371 ( .A(n32382), .B(n32383), .Z(n32095) );
  AND U32372 ( .A(n698), .B(n32384), .Z(n32383) );
  XNOR U32373 ( .A(n32385), .B(n32386), .Z(n32384) );
  XOR U32374 ( .A(n32387), .B(n32388), .Z(n32373) );
  AND U32375 ( .A(n32389), .B(n32390), .Z(n32388) );
  XNOR U32376 ( .A(n32387), .B(n32166), .Z(n32390) );
  XNOR U32377 ( .A(n32391), .B(n32392), .Z(n32166) );
  AND U32378 ( .A(n690), .B(n32393), .Z(n32392) );
  XOR U32379 ( .A(n32394), .B(n32391), .Z(n32393) );
  XNOR U32380 ( .A(n32395), .B(n32387), .Z(n32389) );
  IV U32381 ( .A(n32107), .Z(n32395) );
  XOR U32382 ( .A(n32396), .B(n32397), .Z(n32107) );
  AND U32383 ( .A(n698), .B(n32398), .Z(n32397) );
  XOR U32384 ( .A(n32399), .B(n32400), .Z(n32387) );
  AND U32385 ( .A(n32401), .B(n32402), .Z(n32400) );
  XNOR U32386 ( .A(n32399), .B(n32191), .Z(n32402) );
  XNOR U32387 ( .A(n32403), .B(n32404), .Z(n32191) );
  AND U32388 ( .A(n690), .B(n32405), .Z(n32404) );
  XNOR U32389 ( .A(n32406), .B(n32403), .Z(n32405) );
  XOR U32390 ( .A(n32118), .B(n32399), .Z(n32401) );
  XOR U32391 ( .A(n32407), .B(n32408), .Z(n32118) );
  AND U32392 ( .A(n698), .B(n32409), .Z(n32408) );
  XOR U32393 ( .A(n32367), .B(n32410), .Z(n32399) );
  AND U32394 ( .A(n32411), .B(n32370), .Z(n32410) );
  XNOR U32395 ( .A(n32237), .B(n32367), .Z(n32370) );
  XNOR U32396 ( .A(n32412), .B(n32413), .Z(n32237) );
  AND U32397 ( .A(n690), .B(n32414), .Z(n32413) );
  XOR U32398 ( .A(n32415), .B(n32412), .Z(n32414) );
  XNOR U32399 ( .A(n32416), .B(n32367), .Z(n32411) );
  IV U32400 ( .A(n32128), .Z(n32416) );
  XOR U32401 ( .A(n32417), .B(n32418), .Z(n32128) );
  AND U32402 ( .A(n698), .B(n32419), .Z(n32418) );
  XOR U32403 ( .A(n32420), .B(n32421), .Z(n32367) );
  AND U32404 ( .A(n32422), .B(n32423), .Z(n32421) );
  XNOR U32405 ( .A(n32420), .B(n32331), .Z(n32423) );
  XNOR U32406 ( .A(n32424), .B(n32425), .Z(n32331) );
  AND U32407 ( .A(n690), .B(n32426), .Z(n32425) );
  XNOR U32408 ( .A(n32427), .B(n32424), .Z(n32426) );
  XNOR U32409 ( .A(n32428), .B(n32420), .Z(n32422) );
  IV U32410 ( .A(n32140), .Z(n32428) );
  XOR U32411 ( .A(n32429), .B(n32430), .Z(n32140) );
  AND U32412 ( .A(n698), .B(n32431), .Z(n32430) );
  AND U32413 ( .A(n32371), .B(n32352), .Z(n32420) );
  XNOR U32414 ( .A(n32432), .B(n32433), .Z(n32352) );
  AND U32415 ( .A(n690), .B(n32434), .Z(n32433) );
  XNOR U32416 ( .A(n32435), .B(n32432), .Z(n32434) );
  XNOR U32417 ( .A(n32436), .B(n32437), .Z(n690) );
  AND U32418 ( .A(n32438), .B(n32439), .Z(n32437) );
  XOR U32419 ( .A(n32381), .B(n32436), .Z(n32439) );
  AND U32420 ( .A(n32440), .B(n32441), .Z(n32381) );
  XOR U32421 ( .A(n32436), .B(n32378), .Z(n32438) );
  XOR U32422 ( .A(n32385), .B(n32442), .Z(n32378) );
  AND U32423 ( .A(n694), .B(n32443), .Z(n32442) );
  XOR U32424 ( .A(n32385), .B(n32382), .Z(n32443) );
  XOR U32425 ( .A(n32444), .B(n32445), .Z(n32436) );
  AND U32426 ( .A(n32446), .B(n32447), .Z(n32445) );
  XNOR U32427 ( .A(n32444), .B(n32440), .Z(n32447) );
  IV U32428 ( .A(n32394), .Z(n32440) );
  XOR U32429 ( .A(n32448), .B(n32449), .Z(n32394) );
  XOR U32430 ( .A(n32450), .B(n32441), .Z(n32449) );
  AND U32431 ( .A(n32406), .B(n32451), .Z(n32441) );
  AND U32432 ( .A(n32452), .B(n32453), .Z(n32450) );
  XOR U32433 ( .A(n32454), .B(n32448), .Z(n32452) );
  XNOR U32434 ( .A(n32391), .B(n32444), .Z(n32446) );
  XNOR U32435 ( .A(n32455), .B(n32456), .Z(n32391) );
  AND U32436 ( .A(n694), .B(n32398), .Z(n32456) );
  XOR U32437 ( .A(n32455), .B(n32396), .Z(n32398) );
  XOR U32438 ( .A(n32457), .B(n32458), .Z(n32444) );
  AND U32439 ( .A(n32459), .B(n32460), .Z(n32458) );
  XNOR U32440 ( .A(n32457), .B(n32406), .Z(n32460) );
  XOR U32441 ( .A(n32461), .B(n32453), .Z(n32406) );
  XNOR U32442 ( .A(n32462), .B(n32448), .Z(n32453) );
  XOR U32443 ( .A(n32463), .B(n32464), .Z(n32448) );
  AND U32444 ( .A(n32465), .B(n32466), .Z(n32464) );
  XOR U32445 ( .A(n32467), .B(n32463), .Z(n32465) );
  XNOR U32446 ( .A(n32468), .B(n32469), .Z(n32462) );
  AND U32447 ( .A(n32470), .B(n32471), .Z(n32469) );
  XOR U32448 ( .A(n32468), .B(n32472), .Z(n32470) );
  XNOR U32449 ( .A(n32454), .B(n32451), .Z(n32461) );
  AND U32450 ( .A(n32473), .B(n32474), .Z(n32451) );
  XOR U32451 ( .A(n32475), .B(n32476), .Z(n32454) );
  AND U32452 ( .A(n32477), .B(n32478), .Z(n32476) );
  XOR U32453 ( .A(n32475), .B(n32479), .Z(n32477) );
  XNOR U32454 ( .A(n32403), .B(n32457), .Z(n32459) );
  XNOR U32455 ( .A(n32480), .B(n32481), .Z(n32403) );
  AND U32456 ( .A(n694), .B(n32409), .Z(n32481) );
  XOR U32457 ( .A(n32480), .B(n32407), .Z(n32409) );
  XOR U32458 ( .A(n32482), .B(n32483), .Z(n32457) );
  AND U32459 ( .A(n32484), .B(n32485), .Z(n32483) );
  XNOR U32460 ( .A(n32482), .B(n32473), .Z(n32485) );
  IV U32461 ( .A(n32415), .Z(n32473) );
  XNOR U32462 ( .A(n32486), .B(n32466), .Z(n32415) );
  XNOR U32463 ( .A(n32487), .B(n32472), .Z(n32466) );
  XOR U32464 ( .A(n32488), .B(n32489), .Z(n32472) );
  AND U32465 ( .A(n32490), .B(n32491), .Z(n32489) );
  XOR U32466 ( .A(n32488), .B(n32492), .Z(n32490) );
  XNOR U32467 ( .A(n32471), .B(n32463), .Z(n32487) );
  XOR U32468 ( .A(n32493), .B(n32494), .Z(n32463) );
  AND U32469 ( .A(n32495), .B(n32496), .Z(n32494) );
  XNOR U32470 ( .A(n32497), .B(n32493), .Z(n32495) );
  XNOR U32471 ( .A(n32498), .B(n32468), .Z(n32471) );
  XOR U32472 ( .A(n32499), .B(n32500), .Z(n32468) );
  AND U32473 ( .A(n32501), .B(n32502), .Z(n32500) );
  XOR U32474 ( .A(n32499), .B(n32503), .Z(n32501) );
  XNOR U32475 ( .A(n32504), .B(n32505), .Z(n32498) );
  AND U32476 ( .A(n32506), .B(n32507), .Z(n32505) );
  XNOR U32477 ( .A(n32504), .B(n32508), .Z(n32506) );
  XNOR U32478 ( .A(n32467), .B(n32474), .Z(n32486) );
  AND U32479 ( .A(n32427), .B(n32509), .Z(n32474) );
  XOR U32480 ( .A(n32479), .B(n32478), .Z(n32467) );
  XNOR U32481 ( .A(n32510), .B(n32475), .Z(n32478) );
  XOR U32482 ( .A(n32511), .B(n32512), .Z(n32475) );
  AND U32483 ( .A(n32513), .B(n32514), .Z(n32512) );
  XOR U32484 ( .A(n32511), .B(n32515), .Z(n32513) );
  XNOR U32485 ( .A(n32516), .B(n32517), .Z(n32510) );
  AND U32486 ( .A(n32518), .B(n32519), .Z(n32517) );
  XOR U32487 ( .A(n32516), .B(n32520), .Z(n32518) );
  XOR U32488 ( .A(n32521), .B(n32522), .Z(n32479) );
  AND U32489 ( .A(n32523), .B(n32524), .Z(n32522) );
  XOR U32490 ( .A(n32521), .B(n32525), .Z(n32523) );
  XNOR U32491 ( .A(n32412), .B(n32482), .Z(n32484) );
  XNOR U32492 ( .A(n32526), .B(n32527), .Z(n32412) );
  AND U32493 ( .A(n694), .B(n32419), .Z(n32527) );
  XOR U32494 ( .A(n32526), .B(n32417), .Z(n32419) );
  XOR U32495 ( .A(n32528), .B(n32529), .Z(n32482) );
  AND U32496 ( .A(n32530), .B(n32531), .Z(n32529) );
  XNOR U32497 ( .A(n32528), .B(n32427), .Z(n32531) );
  XOR U32498 ( .A(n32532), .B(n32496), .Z(n32427) );
  XNOR U32499 ( .A(n32533), .B(n32503), .Z(n32496) );
  XOR U32500 ( .A(n32492), .B(n32491), .Z(n32503) );
  XNOR U32501 ( .A(n32534), .B(n32488), .Z(n32491) );
  XOR U32502 ( .A(n32535), .B(n32536), .Z(n32488) );
  AND U32503 ( .A(n32537), .B(n32538), .Z(n32536) );
  XNOR U32504 ( .A(n32539), .B(n32540), .Z(n32537) );
  IV U32505 ( .A(n32535), .Z(n32539) );
  XNOR U32506 ( .A(n32541), .B(n32542), .Z(n32534) );
  NOR U32507 ( .A(n32543), .B(n32544), .Z(n32542) );
  XNOR U32508 ( .A(n32541), .B(n32545), .Z(n32543) );
  XOR U32509 ( .A(n32546), .B(n32547), .Z(n32492) );
  NOR U32510 ( .A(n32548), .B(n32549), .Z(n32547) );
  XNOR U32511 ( .A(n32546), .B(n32550), .Z(n32548) );
  XNOR U32512 ( .A(n32502), .B(n32493), .Z(n32533) );
  XOR U32513 ( .A(n32551), .B(n32552), .Z(n32493) );
  AND U32514 ( .A(n32553), .B(n32554), .Z(n32552) );
  XOR U32515 ( .A(n32551), .B(n32555), .Z(n32553) );
  XOR U32516 ( .A(n32556), .B(n32508), .Z(n32502) );
  XOR U32517 ( .A(n32557), .B(n32558), .Z(n32508) );
  NOR U32518 ( .A(n32559), .B(n32560), .Z(n32558) );
  XOR U32519 ( .A(n32557), .B(n32561), .Z(n32559) );
  XNOR U32520 ( .A(n32507), .B(n32499), .Z(n32556) );
  XOR U32521 ( .A(n32562), .B(n32563), .Z(n32499) );
  AND U32522 ( .A(n32564), .B(n32565), .Z(n32563) );
  XOR U32523 ( .A(n32562), .B(n32566), .Z(n32564) );
  XNOR U32524 ( .A(n32567), .B(n32504), .Z(n32507) );
  XOR U32525 ( .A(n32568), .B(n32569), .Z(n32504) );
  AND U32526 ( .A(n32570), .B(n32571), .Z(n32569) );
  XNOR U32527 ( .A(n32572), .B(n32573), .Z(n32570) );
  IV U32528 ( .A(n32568), .Z(n32572) );
  XNOR U32529 ( .A(n32574), .B(n32575), .Z(n32567) );
  NOR U32530 ( .A(n32576), .B(n32577), .Z(n32575) );
  XNOR U32531 ( .A(n32574), .B(n32578), .Z(n32576) );
  XOR U32532 ( .A(n32497), .B(n32509), .Z(n32532) );
  NOR U32533 ( .A(n32435), .B(n32579), .Z(n32509) );
  XNOR U32534 ( .A(n32515), .B(n32514), .Z(n32497) );
  XNOR U32535 ( .A(n32580), .B(n32520), .Z(n32514) );
  XNOR U32536 ( .A(n32581), .B(n32582), .Z(n32520) );
  NOR U32537 ( .A(n32583), .B(n32584), .Z(n32582) );
  XOR U32538 ( .A(n32581), .B(n32585), .Z(n32583) );
  XNOR U32539 ( .A(n32519), .B(n32511), .Z(n32580) );
  XOR U32540 ( .A(n32586), .B(n32587), .Z(n32511) );
  AND U32541 ( .A(n32588), .B(n32589), .Z(n32587) );
  XOR U32542 ( .A(n32586), .B(n32590), .Z(n32588) );
  XNOR U32543 ( .A(n32591), .B(n32516), .Z(n32519) );
  XOR U32544 ( .A(n32592), .B(n32593), .Z(n32516) );
  AND U32545 ( .A(n32594), .B(n32595), .Z(n32593) );
  XNOR U32546 ( .A(n32596), .B(n32597), .Z(n32594) );
  IV U32547 ( .A(n32592), .Z(n32596) );
  XNOR U32548 ( .A(n32598), .B(n32599), .Z(n32591) );
  NOR U32549 ( .A(n32600), .B(n32601), .Z(n32599) );
  XNOR U32550 ( .A(n32598), .B(n32602), .Z(n32600) );
  XOR U32551 ( .A(n32525), .B(n32524), .Z(n32515) );
  XNOR U32552 ( .A(n32603), .B(n32521), .Z(n32524) );
  XOR U32553 ( .A(n32604), .B(n32605), .Z(n32521) );
  AND U32554 ( .A(n32606), .B(n32607), .Z(n32605) );
  XNOR U32555 ( .A(n32608), .B(n32609), .Z(n32606) );
  IV U32556 ( .A(n32604), .Z(n32608) );
  XNOR U32557 ( .A(n32610), .B(n32611), .Z(n32603) );
  NOR U32558 ( .A(n32612), .B(n32613), .Z(n32611) );
  XNOR U32559 ( .A(n32610), .B(n32614), .Z(n32612) );
  XOR U32560 ( .A(n32615), .B(n32616), .Z(n32525) );
  NOR U32561 ( .A(n32617), .B(n32618), .Z(n32616) );
  XNOR U32562 ( .A(n32615), .B(n32619), .Z(n32617) );
  XNOR U32563 ( .A(n32424), .B(n32528), .Z(n32530) );
  XNOR U32564 ( .A(n32620), .B(n32621), .Z(n32424) );
  AND U32565 ( .A(n694), .B(n32431), .Z(n32621) );
  XOR U32566 ( .A(n32620), .B(n32429), .Z(n32431) );
  AND U32567 ( .A(n32432), .B(n32435), .Z(n32528) );
  XOR U32568 ( .A(n32622), .B(n32579), .Z(n32435) );
  XNOR U32569 ( .A(p_input[1824]), .B(p_input[2048]), .Z(n32579) );
  XNOR U32570 ( .A(n32555), .B(n32554), .Z(n32622) );
  XNOR U32571 ( .A(n32623), .B(n32566), .Z(n32554) );
  XOR U32572 ( .A(n32540), .B(n32538), .Z(n32566) );
  XNOR U32573 ( .A(n32624), .B(n32545), .Z(n32538) );
  XOR U32574 ( .A(p_input[1848]), .B(p_input[2072]), .Z(n32545) );
  XOR U32575 ( .A(n32535), .B(n32544), .Z(n32624) );
  XOR U32576 ( .A(n32625), .B(n32541), .Z(n32544) );
  XOR U32577 ( .A(p_input[1846]), .B(p_input[2070]), .Z(n32541) );
  XOR U32578 ( .A(p_input[1847]), .B(n17295), .Z(n32625) );
  XOR U32579 ( .A(p_input[1842]), .B(p_input[2066]), .Z(n32535) );
  XNOR U32580 ( .A(n32550), .B(n32549), .Z(n32540) );
  XOR U32581 ( .A(n32626), .B(n32546), .Z(n32549) );
  XOR U32582 ( .A(p_input[1843]), .B(p_input[2067]), .Z(n32546) );
  XOR U32583 ( .A(p_input[1844]), .B(n17297), .Z(n32626) );
  XOR U32584 ( .A(p_input[1845]), .B(p_input[2069]), .Z(n32550) );
  XOR U32585 ( .A(n32565), .B(n32627), .Z(n32623) );
  IV U32586 ( .A(n32551), .Z(n32627) );
  XOR U32587 ( .A(p_input[1825]), .B(p_input[2049]), .Z(n32551) );
  XNOR U32588 ( .A(n32628), .B(n32573), .Z(n32565) );
  XNOR U32589 ( .A(n32561), .B(n32560), .Z(n32573) );
  XNOR U32590 ( .A(n32629), .B(n32557), .Z(n32560) );
  XNOR U32591 ( .A(p_input[1850]), .B(p_input[2074]), .Z(n32557) );
  XOR U32592 ( .A(p_input[1851]), .B(n17300), .Z(n32629) );
  XOR U32593 ( .A(p_input[1852]), .B(p_input[2076]), .Z(n32561) );
  XOR U32594 ( .A(n32571), .B(n32630), .Z(n32628) );
  IV U32595 ( .A(n32562), .Z(n32630) );
  XOR U32596 ( .A(p_input[1841]), .B(p_input[2065]), .Z(n32562) );
  XNOR U32597 ( .A(n32631), .B(n32578), .Z(n32571) );
  XNOR U32598 ( .A(p_input[1855]), .B(n17303), .Z(n32578) );
  XOR U32599 ( .A(n32568), .B(n32577), .Z(n32631) );
  XOR U32600 ( .A(n32632), .B(n32574), .Z(n32577) );
  XOR U32601 ( .A(p_input[1853]), .B(p_input[2077]), .Z(n32574) );
  XOR U32602 ( .A(p_input[1854]), .B(n17305), .Z(n32632) );
  XOR U32603 ( .A(p_input[1849]), .B(p_input[2073]), .Z(n32568) );
  XOR U32604 ( .A(n32590), .B(n32589), .Z(n32555) );
  XNOR U32605 ( .A(n32633), .B(n32597), .Z(n32589) );
  XNOR U32606 ( .A(n32585), .B(n32584), .Z(n32597) );
  XNOR U32607 ( .A(n32634), .B(n32581), .Z(n32584) );
  XNOR U32608 ( .A(p_input[1835]), .B(p_input[2059]), .Z(n32581) );
  XOR U32609 ( .A(p_input[1836]), .B(n16451), .Z(n32634) );
  XOR U32610 ( .A(p_input[1837]), .B(p_input[2061]), .Z(n32585) );
  XOR U32611 ( .A(n32595), .B(n32635), .Z(n32633) );
  IV U32612 ( .A(n32586), .Z(n32635) );
  XOR U32613 ( .A(p_input[1826]), .B(p_input[2050]), .Z(n32586) );
  XNOR U32614 ( .A(n32636), .B(n32602), .Z(n32595) );
  XNOR U32615 ( .A(p_input[1840]), .B(n16454), .Z(n32602) );
  XOR U32616 ( .A(n32592), .B(n32601), .Z(n32636) );
  XOR U32617 ( .A(n32637), .B(n32598), .Z(n32601) );
  XOR U32618 ( .A(p_input[1838]), .B(p_input[2062]), .Z(n32598) );
  XOR U32619 ( .A(p_input[1839]), .B(n16456), .Z(n32637) );
  XOR U32620 ( .A(p_input[1834]), .B(p_input[2058]), .Z(n32592) );
  XOR U32621 ( .A(n32609), .B(n32607), .Z(n32590) );
  XNOR U32622 ( .A(n32638), .B(n32614), .Z(n32607) );
  XOR U32623 ( .A(p_input[1833]), .B(p_input[2057]), .Z(n32614) );
  XOR U32624 ( .A(n32604), .B(n32613), .Z(n32638) );
  XOR U32625 ( .A(n32639), .B(n32610), .Z(n32613) );
  XOR U32626 ( .A(p_input[1831]), .B(p_input[2055]), .Z(n32610) );
  XOR U32627 ( .A(p_input[1832]), .B(n17312), .Z(n32639) );
  XOR U32628 ( .A(p_input[1827]), .B(p_input[2051]), .Z(n32604) );
  XNOR U32629 ( .A(n32619), .B(n32618), .Z(n32609) );
  XOR U32630 ( .A(n32640), .B(n32615), .Z(n32618) );
  XOR U32631 ( .A(p_input[1828]), .B(p_input[2052]), .Z(n32615) );
  XOR U32632 ( .A(p_input[1829]), .B(n17314), .Z(n32640) );
  XOR U32633 ( .A(p_input[1830]), .B(p_input[2054]), .Z(n32619) );
  XNOR U32634 ( .A(n32641), .B(n32642), .Z(n32432) );
  AND U32635 ( .A(n694), .B(n32643), .Z(n32642) );
  XNOR U32636 ( .A(n32644), .B(n32645), .Z(n694) );
  AND U32637 ( .A(n32646), .B(n32647), .Z(n32645) );
  XNOR U32638 ( .A(n32644), .B(n32385), .Z(n32647) );
  XOR U32639 ( .A(n32644), .B(n32382), .Z(n32646) );
  XOR U32640 ( .A(n32648), .B(n32649), .Z(n32644) );
  AND U32641 ( .A(n32650), .B(n32651), .Z(n32649) );
  XNOR U32642 ( .A(n32455), .B(n32648), .Z(n32651) );
  XOR U32643 ( .A(n32648), .B(n32396), .Z(n32650) );
  XOR U32644 ( .A(n32652), .B(n32653), .Z(n32648) );
  AND U32645 ( .A(n32654), .B(n32655), .Z(n32653) );
  XNOR U32646 ( .A(n32480), .B(n32652), .Z(n32655) );
  XOR U32647 ( .A(n32652), .B(n32407), .Z(n32654) );
  XOR U32648 ( .A(n32656), .B(n32657), .Z(n32652) );
  AND U32649 ( .A(n32658), .B(n32659), .Z(n32657) );
  XOR U32650 ( .A(n32656), .B(n32417), .Z(n32658) );
  XOR U32651 ( .A(n32660), .B(n32661), .Z(n32371) );
  AND U32652 ( .A(n698), .B(n32643), .Z(n32661) );
  XNOR U32653 ( .A(n32641), .B(n32660), .Z(n32643) );
  XNOR U32654 ( .A(n32662), .B(n32663), .Z(n698) );
  AND U32655 ( .A(n32664), .B(n32665), .Z(n32663) );
  XNOR U32656 ( .A(n32385), .B(n32662), .Z(n32665) );
  XOR U32657 ( .A(n32666), .B(n32667), .Z(n32385) );
  AND U32658 ( .A(n32668), .B(n701), .Z(n32667) );
  NOR U32659 ( .A(n32669), .B(n32666), .Z(n32668) );
  XOR U32660 ( .A(n32662), .B(n32382), .Z(n32664) );
  IV U32661 ( .A(n32386), .Z(n32382) );
  AND U32662 ( .A(n32670), .B(n32671), .Z(n32386) );
  XOR U32663 ( .A(n32672), .B(n32673), .Z(n32662) );
  AND U32664 ( .A(n32674), .B(n32675), .Z(n32673) );
  XNOR U32665 ( .A(n32672), .B(n32455), .Z(n32675) );
  XNOR U32666 ( .A(n32676), .B(n32677), .Z(n32455) );
  AND U32667 ( .A(n701), .B(n32678), .Z(n32677) );
  XOR U32668 ( .A(n32679), .B(n32676), .Z(n32678) );
  XNOR U32669 ( .A(n32680), .B(n32672), .Z(n32674) );
  IV U32670 ( .A(n32396), .Z(n32680) );
  XOR U32671 ( .A(n32681), .B(n32682), .Z(n32396) );
  AND U32672 ( .A(n709), .B(n32683), .Z(n32682) );
  XOR U32673 ( .A(n32684), .B(n32685), .Z(n32672) );
  AND U32674 ( .A(n32686), .B(n32687), .Z(n32685) );
  XNOR U32675 ( .A(n32684), .B(n32480), .Z(n32687) );
  XNOR U32676 ( .A(n32688), .B(n32689), .Z(n32480) );
  AND U32677 ( .A(n701), .B(n32690), .Z(n32689) );
  XNOR U32678 ( .A(n32691), .B(n32688), .Z(n32690) );
  XOR U32679 ( .A(n32407), .B(n32684), .Z(n32686) );
  XOR U32680 ( .A(n32692), .B(n32693), .Z(n32407) );
  AND U32681 ( .A(n709), .B(n32694), .Z(n32693) );
  XOR U32682 ( .A(n32656), .B(n32695), .Z(n32684) );
  AND U32683 ( .A(n32696), .B(n32659), .Z(n32695) );
  XNOR U32684 ( .A(n32526), .B(n32656), .Z(n32659) );
  XNOR U32685 ( .A(n32697), .B(n32698), .Z(n32526) );
  AND U32686 ( .A(n701), .B(n32699), .Z(n32698) );
  XOR U32687 ( .A(n32700), .B(n32697), .Z(n32699) );
  XNOR U32688 ( .A(n32701), .B(n32656), .Z(n32696) );
  IV U32689 ( .A(n32417), .Z(n32701) );
  XOR U32690 ( .A(n32702), .B(n32703), .Z(n32417) );
  AND U32691 ( .A(n709), .B(n32704), .Z(n32703) );
  XOR U32692 ( .A(n32705), .B(n32706), .Z(n32656) );
  AND U32693 ( .A(n32707), .B(n32708), .Z(n32706) );
  XNOR U32694 ( .A(n32705), .B(n32620), .Z(n32708) );
  XNOR U32695 ( .A(n32709), .B(n32710), .Z(n32620) );
  AND U32696 ( .A(n701), .B(n32711), .Z(n32710) );
  XNOR U32697 ( .A(n32712), .B(n32709), .Z(n32711) );
  XNOR U32698 ( .A(n32713), .B(n32705), .Z(n32707) );
  IV U32699 ( .A(n32429), .Z(n32713) );
  XOR U32700 ( .A(n32714), .B(n32715), .Z(n32429) );
  AND U32701 ( .A(n709), .B(n32716), .Z(n32715) );
  AND U32702 ( .A(n32660), .B(n32641), .Z(n32705) );
  XNOR U32703 ( .A(n32717), .B(n32718), .Z(n32641) );
  AND U32704 ( .A(n701), .B(n32719), .Z(n32718) );
  XNOR U32705 ( .A(n32720), .B(n32717), .Z(n32719) );
  XNOR U32706 ( .A(n32721), .B(n32722), .Z(n701) );
  NOR U32707 ( .A(n32723), .B(n32724), .Z(n32722) );
  XNOR U32708 ( .A(n32721), .B(n32666), .Z(n32724) );
  NOR U32709 ( .A(n32670), .B(n32671), .Z(n32666) );
  NOR U32710 ( .A(n32721), .B(n32669), .Z(n32723) );
  AND U32711 ( .A(n32725), .B(n32726), .Z(n32669) );
  XOR U32712 ( .A(n32727), .B(n32728), .Z(n32721) );
  AND U32713 ( .A(n32729), .B(n32730), .Z(n32728) );
  XNOR U32714 ( .A(n32727), .B(n32725), .Z(n32730) );
  IV U32715 ( .A(n32679), .Z(n32725) );
  XOR U32716 ( .A(n32731), .B(n32732), .Z(n32679) );
  XOR U32717 ( .A(n32733), .B(n32726), .Z(n32732) );
  AND U32718 ( .A(n32691), .B(n32734), .Z(n32726) );
  AND U32719 ( .A(n32735), .B(n32736), .Z(n32733) );
  XOR U32720 ( .A(n32737), .B(n32731), .Z(n32735) );
  XNOR U32721 ( .A(n32676), .B(n32727), .Z(n32729) );
  XNOR U32722 ( .A(n32738), .B(n32739), .Z(n32676) );
  AND U32723 ( .A(n705), .B(n32683), .Z(n32739) );
  XOR U32724 ( .A(n32738), .B(n32681), .Z(n32683) );
  XOR U32725 ( .A(n32740), .B(n32741), .Z(n32727) );
  AND U32726 ( .A(n32742), .B(n32743), .Z(n32741) );
  XNOR U32727 ( .A(n32740), .B(n32691), .Z(n32743) );
  XOR U32728 ( .A(n32744), .B(n32736), .Z(n32691) );
  XNOR U32729 ( .A(n32745), .B(n32731), .Z(n32736) );
  XOR U32730 ( .A(n32746), .B(n32747), .Z(n32731) );
  AND U32731 ( .A(n32748), .B(n32749), .Z(n32747) );
  XOR U32732 ( .A(n32750), .B(n32746), .Z(n32748) );
  XNOR U32733 ( .A(n32751), .B(n32752), .Z(n32745) );
  AND U32734 ( .A(n32753), .B(n32754), .Z(n32752) );
  XOR U32735 ( .A(n32751), .B(n32755), .Z(n32753) );
  XNOR U32736 ( .A(n32737), .B(n32734), .Z(n32744) );
  AND U32737 ( .A(n32756), .B(n32757), .Z(n32734) );
  XOR U32738 ( .A(n32758), .B(n32759), .Z(n32737) );
  AND U32739 ( .A(n32760), .B(n32761), .Z(n32759) );
  XOR U32740 ( .A(n32758), .B(n32762), .Z(n32760) );
  XNOR U32741 ( .A(n32688), .B(n32740), .Z(n32742) );
  XNOR U32742 ( .A(n32763), .B(n32764), .Z(n32688) );
  AND U32743 ( .A(n705), .B(n32694), .Z(n32764) );
  XOR U32744 ( .A(n32763), .B(n32692), .Z(n32694) );
  XOR U32745 ( .A(n32765), .B(n32766), .Z(n32740) );
  AND U32746 ( .A(n32767), .B(n32768), .Z(n32766) );
  XNOR U32747 ( .A(n32765), .B(n32756), .Z(n32768) );
  IV U32748 ( .A(n32700), .Z(n32756) );
  XNOR U32749 ( .A(n32769), .B(n32749), .Z(n32700) );
  XNOR U32750 ( .A(n32770), .B(n32755), .Z(n32749) );
  XOR U32751 ( .A(n32771), .B(n32772), .Z(n32755) );
  AND U32752 ( .A(n32773), .B(n32774), .Z(n32772) );
  XOR U32753 ( .A(n32771), .B(n32775), .Z(n32773) );
  XNOR U32754 ( .A(n32754), .B(n32746), .Z(n32770) );
  XOR U32755 ( .A(n32776), .B(n32777), .Z(n32746) );
  AND U32756 ( .A(n32778), .B(n32779), .Z(n32777) );
  XNOR U32757 ( .A(n32780), .B(n32776), .Z(n32778) );
  XNOR U32758 ( .A(n32781), .B(n32751), .Z(n32754) );
  XOR U32759 ( .A(n32782), .B(n32783), .Z(n32751) );
  AND U32760 ( .A(n32784), .B(n32785), .Z(n32783) );
  XOR U32761 ( .A(n32782), .B(n32786), .Z(n32784) );
  XNOR U32762 ( .A(n32787), .B(n32788), .Z(n32781) );
  AND U32763 ( .A(n32789), .B(n32790), .Z(n32788) );
  XNOR U32764 ( .A(n32787), .B(n32791), .Z(n32789) );
  XNOR U32765 ( .A(n32750), .B(n32757), .Z(n32769) );
  AND U32766 ( .A(n32712), .B(n32792), .Z(n32757) );
  XOR U32767 ( .A(n32762), .B(n32761), .Z(n32750) );
  XNOR U32768 ( .A(n32793), .B(n32758), .Z(n32761) );
  XOR U32769 ( .A(n32794), .B(n32795), .Z(n32758) );
  AND U32770 ( .A(n32796), .B(n32797), .Z(n32795) );
  XOR U32771 ( .A(n32794), .B(n32798), .Z(n32796) );
  XNOR U32772 ( .A(n32799), .B(n32800), .Z(n32793) );
  AND U32773 ( .A(n32801), .B(n32802), .Z(n32800) );
  XOR U32774 ( .A(n32799), .B(n32803), .Z(n32801) );
  XOR U32775 ( .A(n32804), .B(n32805), .Z(n32762) );
  AND U32776 ( .A(n32806), .B(n32807), .Z(n32805) );
  XOR U32777 ( .A(n32804), .B(n32808), .Z(n32806) );
  XNOR U32778 ( .A(n32697), .B(n32765), .Z(n32767) );
  XNOR U32779 ( .A(n32809), .B(n32810), .Z(n32697) );
  AND U32780 ( .A(n705), .B(n32704), .Z(n32810) );
  XOR U32781 ( .A(n32809), .B(n32702), .Z(n32704) );
  XOR U32782 ( .A(n32811), .B(n32812), .Z(n32765) );
  AND U32783 ( .A(n32813), .B(n32814), .Z(n32812) );
  XNOR U32784 ( .A(n32811), .B(n32712), .Z(n32814) );
  XOR U32785 ( .A(n32815), .B(n32779), .Z(n32712) );
  XNOR U32786 ( .A(n32816), .B(n32786), .Z(n32779) );
  XOR U32787 ( .A(n32775), .B(n32774), .Z(n32786) );
  XNOR U32788 ( .A(n32817), .B(n32771), .Z(n32774) );
  XOR U32789 ( .A(n32818), .B(n32819), .Z(n32771) );
  AND U32790 ( .A(n32820), .B(n32821), .Z(n32819) );
  XNOR U32791 ( .A(n32822), .B(n32823), .Z(n32820) );
  IV U32792 ( .A(n32818), .Z(n32822) );
  XNOR U32793 ( .A(n32824), .B(n32825), .Z(n32817) );
  NOR U32794 ( .A(n32826), .B(n32827), .Z(n32825) );
  XNOR U32795 ( .A(n32824), .B(n32828), .Z(n32826) );
  XOR U32796 ( .A(n32829), .B(n32830), .Z(n32775) );
  NOR U32797 ( .A(n32831), .B(n32832), .Z(n32830) );
  XNOR U32798 ( .A(n32829), .B(n32833), .Z(n32831) );
  XNOR U32799 ( .A(n32785), .B(n32776), .Z(n32816) );
  XOR U32800 ( .A(n32834), .B(n32835), .Z(n32776) );
  AND U32801 ( .A(n32836), .B(n32837), .Z(n32835) );
  XOR U32802 ( .A(n32834), .B(n32838), .Z(n32836) );
  XOR U32803 ( .A(n32839), .B(n32791), .Z(n32785) );
  XOR U32804 ( .A(n32840), .B(n32841), .Z(n32791) );
  NOR U32805 ( .A(n32842), .B(n32843), .Z(n32841) );
  XOR U32806 ( .A(n32840), .B(n32844), .Z(n32842) );
  XNOR U32807 ( .A(n32790), .B(n32782), .Z(n32839) );
  XOR U32808 ( .A(n32845), .B(n32846), .Z(n32782) );
  AND U32809 ( .A(n32847), .B(n32848), .Z(n32846) );
  XOR U32810 ( .A(n32845), .B(n32849), .Z(n32847) );
  XNOR U32811 ( .A(n32850), .B(n32787), .Z(n32790) );
  XOR U32812 ( .A(n32851), .B(n32852), .Z(n32787) );
  AND U32813 ( .A(n32853), .B(n32854), .Z(n32852) );
  XNOR U32814 ( .A(n32855), .B(n32856), .Z(n32853) );
  IV U32815 ( .A(n32851), .Z(n32855) );
  XNOR U32816 ( .A(n32857), .B(n32858), .Z(n32850) );
  NOR U32817 ( .A(n32859), .B(n32860), .Z(n32858) );
  XNOR U32818 ( .A(n32857), .B(n32861), .Z(n32859) );
  XOR U32819 ( .A(n32780), .B(n32792), .Z(n32815) );
  NOR U32820 ( .A(n32720), .B(n32862), .Z(n32792) );
  XNOR U32821 ( .A(n32798), .B(n32797), .Z(n32780) );
  XNOR U32822 ( .A(n32863), .B(n32803), .Z(n32797) );
  XNOR U32823 ( .A(n32864), .B(n32865), .Z(n32803) );
  NOR U32824 ( .A(n32866), .B(n32867), .Z(n32865) );
  XOR U32825 ( .A(n32864), .B(n32868), .Z(n32866) );
  XNOR U32826 ( .A(n32802), .B(n32794), .Z(n32863) );
  XOR U32827 ( .A(n32869), .B(n32870), .Z(n32794) );
  AND U32828 ( .A(n32871), .B(n32872), .Z(n32870) );
  XOR U32829 ( .A(n32869), .B(n32873), .Z(n32871) );
  XNOR U32830 ( .A(n32874), .B(n32799), .Z(n32802) );
  XOR U32831 ( .A(n32875), .B(n32876), .Z(n32799) );
  AND U32832 ( .A(n32877), .B(n32878), .Z(n32876) );
  XNOR U32833 ( .A(n32879), .B(n32880), .Z(n32877) );
  IV U32834 ( .A(n32875), .Z(n32879) );
  XNOR U32835 ( .A(n32881), .B(n32882), .Z(n32874) );
  NOR U32836 ( .A(n32883), .B(n32884), .Z(n32882) );
  XNOR U32837 ( .A(n32881), .B(n32885), .Z(n32883) );
  XOR U32838 ( .A(n32808), .B(n32807), .Z(n32798) );
  XNOR U32839 ( .A(n32886), .B(n32804), .Z(n32807) );
  XOR U32840 ( .A(n32887), .B(n32888), .Z(n32804) );
  AND U32841 ( .A(n32889), .B(n32890), .Z(n32888) );
  XNOR U32842 ( .A(n32891), .B(n32892), .Z(n32889) );
  IV U32843 ( .A(n32887), .Z(n32891) );
  XNOR U32844 ( .A(n32893), .B(n32894), .Z(n32886) );
  NOR U32845 ( .A(n32895), .B(n32896), .Z(n32894) );
  XNOR U32846 ( .A(n32893), .B(n32897), .Z(n32895) );
  XOR U32847 ( .A(n32898), .B(n32899), .Z(n32808) );
  NOR U32848 ( .A(n32900), .B(n32901), .Z(n32899) );
  XNOR U32849 ( .A(n32898), .B(n32902), .Z(n32900) );
  XNOR U32850 ( .A(n32709), .B(n32811), .Z(n32813) );
  XNOR U32851 ( .A(n32903), .B(n32904), .Z(n32709) );
  AND U32852 ( .A(n705), .B(n32716), .Z(n32904) );
  XOR U32853 ( .A(n32903), .B(n32714), .Z(n32716) );
  AND U32854 ( .A(n32717), .B(n32720), .Z(n32811) );
  XOR U32855 ( .A(n32905), .B(n32862), .Z(n32720) );
  XNOR U32856 ( .A(p_input[1856]), .B(p_input[2048]), .Z(n32862) );
  XNOR U32857 ( .A(n32838), .B(n32837), .Z(n32905) );
  XNOR U32858 ( .A(n32906), .B(n32849), .Z(n32837) );
  XOR U32859 ( .A(n32823), .B(n32821), .Z(n32849) );
  XNOR U32860 ( .A(n32907), .B(n32828), .Z(n32821) );
  XOR U32861 ( .A(p_input[1880]), .B(p_input[2072]), .Z(n32828) );
  XOR U32862 ( .A(n32818), .B(n32827), .Z(n32907) );
  XOR U32863 ( .A(n32908), .B(n32824), .Z(n32827) );
  XOR U32864 ( .A(p_input[1878]), .B(p_input[2070]), .Z(n32824) );
  XOR U32865 ( .A(p_input[1879]), .B(n17295), .Z(n32908) );
  XOR U32866 ( .A(p_input[1874]), .B(p_input[2066]), .Z(n32818) );
  XNOR U32867 ( .A(n32833), .B(n32832), .Z(n32823) );
  XOR U32868 ( .A(n32909), .B(n32829), .Z(n32832) );
  XOR U32869 ( .A(p_input[1875]), .B(p_input[2067]), .Z(n32829) );
  XOR U32870 ( .A(p_input[1876]), .B(n17297), .Z(n32909) );
  XOR U32871 ( .A(p_input[1877]), .B(p_input[2069]), .Z(n32833) );
  XOR U32872 ( .A(n32848), .B(n32910), .Z(n32906) );
  IV U32873 ( .A(n32834), .Z(n32910) );
  XOR U32874 ( .A(p_input[1857]), .B(p_input[2049]), .Z(n32834) );
  XNOR U32875 ( .A(n32911), .B(n32856), .Z(n32848) );
  XNOR U32876 ( .A(n32844), .B(n32843), .Z(n32856) );
  XNOR U32877 ( .A(n32912), .B(n32840), .Z(n32843) );
  XNOR U32878 ( .A(p_input[1882]), .B(p_input[2074]), .Z(n32840) );
  XOR U32879 ( .A(p_input[1883]), .B(n17300), .Z(n32912) );
  XOR U32880 ( .A(p_input[1884]), .B(p_input[2076]), .Z(n32844) );
  XOR U32881 ( .A(n32854), .B(n32913), .Z(n32911) );
  IV U32882 ( .A(n32845), .Z(n32913) );
  XOR U32883 ( .A(p_input[1873]), .B(p_input[2065]), .Z(n32845) );
  XNOR U32884 ( .A(n32914), .B(n32861), .Z(n32854) );
  XNOR U32885 ( .A(p_input[1887]), .B(n17303), .Z(n32861) );
  XOR U32886 ( .A(n32851), .B(n32860), .Z(n32914) );
  XOR U32887 ( .A(n32915), .B(n32857), .Z(n32860) );
  XOR U32888 ( .A(p_input[1885]), .B(p_input[2077]), .Z(n32857) );
  XOR U32889 ( .A(p_input[1886]), .B(n17305), .Z(n32915) );
  XOR U32890 ( .A(p_input[1881]), .B(p_input[2073]), .Z(n32851) );
  XOR U32891 ( .A(n32873), .B(n32872), .Z(n32838) );
  XNOR U32892 ( .A(n32916), .B(n32880), .Z(n32872) );
  XNOR U32893 ( .A(n32868), .B(n32867), .Z(n32880) );
  XNOR U32894 ( .A(n32917), .B(n32864), .Z(n32867) );
  XNOR U32895 ( .A(p_input[1867]), .B(p_input[2059]), .Z(n32864) );
  XOR U32896 ( .A(p_input[1868]), .B(n16451), .Z(n32917) );
  XOR U32897 ( .A(p_input[1869]), .B(p_input[2061]), .Z(n32868) );
  XOR U32898 ( .A(n32878), .B(n32918), .Z(n32916) );
  IV U32899 ( .A(n32869), .Z(n32918) );
  XOR U32900 ( .A(p_input[1858]), .B(p_input[2050]), .Z(n32869) );
  XNOR U32901 ( .A(n32919), .B(n32885), .Z(n32878) );
  XNOR U32902 ( .A(p_input[1872]), .B(n16454), .Z(n32885) );
  XOR U32903 ( .A(n32875), .B(n32884), .Z(n32919) );
  XOR U32904 ( .A(n32920), .B(n32881), .Z(n32884) );
  XOR U32905 ( .A(p_input[1870]), .B(p_input[2062]), .Z(n32881) );
  XOR U32906 ( .A(p_input[1871]), .B(n16456), .Z(n32920) );
  XOR U32907 ( .A(p_input[1866]), .B(p_input[2058]), .Z(n32875) );
  XOR U32908 ( .A(n32892), .B(n32890), .Z(n32873) );
  XNOR U32909 ( .A(n32921), .B(n32897), .Z(n32890) );
  XOR U32910 ( .A(p_input[1865]), .B(p_input[2057]), .Z(n32897) );
  XOR U32911 ( .A(n32887), .B(n32896), .Z(n32921) );
  XOR U32912 ( .A(n32922), .B(n32893), .Z(n32896) );
  XOR U32913 ( .A(p_input[1863]), .B(p_input[2055]), .Z(n32893) );
  XOR U32914 ( .A(p_input[1864]), .B(n17312), .Z(n32922) );
  XOR U32915 ( .A(p_input[1859]), .B(p_input[2051]), .Z(n32887) );
  XNOR U32916 ( .A(n32902), .B(n32901), .Z(n32892) );
  XOR U32917 ( .A(n32923), .B(n32898), .Z(n32901) );
  XOR U32918 ( .A(p_input[1860]), .B(p_input[2052]), .Z(n32898) );
  XOR U32919 ( .A(p_input[1861]), .B(n17314), .Z(n32923) );
  XOR U32920 ( .A(p_input[1862]), .B(p_input[2054]), .Z(n32902) );
  XNOR U32921 ( .A(n32924), .B(n32925), .Z(n32717) );
  AND U32922 ( .A(n705), .B(n32926), .Z(n32925) );
  XNOR U32923 ( .A(n32927), .B(n32928), .Z(n705) );
  NOR U32924 ( .A(n32929), .B(n32930), .Z(n32928) );
  XOR U32925 ( .A(n32671), .B(n32927), .Z(n32930) );
  NOR U32926 ( .A(n32927), .B(n32670), .Z(n32929) );
  XOR U32927 ( .A(n32931), .B(n32932), .Z(n32927) );
  AND U32928 ( .A(n32933), .B(n32934), .Z(n32932) );
  XNOR U32929 ( .A(n32738), .B(n32931), .Z(n32934) );
  XOR U32930 ( .A(n32931), .B(n32681), .Z(n32933) );
  XOR U32931 ( .A(n32935), .B(n32936), .Z(n32931) );
  AND U32932 ( .A(n32937), .B(n32938), .Z(n32936) );
  XNOR U32933 ( .A(n32763), .B(n32935), .Z(n32938) );
  XOR U32934 ( .A(n32935), .B(n32692), .Z(n32937) );
  XOR U32935 ( .A(n32939), .B(n32940), .Z(n32935) );
  AND U32936 ( .A(n32941), .B(n32942), .Z(n32940) );
  XOR U32937 ( .A(n32939), .B(n32702), .Z(n32941) );
  XOR U32938 ( .A(n32943), .B(n32944), .Z(n32660) );
  AND U32939 ( .A(n709), .B(n32926), .Z(n32944) );
  XNOR U32940 ( .A(n32924), .B(n32943), .Z(n32926) );
  XNOR U32941 ( .A(n32945), .B(n32946), .Z(n709) );
  NOR U32942 ( .A(n32947), .B(n32948), .Z(n32946) );
  XNOR U32943 ( .A(n32671), .B(n32949), .Z(n32948) );
  IV U32944 ( .A(n32945), .Z(n32949) );
  AND U32945 ( .A(n32950), .B(n32951), .Z(n32671) );
  NOR U32946 ( .A(n32945), .B(n32670), .Z(n32947) );
  AND U32947 ( .A(n32952), .B(n32953), .Z(n32670) );
  IV U32948 ( .A(n32954), .Z(n32952) );
  XOR U32949 ( .A(n32955), .B(n32956), .Z(n32945) );
  AND U32950 ( .A(n32957), .B(n32958), .Z(n32956) );
  XNOR U32951 ( .A(n32955), .B(n32738), .Z(n32958) );
  XNOR U32952 ( .A(n32959), .B(n32960), .Z(n32738) );
  AND U32953 ( .A(n712), .B(n32961), .Z(n32960) );
  XOR U32954 ( .A(n32962), .B(n32959), .Z(n32961) );
  XNOR U32955 ( .A(n32963), .B(n32955), .Z(n32957) );
  IV U32956 ( .A(n32681), .Z(n32963) );
  XOR U32957 ( .A(n32964), .B(n32965), .Z(n32681) );
  AND U32958 ( .A(n720), .B(n32966), .Z(n32965) );
  XOR U32959 ( .A(n32967), .B(n32968), .Z(n32955) );
  AND U32960 ( .A(n32969), .B(n32970), .Z(n32968) );
  XNOR U32961 ( .A(n32967), .B(n32763), .Z(n32970) );
  XNOR U32962 ( .A(n32971), .B(n32972), .Z(n32763) );
  AND U32963 ( .A(n712), .B(n32973), .Z(n32972) );
  XNOR U32964 ( .A(n32974), .B(n32971), .Z(n32973) );
  XOR U32965 ( .A(n32692), .B(n32967), .Z(n32969) );
  XOR U32966 ( .A(n32975), .B(n32976), .Z(n32692) );
  AND U32967 ( .A(n720), .B(n32977), .Z(n32976) );
  XOR U32968 ( .A(n32939), .B(n32978), .Z(n32967) );
  AND U32969 ( .A(n32979), .B(n32942), .Z(n32978) );
  XNOR U32970 ( .A(n32809), .B(n32939), .Z(n32942) );
  XNOR U32971 ( .A(n32980), .B(n32981), .Z(n32809) );
  AND U32972 ( .A(n712), .B(n32982), .Z(n32981) );
  XOR U32973 ( .A(n32983), .B(n32980), .Z(n32982) );
  XNOR U32974 ( .A(n32984), .B(n32939), .Z(n32979) );
  IV U32975 ( .A(n32702), .Z(n32984) );
  XOR U32976 ( .A(n32985), .B(n32986), .Z(n32702) );
  AND U32977 ( .A(n720), .B(n32987), .Z(n32986) );
  XOR U32978 ( .A(n32988), .B(n32989), .Z(n32939) );
  AND U32979 ( .A(n32990), .B(n32991), .Z(n32989) );
  XNOR U32980 ( .A(n32988), .B(n32903), .Z(n32991) );
  XNOR U32981 ( .A(n32992), .B(n32993), .Z(n32903) );
  AND U32982 ( .A(n712), .B(n32994), .Z(n32993) );
  XNOR U32983 ( .A(n32995), .B(n32992), .Z(n32994) );
  XNOR U32984 ( .A(n32996), .B(n32988), .Z(n32990) );
  IV U32985 ( .A(n32714), .Z(n32996) );
  XOR U32986 ( .A(n32997), .B(n32998), .Z(n32714) );
  AND U32987 ( .A(n720), .B(n32999), .Z(n32998) );
  AND U32988 ( .A(n32943), .B(n32924), .Z(n32988) );
  XNOR U32989 ( .A(n33000), .B(n33001), .Z(n32924) );
  AND U32990 ( .A(n712), .B(n33002), .Z(n33001) );
  XNOR U32991 ( .A(n33003), .B(n33000), .Z(n33002) );
  XNOR U32992 ( .A(n33004), .B(n33005), .Z(n712) );
  NOR U32993 ( .A(n33006), .B(n33007), .Z(n33005) );
  XNOR U32994 ( .A(n33004), .B(n32954), .Z(n33007) );
  NOR U32995 ( .A(n32950), .B(n32951), .Z(n32954) );
  NOR U32996 ( .A(n33004), .B(n32953), .Z(n33006) );
  AND U32997 ( .A(n33008), .B(n33009), .Z(n32953) );
  XOR U32998 ( .A(n33010), .B(n33011), .Z(n33004) );
  AND U32999 ( .A(n33012), .B(n33013), .Z(n33011) );
  XNOR U33000 ( .A(n33010), .B(n33008), .Z(n33013) );
  IV U33001 ( .A(n32962), .Z(n33008) );
  XOR U33002 ( .A(n33014), .B(n33015), .Z(n32962) );
  XOR U33003 ( .A(n33016), .B(n33009), .Z(n33015) );
  AND U33004 ( .A(n32974), .B(n33017), .Z(n33009) );
  AND U33005 ( .A(n33018), .B(n33019), .Z(n33016) );
  XOR U33006 ( .A(n33020), .B(n33014), .Z(n33018) );
  XNOR U33007 ( .A(n32959), .B(n33010), .Z(n33012) );
  XNOR U33008 ( .A(n33021), .B(n33022), .Z(n32959) );
  AND U33009 ( .A(n716), .B(n32966), .Z(n33022) );
  XOR U33010 ( .A(n33021), .B(n32964), .Z(n32966) );
  XOR U33011 ( .A(n33023), .B(n33024), .Z(n33010) );
  AND U33012 ( .A(n33025), .B(n33026), .Z(n33024) );
  XNOR U33013 ( .A(n33023), .B(n32974), .Z(n33026) );
  XOR U33014 ( .A(n33027), .B(n33019), .Z(n32974) );
  XNOR U33015 ( .A(n33028), .B(n33014), .Z(n33019) );
  XOR U33016 ( .A(n33029), .B(n33030), .Z(n33014) );
  AND U33017 ( .A(n33031), .B(n33032), .Z(n33030) );
  XOR U33018 ( .A(n33033), .B(n33029), .Z(n33031) );
  XNOR U33019 ( .A(n33034), .B(n33035), .Z(n33028) );
  AND U33020 ( .A(n33036), .B(n33037), .Z(n33035) );
  XOR U33021 ( .A(n33034), .B(n33038), .Z(n33036) );
  XNOR U33022 ( .A(n33020), .B(n33017), .Z(n33027) );
  AND U33023 ( .A(n33039), .B(n33040), .Z(n33017) );
  XOR U33024 ( .A(n33041), .B(n33042), .Z(n33020) );
  AND U33025 ( .A(n33043), .B(n33044), .Z(n33042) );
  XOR U33026 ( .A(n33041), .B(n33045), .Z(n33043) );
  XNOR U33027 ( .A(n32971), .B(n33023), .Z(n33025) );
  XNOR U33028 ( .A(n33046), .B(n33047), .Z(n32971) );
  AND U33029 ( .A(n716), .B(n32977), .Z(n33047) );
  XOR U33030 ( .A(n33046), .B(n32975), .Z(n32977) );
  XOR U33031 ( .A(n33048), .B(n33049), .Z(n33023) );
  AND U33032 ( .A(n33050), .B(n33051), .Z(n33049) );
  XNOR U33033 ( .A(n33048), .B(n33039), .Z(n33051) );
  IV U33034 ( .A(n32983), .Z(n33039) );
  XNOR U33035 ( .A(n33052), .B(n33032), .Z(n32983) );
  XNOR U33036 ( .A(n33053), .B(n33038), .Z(n33032) );
  XOR U33037 ( .A(n33054), .B(n33055), .Z(n33038) );
  AND U33038 ( .A(n33056), .B(n33057), .Z(n33055) );
  XOR U33039 ( .A(n33054), .B(n33058), .Z(n33056) );
  XNOR U33040 ( .A(n33037), .B(n33029), .Z(n33053) );
  XOR U33041 ( .A(n33059), .B(n33060), .Z(n33029) );
  AND U33042 ( .A(n33061), .B(n33062), .Z(n33060) );
  XNOR U33043 ( .A(n33063), .B(n33059), .Z(n33061) );
  XNOR U33044 ( .A(n33064), .B(n33034), .Z(n33037) );
  XOR U33045 ( .A(n33065), .B(n33066), .Z(n33034) );
  AND U33046 ( .A(n33067), .B(n33068), .Z(n33066) );
  XOR U33047 ( .A(n33065), .B(n33069), .Z(n33067) );
  XNOR U33048 ( .A(n33070), .B(n33071), .Z(n33064) );
  AND U33049 ( .A(n33072), .B(n33073), .Z(n33071) );
  XNOR U33050 ( .A(n33070), .B(n33074), .Z(n33072) );
  XNOR U33051 ( .A(n33033), .B(n33040), .Z(n33052) );
  AND U33052 ( .A(n32995), .B(n33075), .Z(n33040) );
  XOR U33053 ( .A(n33045), .B(n33044), .Z(n33033) );
  XNOR U33054 ( .A(n33076), .B(n33041), .Z(n33044) );
  XOR U33055 ( .A(n33077), .B(n33078), .Z(n33041) );
  AND U33056 ( .A(n33079), .B(n33080), .Z(n33078) );
  XOR U33057 ( .A(n33077), .B(n33081), .Z(n33079) );
  XNOR U33058 ( .A(n33082), .B(n33083), .Z(n33076) );
  AND U33059 ( .A(n33084), .B(n33085), .Z(n33083) );
  XOR U33060 ( .A(n33082), .B(n33086), .Z(n33084) );
  XOR U33061 ( .A(n33087), .B(n33088), .Z(n33045) );
  AND U33062 ( .A(n33089), .B(n33090), .Z(n33088) );
  XOR U33063 ( .A(n33087), .B(n33091), .Z(n33089) );
  XNOR U33064 ( .A(n32980), .B(n33048), .Z(n33050) );
  XNOR U33065 ( .A(n33092), .B(n33093), .Z(n32980) );
  AND U33066 ( .A(n716), .B(n32987), .Z(n33093) );
  XOR U33067 ( .A(n33092), .B(n32985), .Z(n32987) );
  XOR U33068 ( .A(n33094), .B(n33095), .Z(n33048) );
  AND U33069 ( .A(n33096), .B(n33097), .Z(n33095) );
  XNOR U33070 ( .A(n33094), .B(n32995), .Z(n33097) );
  XOR U33071 ( .A(n33098), .B(n33062), .Z(n32995) );
  XNOR U33072 ( .A(n33099), .B(n33069), .Z(n33062) );
  XOR U33073 ( .A(n33058), .B(n33057), .Z(n33069) );
  XNOR U33074 ( .A(n33100), .B(n33054), .Z(n33057) );
  XOR U33075 ( .A(n33101), .B(n33102), .Z(n33054) );
  AND U33076 ( .A(n33103), .B(n33104), .Z(n33102) );
  XNOR U33077 ( .A(n33105), .B(n33106), .Z(n33103) );
  IV U33078 ( .A(n33101), .Z(n33105) );
  XNOR U33079 ( .A(n33107), .B(n33108), .Z(n33100) );
  NOR U33080 ( .A(n33109), .B(n33110), .Z(n33108) );
  XNOR U33081 ( .A(n33107), .B(n33111), .Z(n33109) );
  XOR U33082 ( .A(n33112), .B(n33113), .Z(n33058) );
  NOR U33083 ( .A(n33114), .B(n33115), .Z(n33113) );
  XNOR U33084 ( .A(n33112), .B(n33116), .Z(n33114) );
  XNOR U33085 ( .A(n33068), .B(n33059), .Z(n33099) );
  XOR U33086 ( .A(n33117), .B(n33118), .Z(n33059) );
  AND U33087 ( .A(n33119), .B(n33120), .Z(n33118) );
  XOR U33088 ( .A(n33117), .B(n33121), .Z(n33119) );
  XOR U33089 ( .A(n33122), .B(n33074), .Z(n33068) );
  XOR U33090 ( .A(n33123), .B(n33124), .Z(n33074) );
  NOR U33091 ( .A(n33125), .B(n33126), .Z(n33124) );
  XOR U33092 ( .A(n33123), .B(n33127), .Z(n33125) );
  XNOR U33093 ( .A(n33073), .B(n33065), .Z(n33122) );
  XOR U33094 ( .A(n33128), .B(n33129), .Z(n33065) );
  AND U33095 ( .A(n33130), .B(n33131), .Z(n33129) );
  XOR U33096 ( .A(n33128), .B(n33132), .Z(n33130) );
  XNOR U33097 ( .A(n33133), .B(n33070), .Z(n33073) );
  XOR U33098 ( .A(n33134), .B(n33135), .Z(n33070) );
  AND U33099 ( .A(n33136), .B(n33137), .Z(n33135) );
  XNOR U33100 ( .A(n33138), .B(n33139), .Z(n33136) );
  IV U33101 ( .A(n33134), .Z(n33138) );
  XNOR U33102 ( .A(n33140), .B(n33141), .Z(n33133) );
  NOR U33103 ( .A(n33142), .B(n33143), .Z(n33141) );
  XNOR U33104 ( .A(n33140), .B(n33144), .Z(n33142) );
  XOR U33105 ( .A(n33063), .B(n33075), .Z(n33098) );
  NOR U33106 ( .A(n33003), .B(n33145), .Z(n33075) );
  XNOR U33107 ( .A(n33081), .B(n33080), .Z(n33063) );
  XNOR U33108 ( .A(n33146), .B(n33086), .Z(n33080) );
  XNOR U33109 ( .A(n33147), .B(n33148), .Z(n33086) );
  NOR U33110 ( .A(n33149), .B(n33150), .Z(n33148) );
  XOR U33111 ( .A(n33147), .B(n33151), .Z(n33149) );
  XNOR U33112 ( .A(n33085), .B(n33077), .Z(n33146) );
  XOR U33113 ( .A(n33152), .B(n33153), .Z(n33077) );
  AND U33114 ( .A(n33154), .B(n33155), .Z(n33153) );
  XOR U33115 ( .A(n33152), .B(n33156), .Z(n33154) );
  XNOR U33116 ( .A(n33157), .B(n33082), .Z(n33085) );
  XOR U33117 ( .A(n33158), .B(n33159), .Z(n33082) );
  AND U33118 ( .A(n33160), .B(n33161), .Z(n33159) );
  XNOR U33119 ( .A(n33162), .B(n33163), .Z(n33160) );
  IV U33120 ( .A(n33158), .Z(n33162) );
  XNOR U33121 ( .A(n33164), .B(n33165), .Z(n33157) );
  NOR U33122 ( .A(n33166), .B(n33167), .Z(n33165) );
  XNOR U33123 ( .A(n33164), .B(n33168), .Z(n33166) );
  XOR U33124 ( .A(n33091), .B(n33090), .Z(n33081) );
  XNOR U33125 ( .A(n33169), .B(n33087), .Z(n33090) );
  XOR U33126 ( .A(n33170), .B(n33171), .Z(n33087) );
  AND U33127 ( .A(n33172), .B(n33173), .Z(n33171) );
  XNOR U33128 ( .A(n33174), .B(n33175), .Z(n33172) );
  IV U33129 ( .A(n33170), .Z(n33174) );
  XNOR U33130 ( .A(n33176), .B(n33177), .Z(n33169) );
  NOR U33131 ( .A(n33178), .B(n33179), .Z(n33177) );
  XNOR U33132 ( .A(n33176), .B(n33180), .Z(n33178) );
  XOR U33133 ( .A(n33181), .B(n33182), .Z(n33091) );
  NOR U33134 ( .A(n33183), .B(n33184), .Z(n33182) );
  XNOR U33135 ( .A(n33181), .B(n33185), .Z(n33183) );
  XNOR U33136 ( .A(n32992), .B(n33094), .Z(n33096) );
  XNOR U33137 ( .A(n33186), .B(n33187), .Z(n32992) );
  AND U33138 ( .A(n716), .B(n32999), .Z(n33187) );
  XOR U33139 ( .A(n33186), .B(n32997), .Z(n32999) );
  AND U33140 ( .A(n33000), .B(n33003), .Z(n33094) );
  XOR U33141 ( .A(n33188), .B(n33145), .Z(n33003) );
  XNOR U33142 ( .A(p_input[1888]), .B(p_input[2048]), .Z(n33145) );
  XNOR U33143 ( .A(n33121), .B(n33120), .Z(n33188) );
  XNOR U33144 ( .A(n33189), .B(n33132), .Z(n33120) );
  XOR U33145 ( .A(n33106), .B(n33104), .Z(n33132) );
  XNOR U33146 ( .A(n33190), .B(n33111), .Z(n33104) );
  XOR U33147 ( .A(p_input[1912]), .B(p_input[2072]), .Z(n33111) );
  XOR U33148 ( .A(n33101), .B(n33110), .Z(n33190) );
  XOR U33149 ( .A(n33191), .B(n33107), .Z(n33110) );
  XOR U33150 ( .A(p_input[1910]), .B(p_input[2070]), .Z(n33107) );
  XOR U33151 ( .A(p_input[1911]), .B(n17295), .Z(n33191) );
  XOR U33152 ( .A(p_input[1906]), .B(p_input[2066]), .Z(n33101) );
  XNOR U33153 ( .A(n33116), .B(n33115), .Z(n33106) );
  XOR U33154 ( .A(n33192), .B(n33112), .Z(n33115) );
  XOR U33155 ( .A(p_input[1907]), .B(p_input[2067]), .Z(n33112) );
  XOR U33156 ( .A(p_input[1908]), .B(n17297), .Z(n33192) );
  XOR U33157 ( .A(p_input[1909]), .B(p_input[2069]), .Z(n33116) );
  XOR U33158 ( .A(n33131), .B(n33193), .Z(n33189) );
  IV U33159 ( .A(n33117), .Z(n33193) );
  XOR U33160 ( .A(p_input[1889]), .B(p_input[2049]), .Z(n33117) );
  XNOR U33161 ( .A(n33194), .B(n33139), .Z(n33131) );
  XNOR U33162 ( .A(n33127), .B(n33126), .Z(n33139) );
  XNOR U33163 ( .A(n33195), .B(n33123), .Z(n33126) );
  XNOR U33164 ( .A(p_input[1914]), .B(p_input[2074]), .Z(n33123) );
  XOR U33165 ( .A(p_input[1915]), .B(n17300), .Z(n33195) );
  XOR U33166 ( .A(p_input[1916]), .B(p_input[2076]), .Z(n33127) );
  XOR U33167 ( .A(n33137), .B(n33196), .Z(n33194) );
  IV U33168 ( .A(n33128), .Z(n33196) );
  XOR U33169 ( .A(p_input[1905]), .B(p_input[2065]), .Z(n33128) );
  XNOR U33170 ( .A(n33197), .B(n33144), .Z(n33137) );
  XNOR U33171 ( .A(p_input[1919]), .B(n17303), .Z(n33144) );
  XOR U33172 ( .A(n33134), .B(n33143), .Z(n33197) );
  XOR U33173 ( .A(n33198), .B(n33140), .Z(n33143) );
  XOR U33174 ( .A(p_input[1917]), .B(p_input[2077]), .Z(n33140) );
  XOR U33175 ( .A(p_input[1918]), .B(n17305), .Z(n33198) );
  XOR U33176 ( .A(p_input[1913]), .B(p_input[2073]), .Z(n33134) );
  XOR U33177 ( .A(n33156), .B(n33155), .Z(n33121) );
  XNOR U33178 ( .A(n33199), .B(n33163), .Z(n33155) );
  XNOR U33179 ( .A(n33151), .B(n33150), .Z(n33163) );
  XNOR U33180 ( .A(n33200), .B(n33147), .Z(n33150) );
  XNOR U33181 ( .A(p_input[1899]), .B(p_input[2059]), .Z(n33147) );
  XOR U33182 ( .A(p_input[1900]), .B(n16451), .Z(n33200) );
  XOR U33183 ( .A(p_input[1901]), .B(p_input[2061]), .Z(n33151) );
  XOR U33184 ( .A(n33161), .B(n33201), .Z(n33199) );
  IV U33185 ( .A(n33152), .Z(n33201) );
  XOR U33186 ( .A(p_input[1890]), .B(p_input[2050]), .Z(n33152) );
  XNOR U33187 ( .A(n33202), .B(n33168), .Z(n33161) );
  XNOR U33188 ( .A(p_input[1904]), .B(n16454), .Z(n33168) );
  XOR U33189 ( .A(n33158), .B(n33167), .Z(n33202) );
  XOR U33190 ( .A(n33203), .B(n33164), .Z(n33167) );
  XOR U33191 ( .A(p_input[1902]), .B(p_input[2062]), .Z(n33164) );
  XOR U33192 ( .A(p_input[1903]), .B(n16456), .Z(n33203) );
  XOR U33193 ( .A(p_input[1898]), .B(p_input[2058]), .Z(n33158) );
  XOR U33194 ( .A(n33175), .B(n33173), .Z(n33156) );
  XNOR U33195 ( .A(n33204), .B(n33180), .Z(n33173) );
  XOR U33196 ( .A(p_input[1897]), .B(p_input[2057]), .Z(n33180) );
  XOR U33197 ( .A(n33170), .B(n33179), .Z(n33204) );
  XOR U33198 ( .A(n33205), .B(n33176), .Z(n33179) );
  XOR U33199 ( .A(p_input[1895]), .B(p_input[2055]), .Z(n33176) );
  XOR U33200 ( .A(p_input[1896]), .B(n17312), .Z(n33205) );
  XOR U33201 ( .A(p_input[1891]), .B(p_input[2051]), .Z(n33170) );
  XNOR U33202 ( .A(n33185), .B(n33184), .Z(n33175) );
  XOR U33203 ( .A(n33206), .B(n33181), .Z(n33184) );
  XOR U33204 ( .A(p_input[1892]), .B(p_input[2052]), .Z(n33181) );
  XOR U33205 ( .A(p_input[1893]), .B(n17314), .Z(n33206) );
  XOR U33206 ( .A(p_input[1894]), .B(p_input[2054]), .Z(n33185) );
  XNOR U33207 ( .A(n33207), .B(n33208), .Z(n33000) );
  AND U33208 ( .A(n716), .B(n33209), .Z(n33208) );
  XNOR U33209 ( .A(n33210), .B(n33211), .Z(n716) );
  NOR U33210 ( .A(n33212), .B(n33213), .Z(n33211) );
  XOR U33211 ( .A(n32951), .B(n33210), .Z(n33213) );
  NOR U33212 ( .A(n33210), .B(n32950), .Z(n33212) );
  XOR U33213 ( .A(n33214), .B(n33215), .Z(n33210) );
  AND U33214 ( .A(n33216), .B(n33217), .Z(n33215) );
  XNOR U33215 ( .A(n33021), .B(n33214), .Z(n33217) );
  XOR U33216 ( .A(n33214), .B(n32964), .Z(n33216) );
  XOR U33217 ( .A(n33218), .B(n33219), .Z(n33214) );
  AND U33218 ( .A(n33220), .B(n33221), .Z(n33219) );
  XNOR U33219 ( .A(n33046), .B(n33218), .Z(n33221) );
  XOR U33220 ( .A(n33218), .B(n32975), .Z(n33220) );
  XOR U33221 ( .A(n33222), .B(n33223), .Z(n33218) );
  AND U33222 ( .A(n33224), .B(n33225), .Z(n33223) );
  XOR U33223 ( .A(n33222), .B(n32985), .Z(n33224) );
  XOR U33224 ( .A(n33226), .B(n33227), .Z(n32943) );
  AND U33225 ( .A(n720), .B(n33209), .Z(n33227) );
  XNOR U33226 ( .A(n33207), .B(n33226), .Z(n33209) );
  XNOR U33227 ( .A(n33228), .B(n33229), .Z(n720) );
  NOR U33228 ( .A(n33230), .B(n33231), .Z(n33229) );
  XNOR U33229 ( .A(n32951), .B(n33232), .Z(n33231) );
  IV U33230 ( .A(n33228), .Z(n33232) );
  AND U33231 ( .A(n33233), .B(n33234), .Z(n32951) );
  NOR U33232 ( .A(n33228), .B(n32950), .Z(n33230) );
  AND U33233 ( .A(n33235), .B(n33236), .Z(n32950) );
  IV U33234 ( .A(n33237), .Z(n33235) );
  XOR U33235 ( .A(n33238), .B(n33239), .Z(n33228) );
  AND U33236 ( .A(n33240), .B(n33241), .Z(n33239) );
  XNOR U33237 ( .A(n33238), .B(n33021), .Z(n33241) );
  XNOR U33238 ( .A(n33242), .B(n33243), .Z(n33021) );
  AND U33239 ( .A(n723), .B(n33244), .Z(n33243) );
  XOR U33240 ( .A(n33245), .B(n33242), .Z(n33244) );
  XNOR U33241 ( .A(n33246), .B(n33238), .Z(n33240) );
  IV U33242 ( .A(n32964), .Z(n33246) );
  XOR U33243 ( .A(n33247), .B(n33248), .Z(n32964) );
  AND U33244 ( .A(n731), .B(n33249), .Z(n33248) );
  XOR U33245 ( .A(n33250), .B(n33251), .Z(n33238) );
  AND U33246 ( .A(n33252), .B(n33253), .Z(n33251) );
  XNOR U33247 ( .A(n33250), .B(n33046), .Z(n33253) );
  XNOR U33248 ( .A(n33254), .B(n33255), .Z(n33046) );
  AND U33249 ( .A(n723), .B(n33256), .Z(n33255) );
  XNOR U33250 ( .A(n33257), .B(n33254), .Z(n33256) );
  XOR U33251 ( .A(n32975), .B(n33250), .Z(n33252) );
  XOR U33252 ( .A(n33258), .B(n33259), .Z(n32975) );
  AND U33253 ( .A(n731), .B(n33260), .Z(n33259) );
  XOR U33254 ( .A(n33222), .B(n33261), .Z(n33250) );
  AND U33255 ( .A(n33262), .B(n33225), .Z(n33261) );
  XNOR U33256 ( .A(n33092), .B(n33222), .Z(n33225) );
  XNOR U33257 ( .A(n33263), .B(n33264), .Z(n33092) );
  AND U33258 ( .A(n723), .B(n33265), .Z(n33264) );
  XOR U33259 ( .A(n33266), .B(n33263), .Z(n33265) );
  XNOR U33260 ( .A(n33267), .B(n33222), .Z(n33262) );
  IV U33261 ( .A(n32985), .Z(n33267) );
  XOR U33262 ( .A(n33268), .B(n33269), .Z(n32985) );
  AND U33263 ( .A(n731), .B(n33270), .Z(n33269) );
  XOR U33264 ( .A(n33271), .B(n33272), .Z(n33222) );
  AND U33265 ( .A(n33273), .B(n33274), .Z(n33272) );
  XNOR U33266 ( .A(n33271), .B(n33186), .Z(n33274) );
  XNOR U33267 ( .A(n33275), .B(n33276), .Z(n33186) );
  AND U33268 ( .A(n723), .B(n33277), .Z(n33276) );
  XNOR U33269 ( .A(n33278), .B(n33275), .Z(n33277) );
  XNOR U33270 ( .A(n33279), .B(n33271), .Z(n33273) );
  IV U33271 ( .A(n32997), .Z(n33279) );
  XOR U33272 ( .A(n33280), .B(n33281), .Z(n32997) );
  AND U33273 ( .A(n731), .B(n33282), .Z(n33281) );
  AND U33274 ( .A(n33226), .B(n33207), .Z(n33271) );
  XNOR U33275 ( .A(n33283), .B(n33284), .Z(n33207) );
  AND U33276 ( .A(n723), .B(n33285), .Z(n33284) );
  XNOR U33277 ( .A(n33286), .B(n33283), .Z(n33285) );
  XNOR U33278 ( .A(n33287), .B(n33288), .Z(n723) );
  NOR U33279 ( .A(n33289), .B(n33290), .Z(n33288) );
  XNOR U33280 ( .A(n33287), .B(n33237), .Z(n33290) );
  NOR U33281 ( .A(n33233), .B(n33234), .Z(n33237) );
  NOR U33282 ( .A(n33287), .B(n33236), .Z(n33289) );
  AND U33283 ( .A(n33291), .B(n33292), .Z(n33236) );
  XOR U33284 ( .A(n33293), .B(n33294), .Z(n33287) );
  AND U33285 ( .A(n33295), .B(n33296), .Z(n33294) );
  XNOR U33286 ( .A(n33293), .B(n33291), .Z(n33296) );
  IV U33287 ( .A(n33245), .Z(n33291) );
  XOR U33288 ( .A(n33297), .B(n33298), .Z(n33245) );
  XOR U33289 ( .A(n33299), .B(n33292), .Z(n33298) );
  AND U33290 ( .A(n33257), .B(n33300), .Z(n33292) );
  AND U33291 ( .A(n33301), .B(n33302), .Z(n33299) );
  XOR U33292 ( .A(n33303), .B(n33297), .Z(n33301) );
  XNOR U33293 ( .A(n33242), .B(n33293), .Z(n33295) );
  XNOR U33294 ( .A(n33304), .B(n33305), .Z(n33242) );
  AND U33295 ( .A(n727), .B(n33249), .Z(n33305) );
  XOR U33296 ( .A(n33304), .B(n33247), .Z(n33249) );
  XOR U33297 ( .A(n33306), .B(n33307), .Z(n33293) );
  AND U33298 ( .A(n33308), .B(n33309), .Z(n33307) );
  XNOR U33299 ( .A(n33306), .B(n33257), .Z(n33309) );
  XOR U33300 ( .A(n33310), .B(n33302), .Z(n33257) );
  XNOR U33301 ( .A(n33311), .B(n33297), .Z(n33302) );
  XOR U33302 ( .A(n33312), .B(n33313), .Z(n33297) );
  AND U33303 ( .A(n33314), .B(n33315), .Z(n33313) );
  XOR U33304 ( .A(n33316), .B(n33312), .Z(n33314) );
  XNOR U33305 ( .A(n33317), .B(n33318), .Z(n33311) );
  AND U33306 ( .A(n33319), .B(n33320), .Z(n33318) );
  XOR U33307 ( .A(n33317), .B(n33321), .Z(n33319) );
  XNOR U33308 ( .A(n33303), .B(n33300), .Z(n33310) );
  AND U33309 ( .A(n33322), .B(n33323), .Z(n33300) );
  XOR U33310 ( .A(n33324), .B(n33325), .Z(n33303) );
  AND U33311 ( .A(n33326), .B(n33327), .Z(n33325) );
  XOR U33312 ( .A(n33324), .B(n33328), .Z(n33326) );
  XNOR U33313 ( .A(n33254), .B(n33306), .Z(n33308) );
  XNOR U33314 ( .A(n33329), .B(n33330), .Z(n33254) );
  AND U33315 ( .A(n727), .B(n33260), .Z(n33330) );
  XOR U33316 ( .A(n33329), .B(n33258), .Z(n33260) );
  XOR U33317 ( .A(n33331), .B(n33332), .Z(n33306) );
  AND U33318 ( .A(n33333), .B(n33334), .Z(n33332) );
  XNOR U33319 ( .A(n33331), .B(n33322), .Z(n33334) );
  IV U33320 ( .A(n33266), .Z(n33322) );
  XNOR U33321 ( .A(n33335), .B(n33315), .Z(n33266) );
  XNOR U33322 ( .A(n33336), .B(n33321), .Z(n33315) );
  XOR U33323 ( .A(n33337), .B(n33338), .Z(n33321) );
  AND U33324 ( .A(n33339), .B(n33340), .Z(n33338) );
  XOR U33325 ( .A(n33337), .B(n33341), .Z(n33339) );
  XNOR U33326 ( .A(n33320), .B(n33312), .Z(n33336) );
  XOR U33327 ( .A(n33342), .B(n33343), .Z(n33312) );
  AND U33328 ( .A(n33344), .B(n33345), .Z(n33343) );
  XNOR U33329 ( .A(n33346), .B(n33342), .Z(n33344) );
  XNOR U33330 ( .A(n33347), .B(n33317), .Z(n33320) );
  XOR U33331 ( .A(n33348), .B(n33349), .Z(n33317) );
  AND U33332 ( .A(n33350), .B(n33351), .Z(n33349) );
  XOR U33333 ( .A(n33348), .B(n33352), .Z(n33350) );
  XNOR U33334 ( .A(n33353), .B(n33354), .Z(n33347) );
  AND U33335 ( .A(n33355), .B(n33356), .Z(n33354) );
  XNOR U33336 ( .A(n33353), .B(n33357), .Z(n33355) );
  XNOR U33337 ( .A(n33316), .B(n33323), .Z(n33335) );
  AND U33338 ( .A(n33278), .B(n33358), .Z(n33323) );
  XOR U33339 ( .A(n33328), .B(n33327), .Z(n33316) );
  XNOR U33340 ( .A(n33359), .B(n33324), .Z(n33327) );
  XOR U33341 ( .A(n33360), .B(n33361), .Z(n33324) );
  AND U33342 ( .A(n33362), .B(n33363), .Z(n33361) );
  XOR U33343 ( .A(n33360), .B(n33364), .Z(n33362) );
  XNOR U33344 ( .A(n33365), .B(n33366), .Z(n33359) );
  AND U33345 ( .A(n33367), .B(n33368), .Z(n33366) );
  XOR U33346 ( .A(n33365), .B(n33369), .Z(n33367) );
  XOR U33347 ( .A(n33370), .B(n33371), .Z(n33328) );
  AND U33348 ( .A(n33372), .B(n33373), .Z(n33371) );
  XOR U33349 ( .A(n33370), .B(n33374), .Z(n33372) );
  XNOR U33350 ( .A(n33263), .B(n33331), .Z(n33333) );
  XNOR U33351 ( .A(n33375), .B(n33376), .Z(n33263) );
  AND U33352 ( .A(n727), .B(n33270), .Z(n33376) );
  XOR U33353 ( .A(n33375), .B(n33268), .Z(n33270) );
  XOR U33354 ( .A(n33377), .B(n33378), .Z(n33331) );
  AND U33355 ( .A(n33379), .B(n33380), .Z(n33378) );
  XNOR U33356 ( .A(n33377), .B(n33278), .Z(n33380) );
  XOR U33357 ( .A(n33381), .B(n33345), .Z(n33278) );
  XNOR U33358 ( .A(n33382), .B(n33352), .Z(n33345) );
  XOR U33359 ( .A(n33341), .B(n33340), .Z(n33352) );
  XNOR U33360 ( .A(n33383), .B(n33337), .Z(n33340) );
  XOR U33361 ( .A(n33384), .B(n33385), .Z(n33337) );
  AND U33362 ( .A(n33386), .B(n33387), .Z(n33385) );
  XNOR U33363 ( .A(n33388), .B(n33389), .Z(n33386) );
  IV U33364 ( .A(n33384), .Z(n33388) );
  XNOR U33365 ( .A(n33390), .B(n33391), .Z(n33383) );
  NOR U33366 ( .A(n33392), .B(n33393), .Z(n33391) );
  XNOR U33367 ( .A(n33390), .B(n33394), .Z(n33392) );
  XOR U33368 ( .A(n33395), .B(n33396), .Z(n33341) );
  NOR U33369 ( .A(n33397), .B(n33398), .Z(n33396) );
  XNOR U33370 ( .A(n33395), .B(n33399), .Z(n33397) );
  XNOR U33371 ( .A(n33351), .B(n33342), .Z(n33382) );
  XOR U33372 ( .A(n33400), .B(n33401), .Z(n33342) );
  AND U33373 ( .A(n33402), .B(n33403), .Z(n33401) );
  XOR U33374 ( .A(n33400), .B(n33404), .Z(n33402) );
  XOR U33375 ( .A(n33405), .B(n33357), .Z(n33351) );
  XOR U33376 ( .A(n33406), .B(n33407), .Z(n33357) );
  NOR U33377 ( .A(n33408), .B(n33409), .Z(n33407) );
  XOR U33378 ( .A(n33406), .B(n33410), .Z(n33408) );
  XNOR U33379 ( .A(n33356), .B(n33348), .Z(n33405) );
  XOR U33380 ( .A(n33411), .B(n33412), .Z(n33348) );
  AND U33381 ( .A(n33413), .B(n33414), .Z(n33412) );
  XOR U33382 ( .A(n33411), .B(n33415), .Z(n33413) );
  XNOR U33383 ( .A(n33416), .B(n33353), .Z(n33356) );
  XOR U33384 ( .A(n33417), .B(n33418), .Z(n33353) );
  AND U33385 ( .A(n33419), .B(n33420), .Z(n33418) );
  XNOR U33386 ( .A(n33421), .B(n33422), .Z(n33419) );
  IV U33387 ( .A(n33417), .Z(n33421) );
  XNOR U33388 ( .A(n33423), .B(n33424), .Z(n33416) );
  NOR U33389 ( .A(n33425), .B(n33426), .Z(n33424) );
  XNOR U33390 ( .A(n33423), .B(n33427), .Z(n33425) );
  XOR U33391 ( .A(n33346), .B(n33358), .Z(n33381) );
  NOR U33392 ( .A(n33286), .B(n33428), .Z(n33358) );
  XNOR U33393 ( .A(n33364), .B(n33363), .Z(n33346) );
  XNOR U33394 ( .A(n33429), .B(n33369), .Z(n33363) );
  XNOR U33395 ( .A(n33430), .B(n33431), .Z(n33369) );
  NOR U33396 ( .A(n33432), .B(n33433), .Z(n33431) );
  XOR U33397 ( .A(n33430), .B(n33434), .Z(n33432) );
  XNOR U33398 ( .A(n33368), .B(n33360), .Z(n33429) );
  XOR U33399 ( .A(n33435), .B(n33436), .Z(n33360) );
  AND U33400 ( .A(n33437), .B(n33438), .Z(n33436) );
  XOR U33401 ( .A(n33435), .B(n33439), .Z(n33437) );
  XNOR U33402 ( .A(n33440), .B(n33365), .Z(n33368) );
  XOR U33403 ( .A(n33441), .B(n33442), .Z(n33365) );
  AND U33404 ( .A(n33443), .B(n33444), .Z(n33442) );
  XNOR U33405 ( .A(n33445), .B(n33446), .Z(n33443) );
  IV U33406 ( .A(n33441), .Z(n33445) );
  XNOR U33407 ( .A(n33447), .B(n33448), .Z(n33440) );
  NOR U33408 ( .A(n33449), .B(n33450), .Z(n33448) );
  XNOR U33409 ( .A(n33447), .B(n33451), .Z(n33449) );
  XOR U33410 ( .A(n33374), .B(n33373), .Z(n33364) );
  XNOR U33411 ( .A(n33452), .B(n33370), .Z(n33373) );
  XOR U33412 ( .A(n33453), .B(n33454), .Z(n33370) );
  AND U33413 ( .A(n33455), .B(n33456), .Z(n33454) );
  XNOR U33414 ( .A(n33457), .B(n33458), .Z(n33455) );
  IV U33415 ( .A(n33453), .Z(n33457) );
  XNOR U33416 ( .A(n33459), .B(n33460), .Z(n33452) );
  NOR U33417 ( .A(n33461), .B(n33462), .Z(n33460) );
  XNOR U33418 ( .A(n33459), .B(n33463), .Z(n33461) );
  XOR U33419 ( .A(n33464), .B(n33465), .Z(n33374) );
  NOR U33420 ( .A(n33466), .B(n33467), .Z(n33465) );
  XNOR U33421 ( .A(n33464), .B(n33468), .Z(n33466) );
  XNOR U33422 ( .A(n33275), .B(n33377), .Z(n33379) );
  XNOR U33423 ( .A(n33469), .B(n33470), .Z(n33275) );
  AND U33424 ( .A(n727), .B(n33282), .Z(n33470) );
  XOR U33425 ( .A(n33469), .B(n33280), .Z(n33282) );
  AND U33426 ( .A(n33283), .B(n33286), .Z(n33377) );
  XOR U33427 ( .A(n33471), .B(n33428), .Z(n33286) );
  XNOR U33428 ( .A(p_input[1920]), .B(p_input[2048]), .Z(n33428) );
  XNOR U33429 ( .A(n33404), .B(n33403), .Z(n33471) );
  XNOR U33430 ( .A(n33472), .B(n33415), .Z(n33403) );
  XOR U33431 ( .A(n33389), .B(n33387), .Z(n33415) );
  XNOR U33432 ( .A(n33473), .B(n33394), .Z(n33387) );
  XOR U33433 ( .A(p_input[1944]), .B(p_input[2072]), .Z(n33394) );
  XOR U33434 ( .A(n33384), .B(n33393), .Z(n33473) );
  XOR U33435 ( .A(n33474), .B(n33390), .Z(n33393) );
  XOR U33436 ( .A(p_input[1942]), .B(p_input[2070]), .Z(n33390) );
  XOR U33437 ( .A(p_input[1943]), .B(n17295), .Z(n33474) );
  XOR U33438 ( .A(p_input[1938]), .B(p_input[2066]), .Z(n33384) );
  XNOR U33439 ( .A(n33399), .B(n33398), .Z(n33389) );
  XOR U33440 ( .A(n33475), .B(n33395), .Z(n33398) );
  XOR U33441 ( .A(p_input[1939]), .B(p_input[2067]), .Z(n33395) );
  XOR U33442 ( .A(p_input[1940]), .B(n17297), .Z(n33475) );
  XOR U33443 ( .A(p_input[1941]), .B(p_input[2069]), .Z(n33399) );
  XOR U33444 ( .A(n33414), .B(n33476), .Z(n33472) );
  IV U33445 ( .A(n33400), .Z(n33476) );
  XOR U33446 ( .A(p_input[1921]), .B(p_input[2049]), .Z(n33400) );
  XNOR U33447 ( .A(n33477), .B(n33422), .Z(n33414) );
  XNOR U33448 ( .A(n33410), .B(n33409), .Z(n33422) );
  XNOR U33449 ( .A(n33478), .B(n33406), .Z(n33409) );
  XNOR U33450 ( .A(p_input[1946]), .B(p_input[2074]), .Z(n33406) );
  XOR U33451 ( .A(p_input[1947]), .B(n17300), .Z(n33478) );
  XOR U33452 ( .A(p_input[1948]), .B(p_input[2076]), .Z(n33410) );
  XOR U33453 ( .A(n33420), .B(n33479), .Z(n33477) );
  IV U33454 ( .A(n33411), .Z(n33479) );
  XOR U33455 ( .A(p_input[1937]), .B(p_input[2065]), .Z(n33411) );
  XNOR U33456 ( .A(n33480), .B(n33427), .Z(n33420) );
  XNOR U33457 ( .A(p_input[1951]), .B(n17303), .Z(n33427) );
  XOR U33458 ( .A(n33417), .B(n33426), .Z(n33480) );
  XOR U33459 ( .A(n33481), .B(n33423), .Z(n33426) );
  XOR U33460 ( .A(p_input[1949]), .B(p_input[2077]), .Z(n33423) );
  XOR U33461 ( .A(p_input[1950]), .B(n17305), .Z(n33481) );
  XOR U33462 ( .A(p_input[1945]), .B(p_input[2073]), .Z(n33417) );
  XOR U33463 ( .A(n33439), .B(n33438), .Z(n33404) );
  XNOR U33464 ( .A(n33482), .B(n33446), .Z(n33438) );
  XNOR U33465 ( .A(n33434), .B(n33433), .Z(n33446) );
  XNOR U33466 ( .A(n33483), .B(n33430), .Z(n33433) );
  XNOR U33467 ( .A(p_input[1931]), .B(p_input[2059]), .Z(n33430) );
  XOR U33468 ( .A(p_input[1932]), .B(n16451), .Z(n33483) );
  XOR U33469 ( .A(p_input[1933]), .B(p_input[2061]), .Z(n33434) );
  XOR U33470 ( .A(n33444), .B(n33484), .Z(n33482) );
  IV U33471 ( .A(n33435), .Z(n33484) );
  XOR U33472 ( .A(p_input[1922]), .B(p_input[2050]), .Z(n33435) );
  XNOR U33473 ( .A(n33485), .B(n33451), .Z(n33444) );
  XNOR U33474 ( .A(p_input[1936]), .B(n16454), .Z(n33451) );
  XOR U33475 ( .A(n33441), .B(n33450), .Z(n33485) );
  XOR U33476 ( .A(n33486), .B(n33447), .Z(n33450) );
  XOR U33477 ( .A(p_input[1934]), .B(p_input[2062]), .Z(n33447) );
  XOR U33478 ( .A(p_input[1935]), .B(n16456), .Z(n33486) );
  XOR U33479 ( .A(p_input[1930]), .B(p_input[2058]), .Z(n33441) );
  XOR U33480 ( .A(n33458), .B(n33456), .Z(n33439) );
  XNOR U33481 ( .A(n33487), .B(n33463), .Z(n33456) );
  XOR U33482 ( .A(p_input[1929]), .B(p_input[2057]), .Z(n33463) );
  XOR U33483 ( .A(n33453), .B(n33462), .Z(n33487) );
  XOR U33484 ( .A(n33488), .B(n33459), .Z(n33462) );
  XOR U33485 ( .A(p_input[1927]), .B(p_input[2055]), .Z(n33459) );
  XOR U33486 ( .A(p_input[1928]), .B(n17312), .Z(n33488) );
  XOR U33487 ( .A(p_input[1923]), .B(p_input[2051]), .Z(n33453) );
  XNOR U33488 ( .A(n33468), .B(n33467), .Z(n33458) );
  XOR U33489 ( .A(n33489), .B(n33464), .Z(n33467) );
  XOR U33490 ( .A(p_input[1924]), .B(p_input[2052]), .Z(n33464) );
  XOR U33491 ( .A(p_input[1925]), .B(n17314), .Z(n33489) );
  XOR U33492 ( .A(p_input[1926]), .B(p_input[2054]), .Z(n33468) );
  XNOR U33493 ( .A(n33490), .B(n33491), .Z(n33283) );
  AND U33494 ( .A(n727), .B(n33492), .Z(n33491) );
  XNOR U33495 ( .A(n33493), .B(n33494), .Z(n727) );
  NOR U33496 ( .A(n33495), .B(n33496), .Z(n33494) );
  XOR U33497 ( .A(n33234), .B(n33493), .Z(n33496) );
  NOR U33498 ( .A(n33493), .B(n33233), .Z(n33495) );
  XOR U33499 ( .A(n33497), .B(n33498), .Z(n33493) );
  AND U33500 ( .A(n33499), .B(n33500), .Z(n33498) );
  XNOR U33501 ( .A(n33304), .B(n33497), .Z(n33500) );
  XOR U33502 ( .A(n33497), .B(n33247), .Z(n33499) );
  XOR U33503 ( .A(n33501), .B(n33502), .Z(n33497) );
  AND U33504 ( .A(n33503), .B(n33504), .Z(n33502) );
  XNOR U33505 ( .A(n33329), .B(n33501), .Z(n33504) );
  XOR U33506 ( .A(n33501), .B(n33258), .Z(n33503) );
  XOR U33507 ( .A(n33505), .B(n33506), .Z(n33501) );
  AND U33508 ( .A(n33507), .B(n33508), .Z(n33506) );
  XOR U33509 ( .A(n33505), .B(n33268), .Z(n33507) );
  XOR U33510 ( .A(n33509), .B(n33510), .Z(n33226) );
  AND U33511 ( .A(n731), .B(n33492), .Z(n33510) );
  XNOR U33512 ( .A(n33490), .B(n33509), .Z(n33492) );
  XNOR U33513 ( .A(n33511), .B(n33512), .Z(n731) );
  NOR U33514 ( .A(n33513), .B(n33514), .Z(n33512) );
  XNOR U33515 ( .A(n33234), .B(n33515), .Z(n33514) );
  IV U33516 ( .A(n33511), .Z(n33515) );
  AND U33517 ( .A(n33516), .B(n33517), .Z(n33234) );
  NOR U33518 ( .A(n33511), .B(n33233), .Z(n33513) );
  AND U33519 ( .A(n33518), .B(n33519), .Z(n33233) );
  IV U33520 ( .A(n33520), .Z(n33518) );
  XOR U33521 ( .A(n33521), .B(n33522), .Z(n33511) );
  AND U33522 ( .A(n33523), .B(n33524), .Z(n33522) );
  XNOR U33523 ( .A(n33521), .B(n33304), .Z(n33524) );
  XNOR U33524 ( .A(n33525), .B(n33526), .Z(n33304) );
  AND U33525 ( .A(n734), .B(n33527), .Z(n33526) );
  XOR U33526 ( .A(n33528), .B(n33525), .Z(n33527) );
  XNOR U33527 ( .A(n33529), .B(n33521), .Z(n33523) );
  IV U33528 ( .A(n33247), .Z(n33529) );
  XOR U33529 ( .A(n33530), .B(n33531), .Z(n33247) );
  AND U33530 ( .A(n741), .B(n33532), .Z(n33531) );
  XOR U33531 ( .A(n33533), .B(n33534), .Z(n33521) );
  AND U33532 ( .A(n33535), .B(n33536), .Z(n33534) );
  XNOR U33533 ( .A(n33533), .B(n33329), .Z(n33536) );
  XNOR U33534 ( .A(n33537), .B(n33538), .Z(n33329) );
  AND U33535 ( .A(n734), .B(n33539), .Z(n33538) );
  XNOR U33536 ( .A(n33540), .B(n33537), .Z(n33539) );
  XOR U33537 ( .A(n33258), .B(n33533), .Z(n33535) );
  XOR U33538 ( .A(n33541), .B(n33542), .Z(n33258) );
  AND U33539 ( .A(n741), .B(n33543), .Z(n33542) );
  XOR U33540 ( .A(n33505), .B(n33544), .Z(n33533) );
  AND U33541 ( .A(n33545), .B(n33508), .Z(n33544) );
  XNOR U33542 ( .A(n33375), .B(n33505), .Z(n33508) );
  XNOR U33543 ( .A(n33546), .B(n33547), .Z(n33375) );
  AND U33544 ( .A(n734), .B(n33548), .Z(n33547) );
  XOR U33545 ( .A(n33549), .B(n33546), .Z(n33548) );
  XNOR U33546 ( .A(n33550), .B(n33505), .Z(n33545) );
  IV U33547 ( .A(n33268), .Z(n33550) );
  XOR U33548 ( .A(n33551), .B(n33552), .Z(n33268) );
  AND U33549 ( .A(n741), .B(n33553), .Z(n33552) );
  XOR U33550 ( .A(n33554), .B(n33555), .Z(n33505) );
  AND U33551 ( .A(n33556), .B(n33557), .Z(n33555) );
  XNOR U33552 ( .A(n33554), .B(n33469), .Z(n33557) );
  XNOR U33553 ( .A(n33558), .B(n33559), .Z(n33469) );
  AND U33554 ( .A(n734), .B(n33560), .Z(n33559) );
  XNOR U33555 ( .A(n33561), .B(n33558), .Z(n33560) );
  XNOR U33556 ( .A(n33562), .B(n33554), .Z(n33556) );
  IV U33557 ( .A(n33280), .Z(n33562) );
  XOR U33558 ( .A(n33563), .B(n33564), .Z(n33280) );
  AND U33559 ( .A(n741), .B(n33565), .Z(n33564) );
  AND U33560 ( .A(n33509), .B(n33490), .Z(n33554) );
  XNOR U33561 ( .A(n33566), .B(n33567), .Z(n33490) );
  AND U33562 ( .A(n734), .B(n33568), .Z(n33567) );
  XNOR U33563 ( .A(n33569), .B(n33566), .Z(n33568) );
  XNOR U33564 ( .A(n33570), .B(n33571), .Z(n734) );
  NOR U33565 ( .A(n33572), .B(n33573), .Z(n33571) );
  XNOR U33566 ( .A(n33570), .B(n33520), .Z(n33573) );
  NOR U33567 ( .A(n33516), .B(n33517), .Z(n33520) );
  NOR U33568 ( .A(n33570), .B(n33519), .Z(n33572) );
  AND U33569 ( .A(n33574), .B(n33575), .Z(n33519) );
  XOR U33570 ( .A(n33576), .B(n33577), .Z(n33570) );
  AND U33571 ( .A(n33578), .B(n33579), .Z(n33577) );
  XNOR U33572 ( .A(n33576), .B(n33574), .Z(n33579) );
  IV U33573 ( .A(n33528), .Z(n33574) );
  XOR U33574 ( .A(n33580), .B(n33581), .Z(n33528) );
  XOR U33575 ( .A(n33582), .B(n33575), .Z(n33581) );
  AND U33576 ( .A(n33540), .B(n33583), .Z(n33575) );
  AND U33577 ( .A(n33584), .B(n33585), .Z(n33582) );
  XOR U33578 ( .A(n33586), .B(n33580), .Z(n33584) );
  XNOR U33579 ( .A(n33525), .B(n33576), .Z(n33578) );
  XNOR U33580 ( .A(n33587), .B(n33588), .Z(n33525) );
  AND U33581 ( .A(n738), .B(n33532), .Z(n33588) );
  XOR U33582 ( .A(n33587), .B(n33530), .Z(n33532) );
  XOR U33583 ( .A(n33589), .B(n33590), .Z(n33576) );
  AND U33584 ( .A(n33591), .B(n33592), .Z(n33590) );
  XNOR U33585 ( .A(n33589), .B(n33540), .Z(n33592) );
  XOR U33586 ( .A(n33593), .B(n33585), .Z(n33540) );
  XNOR U33587 ( .A(n33594), .B(n33580), .Z(n33585) );
  XOR U33588 ( .A(n33595), .B(n33596), .Z(n33580) );
  AND U33589 ( .A(n33597), .B(n33598), .Z(n33596) );
  XOR U33590 ( .A(n33599), .B(n33595), .Z(n33597) );
  XNOR U33591 ( .A(n33600), .B(n33601), .Z(n33594) );
  AND U33592 ( .A(n33602), .B(n33603), .Z(n33601) );
  XOR U33593 ( .A(n33600), .B(n33604), .Z(n33602) );
  XNOR U33594 ( .A(n33586), .B(n33583), .Z(n33593) );
  AND U33595 ( .A(n33605), .B(n33606), .Z(n33583) );
  XOR U33596 ( .A(n33607), .B(n33608), .Z(n33586) );
  AND U33597 ( .A(n33609), .B(n33610), .Z(n33608) );
  XOR U33598 ( .A(n33607), .B(n33611), .Z(n33609) );
  XNOR U33599 ( .A(n33537), .B(n33589), .Z(n33591) );
  XNOR U33600 ( .A(n33612), .B(n33613), .Z(n33537) );
  AND U33601 ( .A(n738), .B(n33543), .Z(n33613) );
  XOR U33602 ( .A(n33612), .B(n33541), .Z(n33543) );
  XOR U33603 ( .A(n33614), .B(n33615), .Z(n33589) );
  AND U33604 ( .A(n33616), .B(n33617), .Z(n33615) );
  XNOR U33605 ( .A(n33614), .B(n33605), .Z(n33617) );
  IV U33606 ( .A(n33549), .Z(n33605) );
  XNOR U33607 ( .A(n33618), .B(n33598), .Z(n33549) );
  XNOR U33608 ( .A(n33619), .B(n33604), .Z(n33598) );
  XOR U33609 ( .A(n33620), .B(n33621), .Z(n33604) );
  AND U33610 ( .A(n33622), .B(n33623), .Z(n33621) );
  XOR U33611 ( .A(n33620), .B(n33624), .Z(n33622) );
  XNOR U33612 ( .A(n33603), .B(n33595), .Z(n33619) );
  XOR U33613 ( .A(n33625), .B(n33626), .Z(n33595) );
  AND U33614 ( .A(n33627), .B(n33628), .Z(n33626) );
  XNOR U33615 ( .A(n33629), .B(n33625), .Z(n33627) );
  XNOR U33616 ( .A(n33630), .B(n33600), .Z(n33603) );
  XOR U33617 ( .A(n33631), .B(n33632), .Z(n33600) );
  AND U33618 ( .A(n33633), .B(n33634), .Z(n33632) );
  XOR U33619 ( .A(n33631), .B(n33635), .Z(n33633) );
  XNOR U33620 ( .A(n33636), .B(n33637), .Z(n33630) );
  AND U33621 ( .A(n33638), .B(n33639), .Z(n33637) );
  XNOR U33622 ( .A(n33636), .B(n33640), .Z(n33638) );
  XNOR U33623 ( .A(n33599), .B(n33606), .Z(n33618) );
  AND U33624 ( .A(n33561), .B(n33641), .Z(n33606) );
  XOR U33625 ( .A(n33611), .B(n33610), .Z(n33599) );
  XNOR U33626 ( .A(n33642), .B(n33607), .Z(n33610) );
  XOR U33627 ( .A(n33643), .B(n33644), .Z(n33607) );
  AND U33628 ( .A(n33645), .B(n33646), .Z(n33644) );
  XOR U33629 ( .A(n33643), .B(n33647), .Z(n33645) );
  XNOR U33630 ( .A(n33648), .B(n33649), .Z(n33642) );
  AND U33631 ( .A(n33650), .B(n33651), .Z(n33649) );
  XOR U33632 ( .A(n33648), .B(n33652), .Z(n33650) );
  XOR U33633 ( .A(n33653), .B(n33654), .Z(n33611) );
  AND U33634 ( .A(n33655), .B(n33656), .Z(n33654) );
  XOR U33635 ( .A(n33653), .B(n33657), .Z(n33655) );
  XNOR U33636 ( .A(n33546), .B(n33614), .Z(n33616) );
  XNOR U33637 ( .A(n33658), .B(n33659), .Z(n33546) );
  AND U33638 ( .A(n738), .B(n33553), .Z(n33659) );
  XOR U33639 ( .A(n33658), .B(n33551), .Z(n33553) );
  XOR U33640 ( .A(n33660), .B(n33661), .Z(n33614) );
  AND U33641 ( .A(n33662), .B(n33663), .Z(n33661) );
  XNOR U33642 ( .A(n33660), .B(n33561), .Z(n33663) );
  XOR U33643 ( .A(n33664), .B(n33628), .Z(n33561) );
  XNOR U33644 ( .A(n33665), .B(n33635), .Z(n33628) );
  XOR U33645 ( .A(n33624), .B(n33623), .Z(n33635) );
  XNOR U33646 ( .A(n33666), .B(n33620), .Z(n33623) );
  XOR U33647 ( .A(n33667), .B(n33668), .Z(n33620) );
  AND U33648 ( .A(n33669), .B(n33670), .Z(n33668) );
  XNOR U33649 ( .A(n33671), .B(n33672), .Z(n33669) );
  IV U33650 ( .A(n33667), .Z(n33671) );
  XNOR U33651 ( .A(n33673), .B(n33674), .Z(n33666) );
  NOR U33652 ( .A(n33675), .B(n33676), .Z(n33674) );
  XNOR U33653 ( .A(n33673), .B(n33677), .Z(n33675) );
  XOR U33654 ( .A(n33678), .B(n33679), .Z(n33624) );
  NOR U33655 ( .A(n33680), .B(n33681), .Z(n33679) );
  XNOR U33656 ( .A(n33678), .B(n33682), .Z(n33680) );
  XNOR U33657 ( .A(n33634), .B(n33625), .Z(n33665) );
  XOR U33658 ( .A(n33683), .B(n33684), .Z(n33625) );
  AND U33659 ( .A(n33685), .B(n33686), .Z(n33684) );
  XOR U33660 ( .A(n33683), .B(n33687), .Z(n33685) );
  XOR U33661 ( .A(n33688), .B(n33640), .Z(n33634) );
  XOR U33662 ( .A(n33689), .B(n33690), .Z(n33640) );
  NOR U33663 ( .A(n33691), .B(n33692), .Z(n33690) );
  XOR U33664 ( .A(n33689), .B(n33693), .Z(n33691) );
  XNOR U33665 ( .A(n33639), .B(n33631), .Z(n33688) );
  XOR U33666 ( .A(n33694), .B(n33695), .Z(n33631) );
  AND U33667 ( .A(n33696), .B(n33697), .Z(n33695) );
  XOR U33668 ( .A(n33694), .B(n33698), .Z(n33696) );
  XNOR U33669 ( .A(n33699), .B(n33636), .Z(n33639) );
  XOR U33670 ( .A(n33700), .B(n33701), .Z(n33636) );
  AND U33671 ( .A(n33702), .B(n33703), .Z(n33701) );
  XNOR U33672 ( .A(n33704), .B(n33705), .Z(n33702) );
  IV U33673 ( .A(n33700), .Z(n33704) );
  XNOR U33674 ( .A(n33706), .B(n33707), .Z(n33699) );
  NOR U33675 ( .A(n33708), .B(n33709), .Z(n33707) );
  XNOR U33676 ( .A(n33706), .B(n33710), .Z(n33708) );
  XOR U33677 ( .A(n33629), .B(n33641), .Z(n33664) );
  NOR U33678 ( .A(n33569), .B(n33711), .Z(n33641) );
  XNOR U33679 ( .A(n33647), .B(n33646), .Z(n33629) );
  XNOR U33680 ( .A(n33712), .B(n33652), .Z(n33646) );
  XNOR U33681 ( .A(n33713), .B(n33714), .Z(n33652) );
  NOR U33682 ( .A(n33715), .B(n33716), .Z(n33714) );
  XOR U33683 ( .A(n33713), .B(n33717), .Z(n33715) );
  XNOR U33684 ( .A(n33651), .B(n33643), .Z(n33712) );
  XOR U33685 ( .A(n33718), .B(n33719), .Z(n33643) );
  AND U33686 ( .A(n33720), .B(n33721), .Z(n33719) );
  XOR U33687 ( .A(n33718), .B(n33722), .Z(n33720) );
  XNOR U33688 ( .A(n33723), .B(n33648), .Z(n33651) );
  XOR U33689 ( .A(n33724), .B(n33725), .Z(n33648) );
  AND U33690 ( .A(n33726), .B(n33727), .Z(n33725) );
  XNOR U33691 ( .A(n33728), .B(n33729), .Z(n33726) );
  IV U33692 ( .A(n33724), .Z(n33728) );
  XNOR U33693 ( .A(n33730), .B(n33731), .Z(n33723) );
  NOR U33694 ( .A(n33732), .B(n33733), .Z(n33731) );
  XNOR U33695 ( .A(n33730), .B(n33734), .Z(n33732) );
  XOR U33696 ( .A(n33657), .B(n33656), .Z(n33647) );
  XNOR U33697 ( .A(n33735), .B(n33653), .Z(n33656) );
  XOR U33698 ( .A(n33736), .B(n33737), .Z(n33653) );
  AND U33699 ( .A(n33738), .B(n33739), .Z(n33737) );
  XNOR U33700 ( .A(n33740), .B(n33741), .Z(n33738) );
  IV U33701 ( .A(n33736), .Z(n33740) );
  XNOR U33702 ( .A(n33742), .B(n33743), .Z(n33735) );
  NOR U33703 ( .A(n33744), .B(n33745), .Z(n33743) );
  XNOR U33704 ( .A(n33742), .B(n33746), .Z(n33744) );
  XOR U33705 ( .A(n33747), .B(n33748), .Z(n33657) );
  NOR U33706 ( .A(n33749), .B(n33750), .Z(n33748) );
  XNOR U33707 ( .A(n33747), .B(n33751), .Z(n33749) );
  XNOR U33708 ( .A(n33558), .B(n33660), .Z(n33662) );
  XNOR U33709 ( .A(n33752), .B(n33753), .Z(n33558) );
  AND U33710 ( .A(n738), .B(n33565), .Z(n33753) );
  XOR U33711 ( .A(n33752), .B(n33563), .Z(n33565) );
  AND U33712 ( .A(n33566), .B(n33569), .Z(n33660) );
  XOR U33713 ( .A(n33754), .B(n33711), .Z(n33569) );
  XNOR U33714 ( .A(p_input[1952]), .B(p_input[2048]), .Z(n33711) );
  XNOR U33715 ( .A(n33687), .B(n33686), .Z(n33754) );
  XNOR U33716 ( .A(n33755), .B(n33698), .Z(n33686) );
  XOR U33717 ( .A(n33672), .B(n33670), .Z(n33698) );
  XNOR U33718 ( .A(n33756), .B(n33677), .Z(n33670) );
  XOR U33719 ( .A(p_input[1976]), .B(p_input[2072]), .Z(n33677) );
  XOR U33720 ( .A(n33667), .B(n33676), .Z(n33756) );
  XOR U33721 ( .A(n33757), .B(n33673), .Z(n33676) );
  XOR U33722 ( .A(p_input[1974]), .B(p_input[2070]), .Z(n33673) );
  XOR U33723 ( .A(p_input[1975]), .B(n17295), .Z(n33757) );
  XOR U33724 ( .A(p_input[1970]), .B(p_input[2066]), .Z(n33667) );
  XNOR U33725 ( .A(n33682), .B(n33681), .Z(n33672) );
  XOR U33726 ( .A(n33758), .B(n33678), .Z(n33681) );
  XOR U33727 ( .A(p_input[1971]), .B(p_input[2067]), .Z(n33678) );
  XOR U33728 ( .A(p_input[1972]), .B(n17297), .Z(n33758) );
  XOR U33729 ( .A(p_input[1973]), .B(p_input[2069]), .Z(n33682) );
  XOR U33730 ( .A(n33697), .B(n33759), .Z(n33755) );
  IV U33731 ( .A(n33683), .Z(n33759) );
  XOR U33732 ( .A(p_input[1953]), .B(p_input[2049]), .Z(n33683) );
  XNOR U33733 ( .A(n33760), .B(n33705), .Z(n33697) );
  XNOR U33734 ( .A(n33693), .B(n33692), .Z(n33705) );
  XNOR U33735 ( .A(n33761), .B(n33689), .Z(n33692) );
  XNOR U33736 ( .A(p_input[1978]), .B(p_input[2074]), .Z(n33689) );
  XOR U33737 ( .A(p_input[1979]), .B(n17300), .Z(n33761) );
  XOR U33738 ( .A(p_input[1980]), .B(p_input[2076]), .Z(n33693) );
  XOR U33739 ( .A(n33703), .B(n33762), .Z(n33760) );
  IV U33740 ( .A(n33694), .Z(n33762) );
  XOR U33741 ( .A(p_input[1969]), .B(p_input[2065]), .Z(n33694) );
  XNOR U33742 ( .A(n33763), .B(n33710), .Z(n33703) );
  XNOR U33743 ( .A(p_input[1983]), .B(n17303), .Z(n33710) );
  IV U33744 ( .A(p_input[2079]), .Z(n17303) );
  XOR U33745 ( .A(n33700), .B(n33709), .Z(n33763) );
  XOR U33746 ( .A(n33764), .B(n33706), .Z(n33709) );
  XOR U33747 ( .A(p_input[1981]), .B(p_input[2077]), .Z(n33706) );
  XOR U33748 ( .A(p_input[1982]), .B(n17305), .Z(n33764) );
  XOR U33749 ( .A(p_input[1977]), .B(p_input[2073]), .Z(n33700) );
  XOR U33750 ( .A(n33722), .B(n33721), .Z(n33687) );
  XNOR U33751 ( .A(n33765), .B(n33729), .Z(n33721) );
  XNOR U33752 ( .A(n33717), .B(n33716), .Z(n33729) );
  XNOR U33753 ( .A(n33766), .B(n33713), .Z(n33716) );
  XNOR U33754 ( .A(p_input[1963]), .B(p_input[2059]), .Z(n33713) );
  XOR U33755 ( .A(p_input[1964]), .B(n16451), .Z(n33766) );
  XOR U33756 ( .A(p_input[1965]), .B(p_input[2061]), .Z(n33717) );
  XOR U33757 ( .A(n33727), .B(n33767), .Z(n33765) );
  IV U33758 ( .A(n33718), .Z(n33767) );
  XOR U33759 ( .A(p_input[1954]), .B(p_input[2050]), .Z(n33718) );
  XNOR U33760 ( .A(n33768), .B(n33734), .Z(n33727) );
  XNOR U33761 ( .A(p_input[1968]), .B(n16454), .Z(n33734) );
  IV U33762 ( .A(p_input[2064]), .Z(n16454) );
  XOR U33763 ( .A(n33724), .B(n33733), .Z(n33768) );
  XOR U33764 ( .A(n33769), .B(n33730), .Z(n33733) );
  XOR U33765 ( .A(p_input[1966]), .B(p_input[2062]), .Z(n33730) );
  XOR U33766 ( .A(p_input[1967]), .B(n16456), .Z(n33769) );
  XOR U33767 ( .A(p_input[1962]), .B(p_input[2058]), .Z(n33724) );
  XOR U33768 ( .A(n33741), .B(n33739), .Z(n33722) );
  XNOR U33769 ( .A(n33770), .B(n33746), .Z(n33739) );
  XOR U33770 ( .A(p_input[1961]), .B(p_input[2057]), .Z(n33746) );
  XOR U33771 ( .A(n33736), .B(n33745), .Z(n33770) );
  XOR U33772 ( .A(n33771), .B(n33742), .Z(n33745) );
  XOR U33773 ( .A(p_input[1959]), .B(p_input[2055]), .Z(n33742) );
  XOR U33774 ( .A(p_input[1960]), .B(n17312), .Z(n33771) );
  XOR U33775 ( .A(p_input[1955]), .B(p_input[2051]), .Z(n33736) );
  XNOR U33776 ( .A(n33751), .B(n33750), .Z(n33741) );
  XOR U33777 ( .A(n33772), .B(n33747), .Z(n33750) );
  XOR U33778 ( .A(p_input[1956]), .B(p_input[2052]), .Z(n33747) );
  XOR U33779 ( .A(p_input[1957]), .B(n17314), .Z(n33772) );
  XOR U33780 ( .A(p_input[1958]), .B(p_input[2054]), .Z(n33751) );
  XNOR U33781 ( .A(n33773), .B(n33774), .Z(n33566) );
  AND U33782 ( .A(n738), .B(n33775), .Z(n33774) );
  XNOR U33783 ( .A(n33776), .B(n33777), .Z(n738) );
  NOR U33784 ( .A(n33778), .B(n33779), .Z(n33777) );
  XOR U33785 ( .A(n33517), .B(n33776), .Z(n33779) );
  NOR U33786 ( .A(n33776), .B(n33516), .Z(n33778) );
  XOR U33787 ( .A(n33780), .B(n33781), .Z(n33776) );
  AND U33788 ( .A(n33782), .B(n33783), .Z(n33781) );
  XNOR U33789 ( .A(n33587), .B(n33780), .Z(n33783) );
  XOR U33790 ( .A(n33780), .B(n33530), .Z(n33782) );
  XOR U33791 ( .A(n33784), .B(n33785), .Z(n33780) );
  AND U33792 ( .A(n33786), .B(n33787), .Z(n33785) );
  XNOR U33793 ( .A(n33612), .B(n33784), .Z(n33787) );
  XOR U33794 ( .A(n33784), .B(n33541), .Z(n33786) );
  XOR U33795 ( .A(n33788), .B(n33789), .Z(n33784) );
  AND U33796 ( .A(n33790), .B(n33791), .Z(n33789) );
  XOR U33797 ( .A(n33788), .B(n33551), .Z(n33790) );
  XOR U33798 ( .A(n33792), .B(n33793), .Z(n33509) );
  AND U33799 ( .A(n741), .B(n33775), .Z(n33793) );
  XOR U33800 ( .A(n33794), .B(n33792), .Z(n33775) );
  XNOR U33801 ( .A(n33795), .B(n33796), .Z(n741) );
  NOR U33802 ( .A(n33797), .B(n33798), .Z(n33796) );
  XNOR U33803 ( .A(n33517), .B(n33799), .Z(n33798) );
  IV U33804 ( .A(n33795), .Z(n33799) );
  AND U33805 ( .A(n33530), .B(n33800), .Z(n33517) );
  NOR U33806 ( .A(n33795), .B(n33516), .Z(n33797) );
  AND U33807 ( .A(n33587), .B(n33801), .Z(n33516) );
  XOR U33808 ( .A(n33802), .B(n33803), .Z(n33795) );
  AND U33809 ( .A(n33804), .B(n33805), .Z(n33803) );
  XNOR U33810 ( .A(n33802), .B(n33587), .Z(n33805) );
  XNOR U33811 ( .A(n33806), .B(n33807), .Z(n33587) );
  XOR U33812 ( .A(n33808), .B(n33801), .Z(n33807) );
  AND U33813 ( .A(n33612), .B(n33809), .Z(n33801) );
  AND U33814 ( .A(n33810), .B(n33811), .Z(n33808) );
  XOR U33815 ( .A(n33812), .B(n33806), .Z(n33810) );
  XNOR U33816 ( .A(n33813), .B(n33802), .Z(n33804) );
  IV U33817 ( .A(n33530), .Z(n33813) );
  XNOR U33818 ( .A(n33814), .B(n33815), .Z(n33530) );
  XOR U33819 ( .A(n33816), .B(n33800), .Z(n33815) );
  AND U33820 ( .A(n33541), .B(n33817), .Z(n33800) );
  AND U33821 ( .A(n33818), .B(n33819), .Z(n33816) );
  XNOR U33822 ( .A(n33814), .B(n33820), .Z(n33818) );
  XOR U33823 ( .A(n33821), .B(n33822), .Z(n33802) );
  AND U33824 ( .A(n33823), .B(n33824), .Z(n33822) );
  XNOR U33825 ( .A(n33821), .B(n33612), .Z(n33824) );
  XOR U33826 ( .A(n33825), .B(n33811), .Z(n33612) );
  XNOR U33827 ( .A(n33826), .B(n33806), .Z(n33811) );
  XOR U33828 ( .A(n33827), .B(n33828), .Z(n33806) );
  AND U33829 ( .A(n33829), .B(n33830), .Z(n33828) );
  XOR U33830 ( .A(n33831), .B(n33827), .Z(n33829) );
  XNOR U33831 ( .A(n33832), .B(n33833), .Z(n33826) );
  AND U33832 ( .A(n33834), .B(n33835), .Z(n33833) );
  XOR U33833 ( .A(n33832), .B(n33836), .Z(n33834) );
  XNOR U33834 ( .A(n33812), .B(n33809), .Z(n33825) );
  AND U33835 ( .A(n33658), .B(n33837), .Z(n33809) );
  XOR U33836 ( .A(n33838), .B(n33839), .Z(n33812) );
  AND U33837 ( .A(n33840), .B(n33841), .Z(n33839) );
  XOR U33838 ( .A(n33838), .B(n33842), .Z(n33840) );
  XOR U33839 ( .A(n33541), .B(n33821), .Z(n33823) );
  XNOR U33840 ( .A(n33843), .B(n33820), .Z(n33541) );
  XNOR U33841 ( .A(n33844), .B(n33845), .Z(n33820) );
  AND U33842 ( .A(n33846), .B(n33847), .Z(n33845) );
  XOR U33843 ( .A(n33844), .B(n33848), .Z(n33846) );
  XNOR U33844 ( .A(n33819), .B(n33817), .Z(n33843) );
  AND U33845 ( .A(n33551), .B(n33849), .Z(n33817) );
  XNOR U33846 ( .A(n33850), .B(n33814), .Z(n33819) );
  XOR U33847 ( .A(n33851), .B(n33852), .Z(n33814) );
  AND U33848 ( .A(n33853), .B(n33854), .Z(n33852) );
  XOR U33849 ( .A(n33851), .B(n33855), .Z(n33853) );
  XNOR U33850 ( .A(n33856), .B(n33857), .Z(n33850) );
  AND U33851 ( .A(n33858), .B(n33859), .Z(n33857) );
  XNOR U33852 ( .A(n33856), .B(n33860), .Z(n33858) );
  XOR U33853 ( .A(n33788), .B(n33861), .Z(n33821) );
  AND U33854 ( .A(n33862), .B(n33791), .Z(n33861) );
  XNOR U33855 ( .A(n33658), .B(n33788), .Z(n33791) );
  XOR U33856 ( .A(n33863), .B(n33830), .Z(n33658) );
  XNOR U33857 ( .A(n33864), .B(n33836), .Z(n33830) );
  XOR U33858 ( .A(n33865), .B(n33866), .Z(n33836) );
  AND U33859 ( .A(n33867), .B(n33868), .Z(n33866) );
  XOR U33860 ( .A(n33865), .B(n33869), .Z(n33867) );
  XNOR U33861 ( .A(n33835), .B(n33827), .Z(n33864) );
  XOR U33862 ( .A(n33870), .B(n33871), .Z(n33827) );
  AND U33863 ( .A(n33872), .B(n33873), .Z(n33871) );
  XNOR U33864 ( .A(n33874), .B(n33870), .Z(n33872) );
  XNOR U33865 ( .A(n33875), .B(n33832), .Z(n33835) );
  XOR U33866 ( .A(n33876), .B(n33877), .Z(n33832) );
  AND U33867 ( .A(n33878), .B(n33879), .Z(n33877) );
  XOR U33868 ( .A(n33876), .B(n33880), .Z(n33878) );
  XNOR U33869 ( .A(n33881), .B(n33882), .Z(n33875) );
  AND U33870 ( .A(n33883), .B(n33884), .Z(n33882) );
  XNOR U33871 ( .A(n33881), .B(n33885), .Z(n33883) );
  XNOR U33872 ( .A(n33831), .B(n33837), .Z(n33863) );
  AND U33873 ( .A(n33752), .B(n33886), .Z(n33837) );
  XOR U33874 ( .A(n33842), .B(n33841), .Z(n33831) );
  XNOR U33875 ( .A(n33887), .B(n33838), .Z(n33841) );
  XOR U33876 ( .A(n33888), .B(n33889), .Z(n33838) );
  AND U33877 ( .A(n33890), .B(n33891), .Z(n33889) );
  XOR U33878 ( .A(n33888), .B(n33892), .Z(n33890) );
  XNOR U33879 ( .A(n33893), .B(n33894), .Z(n33887) );
  AND U33880 ( .A(n33895), .B(n33896), .Z(n33894) );
  XOR U33881 ( .A(n33893), .B(n33897), .Z(n33895) );
  XOR U33882 ( .A(n33898), .B(n33899), .Z(n33842) );
  AND U33883 ( .A(n33900), .B(n33901), .Z(n33899) );
  XOR U33884 ( .A(n33898), .B(n33902), .Z(n33900) );
  XNOR U33885 ( .A(n33903), .B(n33788), .Z(n33862) );
  IV U33886 ( .A(n33551), .Z(n33903) );
  XOR U33887 ( .A(n33904), .B(n33855), .Z(n33551) );
  XOR U33888 ( .A(n33848), .B(n33847), .Z(n33855) );
  XNOR U33889 ( .A(n33905), .B(n33844), .Z(n33847) );
  XOR U33890 ( .A(n33906), .B(n33907), .Z(n33844) );
  AND U33891 ( .A(n33908), .B(n33909), .Z(n33907) );
  XOR U33892 ( .A(n33906), .B(n33910), .Z(n33908) );
  XNOR U33893 ( .A(n33911), .B(n33912), .Z(n33905) );
  AND U33894 ( .A(n33913), .B(n33914), .Z(n33912) );
  XOR U33895 ( .A(n33911), .B(n33915), .Z(n33913) );
  XOR U33896 ( .A(n33916), .B(n33917), .Z(n33848) );
  AND U33897 ( .A(n33918), .B(n33919), .Z(n33917) );
  XOR U33898 ( .A(n33916), .B(n33920), .Z(n33918) );
  XNOR U33899 ( .A(n33854), .B(n33849), .Z(n33904) );
  AND U33900 ( .A(n33563), .B(n33921), .Z(n33849) );
  XOR U33901 ( .A(n33922), .B(n33860), .Z(n33854) );
  XNOR U33902 ( .A(n33923), .B(n33924), .Z(n33860) );
  AND U33903 ( .A(n33925), .B(n33926), .Z(n33924) );
  XOR U33904 ( .A(n33923), .B(n33927), .Z(n33925) );
  XNOR U33905 ( .A(n33859), .B(n33851), .Z(n33922) );
  XOR U33906 ( .A(n33928), .B(n33929), .Z(n33851) );
  AND U33907 ( .A(n33930), .B(n33931), .Z(n33929) );
  XOR U33908 ( .A(n33928), .B(n33932), .Z(n33930) );
  XNOR U33909 ( .A(n33933), .B(n33856), .Z(n33859) );
  XOR U33910 ( .A(n33934), .B(n33935), .Z(n33856) );
  AND U33911 ( .A(n33936), .B(n33937), .Z(n33935) );
  XOR U33912 ( .A(n33934), .B(n33938), .Z(n33936) );
  XNOR U33913 ( .A(n33939), .B(n33940), .Z(n33933) );
  AND U33914 ( .A(n33941), .B(n33942), .Z(n33940) );
  XNOR U33915 ( .A(n33939), .B(n33943), .Z(n33941) );
  XOR U33916 ( .A(n33944), .B(n33945), .Z(n33788) );
  AND U33917 ( .A(n33946), .B(n33947), .Z(n33945) );
  XNOR U33918 ( .A(n33944), .B(n33752), .Z(n33947) );
  XOR U33919 ( .A(n33948), .B(n33873), .Z(n33752) );
  XNOR U33920 ( .A(n33949), .B(n33880), .Z(n33873) );
  XOR U33921 ( .A(n33869), .B(n33868), .Z(n33880) );
  XNOR U33922 ( .A(n33950), .B(n33865), .Z(n33868) );
  XOR U33923 ( .A(n33951), .B(n33952), .Z(n33865) );
  AND U33924 ( .A(n33953), .B(n33954), .Z(n33952) );
  XOR U33925 ( .A(n33951), .B(n33955), .Z(n33953) );
  XNOR U33926 ( .A(n33956), .B(n33957), .Z(n33950) );
  NOR U33927 ( .A(n33958), .B(n33959), .Z(n33957) );
  XNOR U33928 ( .A(n33956), .B(n33960), .Z(n33958) );
  XOR U33929 ( .A(n33961), .B(n33962), .Z(n33869) );
  NOR U33930 ( .A(n33963), .B(n33964), .Z(n33962) );
  XNOR U33931 ( .A(n33961), .B(n33965), .Z(n33963) );
  XNOR U33932 ( .A(n33879), .B(n33870), .Z(n33949) );
  XOR U33933 ( .A(n33966), .B(n33967), .Z(n33870) );
  NOR U33934 ( .A(n33968), .B(n33969), .Z(n33967) );
  XNOR U33935 ( .A(n33966), .B(n33970), .Z(n33968) );
  XOR U33936 ( .A(n33971), .B(n33885), .Z(n33879) );
  XNOR U33937 ( .A(n33972), .B(n33973), .Z(n33885) );
  NOR U33938 ( .A(n33974), .B(n33975), .Z(n33973) );
  XNOR U33939 ( .A(n33972), .B(n33976), .Z(n33974) );
  XNOR U33940 ( .A(n33884), .B(n33876), .Z(n33971) );
  XOR U33941 ( .A(n33977), .B(n33978), .Z(n33876) );
  AND U33942 ( .A(n33979), .B(n33980), .Z(n33978) );
  XOR U33943 ( .A(n33977), .B(n33981), .Z(n33979) );
  XNOR U33944 ( .A(n33982), .B(n33881), .Z(n33884) );
  XOR U33945 ( .A(n33983), .B(n33984), .Z(n33881) );
  AND U33946 ( .A(n33985), .B(n33986), .Z(n33984) );
  XOR U33947 ( .A(n33983), .B(n33987), .Z(n33985) );
  XNOR U33948 ( .A(n33988), .B(n33989), .Z(n33982) );
  NOR U33949 ( .A(n33990), .B(n33991), .Z(n33989) );
  XOR U33950 ( .A(n33988), .B(n33992), .Z(n33990) );
  XOR U33951 ( .A(n33874), .B(n33886), .Z(n33948) );
  AND U33952 ( .A(n33794), .B(n33993), .Z(n33886) );
  IV U33953 ( .A(n33773), .Z(n33794) );
  XNOR U33954 ( .A(n33892), .B(n33891), .Z(n33874) );
  XNOR U33955 ( .A(n33994), .B(n33897), .Z(n33891) );
  XOR U33956 ( .A(n33995), .B(n33996), .Z(n33897) );
  NOR U33957 ( .A(n33997), .B(n33998), .Z(n33996) );
  XNOR U33958 ( .A(n33995), .B(n33999), .Z(n33997) );
  XNOR U33959 ( .A(n33896), .B(n33888), .Z(n33994) );
  XOR U33960 ( .A(n34000), .B(n34001), .Z(n33888) );
  AND U33961 ( .A(n34002), .B(n34003), .Z(n34001) );
  XNOR U33962 ( .A(n34000), .B(n34004), .Z(n34002) );
  XNOR U33963 ( .A(n34005), .B(n33893), .Z(n33896) );
  XOR U33964 ( .A(n34006), .B(n34007), .Z(n33893) );
  AND U33965 ( .A(n34008), .B(n34009), .Z(n34007) );
  XOR U33966 ( .A(n34006), .B(n34010), .Z(n34008) );
  XNOR U33967 ( .A(n34011), .B(n34012), .Z(n34005) );
  NOR U33968 ( .A(n34013), .B(n34014), .Z(n34012) );
  XOR U33969 ( .A(n34011), .B(n34015), .Z(n34013) );
  XOR U33970 ( .A(n33902), .B(n33901), .Z(n33892) );
  XNOR U33971 ( .A(n34016), .B(n33898), .Z(n33901) );
  XOR U33972 ( .A(n34017), .B(n34018), .Z(n33898) );
  AND U33973 ( .A(n34019), .B(n34020), .Z(n34018) );
  XOR U33974 ( .A(n34017), .B(n34021), .Z(n34019) );
  XNOR U33975 ( .A(n34022), .B(n34023), .Z(n34016) );
  NOR U33976 ( .A(n34024), .B(n34025), .Z(n34023) );
  XNOR U33977 ( .A(n34022), .B(n34026), .Z(n34024) );
  XOR U33978 ( .A(n34027), .B(n34028), .Z(n33902) );
  NOR U33979 ( .A(n34029), .B(n34030), .Z(n34028) );
  XNOR U33980 ( .A(n34027), .B(n34031), .Z(n34029) );
  XNOR U33981 ( .A(n34032), .B(n33944), .Z(n33946) );
  IV U33982 ( .A(n33563), .Z(n34032) );
  XOR U33983 ( .A(n34033), .B(n33932), .Z(n33563) );
  XOR U33984 ( .A(n33910), .B(n33909), .Z(n33932) );
  XNOR U33985 ( .A(n34034), .B(n33915), .Z(n33909) );
  XOR U33986 ( .A(n34035), .B(n34036), .Z(n33915) );
  NOR U33987 ( .A(n34037), .B(n34038), .Z(n34036) );
  XNOR U33988 ( .A(n34035), .B(n34039), .Z(n34037) );
  XNOR U33989 ( .A(n33914), .B(n33906), .Z(n34034) );
  XOR U33990 ( .A(n34040), .B(n34041), .Z(n33906) );
  AND U33991 ( .A(n34042), .B(n34043), .Z(n34041) );
  XNOR U33992 ( .A(n34040), .B(n34044), .Z(n34042) );
  XNOR U33993 ( .A(n34045), .B(n33911), .Z(n33914) );
  XOR U33994 ( .A(n34046), .B(n34047), .Z(n33911) );
  AND U33995 ( .A(n34048), .B(n34049), .Z(n34047) );
  XOR U33996 ( .A(n34046), .B(n34050), .Z(n34048) );
  XNOR U33997 ( .A(n34051), .B(n34052), .Z(n34045) );
  NOR U33998 ( .A(n34053), .B(n34054), .Z(n34052) );
  XOR U33999 ( .A(n34051), .B(n34055), .Z(n34053) );
  XOR U34000 ( .A(n33920), .B(n33919), .Z(n33910) );
  XNOR U34001 ( .A(n34056), .B(n33916), .Z(n33919) );
  XOR U34002 ( .A(n34057), .B(n34058), .Z(n33916) );
  AND U34003 ( .A(n34059), .B(n34060), .Z(n34058) );
  XOR U34004 ( .A(n34057), .B(n34061), .Z(n34059) );
  XNOR U34005 ( .A(n34062), .B(n34063), .Z(n34056) );
  NOR U34006 ( .A(n34064), .B(n34065), .Z(n34063) );
  XNOR U34007 ( .A(n34062), .B(n34066), .Z(n34064) );
  XOR U34008 ( .A(n34067), .B(n34068), .Z(n33920) );
  NOR U34009 ( .A(n34069), .B(n34070), .Z(n34068) );
  XNOR U34010 ( .A(n34067), .B(n34071), .Z(n34069) );
  XNOR U34011 ( .A(n33931), .B(n33921), .Z(n34033) );
  AND U34012 ( .A(n33792), .B(n34072), .Z(n33921) );
  XNOR U34013 ( .A(n34073), .B(n33938), .Z(n33931) );
  XOR U34014 ( .A(n33927), .B(n33926), .Z(n33938) );
  XNOR U34015 ( .A(n34074), .B(n33923), .Z(n33926) );
  XOR U34016 ( .A(n34075), .B(n34076), .Z(n33923) );
  AND U34017 ( .A(n34077), .B(n34078), .Z(n34076) );
  XOR U34018 ( .A(n34075), .B(n34079), .Z(n34077) );
  XNOR U34019 ( .A(n34080), .B(n34081), .Z(n34074) );
  NOR U34020 ( .A(n34082), .B(n34083), .Z(n34081) );
  XNOR U34021 ( .A(n34080), .B(n34084), .Z(n34082) );
  XOR U34022 ( .A(n34085), .B(n34086), .Z(n33927) );
  NOR U34023 ( .A(n34087), .B(n34088), .Z(n34086) );
  XNOR U34024 ( .A(n34085), .B(n34089), .Z(n34087) );
  XNOR U34025 ( .A(n33937), .B(n33928), .Z(n34073) );
  XOR U34026 ( .A(n34090), .B(n34091), .Z(n33928) );
  NOR U34027 ( .A(n34092), .B(n34093), .Z(n34091) );
  XNOR U34028 ( .A(n34090), .B(n34094), .Z(n34092) );
  XOR U34029 ( .A(n34095), .B(n33943), .Z(n33937) );
  XNOR U34030 ( .A(n34096), .B(n34097), .Z(n33943) );
  NOR U34031 ( .A(n34098), .B(n34099), .Z(n34097) );
  XNOR U34032 ( .A(n34096), .B(n34100), .Z(n34098) );
  XNOR U34033 ( .A(n33942), .B(n33934), .Z(n34095) );
  XOR U34034 ( .A(n34101), .B(n34102), .Z(n33934) );
  AND U34035 ( .A(n34103), .B(n34104), .Z(n34102) );
  XOR U34036 ( .A(n34101), .B(n34105), .Z(n34103) );
  XNOR U34037 ( .A(n34106), .B(n33939), .Z(n33942) );
  XOR U34038 ( .A(n34107), .B(n34108), .Z(n33939) );
  AND U34039 ( .A(n34109), .B(n34110), .Z(n34108) );
  XOR U34040 ( .A(n34107), .B(n34111), .Z(n34109) );
  XNOR U34041 ( .A(n34112), .B(n34113), .Z(n34106) );
  NOR U34042 ( .A(n34114), .B(n34115), .Z(n34113) );
  XOR U34043 ( .A(n34112), .B(n34116), .Z(n34114) );
  AND U34044 ( .A(n33792), .B(n33773), .Z(n33944) );
  XNOR U34045 ( .A(n34117), .B(n33993), .Z(n33773) );
  XOR U34046 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(
        p_input[2048]), .Z(n33993) );
  XOR U34047 ( .A(n33970), .B(n33969), .Z(n34117) );
  XOR U34048 ( .A(n34118), .B(n33981), .Z(n33969) );
  XOR U34049 ( .A(n33955), .B(n33954), .Z(n33981) );
  XNOR U34050 ( .A(n34119), .B(n33960), .Z(n33954) );
  XNOR U34051 ( .A(n8219), .B(p_input[2072]), .Z(n33960) );
  IV U34052 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .Z(n8219) );
  XOR U34053 ( .A(n33951), .B(n33959), .Z(n34119) );
  XOR U34054 ( .A(n34120), .B(n33956), .Z(n33959) );
  XNOR U34055 ( .A(n9214), .B(p_input[2070]), .Z(n33956) );
  IV U34056 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .Z(n9214) );
  XOR U34057 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .B(n17295), 
        .Z(n34120) );
  XNOR U34058 ( .A(n11700), .B(p_input[2066]), .Z(n33951) );
  IV U34059 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .Z(n11700)
         );
  XNOR U34060 ( .A(n33965), .B(n33964), .Z(n33955) );
  XOR U34061 ( .A(n34121), .B(n33961), .Z(n33964) );
  XNOR U34062 ( .A(n11203), .B(p_input[2067]), .Z(n33961) );
  IV U34063 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .Z(n11203)
         );
  XOR U34064 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .B(n17297), 
        .Z(n34121) );
  XNOR U34065 ( .A(n9711), .B(p_input[2069]), .Z(n33965) );
  IV U34066 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .Z(n9711) );
  XNOR U34067 ( .A(n33980), .B(n33966), .Z(n34118) );
  XNOR U34068 ( .A(n10706), .B(p_input[2049]), .Z(n33966) );
  IV U34069 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n10706) );
  XNOR U34070 ( .A(n34122), .B(n33987), .Z(n33980) );
  XNOR U34071 ( .A(n33976), .B(n33975), .Z(n33987) );
  XOR U34072 ( .A(n34123), .B(n33972), .Z(n33975) );
  XNOR U34073 ( .A(n7225), .B(p_input[2074]), .Z(n33972) );
  IV U34074 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .Z(n7225) );
  XOR U34075 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .B(n17300), 
        .Z(n34123) );
  XNOR U34076 ( .A(n6230), .B(p_input[2076]), .Z(n33976) );
  IV U34077 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .Z(n6230) );
  XNOR U34078 ( .A(n33986), .B(n33977), .Z(n34122) );
  XNOR U34079 ( .A(n12197), .B(p_input[2065]), .Z(n33977) );
  IV U34080 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .Z(n12197)
         );
  XOR U34081 ( .A(n34124), .B(n33992), .Z(n33986) );
  XNOR U34082 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .B(
        p_input[2079]), .Z(n33992) );
  XOR U34083 ( .A(n33983), .B(n33991), .Z(n34124) );
  XOR U34084 ( .A(n34125), .B(n33988), .Z(n33991) );
  XNOR U34085 ( .A(n5733), .B(p_input[2077]), .Z(n33988) );
  IV U34086 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .Z(n5733) );
  XOR U34087 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .B(n17305), 
        .Z(n34125) );
  XNOR U34088 ( .A(n7722), .B(p_input[2073]), .Z(n33983) );
  IV U34089 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .Z(n7722) );
  XNOR U34090 ( .A(n34004), .B(n34003), .Z(n33970) );
  XNOR U34091 ( .A(n34126), .B(n34010), .Z(n34003) );
  XNOR U34092 ( .A(n33999), .B(n33998), .Z(n34010) );
  XOR U34093 ( .A(n34127), .B(n33995), .Z(n33998) );
  XNOR U34094 ( .A(n15182), .B(p_input[2059]), .Z(n33995) );
  IV U34095 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n15182)
         );
  XOR U34096 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(n16451), 
        .Z(n34127) );
  XNOR U34097 ( .A(n14187), .B(p_input[2061]), .Z(n33999) );
  IV U34098 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n14187)
         );
  XNOR U34099 ( .A(n34009), .B(n34000), .Z(n34126) );
  XNOR U34100 ( .A(n5236), .B(p_input[2050]), .Z(n34000) );
  IV U34101 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n5236) );
  XOR U34102 ( .A(n34128), .B(n34015), .Z(n34009) );
  XNOR U34103 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .B(
        p_input[2064]), .Z(n34015) );
  XOR U34104 ( .A(n34006), .B(n34014), .Z(n34128) );
  XOR U34105 ( .A(n34129), .B(n34011), .Z(n34014) );
  XNOR U34106 ( .A(n13690), .B(p_input[2062]), .Z(n34011) );
  IV U34107 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n13690)
         );
  XOR U34108 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(n16456), 
        .Z(n34129) );
  XNOR U34109 ( .A(n15679), .B(p_input[2058]), .Z(n34006) );
  IV U34110 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n15679)
         );
  XNOR U34111 ( .A(n34021), .B(n34020), .Z(n34004) );
  XNOR U34112 ( .A(n34130), .B(n34026), .Z(n34020) );
  XNOR U34113 ( .A(n736), .B(p_input[2057]), .Z(n34026) );
  IV U34114 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .Z(n736) );
  XOR U34115 ( .A(n34017), .B(n34025), .Z(n34130) );
  XOR U34116 ( .A(n34131), .B(n34022), .Z(n34025) );
  XNOR U34117 ( .A(n1738), .B(p_input[2055]), .Z(n34022) );
  IV U34118 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .Z(n1738) );
  XOR U34119 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(n17312), 
        .Z(n34131) );
  XNOR U34120 ( .A(n3734), .B(p_input[2051]), .Z(n34017) );
  IV U34121 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .Z(n3734) );
  XNOR U34122 ( .A(n34031), .B(n34030), .Z(n34021) );
  XOR U34123 ( .A(n34132), .B(n34027), .Z(n34030) );
  XNOR U34124 ( .A(n3235), .B(p_input[2052]), .Z(n34027) );
  IV U34125 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .Z(n3235) );
  XOR U34126 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(n17314), 
        .Z(n34132) );
  XNOR U34127 ( .A(n2237), .B(p_input[2054]), .Z(n34031) );
  IV U34128 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .Z(n2237) );
  XOR U34129 ( .A(n34133), .B(n34094), .Z(n33792) );
  XNOR U34130 ( .A(n34044), .B(n34043), .Z(n34094) );
  XNOR U34131 ( .A(n34134), .B(n34050), .Z(n34043) );
  XNOR U34132 ( .A(n34039), .B(n34038), .Z(n34050) );
  XOR U34133 ( .A(n34135), .B(n34035), .Z(n34038) );
  XNOR U34134 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n16737), .Z(n34035) );
  IV U34135 ( .A(p_input[2059]), .Z(n16737) );
  XOR U34136 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n16451), .Z(n34135) );
  IV U34137 ( .A(p_input[2060]), .Z(n16451) );
  XOR U34138 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[2061]), .Z(
        n34039) );
  XNOR U34139 ( .A(n34049), .B(n34040), .Z(n34134) );
  XNOR U34140 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n16452), .Z(n34040) );
  IV U34141 ( .A(p_input[2050]), .Z(n16452) );
  XOR U34142 ( .A(n34136), .B(n34055), .Z(n34049) );
  XNOR U34143 ( .A(\knn_comb_/min_val_out[0][16] ), .B(p_input[2064]), .Z(
        n34055) );
  XOR U34144 ( .A(n34046), .B(n34054), .Z(n34136) );
  XOR U34145 ( .A(n34137), .B(n34051), .Z(n34054) );
  XOR U34146 ( .A(\knn_comb_/min_val_out[0][14] ), .B(p_input[2062]), .Z(
        n34051) );
  XOR U34147 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n16456), .Z(n34137) );
  IV U34148 ( .A(p_input[2063]), .Z(n16456) );
  XNOR U34149 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n16740), .Z(n34046) );
  IV U34150 ( .A(p_input[2058]), .Z(n16740) );
  XNOR U34151 ( .A(n34061), .B(n34060), .Z(n34044) );
  XNOR U34152 ( .A(n34138), .B(n34066), .Z(n34060) );
  XNOR U34153 ( .A(n742), .B(p_input[2057]), .Z(n34066) );
  IV U34154 ( .A(\knn_comb_/min_val_out[0][9] ), .Z(n742) );
  XOR U34155 ( .A(n34057), .B(n34065), .Z(n34138) );
  XOR U34156 ( .A(n34139), .B(n34062), .Z(n34065) );
  XNOR U34157 ( .A(n1742), .B(p_input[2055]), .Z(n34062) );
  IV U34158 ( .A(\knn_comb_/min_val_out[0][7] ), .Z(n1742) );
  XOR U34159 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n17312), .Z(n34139) );
  IV U34160 ( .A(p_input[2056]), .Z(n17312) );
  XNOR U34161 ( .A(n3738), .B(p_input[2051]), .Z(n34057) );
  IV U34162 ( .A(\knn_comb_/min_val_out[0][3] ), .Z(n3738) );
  XNOR U34163 ( .A(n34071), .B(n34070), .Z(n34061) );
  XOR U34164 ( .A(n34140), .B(n34067), .Z(n34070) );
  XNOR U34165 ( .A(n3239), .B(p_input[2052]), .Z(n34067) );
  IV U34166 ( .A(\knn_comb_/min_val_out[0][4] ), .Z(n3239) );
  XOR U34167 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n17314), .Z(n34140) );
  IV U34168 ( .A(p_input[2053]), .Z(n17314) );
  XNOR U34169 ( .A(n2241), .B(p_input[2054]), .Z(n34071) );
  IV U34170 ( .A(\knn_comb_/min_val_out[0][6] ), .Z(n2241) );
  XOR U34171 ( .A(n34093), .B(n34072), .Z(n34133) );
  XOR U34172 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[2048]), .Z(n34072) );
  XOR U34173 ( .A(n34141), .B(n34105), .Z(n34093) );
  XOR U34174 ( .A(n34079), .B(n34078), .Z(n34105) );
  XNOR U34175 ( .A(n34142), .B(n34084), .Z(n34078) );
  XOR U34176 ( .A(\knn_comb_/min_val_out[0][24] ), .B(p_input[2072]), .Z(
        n34084) );
  XOR U34177 ( .A(n34075), .B(n34083), .Z(n34142) );
  XOR U34178 ( .A(n34143), .B(n34080), .Z(n34083) );
  XOR U34179 ( .A(\knn_comb_/min_val_out[0][22] ), .B(p_input[2070]), .Z(
        n34080) );
  XOR U34180 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n17295), .Z(n34143) );
  IV U34181 ( .A(p_input[2071]), .Z(n17295) );
  XNOR U34182 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n16727), .Z(n34075) );
  IV U34183 ( .A(p_input[2066]), .Z(n16727) );
  XNOR U34184 ( .A(n34089), .B(n34088), .Z(n34079) );
  XOR U34185 ( .A(n34144), .B(n34085), .Z(n34088) );
  XOR U34186 ( .A(\knn_comb_/min_val_out[0][19] ), .B(p_input[2067]), .Z(
        n34085) );
  XOR U34187 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n17297), .Z(n34144) );
  IV U34188 ( .A(p_input[2068]), .Z(n17297) );
  XOR U34189 ( .A(\knn_comb_/min_val_out[0][21] ), .B(p_input[2069]), .Z(
        n34089) );
  XNOR U34190 ( .A(n34104), .B(n34090), .Z(n34141) );
  XNOR U34191 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n16729), .Z(n34090) );
  IV U34192 ( .A(p_input[2049]), .Z(n16729) );
  XNOR U34193 ( .A(n34145), .B(n34111), .Z(n34104) );
  XNOR U34194 ( .A(n34100), .B(n34099), .Z(n34111) );
  XOR U34195 ( .A(n34146), .B(n34096), .Z(n34099) );
  XNOR U34196 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n16444), .Z(n34096) );
  IV U34197 ( .A(p_input[2074]), .Z(n16444) );
  XOR U34198 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n17300), .Z(n34146) );
  IV U34199 ( .A(p_input[2075]), .Z(n17300) );
  XOR U34200 ( .A(\knn_comb_/min_val_out[0][28] ), .B(p_input[2076]), .Z(
        n34100) );
  XNOR U34201 ( .A(n34110), .B(n34101), .Z(n34145) );
  XNOR U34202 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n16732), .Z(n34101) );
  IV U34203 ( .A(p_input[2065]), .Z(n16732) );
  XOR U34204 ( .A(n34147), .B(n34116), .Z(n34110) );
  XNOR U34205 ( .A(\knn_comb_/min_val_out[0][31] ), .B(p_input[2079]), .Z(
        n34116) );
  XOR U34206 ( .A(n34107), .B(n34115), .Z(n34147) );
  XOR U34207 ( .A(n34148), .B(n34112), .Z(n34115) );
  XOR U34208 ( .A(\knn_comb_/min_val_out[0][29] ), .B(p_input[2077]), .Z(
        n34112) );
  XOR U34209 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n17305), .Z(n34148) );
  IV U34210 ( .A(p_input[2078]), .Z(n17305) );
  XNOR U34211 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n16448), .Z(n34107) );
  IV U34212 ( .A(p_input[2073]), .Z(n16448) );
endmodule

