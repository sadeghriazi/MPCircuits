
module knn_comb_BMR_W16_K1_N16 ( p_input, o );
  input [271:0] p_input;
  output [15:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485;
  assign \knn_comb_/min_val_out[0][0]  = p_input[240];
  assign \knn_comb_/min_val_out[0][1]  = p_input[241];
  assign \knn_comb_/min_val_out[0][2]  = p_input[242];
  assign \knn_comb_/min_val_out[0][3]  = p_input[243];
  assign \knn_comb_/min_val_out[0][4]  = p_input[244];
  assign \knn_comb_/min_val_out[0][5]  = p_input[245];
  assign \knn_comb_/min_val_out[0][6]  = p_input[246];
  assign \knn_comb_/min_val_out[0][7]  = p_input[247];
  assign \knn_comb_/min_val_out[0][8]  = p_input[248];
  assign \knn_comb_/min_val_out[0][9]  = p_input[249];
  assign \knn_comb_/min_val_out[0][10]  = p_input[250];
  assign \knn_comb_/min_val_out[0][11]  = p_input[251];
  assign \knn_comb_/min_val_out[0][12]  = p_input[252];
  assign \knn_comb_/min_val_out[0][13]  = p_input[253];
  assign \knn_comb_/min_val_out[0][14]  = p_input[254];
  assign \knn_comb_/min_val_out[0][15]  = p_input[255];

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(n3), .B(n4), .Z(n1) );
  XNOR U3 ( .A(p_input[9]), .B(n2), .Z(n4) );
  XOR U4 ( .A(n5), .B(n6), .Z(n2) );
  AND U5 ( .A(n7), .B(n8), .Z(n6) );
  XNOR U6 ( .A(p_input[25]), .B(n5), .Z(n8) );
  XOR U7 ( .A(n9), .B(n10), .Z(n5) );
  AND U8 ( .A(n11), .B(n12), .Z(n10) );
  XNOR U9 ( .A(p_input[41]), .B(n9), .Z(n12) );
  XOR U10 ( .A(n13), .B(n14), .Z(n9) );
  AND U11 ( .A(n15), .B(n16), .Z(n14) );
  XNOR U12 ( .A(p_input[57]), .B(n13), .Z(n16) );
  XOR U13 ( .A(n17), .B(n18), .Z(n13) );
  AND U14 ( .A(n19), .B(n20), .Z(n18) );
  XNOR U15 ( .A(p_input[73]), .B(n17), .Z(n20) );
  XOR U16 ( .A(n21), .B(n22), .Z(n17) );
  AND U17 ( .A(n23), .B(n24), .Z(n22) );
  XNOR U18 ( .A(p_input[89]), .B(n21), .Z(n24) );
  XOR U19 ( .A(n25), .B(n26), .Z(n21) );
  AND U20 ( .A(n27), .B(n28), .Z(n26) );
  XNOR U21 ( .A(p_input[105]), .B(n25), .Z(n28) );
  XOR U22 ( .A(n29), .B(n30), .Z(n25) );
  AND U23 ( .A(n31), .B(n32), .Z(n30) );
  XNOR U24 ( .A(p_input[121]), .B(n29), .Z(n32) );
  XOR U25 ( .A(n33), .B(n34), .Z(n29) );
  AND U26 ( .A(n35), .B(n36), .Z(n34) );
  XNOR U27 ( .A(p_input[137]), .B(n33), .Z(n36) );
  XOR U28 ( .A(n37), .B(n38), .Z(n33) );
  AND U29 ( .A(n39), .B(n40), .Z(n38) );
  XNOR U30 ( .A(p_input[153]), .B(n37), .Z(n40) );
  XOR U31 ( .A(n41), .B(n42), .Z(n37) );
  AND U32 ( .A(n43), .B(n44), .Z(n42) );
  XNOR U33 ( .A(p_input[169]), .B(n41), .Z(n44) );
  XOR U34 ( .A(n45), .B(n46), .Z(n41) );
  AND U35 ( .A(n47), .B(n48), .Z(n46) );
  XNOR U36 ( .A(p_input[185]), .B(n45), .Z(n48) );
  XOR U37 ( .A(n49), .B(n50), .Z(n45) );
  AND U38 ( .A(n51), .B(n52), .Z(n50) );
  XNOR U39 ( .A(p_input[201]), .B(n49), .Z(n52) );
  XNOR U40 ( .A(n53), .B(n54), .Z(n49) );
  AND U41 ( .A(n55), .B(n56), .Z(n54) );
  XOR U42 ( .A(p_input[217]), .B(n53), .Z(n56) );
  XOR U43 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n57), .Z(n53) );
  AND U44 ( .A(n58), .B(n59), .Z(n57) );
  XOR U45 ( .A(p_input[233]), .B(\knn_comb_/min_val_out[0][9] ), .Z(n59) );
  XNOR U46 ( .A(n60), .B(n61), .Z(o[8]) );
  AND U47 ( .A(n3), .B(n62), .Z(n60) );
  XNOR U48 ( .A(p_input[8]), .B(n61), .Z(n62) );
  XOR U49 ( .A(n63), .B(n64), .Z(n61) );
  AND U50 ( .A(n7), .B(n65), .Z(n64) );
  XNOR U51 ( .A(p_input[24]), .B(n63), .Z(n65) );
  XOR U52 ( .A(n66), .B(n67), .Z(n63) );
  AND U53 ( .A(n11), .B(n68), .Z(n67) );
  XNOR U54 ( .A(p_input[40]), .B(n66), .Z(n68) );
  XOR U55 ( .A(n69), .B(n70), .Z(n66) );
  AND U56 ( .A(n15), .B(n71), .Z(n70) );
  XNOR U57 ( .A(p_input[56]), .B(n69), .Z(n71) );
  XOR U58 ( .A(n72), .B(n73), .Z(n69) );
  AND U59 ( .A(n19), .B(n74), .Z(n73) );
  XNOR U60 ( .A(p_input[72]), .B(n72), .Z(n74) );
  XOR U61 ( .A(n75), .B(n76), .Z(n72) );
  AND U62 ( .A(n23), .B(n77), .Z(n76) );
  XNOR U63 ( .A(p_input[88]), .B(n75), .Z(n77) );
  XOR U64 ( .A(n78), .B(n79), .Z(n75) );
  AND U65 ( .A(n27), .B(n80), .Z(n79) );
  XNOR U66 ( .A(p_input[104]), .B(n78), .Z(n80) );
  XOR U67 ( .A(n81), .B(n82), .Z(n78) );
  AND U68 ( .A(n31), .B(n83), .Z(n82) );
  XNOR U69 ( .A(p_input[120]), .B(n81), .Z(n83) );
  XOR U70 ( .A(n84), .B(n85), .Z(n81) );
  AND U71 ( .A(n35), .B(n86), .Z(n85) );
  XNOR U72 ( .A(p_input[136]), .B(n84), .Z(n86) );
  XOR U73 ( .A(n87), .B(n88), .Z(n84) );
  AND U74 ( .A(n39), .B(n89), .Z(n88) );
  XNOR U75 ( .A(p_input[152]), .B(n87), .Z(n89) );
  XOR U76 ( .A(n90), .B(n91), .Z(n87) );
  AND U77 ( .A(n43), .B(n92), .Z(n91) );
  XNOR U78 ( .A(p_input[168]), .B(n90), .Z(n92) );
  XOR U79 ( .A(n93), .B(n94), .Z(n90) );
  AND U80 ( .A(n47), .B(n95), .Z(n94) );
  XNOR U81 ( .A(p_input[184]), .B(n93), .Z(n95) );
  XOR U82 ( .A(n96), .B(n97), .Z(n93) );
  AND U83 ( .A(n51), .B(n98), .Z(n97) );
  XNOR U84 ( .A(p_input[200]), .B(n96), .Z(n98) );
  XNOR U85 ( .A(n99), .B(n100), .Z(n96) );
  AND U86 ( .A(n55), .B(n101), .Z(n100) );
  XOR U87 ( .A(p_input[216]), .B(n99), .Z(n101) );
  XOR U88 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n102), .Z(n99) );
  AND U89 ( .A(n58), .B(n103), .Z(n102) );
  XOR U90 ( .A(p_input[232]), .B(\knn_comb_/min_val_out[0][8] ), .Z(n103) );
  XNOR U91 ( .A(n104), .B(n105), .Z(o[7]) );
  AND U92 ( .A(n3), .B(n106), .Z(n104) );
  XNOR U93 ( .A(p_input[7]), .B(n105), .Z(n106) );
  XOR U94 ( .A(n107), .B(n108), .Z(n105) );
  AND U95 ( .A(n7), .B(n109), .Z(n108) );
  XNOR U96 ( .A(p_input[23]), .B(n107), .Z(n109) );
  XOR U97 ( .A(n110), .B(n111), .Z(n107) );
  AND U98 ( .A(n11), .B(n112), .Z(n111) );
  XNOR U99 ( .A(p_input[39]), .B(n110), .Z(n112) );
  XOR U100 ( .A(n113), .B(n114), .Z(n110) );
  AND U101 ( .A(n15), .B(n115), .Z(n114) );
  XNOR U102 ( .A(p_input[55]), .B(n113), .Z(n115) );
  XOR U103 ( .A(n116), .B(n117), .Z(n113) );
  AND U104 ( .A(n19), .B(n118), .Z(n117) );
  XNOR U105 ( .A(p_input[71]), .B(n116), .Z(n118) );
  XOR U106 ( .A(n119), .B(n120), .Z(n116) );
  AND U107 ( .A(n23), .B(n121), .Z(n120) );
  XNOR U108 ( .A(p_input[87]), .B(n119), .Z(n121) );
  XOR U109 ( .A(n122), .B(n123), .Z(n119) );
  AND U110 ( .A(n27), .B(n124), .Z(n123) );
  XNOR U111 ( .A(p_input[103]), .B(n122), .Z(n124) );
  XOR U112 ( .A(n125), .B(n126), .Z(n122) );
  AND U113 ( .A(n31), .B(n127), .Z(n126) );
  XNOR U114 ( .A(p_input[119]), .B(n125), .Z(n127) );
  XOR U115 ( .A(n128), .B(n129), .Z(n125) );
  AND U116 ( .A(n35), .B(n130), .Z(n129) );
  XNOR U117 ( .A(p_input[135]), .B(n128), .Z(n130) );
  XOR U118 ( .A(n131), .B(n132), .Z(n128) );
  AND U119 ( .A(n39), .B(n133), .Z(n132) );
  XNOR U120 ( .A(p_input[151]), .B(n131), .Z(n133) );
  XOR U121 ( .A(n134), .B(n135), .Z(n131) );
  AND U122 ( .A(n43), .B(n136), .Z(n135) );
  XNOR U123 ( .A(p_input[167]), .B(n134), .Z(n136) );
  XOR U124 ( .A(n137), .B(n138), .Z(n134) );
  AND U125 ( .A(n47), .B(n139), .Z(n138) );
  XNOR U126 ( .A(p_input[183]), .B(n137), .Z(n139) );
  XOR U127 ( .A(n140), .B(n141), .Z(n137) );
  AND U128 ( .A(n51), .B(n142), .Z(n141) );
  XNOR U129 ( .A(p_input[199]), .B(n140), .Z(n142) );
  XNOR U130 ( .A(n143), .B(n144), .Z(n140) );
  AND U131 ( .A(n55), .B(n145), .Z(n144) );
  XOR U132 ( .A(p_input[215]), .B(n143), .Z(n145) );
  XOR U133 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n146), .Z(n143) );
  AND U134 ( .A(n58), .B(n147), .Z(n146) );
  XOR U135 ( .A(p_input[231]), .B(\knn_comb_/min_val_out[0][7] ), .Z(n147) );
  XNOR U136 ( .A(n148), .B(n149), .Z(o[6]) );
  AND U137 ( .A(n3), .B(n150), .Z(n148) );
  XNOR U138 ( .A(p_input[6]), .B(n149), .Z(n150) );
  XOR U139 ( .A(n151), .B(n152), .Z(n149) );
  AND U140 ( .A(n7), .B(n153), .Z(n152) );
  XNOR U141 ( .A(p_input[22]), .B(n151), .Z(n153) );
  XOR U142 ( .A(n154), .B(n155), .Z(n151) );
  AND U143 ( .A(n11), .B(n156), .Z(n155) );
  XNOR U144 ( .A(p_input[38]), .B(n154), .Z(n156) );
  XOR U145 ( .A(n157), .B(n158), .Z(n154) );
  AND U146 ( .A(n15), .B(n159), .Z(n158) );
  XNOR U147 ( .A(p_input[54]), .B(n157), .Z(n159) );
  XOR U148 ( .A(n160), .B(n161), .Z(n157) );
  AND U149 ( .A(n19), .B(n162), .Z(n161) );
  XNOR U150 ( .A(p_input[70]), .B(n160), .Z(n162) );
  XOR U151 ( .A(n163), .B(n164), .Z(n160) );
  AND U152 ( .A(n23), .B(n165), .Z(n164) );
  XNOR U153 ( .A(p_input[86]), .B(n163), .Z(n165) );
  XOR U154 ( .A(n166), .B(n167), .Z(n163) );
  AND U155 ( .A(n27), .B(n168), .Z(n167) );
  XNOR U156 ( .A(p_input[102]), .B(n166), .Z(n168) );
  XOR U157 ( .A(n169), .B(n170), .Z(n166) );
  AND U158 ( .A(n31), .B(n171), .Z(n170) );
  XNOR U159 ( .A(p_input[118]), .B(n169), .Z(n171) );
  XOR U160 ( .A(n172), .B(n173), .Z(n169) );
  AND U161 ( .A(n35), .B(n174), .Z(n173) );
  XNOR U162 ( .A(p_input[134]), .B(n172), .Z(n174) );
  XOR U163 ( .A(n175), .B(n176), .Z(n172) );
  AND U164 ( .A(n39), .B(n177), .Z(n176) );
  XNOR U165 ( .A(p_input[150]), .B(n175), .Z(n177) );
  XOR U166 ( .A(n178), .B(n179), .Z(n175) );
  AND U167 ( .A(n43), .B(n180), .Z(n179) );
  XNOR U168 ( .A(p_input[166]), .B(n178), .Z(n180) );
  XOR U169 ( .A(n181), .B(n182), .Z(n178) );
  AND U170 ( .A(n47), .B(n183), .Z(n182) );
  XNOR U171 ( .A(p_input[182]), .B(n181), .Z(n183) );
  XOR U172 ( .A(n184), .B(n185), .Z(n181) );
  AND U173 ( .A(n51), .B(n186), .Z(n185) );
  XNOR U174 ( .A(p_input[198]), .B(n184), .Z(n186) );
  XNOR U175 ( .A(n187), .B(n188), .Z(n184) );
  AND U176 ( .A(n55), .B(n189), .Z(n188) );
  XOR U177 ( .A(p_input[214]), .B(n187), .Z(n189) );
  XOR U178 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n190), .Z(n187) );
  AND U179 ( .A(n58), .B(n191), .Z(n190) );
  XOR U180 ( .A(p_input[230]), .B(\knn_comb_/min_val_out[0][6] ), .Z(n191) );
  XNOR U181 ( .A(n192), .B(n193), .Z(o[5]) );
  AND U182 ( .A(n3), .B(n194), .Z(n192) );
  XNOR U183 ( .A(p_input[5]), .B(n193), .Z(n194) );
  XOR U184 ( .A(n195), .B(n196), .Z(n193) );
  AND U185 ( .A(n7), .B(n197), .Z(n196) );
  XNOR U186 ( .A(p_input[21]), .B(n195), .Z(n197) );
  XOR U187 ( .A(n198), .B(n199), .Z(n195) );
  AND U188 ( .A(n11), .B(n200), .Z(n199) );
  XNOR U189 ( .A(p_input[37]), .B(n198), .Z(n200) );
  XOR U190 ( .A(n201), .B(n202), .Z(n198) );
  AND U191 ( .A(n15), .B(n203), .Z(n202) );
  XNOR U192 ( .A(p_input[53]), .B(n201), .Z(n203) );
  XOR U193 ( .A(n204), .B(n205), .Z(n201) );
  AND U194 ( .A(n19), .B(n206), .Z(n205) );
  XNOR U195 ( .A(p_input[69]), .B(n204), .Z(n206) );
  XOR U196 ( .A(n207), .B(n208), .Z(n204) );
  AND U197 ( .A(n23), .B(n209), .Z(n208) );
  XNOR U198 ( .A(p_input[85]), .B(n207), .Z(n209) );
  XOR U199 ( .A(n210), .B(n211), .Z(n207) );
  AND U200 ( .A(n27), .B(n212), .Z(n211) );
  XNOR U201 ( .A(p_input[101]), .B(n210), .Z(n212) );
  XOR U202 ( .A(n213), .B(n214), .Z(n210) );
  AND U203 ( .A(n31), .B(n215), .Z(n214) );
  XNOR U204 ( .A(p_input[117]), .B(n213), .Z(n215) );
  XOR U205 ( .A(n216), .B(n217), .Z(n213) );
  AND U206 ( .A(n35), .B(n218), .Z(n217) );
  XNOR U207 ( .A(p_input[133]), .B(n216), .Z(n218) );
  XOR U208 ( .A(n219), .B(n220), .Z(n216) );
  AND U209 ( .A(n39), .B(n221), .Z(n220) );
  XNOR U210 ( .A(p_input[149]), .B(n219), .Z(n221) );
  XOR U211 ( .A(n222), .B(n223), .Z(n219) );
  AND U212 ( .A(n43), .B(n224), .Z(n223) );
  XNOR U213 ( .A(p_input[165]), .B(n222), .Z(n224) );
  XOR U214 ( .A(n225), .B(n226), .Z(n222) );
  AND U215 ( .A(n47), .B(n227), .Z(n226) );
  XNOR U216 ( .A(p_input[181]), .B(n225), .Z(n227) );
  XOR U217 ( .A(n228), .B(n229), .Z(n225) );
  AND U218 ( .A(n51), .B(n230), .Z(n229) );
  XNOR U219 ( .A(p_input[197]), .B(n228), .Z(n230) );
  XNOR U220 ( .A(n231), .B(n232), .Z(n228) );
  AND U221 ( .A(n55), .B(n233), .Z(n232) );
  XOR U222 ( .A(p_input[213]), .B(n231), .Z(n233) );
  XOR U223 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n234), .Z(n231) );
  AND U224 ( .A(n58), .B(n235), .Z(n234) );
  XOR U225 ( .A(p_input[229]), .B(\knn_comb_/min_val_out[0][5] ), .Z(n235) );
  XNOR U226 ( .A(n236), .B(n237), .Z(o[4]) );
  AND U227 ( .A(n3), .B(n238), .Z(n236) );
  XNOR U228 ( .A(p_input[4]), .B(n237), .Z(n238) );
  XOR U229 ( .A(n239), .B(n240), .Z(n237) );
  AND U230 ( .A(n7), .B(n241), .Z(n240) );
  XNOR U231 ( .A(p_input[20]), .B(n239), .Z(n241) );
  XOR U232 ( .A(n242), .B(n243), .Z(n239) );
  AND U233 ( .A(n11), .B(n244), .Z(n243) );
  XNOR U234 ( .A(p_input[36]), .B(n242), .Z(n244) );
  XOR U235 ( .A(n245), .B(n246), .Z(n242) );
  AND U236 ( .A(n15), .B(n247), .Z(n246) );
  XNOR U237 ( .A(p_input[52]), .B(n245), .Z(n247) );
  XOR U238 ( .A(n248), .B(n249), .Z(n245) );
  AND U239 ( .A(n19), .B(n250), .Z(n249) );
  XNOR U240 ( .A(p_input[68]), .B(n248), .Z(n250) );
  XOR U241 ( .A(n251), .B(n252), .Z(n248) );
  AND U242 ( .A(n23), .B(n253), .Z(n252) );
  XNOR U243 ( .A(p_input[84]), .B(n251), .Z(n253) );
  XOR U244 ( .A(n254), .B(n255), .Z(n251) );
  AND U245 ( .A(n27), .B(n256), .Z(n255) );
  XNOR U246 ( .A(p_input[100]), .B(n254), .Z(n256) );
  XOR U247 ( .A(n257), .B(n258), .Z(n254) );
  AND U248 ( .A(n31), .B(n259), .Z(n258) );
  XNOR U249 ( .A(p_input[116]), .B(n257), .Z(n259) );
  XOR U250 ( .A(n260), .B(n261), .Z(n257) );
  AND U251 ( .A(n35), .B(n262), .Z(n261) );
  XNOR U252 ( .A(p_input[132]), .B(n260), .Z(n262) );
  XOR U253 ( .A(n263), .B(n264), .Z(n260) );
  AND U254 ( .A(n39), .B(n265), .Z(n264) );
  XNOR U255 ( .A(p_input[148]), .B(n263), .Z(n265) );
  XOR U256 ( .A(n266), .B(n267), .Z(n263) );
  AND U257 ( .A(n43), .B(n268), .Z(n267) );
  XNOR U258 ( .A(p_input[164]), .B(n266), .Z(n268) );
  XOR U259 ( .A(n269), .B(n270), .Z(n266) );
  AND U260 ( .A(n47), .B(n271), .Z(n270) );
  XNOR U261 ( .A(p_input[180]), .B(n269), .Z(n271) );
  XOR U262 ( .A(n272), .B(n273), .Z(n269) );
  AND U263 ( .A(n51), .B(n274), .Z(n273) );
  XNOR U264 ( .A(p_input[196]), .B(n272), .Z(n274) );
  XNOR U265 ( .A(n275), .B(n276), .Z(n272) );
  AND U266 ( .A(n55), .B(n277), .Z(n276) );
  XOR U267 ( .A(p_input[212]), .B(n275), .Z(n277) );
  XOR U268 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n278), .Z(n275) );
  AND U269 ( .A(n58), .B(n279), .Z(n278) );
  XOR U270 ( .A(p_input[228]), .B(\knn_comb_/min_val_out[0][4] ), .Z(n279) );
  XNOR U271 ( .A(n280), .B(n281), .Z(o[3]) );
  AND U272 ( .A(n3), .B(n282), .Z(n280) );
  XNOR U273 ( .A(p_input[3]), .B(n281), .Z(n282) );
  XOR U274 ( .A(n283), .B(n284), .Z(n281) );
  AND U275 ( .A(n7), .B(n285), .Z(n284) );
  XNOR U276 ( .A(p_input[19]), .B(n283), .Z(n285) );
  XOR U277 ( .A(n286), .B(n287), .Z(n283) );
  AND U278 ( .A(n11), .B(n288), .Z(n287) );
  XNOR U279 ( .A(p_input[35]), .B(n286), .Z(n288) );
  XOR U280 ( .A(n289), .B(n290), .Z(n286) );
  AND U281 ( .A(n15), .B(n291), .Z(n290) );
  XNOR U282 ( .A(p_input[51]), .B(n289), .Z(n291) );
  XOR U283 ( .A(n292), .B(n293), .Z(n289) );
  AND U284 ( .A(n19), .B(n294), .Z(n293) );
  XNOR U285 ( .A(p_input[67]), .B(n292), .Z(n294) );
  XOR U286 ( .A(n295), .B(n296), .Z(n292) );
  AND U287 ( .A(n23), .B(n297), .Z(n296) );
  XNOR U288 ( .A(p_input[83]), .B(n295), .Z(n297) );
  XOR U289 ( .A(n298), .B(n299), .Z(n295) );
  AND U290 ( .A(n27), .B(n300), .Z(n299) );
  XNOR U291 ( .A(p_input[99]), .B(n298), .Z(n300) );
  XOR U292 ( .A(n301), .B(n302), .Z(n298) );
  AND U293 ( .A(n31), .B(n303), .Z(n302) );
  XNOR U294 ( .A(p_input[115]), .B(n301), .Z(n303) );
  XOR U295 ( .A(n304), .B(n305), .Z(n301) );
  AND U296 ( .A(n35), .B(n306), .Z(n305) );
  XNOR U297 ( .A(p_input[131]), .B(n304), .Z(n306) );
  XOR U298 ( .A(n307), .B(n308), .Z(n304) );
  AND U299 ( .A(n39), .B(n309), .Z(n308) );
  XNOR U300 ( .A(p_input[147]), .B(n307), .Z(n309) );
  XOR U301 ( .A(n310), .B(n311), .Z(n307) );
  AND U302 ( .A(n43), .B(n312), .Z(n311) );
  XNOR U303 ( .A(p_input[163]), .B(n310), .Z(n312) );
  XOR U304 ( .A(n313), .B(n314), .Z(n310) );
  AND U305 ( .A(n47), .B(n315), .Z(n314) );
  XNOR U306 ( .A(p_input[179]), .B(n313), .Z(n315) );
  XOR U307 ( .A(n316), .B(n317), .Z(n313) );
  AND U308 ( .A(n51), .B(n318), .Z(n317) );
  XNOR U309 ( .A(p_input[195]), .B(n316), .Z(n318) );
  XNOR U310 ( .A(n319), .B(n320), .Z(n316) );
  AND U311 ( .A(n55), .B(n321), .Z(n320) );
  XOR U312 ( .A(p_input[211]), .B(n319), .Z(n321) );
  XOR U313 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n322), .Z(n319) );
  AND U314 ( .A(n58), .B(n323), .Z(n322) );
  XOR U315 ( .A(p_input[227]), .B(\knn_comb_/min_val_out[0][3] ), .Z(n323) );
  XNOR U316 ( .A(n324), .B(n325), .Z(o[2]) );
  AND U317 ( .A(n3), .B(n326), .Z(n324) );
  XNOR U318 ( .A(p_input[2]), .B(n325), .Z(n326) );
  XOR U319 ( .A(n327), .B(n328), .Z(n325) );
  AND U320 ( .A(n7), .B(n329), .Z(n328) );
  XNOR U321 ( .A(p_input[18]), .B(n327), .Z(n329) );
  XOR U322 ( .A(n330), .B(n331), .Z(n327) );
  AND U323 ( .A(n11), .B(n332), .Z(n331) );
  XNOR U324 ( .A(p_input[34]), .B(n330), .Z(n332) );
  XOR U325 ( .A(n333), .B(n334), .Z(n330) );
  AND U326 ( .A(n15), .B(n335), .Z(n334) );
  XNOR U327 ( .A(p_input[50]), .B(n333), .Z(n335) );
  XOR U328 ( .A(n336), .B(n337), .Z(n333) );
  AND U329 ( .A(n19), .B(n338), .Z(n337) );
  XNOR U330 ( .A(p_input[66]), .B(n336), .Z(n338) );
  XOR U331 ( .A(n339), .B(n340), .Z(n336) );
  AND U332 ( .A(n23), .B(n341), .Z(n340) );
  XNOR U333 ( .A(p_input[82]), .B(n339), .Z(n341) );
  XOR U334 ( .A(n342), .B(n343), .Z(n339) );
  AND U335 ( .A(n27), .B(n344), .Z(n343) );
  XNOR U336 ( .A(p_input[98]), .B(n342), .Z(n344) );
  XOR U337 ( .A(n345), .B(n346), .Z(n342) );
  AND U338 ( .A(n31), .B(n347), .Z(n346) );
  XNOR U339 ( .A(p_input[114]), .B(n345), .Z(n347) );
  XOR U340 ( .A(n348), .B(n349), .Z(n345) );
  AND U341 ( .A(n35), .B(n350), .Z(n349) );
  XNOR U342 ( .A(p_input[130]), .B(n348), .Z(n350) );
  XOR U343 ( .A(n351), .B(n352), .Z(n348) );
  AND U344 ( .A(n39), .B(n353), .Z(n352) );
  XNOR U345 ( .A(p_input[146]), .B(n351), .Z(n353) );
  XOR U346 ( .A(n354), .B(n355), .Z(n351) );
  AND U347 ( .A(n43), .B(n356), .Z(n355) );
  XNOR U348 ( .A(p_input[162]), .B(n354), .Z(n356) );
  XOR U349 ( .A(n357), .B(n358), .Z(n354) );
  AND U350 ( .A(n47), .B(n359), .Z(n358) );
  XNOR U351 ( .A(p_input[178]), .B(n357), .Z(n359) );
  XOR U352 ( .A(n360), .B(n361), .Z(n357) );
  AND U353 ( .A(n51), .B(n362), .Z(n361) );
  XNOR U354 ( .A(p_input[194]), .B(n360), .Z(n362) );
  XNOR U355 ( .A(n363), .B(n364), .Z(n360) );
  AND U356 ( .A(n55), .B(n365), .Z(n364) );
  XOR U357 ( .A(p_input[210]), .B(n363), .Z(n365) );
  XOR U358 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n366), .Z(n363) );
  AND U359 ( .A(n58), .B(n367), .Z(n366) );
  XOR U360 ( .A(p_input[226]), .B(\knn_comb_/min_val_out[0][2] ), .Z(n367) );
  XNOR U361 ( .A(n368), .B(n369), .Z(o[1]) );
  AND U362 ( .A(n3), .B(n370), .Z(n368) );
  XNOR U363 ( .A(p_input[1]), .B(n369), .Z(n370) );
  XOR U364 ( .A(n371), .B(n372), .Z(n369) );
  AND U365 ( .A(n7), .B(n373), .Z(n372) );
  XNOR U366 ( .A(p_input[17]), .B(n371), .Z(n373) );
  XOR U367 ( .A(n374), .B(n375), .Z(n371) );
  AND U368 ( .A(n11), .B(n376), .Z(n375) );
  XNOR U369 ( .A(p_input[33]), .B(n374), .Z(n376) );
  XOR U370 ( .A(n377), .B(n378), .Z(n374) );
  AND U371 ( .A(n15), .B(n379), .Z(n378) );
  XNOR U372 ( .A(p_input[49]), .B(n377), .Z(n379) );
  XOR U373 ( .A(n380), .B(n381), .Z(n377) );
  AND U374 ( .A(n19), .B(n382), .Z(n381) );
  XNOR U375 ( .A(p_input[65]), .B(n380), .Z(n382) );
  XOR U376 ( .A(n383), .B(n384), .Z(n380) );
  AND U377 ( .A(n23), .B(n385), .Z(n384) );
  XNOR U378 ( .A(p_input[81]), .B(n383), .Z(n385) );
  XOR U379 ( .A(n386), .B(n387), .Z(n383) );
  AND U380 ( .A(n27), .B(n388), .Z(n387) );
  XNOR U381 ( .A(p_input[97]), .B(n386), .Z(n388) );
  XOR U382 ( .A(n389), .B(n390), .Z(n386) );
  AND U383 ( .A(n31), .B(n391), .Z(n390) );
  XNOR U384 ( .A(p_input[113]), .B(n389), .Z(n391) );
  XOR U385 ( .A(n392), .B(n393), .Z(n389) );
  AND U386 ( .A(n35), .B(n394), .Z(n393) );
  XNOR U387 ( .A(p_input[129]), .B(n392), .Z(n394) );
  XOR U388 ( .A(n395), .B(n396), .Z(n392) );
  AND U389 ( .A(n39), .B(n397), .Z(n396) );
  XNOR U390 ( .A(p_input[145]), .B(n395), .Z(n397) );
  XOR U391 ( .A(n398), .B(n399), .Z(n395) );
  AND U392 ( .A(n43), .B(n400), .Z(n399) );
  XNOR U393 ( .A(p_input[161]), .B(n398), .Z(n400) );
  XOR U394 ( .A(n401), .B(n402), .Z(n398) );
  AND U395 ( .A(n47), .B(n403), .Z(n402) );
  XNOR U396 ( .A(p_input[177]), .B(n401), .Z(n403) );
  XOR U397 ( .A(n404), .B(n405), .Z(n401) );
  AND U398 ( .A(n51), .B(n406), .Z(n405) );
  XNOR U399 ( .A(p_input[193]), .B(n404), .Z(n406) );
  XNOR U400 ( .A(n407), .B(n408), .Z(n404) );
  AND U401 ( .A(n55), .B(n409), .Z(n408) );
  XOR U402 ( .A(p_input[209]), .B(n407), .Z(n409) );
  XOR U403 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n410), .Z(n407) );
  AND U404 ( .A(n58), .B(n411), .Z(n410) );
  XOR U405 ( .A(p_input[225]), .B(\knn_comb_/min_val_out[0][1] ), .Z(n411) );
  XNOR U406 ( .A(n412), .B(n413), .Z(o[15]) );
  AND U407 ( .A(n3), .B(n414), .Z(n412) );
  XNOR U408 ( .A(p_input[15]), .B(n413), .Z(n414) );
  XOR U409 ( .A(n415), .B(n416), .Z(n413) );
  AND U410 ( .A(n7), .B(n417), .Z(n416) );
  XNOR U411 ( .A(p_input[31]), .B(n415), .Z(n417) );
  XOR U412 ( .A(n418), .B(n419), .Z(n415) );
  AND U413 ( .A(n11), .B(n420), .Z(n419) );
  XNOR U414 ( .A(p_input[47]), .B(n418), .Z(n420) );
  XOR U415 ( .A(n421), .B(n422), .Z(n418) );
  AND U416 ( .A(n15), .B(n423), .Z(n422) );
  XNOR U417 ( .A(p_input[63]), .B(n421), .Z(n423) );
  XOR U418 ( .A(n424), .B(n425), .Z(n421) );
  AND U419 ( .A(n19), .B(n426), .Z(n425) );
  XNOR U420 ( .A(p_input[79]), .B(n424), .Z(n426) );
  XOR U421 ( .A(n427), .B(n428), .Z(n424) );
  AND U422 ( .A(n23), .B(n429), .Z(n428) );
  XNOR U423 ( .A(p_input[95]), .B(n427), .Z(n429) );
  XOR U424 ( .A(n430), .B(n431), .Z(n427) );
  AND U425 ( .A(n27), .B(n432), .Z(n431) );
  XNOR U426 ( .A(p_input[111]), .B(n430), .Z(n432) );
  XOR U427 ( .A(n433), .B(n434), .Z(n430) );
  AND U428 ( .A(n31), .B(n435), .Z(n434) );
  XNOR U429 ( .A(p_input[127]), .B(n433), .Z(n435) );
  XOR U430 ( .A(n436), .B(n437), .Z(n433) );
  AND U431 ( .A(n35), .B(n438), .Z(n437) );
  XNOR U432 ( .A(p_input[143]), .B(n436), .Z(n438) );
  XOR U433 ( .A(n439), .B(n440), .Z(n436) );
  AND U434 ( .A(n39), .B(n441), .Z(n440) );
  XNOR U435 ( .A(p_input[159]), .B(n439), .Z(n441) );
  XOR U436 ( .A(n442), .B(n443), .Z(n439) );
  AND U437 ( .A(n43), .B(n444), .Z(n443) );
  XNOR U438 ( .A(p_input[175]), .B(n442), .Z(n444) );
  XOR U439 ( .A(n445), .B(n446), .Z(n442) );
  AND U440 ( .A(n47), .B(n447), .Z(n446) );
  XNOR U441 ( .A(p_input[191]), .B(n445), .Z(n447) );
  XOR U442 ( .A(n448), .B(n449), .Z(n445) );
  AND U443 ( .A(n51), .B(n450), .Z(n449) );
  XNOR U444 ( .A(p_input[207]), .B(n448), .Z(n450) );
  XNOR U445 ( .A(n451), .B(n452), .Z(n448) );
  AND U446 ( .A(n55), .B(n453), .Z(n452) );
  XOR U447 ( .A(p_input[223]), .B(n451), .Z(n453) );
  XOR U448 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n454), .Z(n451) );
  AND U449 ( .A(n58), .B(n455), .Z(n454) );
  XOR U450 ( .A(p_input[239]), .B(\knn_comb_/min_val_out[0][15] ), .Z(n455) );
  XNOR U451 ( .A(n456), .B(n457), .Z(o[14]) );
  AND U452 ( .A(n3), .B(n458), .Z(n456) );
  XNOR U453 ( .A(p_input[14]), .B(n457), .Z(n458) );
  XOR U454 ( .A(n459), .B(n460), .Z(n457) );
  AND U455 ( .A(n7), .B(n461), .Z(n460) );
  XNOR U456 ( .A(p_input[30]), .B(n459), .Z(n461) );
  XOR U457 ( .A(n462), .B(n463), .Z(n459) );
  AND U458 ( .A(n11), .B(n464), .Z(n463) );
  XNOR U459 ( .A(p_input[46]), .B(n462), .Z(n464) );
  XOR U460 ( .A(n465), .B(n466), .Z(n462) );
  AND U461 ( .A(n15), .B(n467), .Z(n466) );
  XNOR U462 ( .A(p_input[62]), .B(n465), .Z(n467) );
  XOR U463 ( .A(n468), .B(n469), .Z(n465) );
  AND U464 ( .A(n19), .B(n470), .Z(n469) );
  XNOR U465 ( .A(p_input[78]), .B(n468), .Z(n470) );
  XOR U466 ( .A(n471), .B(n472), .Z(n468) );
  AND U467 ( .A(n23), .B(n473), .Z(n472) );
  XNOR U468 ( .A(p_input[94]), .B(n471), .Z(n473) );
  XOR U469 ( .A(n474), .B(n475), .Z(n471) );
  AND U470 ( .A(n27), .B(n476), .Z(n475) );
  XNOR U471 ( .A(p_input[110]), .B(n474), .Z(n476) );
  XOR U472 ( .A(n477), .B(n478), .Z(n474) );
  AND U473 ( .A(n31), .B(n479), .Z(n478) );
  XNOR U474 ( .A(p_input[126]), .B(n477), .Z(n479) );
  XOR U475 ( .A(n480), .B(n481), .Z(n477) );
  AND U476 ( .A(n35), .B(n482), .Z(n481) );
  XNOR U477 ( .A(p_input[142]), .B(n480), .Z(n482) );
  XOR U478 ( .A(n483), .B(n484), .Z(n480) );
  AND U479 ( .A(n39), .B(n485), .Z(n484) );
  XNOR U480 ( .A(p_input[158]), .B(n483), .Z(n485) );
  XOR U481 ( .A(n486), .B(n487), .Z(n483) );
  AND U482 ( .A(n43), .B(n488), .Z(n487) );
  XNOR U483 ( .A(p_input[174]), .B(n486), .Z(n488) );
  XOR U484 ( .A(n489), .B(n490), .Z(n486) );
  AND U485 ( .A(n47), .B(n491), .Z(n490) );
  XNOR U486 ( .A(p_input[190]), .B(n489), .Z(n491) );
  XOR U487 ( .A(n492), .B(n493), .Z(n489) );
  AND U488 ( .A(n51), .B(n494), .Z(n493) );
  XNOR U489 ( .A(p_input[206]), .B(n492), .Z(n494) );
  XNOR U490 ( .A(n495), .B(n496), .Z(n492) );
  AND U491 ( .A(n55), .B(n497), .Z(n496) );
  XOR U492 ( .A(p_input[222]), .B(n495), .Z(n497) );
  XOR U493 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n498), .Z(n495) );
  AND U494 ( .A(n58), .B(n499), .Z(n498) );
  XOR U495 ( .A(p_input[238]), .B(\knn_comb_/min_val_out[0][14] ), .Z(n499) );
  XNOR U496 ( .A(n500), .B(n501), .Z(o[13]) );
  AND U497 ( .A(n3), .B(n502), .Z(n500) );
  XNOR U498 ( .A(p_input[13]), .B(n501), .Z(n502) );
  XOR U499 ( .A(n503), .B(n504), .Z(n501) );
  AND U500 ( .A(n7), .B(n505), .Z(n504) );
  XNOR U501 ( .A(p_input[29]), .B(n503), .Z(n505) );
  XOR U502 ( .A(n506), .B(n507), .Z(n503) );
  AND U503 ( .A(n11), .B(n508), .Z(n507) );
  XNOR U504 ( .A(p_input[45]), .B(n506), .Z(n508) );
  XOR U505 ( .A(n509), .B(n510), .Z(n506) );
  AND U506 ( .A(n15), .B(n511), .Z(n510) );
  XNOR U507 ( .A(p_input[61]), .B(n509), .Z(n511) );
  XOR U508 ( .A(n512), .B(n513), .Z(n509) );
  AND U509 ( .A(n19), .B(n514), .Z(n513) );
  XNOR U510 ( .A(p_input[77]), .B(n512), .Z(n514) );
  XOR U511 ( .A(n515), .B(n516), .Z(n512) );
  AND U512 ( .A(n23), .B(n517), .Z(n516) );
  XNOR U513 ( .A(p_input[93]), .B(n515), .Z(n517) );
  XOR U514 ( .A(n518), .B(n519), .Z(n515) );
  AND U515 ( .A(n27), .B(n520), .Z(n519) );
  XNOR U516 ( .A(p_input[109]), .B(n518), .Z(n520) );
  XOR U517 ( .A(n521), .B(n522), .Z(n518) );
  AND U518 ( .A(n31), .B(n523), .Z(n522) );
  XNOR U519 ( .A(p_input[125]), .B(n521), .Z(n523) );
  XOR U520 ( .A(n524), .B(n525), .Z(n521) );
  AND U521 ( .A(n35), .B(n526), .Z(n525) );
  XNOR U522 ( .A(p_input[141]), .B(n524), .Z(n526) );
  XOR U523 ( .A(n527), .B(n528), .Z(n524) );
  AND U524 ( .A(n39), .B(n529), .Z(n528) );
  XNOR U525 ( .A(p_input[157]), .B(n527), .Z(n529) );
  XOR U526 ( .A(n530), .B(n531), .Z(n527) );
  AND U527 ( .A(n43), .B(n532), .Z(n531) );
  XNOR U528 ( .A(p_input[173]), .B(n530), .Z(n532) );
  XOR U529 ( .A(n533), .B(n534), .Z(n530) );
  AND U530 ( .A(n47), .B(n535), .Z(n534) );
  XNOR U531 ( .A(p_input[189]), .B(n533), .Z(n535) );
  XOR U532 ( .A(n536), .B(n537), .Z(n533) );
  AND U533 ( .A(n51), .B(n538), .Z(n537) );
  XNOR U534 ( .A(p_input[205]), .B(n536), .Z(n538) );
  XNOR U535 ( .A(n539), .B(n540), .Z(n536) );
  AND U536 ( .A(n55), .B(n541), .Z(n540) );
  XOR U537 ( .A(p_input[221]), .B(n539), .Z(n541) );
  XOR U538 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n542), .Z(n539) );
  AND U539 ( .A(n58), .B(n543), .Z(n542) );
  XOR U540 ( .A(p_input[237]), .B(\knn_comb_/min_val_out[0][13] ), .Z(n543) );
  XNOR U541 ( .A(n544), .B(n545), .Z(o[12]) );
  AND U542 ( .A(n3), .B(n546), .Z(n544) );
  XNOR U543 ( .A(p_input[12]), .B(n545), .Z(n546) );
  XOR U544 ( .A(n547), .B(n548), .Z(n545) );
  AND U545 ( .A(n7), .B(n549), .Z(n548) );
  XNOR U546 ( .A(p_input[28]), .B(n547), .Z(n549) );
  XOR U547 ( .A(n550), .B(n551), .Z(n547) );
  AND U548 ( .A(n11), .B(n552), .Z(n551) );
  XNOR U549 ( .A(p_input[44]), .B(n550), .Z(n552) );
  XOR U550 ( .A(n553), .B(n554), .Z(n550) );
  AND U551 ( .A(n15), .B(n555), .Z(n554) );
  XNOR U552 ( .A(p_input[60]), .B(n553), .Z(n555) );
  XOR U553 ( .A(n556), .B(n557), .Z(n553) );
  AND U554 ( .A(n19), .B(n558), .Z(n557) );
  XNOR U555 ( .A(p_input[76]), .B(n556), .Z(n558) );
  XOR U556 ( .A(n559), .B(n560), .Z(n556) );
  AND U557 ( .A(n23), .B(n561), .Z(n560) );
  XNOR U558 ( .A(p_input[92]), .B(n559), .Z(n561) );
  XOR U559 ( .A(n562), .B(n563), .Z(n559) );
  AND U560 ( .A(n27), .B(n564), .Z(n563) );
  XNOR U561 ( .A(p_input[108]), .B(n562), .Z(n564) );
  XOR U562 ( .A(n565), .B(n566), .Z(n562) );
  AND U563 ( .A(n31), .B(n567), .Z(n566) );
  XNOR U564 ( .A(p_input[124]), .B(n565), .Z(n567) );
  XOR U565 ( .A(n568), .B(n569), .Z(n565) );
  AND U566 ( .A(n35), .B(n570), .Z(n569) );
  XNOR U567 ( .A(p_input[140]), .B(n568), .Z(n570) );
  XOR U568 ( .A(n571), .B(n572), .Z(n568) );
  AND U569 ( .A(n39), .B(n573), .Z(n572) );
  XNOR U570 ( .A(p_input[156]), .B(n571), .Z(n573) );
  XOR U571 ( .A(n574), .B(n575), .Z(n571) );
  AND U572 ( .A(n43), .B(n576), .Z(n575) );
  XNOR U573 ( .A(p_input[172]), .B(n574), .Z(n576) );
  XOR U574 ( .A(n577), .B(n578), .Z(n574) );
  AND U575 ( .A(n47), .B(n579), .Z(n578) );
  XNOR U576 ( .A(p_input[188]), .B(n577), .Z(n579) );
  XOR U577 ( .A(n580), .B(n581), .Z(n577) );
  AND U578 ( .A(n51), .B(n582), .Z(n581) );
  XNOR U579 ( .A(p_input[204]), .B(n580), .Z(n582) );
  XNOR U580 ( .A(n583), .B(n584), .Z(n580) );
  AND U581 ( .A(n55), .B(n585), .Z(n584) );
  XOR U582 ( .A(p_input[220]), .B(n583), .Z(n585) );
  XOR U583 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n586), .Z(n583) );
  AND U584 ( .A(n58), .B(n587), .Z(n586) );
  XOR U585 ( .A(p_input[236]), .B(\knn_comb_/min_val_out[0][12] ), .Z(n587) );
  XNOR U586 ( .A(n588), .B(n589), .Z(o[11]) );
  AND U587 ( .A(n3), .B(n590), .Z(n588) );
  XNOR U588 ( .A(p_input[11]), .B(n589), .Z(n590) );
  XOR U589 ( .A(n591), .B(n592), .Z(n589) );
  AND U590 ( .A(n7), .B(n593), .Z(n592) );
  XNOR U591 ( .A(p_input[27]), .B(n591), .Z(n593) );
  XOR U592 ( .A(n594), .B(n595), .Z(n591) );
  AND U593 ( .A(n11), .B(n596), .Z(n595) );
  XNOR U594 ( .A(p_input[43]), .B(n594), .Z(n596) );
  XOR U595 ( .A(n597), .B(n598), .Z(n594) );
  AND U596 ( .A(n15), .B(n599), .Z(n598) );
  XNOR U597 ( .A(p_input[59]), .B(n597), .Z(n599) );
  XOR U598 ( .A(n600), .B(n601), .Z(n597) );
  AND U599 ( .A(n19), .B(n602), .Z(n601) );
  XNOR U600 ( .A(p_input[75]), .B(n600), .Z(n602) );
  XOR U601 ( .A(n603), .B(n604), .Z(n600) );
  AND U602 ( .A(n23), .B(n605), .Z(n604) );
  XNOR U603 ( .A(p_input[91]), .B(n603), .Z(n605) );
  XOR U604 ( .A(n606), .B(n607), .Z(n603) );
  AND U605 ( .A(n27), .B(n608), .Z(n607) );
  XNOR U606 ( .A(p_input[107]), .B(n606), .Z(n608) );
  XOR U607 ( .A(n609), .B(n610), .Z(n606) );
  AND U608 ( .A(n31), .B(n611), .Z(n610) );
  XNOR U609 ( .A(p_input[123]), .B(n609), .Z(n611) );
  XOR U610 ( .A(n612), .B(n613), .Z(n609) );
  AND U611 ( .A(n35), .B(n614), .Z(n613) );
  XNOR U612 ( .A(p_input[139]), .B(n612), .Z(n614) );
  XOR U613 ( .A(n615), .B(n616), .Z(n612) );
  AND U614 ( .A(n39), .B(n617), .Z(n616) );
  XNOR U615 ( .A(p_input[155]), .B(n615), .Z(n617) );
  XOR U616 ( .A(n618), .B(n619), .Z(n615) );
  AND U617 ( .A(n43), .B(n620), .Z(n619) );
  XNOR U618 ( .A(p_input[171]), .B(n618), .Z(n620) );
  XOR U619 ( .A(n621), .B(n622), .Z(n618) );
  AND U620 ( .A(n47), .B(n623), .Z(n622) );
  XNOR U621 ( .A(p_input[187]), .B(n621), .Z(n623) );
  XOR U622 ( .A(n624), .B(n625), .Z(n621) );
  AND U623 ( .A(n51), .B(n626), .Z(n625) );
  XNOR U624 ( .A(p_input[203]), .B(n624), .Z(n626) );
  XNOR U625 ( .A(n627), .B(n628), .Z(n624) );
  AND U626 ( .A(n55), .B(n629), .Z(n628) );
  XOR U627 ( .A(p_input[219]), .B(n627), .Z(n629) );
  XOR U628 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n630), .Z(n627) );
  AND U629 ( .A(n58), .B(n631), .Z(n630) );
  XOR U630 ( .A(p_input[235]), .B(\knn_comb_/min_val_out[0][11] ), .Z(n631) );
  XNOR U631 ( .A(n632), .B(n633), .Z(o[10]) );
  AND U632 ( .A(n3), .B(n634), .Z(n632) );
  XNOR U633 ( .A(p_input[10]), .B(n633), .Z(n634) );
  XOR U634 ( .A(n635), .B(n636), .Z(n633) );
  AND U635 ( .A(n7), .B(n637), .Z(n636) );
  XNOR U636 ( .A(p_input[26]), .B(n635), .Z(n637) );
  XOR U637 ( .A(n638), .B(n639), .Z(n635) );
  AND U638 ( .A(n11), .B(n640), .Z(n639) );
  XNOR U639 ( .A(p_input[42]), .B(n638), .Z(n640) );
  XOR U640 ( .A(n641), .B(n642), .Z(n638) );
  AND U641 ( .A(n15), .B(n643), .Z(n642) );
  XNOR U642 ( .A(p_input[58]), .B(n641), .Z(n643) );
  XOR U643 ( .A(n644), .B(n645), .Z(n641) );
  AND U644 ( .A(n19), .B(n646), .Z(n645) );
  XNOR U645 ( .A(p_input[74]), .B(n644), .Z(n646) );
  XOR U646 ( .A(n647), .B(n648), .Z(n644) );
  AND U647 ( .A(n23), .B(n649), .Z(n648) );
  XNOR U648 ( .A(p_input[90]), .B(n647), .Z(n649) );
  XOR U649 ( .A(n650), .B(n651), .Z(n647) );
  AND U650 ( .A(n27), .B(n652), .Z(n651) );
  XNOR U651 ( .A(p_input[106]), .B(n650), .Z(n652) );
  XOR U652 ( .A(n653), .B(n654), .Z(n650) );
  AND U653 ( .A(n31), .B(n655), .Z(n654) );
  XNOR U654 ( .A(p_input[122]), .B(n653), .Z(n655) );
  XOR U655 ( .A(n656), .B(n657), .Z(n653) );
  AND U656 ( .A(n35), .B(n658), .Z(n657) );
  XNOR U657 ( .A(p_input[138]), .B(n656), .Z(n658) );
  XOR U658 ( .A(n659), .B(n660), .Z(n656) );
  AND U659 ( .A(n39), .B(n661), .Z(n660) );
  XNOR U660 ( .A(p_input[154]), .B(n659), .Z(n661) );
  XOR U661 ( .A(n662), .B(n663), .Z(n659) );
  AND U662 ( .A(n43), .B(n664), .Z(n663) );
  XNOR U663 ( .A(p_input[170]), .B(n662), .Z(n664) );
  XOR U664 ( .A(n665), .B(n666), .Z(n662) );
  AND U665 ( .A(n47), .B(n667), .Z(n666) );
  XNOR U666 ( .A(p_input[186]), .B(n665), .Z(n667) );
  XOR U667 ( .A(n668), .B(n669), .Z(n665) );
  AND U668 ( .A(n51), .B(n670), .Z(n669) );
  XNOR U669 ( .A(p_input[202]), .B(n668), .Z(n670) );
  XNOR U670 ( .A(n671), .B(n672), .Z(n668) );
  AND U671 ( .A(n55), .B(n673), .Z(n672) );
  XOR U672 ( .A(p_input[218]), .B(n671), .Z(n673) );
  XOR U673 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n674), .Z(n671) );
  AND U674 ( .A(n58), .B(n675), .Z(n674) );
  XOR U675 ( .A(p_input[234]), .B(\knn_comb_/min_val_out[0][10] ), .Z(n675) );
  XNOR U676 ( .A(n676), .B(n677), .Z(o[0]) );
  AND U677 ( .A(n3), .B(n678), .Z(n676) );
  XNOR U678 ( .A(p_input[0]), .B(n677), .Z(n678) );
  XOR U679 ( .A(n679), .B(n680), .Z(n677) );
  AND U680 ( .A(n7), .B(n681), .Z(n680) );
  XNOR U681 ( .A(p_input[16]), .B(n679), .Z(n681) );
  XOR U682 ( .A(n682), .B(n683), .Z(n679) );
  AND U683 ( .A(n11), .B(n684), .Z(n683) );
  XNOR U684 ( .A(p_input[32]), .B(n682), .Z(n684) );
  XOR U685 ( .A(n685), .B(n686), .Z(n682) );
  AND U686 ( .A(n15), .B(n687), .Z(n686) );
  XNOR U687 ( .A(p_input[48]), .B(n685), .Z(n687) );
  XOR U688 ( .A(n688), .B(n689), .Z(n685) );
  AND U689 ( .A(n19), .B(n690), .Z(n689) );
  XNOR U690 ( .A(p_input[64]), .B(n688), .Z(n690) );
  XOR U691 ( .A(n691), .B(n692), .Z(n688) );
  AND U692 ( .A(n23), .B(n693), .Z(n692) );
  XNOR U693 ( .A(p_input[80]), .B(n691), .Z(n693) );
  XOR U694 ( .A(n694), .B(n695), .Z(n691) );
  AND U695 ( .A(n27), .B(n696), .Z(n695) );
  XNOR U696 ( .A(p_input[96]), .B(n694), .Z(n696) );
  XOR U697 ( .A(n697), .B(n698), .Z(n694) );
  AND U698 ( .A(n31), .B(n699), .Z(n698) );
  XNOR U699 ( .A(p_input[112]), .B(n697), .Z(n699) );
  XOR U700 ( .A(n700), .B(n701), .Z(n697) );
  AND U701 ( .A(n35), .B(n702), .Z(n701) );
  XNOR U702 ( .A(p_input[128]), .B(n700), .Z(n702) );
  XOR U703 ( .A(n703), .B(n704), .Z(n700) );
  AND U704 ( .A(n39), .B(n705), .Z(n704) );
  XNOR U705 ( .A(p_input[144]), .B(n703), .Z(n705) );
  XOR U706 ( .A(n706), .B(n707), .Z(n703) );
  AND U707 ( .A(n43), .B(n708), .Z(n707) );
  XNOR U708 ( .A(p_input[160]), .B(n706), .Z(n708) );
  XOR U709 ( .A(n709), .B(n710), .Z(n706) );
  AND U710 ( .A(n47), .B(n711), .Z(n710) );
  XNOR U711 ( .A(p_input[176]), .B(n709), .Z(n711) );
  XOR U712 ( .A(n712), .B(n713), .Z(n709) );
  AND U713 ( .A(n51), .B(n714), .Z(n713) );
  XNOR U714 ( .A(p_input[192]), .B(n712), .Z(n714) );
  XNOR U715 ( .A(n715), .B(n716), .Z(n712) );
  AND U716 ( .A(n55), .B(n717), .Z(n716) );
  XOR U717 ( .A(p_input[208]), .B(n715), .Z(n717) );
  XOR U718 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n718), .Z(n715) );
  AND U719 ( .A(n58), .B(n719), .Z(n718) );
  XOR U720 ( .A(p_input[224]), .B(\knn_comb_/min_val_out[0][0] ), .Z(n719) );
  XNOR U721 ( .A(n720), .B(n721), .Z(n3) );
  AND U722 ( .A(n722), .B(n723), .Z(n721) );
  XOR U723 ( .A(n724), .B(n720), .Z(n723) );
  AND U724 ( .A(n725), .B(n726), .Z(n724) );
  XOR U725 ( .A(n727), .B(n720), .Z(n722) );
  XNOR U726 ( .A(n728), .B(n729), .Z(n727) );
  AND U727 ( .A(n7), .B(n730), .Z(n729) );
  XOR U728 ( .A(n731), .B(n728), .Z(n730) );
  XOR U729 ( .A(n732), .B(n733), .Z(n720) );
  AND U730 ( .A(n734), .B(n735), .Z(n733) );
  XNOR U731 ( .A(n732), .B(n725), .Z(n735) );
  XNOR U732 ( .A(n736), .B(n737), .Z(n725) );
  XOR U733 ( .A(n738), .B(n726), .Z(n737) );
  AND U734 ( .A(n739), .B(n740), .Z(n726) );
  AND U735 ( .A(n741), .B(n742), .Z(n738) );
  XOR U736 ( .A(n743), .B(n736), .Z(n741) );
  XOR U737 ( .A(n744), .B(n732), .Z(n734) );
  XNOR U738 ( .A(n745), .B(n746), .Z(n744) );
  AND U739 ( .A(n7), .B(n747), .Z(n746) );
  XOR U740 ( .A(n748), .B(n745), .Z(n747) );
  XOR U741 ( .A(n749), .B(n750), .Z(n732) );
  AND U742 ( .A(n751), .B(n752), .Z(n750) );
  XNOR U743 ( .A(n749), .B(n739), .Z(n752) );
  XOR U744 ( .A(n753), .B(n742), .Z(n739) );
  XNOR U745 ( .A(n754), .B(n736), .Z(n742) );
  XOR U746 ( .A(n755), .B(n756), .Z(n736) );
  AND U747 ( .A(n757), .B(n758), .Z(n756) );
  XOR U748 ( .A(n759), .B(n755), .Z(n757) );
  XNOR U749 ( .A(n760), .B(n761), .Z(n754) );
  AND U750 ( .A(n762), .B(n763), .Z(n761) );
  XOR U751 ( .A(n760), .B(n764), .Z(n762) );
  XNOR U752 ( .A(n743), .B(n740), .Z(n753) );
  AND U753 ( .A(n765), .B(n766), .Z(n740) );
  XOR U754 ( .A(n767), .B(n768), .Z(n743) );
  AND U755 ( .A(n769), .B(n770), .Z(n768) );
  XOR U756 ( .A(n767), .B(n771), .Z(n769) );
  XOR U757 ( .A(n772), .B(n749), .Z(n751) );
  XNOR U758 ( .A(n773), .B(n774), .Z(n772) );
  AND U759 ( .A(n7), .B(n775), .Z(n774) );
  XNOR U760 ( .A(n776), .B(n773), .Z(n775) );
  XOR U761 ( .A(n777), .B(n778), .Z(n749) );
  AND U762 ( .A(n779), .B(n780), .Z(n778) );
  XNOR U763 ( .A(n777), .B(n765), .Z(n780) );
  XOR U764 ( .A(n781), .B(n758), .Z(n765) );
  XNOR U765 ( .A(n782), .B(n764), .Z(n758) );
  XNOR U766 ( .A(n783), .B(n784), .Z(n764) );
  NOR U767 ( .A(n785), .B(n786), .Z(n784) );
  XOR U768 ( .A(n783), .B(n787), .Z(n785) );
  XNOR U769 ( .A(n763), .B(n755), .Z(n782) );
  XOR U770 ( .A(n788), .B(n789), .Z(n755) );
  AND U771 ( .A(n790), .B(n791), .Z(n789) );
  XNOR U772 ( .A(n788), .B(n792), .Z(n790) );
  XNOR U773 ( .A(n793), .B(n760), .Z(n763) );
  XOR U774 ( .A(n794), .B(n795), .Z(n760) );
  AND U775 ( .A(n796), .B(n797), .Z(n795) );
  XOR U776 ( .A(n794), .B(n798), .Z(n796) );
  XNOR U777 ( .A(n799), .B(n800), .Z(n793) );
  NOR U778 ( .A(n801), .B(n802), .Z(n800) );
  XNOR U779 ( .A(n799), .B(n803), .Z(n801) );
  XNOR U780 ( .A(n759), .B(n766), .Z(n781) );
  NOR U781 ( .A(n804), .B(n805), .Z(n766) );
  XOR U782 ( .A(n771), .B(n770), .Z(n759) );
  XNOR U783 ( .A(n806), .B(n767), .Z(n770) );
  XOR U784 ( .A(n807), .B(n808), .Z(n767) );
  AND U785 ( .A(n809), .B(n810), .Z(n808) );
  XOR U786 ( .A(n807), .B(n811), .Z(n809) );
  XNOR U787 ( .A(n812), .B(n813), .Z(n806) );
  NOR U788 ( .A(n814), .B(n815), .Z(n813) );
  XNOR U789 ( .A(n812), .B(n816), .Z(n814) );
  XOR U790 ( .A(n817), .B(n818), .Z(n771) );
  NOR U791 ( .A(n819), .B(n820), .Z(n818) );
  XNOR U792 ( .A(n817), .B(n821), .Z(n819) );
  XNOR U793 ( .A(n822), .B(n823), .Z(n779) );
  XOR U794 ( .A(n777), .B(n824), .Z(n823) );
  AND U795 ( .A(n7), .B(n825), .Z(n824) );
  XOR U796 ( .A(n826), .B(n822), .Z(n825) );
  AND U797 ( .A(n827), .B(n804), .Z(n777) );
  XOR U798 ( .A(n828), .B(n805), .Z(n804) );
  XNOR U799 ( .A(p_input[0]), .B(p_input[256]), .Z(n805) );
  XOR U800 ( .A(n792), .B(n791), .Z(n828) );
  XNOR U801 ( .A(n829), .B(n798), .Z(n791) );
  XNOR U802 ( .A(n787), .B(n786), .Z(n798) );
  XNOR U803 ( .A(n830), .B(n783), .Z(n786) );
  XNOR U804 ( .A(p_input[10]), .B(p_input[266]), .Z(n783) );
  XOR U805 ( .A(p_input[11]), .B(n831), .Z(n830) );
  XOR U806 ( .A(p_input[12]), .B(p_input[268]), .Z(n787) );
  XOR U807 ( .A(n797), .B(n832), .Z(n829) );
  IV U808 ( .A(n788), .Z(n832) );
  XOR U809 ( .A(p_input[1]), .B(p_input[257]), .Z(n788) );
  XNOR U810 ( .A(n833), .B(n803), .Z(n797) );
  XNOR U811 ( .A(p_input[15]), .B(n834), .Z(n803) );
  XOR U812 ( .A(n794), .B(n802), .Z(n833) );
  XOR U813 ( .A(n835), .B(n799), .Z(n802) );
  XOR U814 ( .A(p_input[13]), .B(p_input[269]), .Z(n799) );
  XOR U815 ( .A(p_input[14]), .B(n836), .Z(n835) );
  XNOR U816 ( .A(n837), .B(p_input[9]), .Z(n794) );
  XNOR U817 ( .A(n811), .B(n810), .Z(n792) );
  XNOR U818 ( .A(n838), .B(n816), .Z(n810) );
  XOR U819 ( .A(p_input[264]), .B(p_input[8]), .Z(n816) );
  XOR U820 ( .A(n807), .B(n815), .Z(n838) );
  XOR U821 ( .A(n839), .B(n812), .Z(n815) );
  XOR U822 ( .A(p_input[262]), .B(p_input[6]), .Z(n812) );
  XNOR U823 ( .A(p_input[263]), .B(p_input[7]), .Z(n839) );
  XNOR U824 ( .A(n840), .B(p_input[2]), .Z(n807) );
  XNOR U825 ( .A(n821), .B(n820), .Z(n811) );
  XOR U826 ( .A(n841), .B(n817), .Z(n820) );
  XOR U827 ( .A(p_input[259]), .B(p_input[3]), .Z(n817) );
  XNOR U828 ( .A(p_input[260]), .B(p_input[4]), .Z(n841) );
  XOR U829 ( .A(p_input[261]), .B(p_input[5]), .Z(n821) );
  XNOR U830 ( .A(n842), .B(n843), .Z(n827) );
  AND U831 ( .A(n7), .B(n844), .Z(n843) );
  XNOR U832 ( .A(n845), .B(n846), .Z(n844) );
  XNOR U833 ( .A(n847), .B(n848), .Z(n7) );
  AND U834 ( .A(n849), .B(n850), .Z(n848) );
  XOR U835 ( .A(n731), .B(n847), .Z(n850) );
  AND U836 ( .A(n851), .B(n852), .Z(n731) );
  XNOR U837 ( .A(n728), .B(n847), .Z(n849) );
  XOR U838 ( .A(n853), .B(n854), .Z(n728) );
  AND U839 ( .A(n11), .B(n855), .Z(n854) );
  XOR U840 ( .A(n856), .B(n853), .Z(n855) );
  XOR U841 ( .A(n857), .B(n858), .Z(n847) );
  AND U842 ( .A(n859), .B(n860), .Z(n858) );
  XNOR U843 ( .A(n857), .B(n851), .Z(n860) );
  IV U844 ( .A(n748), .Z(n851) );
  XOR U845 ( .A(n861), .B(n862), .Z(n748) );
  XOR U846 ( .A(n863), .B(n852), .Z(n862) );
  AND U847 ( .A(n776), .B(n864), .Z(n852) );
  AND U848 ( .A(n865), .B(n866), .Z(n863) );
  XOR U849 ( .A(n867), .B(n861), .Z(n865) );
  XNOR U850 ( .A(n745), .B(n857), .Z(n859) );
  XOR U851 ( .A(n868), .B(n869), .Z(n745) );
  AND U852 ( .A(n11), .B(n870), .Z(n869) );
  XOR U853 ( .A(n871), .B(n868), .Z(n870) );
  XOR U854 ( .A(n872), .B(n873), .Z(n857) );
  AND U855 ( .A(n874), .B(n875), .Z(n873) );
  XNOR U856 ( .A(n872), .B(n776), .Z(n875) );
  XOR U857 ( .A(n876), .B(n866), .Z(n776) );
  XNOR U858 ( .A(n877), .B(n861), .Z(n866) );
  XOR U859 ( .A(n878), .B(n879), .Z(n861) );
  AND U860 ( .A(n880), .B(n881), .Z(n879) );
  XOR U861 ( .A(n882), .B(n878), .Z(n880) );
  XNOR U862 ( .A(n883), .B(n884), .Z(n877) );
  AND U863 ( .A(n885), .B(n886), .Z(n884) );
  XOR U864 ( .A(n883), .B(n887), .Z(n885) );
  XNOR U865 ( .A(n867), .B(n864), .Z(n876) );
  AND U866 ( .A(n888), .B(n889), .Z(n864) );
  XOR U867 ( .A(n890), .B(n891), .Z(n867) );
  AND U868 ( .A(n892), .B(n893), .Z(n891) );
  XOR U869 ( .A(n890), .B(n894), .Z(n892) );
  XNOR U870 ( .A(n773), .B(n872), .Z(n874) );
  XOR U871 ( .A(n895), .B(n896), .Z(n773) );
  AND U872 ( .A(n11), .B(n897), .Z(n896) );
  XNOR U873 ( .A(n898), .B(n895), .Z(n897) );
  XOR U874 ( .A(n899), .B(n900), .Z(n872) );
  AND U875 ( .A(n901), .B(n902), .Z(n900) );
  XNOR U876 ( .A(n899), .B(n888), .Z(n902) );
  IV U877 ( .A(n826), .Z(n888) );
  XNOR U878 ( .A(n903), .B(n881), .Z(n826) );
  XNOR U879 ( .A(n904), .B(n887), .Z(n881) );
  XOR U880 ( .A(n905), .B(n906), .Z(n887) );
  NOR U881 ( .A(n907), .B(n908), .Z(n906) );
  XNOR U882 ( .A(n905), .B(n909), .Z(n907) );
  XNOR U883 ( .A(n886), .B(n878), .Z(n904) );
  XOR U884 ( .A(n910), .B(n911), .Z(n878) );
  AND U885 ( .A(n912), .B(n913), .Z(n911) );
  XOR U886 ( .A(n910), .B(n914), .Z(n912) );
  XNOR U887 ( .A(n915), .B(n883), .Z(n886) );
  XOR U888 ( .A(n916), .B(n917), .Z(n883) );
  AND U889 ( .A(n918), .B(n919), .Z(n917) );
  XNOR U890 ( .A(n920), .B(n921), .Z(n918) );
  IV U891 ( .A(n916), .Z(n920) );
  XNOR U892 ( .A(n922), .B(n923), .Z(n915) );
  NOR U893 ( .A(n924), .B(n925), .Z(n923) );
  XOR U894 ( .A(n922), .B(n926), .Z(n924) );
  XNOR U895 ( .A(n882), .B(n889), .Z(n903) );
  NOR U896 ( .A(n845), .B(n927), .Z(n889) );
  XOR U897 ( .A(n894), .B(n893), .Z(n882) );
  XNOR U898 ( .A(n928), .B(n890), .Z(n893) );
  XOR U899 ( .A(n929), .B(n930), .Z(n890) );
  AND U900 ( .A(n931), .B(n932), .Z(n930) );
  XNOR U901 ( .A(n933), .B(n934), .Z(n931) );
  IV U902 ( .A(n929), .Z(n933) );
  XNOR U903 ( .A(n935), .B(n936), .Z(n928) );
  NOR U904 ( .A(n937), .B(n938), .Z(n936) );
  XNOR U905 ( .A(n935), .B(n939), .Z(n937) );
  XOR U906 ( .A(n940), .B(n941), .Z(n894) );
  NOR U907 ( .A(n942), .B(n943), .Z(n941) );
  XNOR U908 ( .A(n940), .B(n944), .Z(n942) );
  XNOR U909 ( .A(n822), .B(n899), .Z(n901) );
  XOR U910 ( .A(n945), .B(n946), .Z(n822) );
  AND U911 ( .A(n11), .B(n947), .Z(n946) );
  XOR U912 ( .A(n948), .B(n945), .Z(n947) );
  AND U913 ( .A(n846), .B(n845), .Z(n899) );
  XOR U914 ( .A(n949), .B(n927), .Z(n845) );
  XNOR U915 ( .A(p_input[16]), .B(p_input[256]), .Z(n927) );
  XNOR U916 ( .A(n914), .B(n913), .Z(n949) );
  XNOR U917 ( .A(n950), .B(n921), .Z(n913) );
  XNOR U918 ( .A(n909), .B(n908), .Z(n921) );
  XOR U919 ( .A(n951), .B(n905), .Z(n908) );
  XNOR U920 ( .A(n952), .B(p_input[26]), .Z(n905) );
  XNOR U921 ( .A(p_input[267]), .B(p_input[27]), .Z(n951) );
  XOR U922 ( .A(p_input[268]), .B(p_input[28]), .Z(n909) );
  XOR U923 ( .A(n919), .B(n953), .Z(n950) );
  IV U924 ( .A(n910), .Z(n953) );
  XOR U925 ( .A(p_input[17]), .B(p_input[257]), .Z(n910) );
  XOR U926 ( .A(n954), .B(n926), .Z(n919) );
  XNOR U927 ( .A(p_input[271]), .B(p_input[31]), .Z(n926) );
  XOR U928 ( .A(n916), .B(n925), .Z(n954) );
  XOR U929 ( .A(n955), .B(n922), .Z(n925) );
  XOR U930 ( .A(p_input[269]), .B(p_input[29]), .Z(n922) );
  XNOR U931 ( .A(p_input[270]), .B(p_input[30]), .Z(n955) );
  XOR U932 ( .A(p_input[25]), .B(p_input[265]), .Z(n916) );
  XOR U933 ( .A(n934), .B(n932), .Z(n914) );
  XNOR U934 ( .A(n956), .B(n939), .Z(n932) );
  XOR U935 ( .A(p_input[24]), .B(p_input[264]), .Z(n939) );
  XOR U936 ( .A(n929), .B(n938), .Z(n956) );
  XOR U937 ( .A(n957), .B(n935), .Z(n938) );
  XOR U938 ( .A(p_input[22]), .B(p_input[262]), .Z(n935) );
  XOR U939 ( .A(p_input[23]), .B(n958), .Z(n957) );
  XOR U940 ( .A(p_input[18]), .B(p_input[258]), .Z(n929) );
  XNOR U941 ( .A(n944), .B(n943), .Z(n934) );
  XOR U942 ( .A(n959), .B(n940), .Z(n943) );
  XOR U943 ( .A(p_input[19]), .B(p_input[259]), .Z(n940) );
  XOR U944 ( .A(p_input[20]), .B(n960), .Z(n959) );
  XOR U945 ( .A(p_input[21]), .B(p_input[261]), .Z(n944) );
  IV U946 ( .A(n842), .Z(n846) );
  XNOR U947 ( .A(n961), .B(n962), .Z(n842) );
  AND U948 ( .A(n11), .B(n963), .Z(n962) );
  XNOR U949 ( .A(n964), .B(n961), .Z(n963) );
  XNOR U950 ( .A(n965), .B(n966), .Z(n11) );
  AND U951 ( .A(n967), .B(n968), .Z(n966) );
  XOR U952 ( .A(n856), .B(n965), .Z(n968) );
  AND U953 ( .A(n969), .B(n970), .Z(n856) );
  XNOR U954 ( .A(n853), .B(n965), .Z(n967) );
  XOR U955 ( .A(n971), .B(n972), .Z(n853) );
  AND U956 ( .A(n15), .B(n973), .Z(n972) );
  XOR U957 ( .A(n974), .B(n971), .Z(n973) );
  XOR U958 ( .A(n975), .B(n976), .Z(n965) );
  AND U959 ( .A(n977), .B(n978), .Z(n976) );
  XNOR U960 ( .A(n975), .B(n969), .Z(n978) );
  IV U961 ( .A(n871), .Z(n969) );
  XOR U962 ( .A(n979), .B(n980), .Z(n871) );
  XOR U963 ( .A(n981), .B(n970), .Z(n980) );
  AND U964 ( .A(n898), .B(n982), .Z(n970) );
  AND U965 ( .A(n983), .B(n984), .Z(n981) );
  XOR U966 ( .A(n985), .B(n979), .Z(n983) );
  XNOR U967 ( .A(n868), .B(n975), .Z(n977) );
  XOR U968 ( .A(n986), .B(n987), .Z(n868) );
  AND U969 ( .A(n15), .B(n988), .Z(n987) );
  XOR U970 ( .A(n989), .B(n986), .Z(n988) );
  XOR U971 ( .A(n990), .B(n991), .Z(n975) );
  AND U972 ( .A(n992), .B(n993), .Z(n991) );
  XNOR U973 ( .A(n990), .B(n898), .Z(n993) );
  XOR U974 ( .A(n994), .B(n984), .Z(n898) );
  XNOR U975 ( .A(n995), .B(n979), .Z(n984) );
  XOR U976 ( .A(n996), .B(n997), .Z(n979) );
  AND U977 ( .A(n998), .B(n999), .Z(n997) );
  XOR U978 ( .A(n1000), .B(n996), .Z(n998) );
  XNOR U979 ( .A(n1001), .B(n1002), .Z(n995) );
  AND U980 ( .A(n1003), .B(n1004), .Z(n1002) );
  XOR U981 ( .A(n1001), .B(n1005), .Z(n1003) );
  XNOR U982 ( .A(n985), .B(n982), .Z(n994) );
  AND U983 ( .A(n1006), .B(n1007), .Z(n982) );
  XOR U984 ( .A(n1008), .B(n1009), .Z(n985) );
  AND U985 ( .A(n1010), .B(n1011), .Z(n1009) );
  XOR U986 ( .A(n1008), .B(n1012), .Z(n1010) );
  XNOR U987 ( .A(n895), .B(n990), .Z(n992) );
  XOR U988 ( .A(n1013), .B(n1014), .Z(n895) );
  AND U989 ( .A(n15), .B(n1015), .Z(n1014) );
  XNOR U990 ( .A(n1016), .B(n1013), .Z(n1015) );
  XOR U991 ( .A(n1017), .B(n1018), .Z(n990) );
  AND U992 ( .A(n1019), .B(n1020), .Z(n1018) );
  XNOR U993 ( .A(n1017), .B(n1006), .Z(n1020) );
  IV U994 ( .A(n948), .Z(n1006) );
  XNOR U995 ( .A(n1021), .B(n999), .Z(n948) );
  XNOR U996 ( .A(n1022), .B(n1005), .Z(n999) );
  XOR U997 ( .A(n1023), .B(n1024), .Z(n1005) );
  NOR U998 ( .A(n1025), .B(n1026), .Z(n1024) );
  XNOR U999 ( .A(n1023), .B(n1027), .Z(n1025) );
  XNOR U1000 ( .A(n1004), .B(n996), .Z(n1022) );
  XOR U1001 ( .A(n1028), .B(n1029), .Z(n996) );
  AND U1002 ( .A(n1030), .B(n1031), .Z(n1029) );
  XNOR U1003 ( .A(n1028), .B(n1032), .Z(n1030) );
  XNOR U1004 ( .A(n1033), .B(n1001), .Z(n1004) );
  XOR U1005 ( .A(n1034), .B(n1035), .Z(n1001) );
  AND U1006 ( .A(n1036), .B(n1037), .Z(n1035) );
  XOR U1007 ( .A(n1034), .B(n1038), .Z(n1036) );
  XNOR U1008 ( .A(n1039), .B(n1040), .Z(n1033) );
  NOR U1009 ( .A(n1041), .B(n1042), .Z(n1040) );
  XOR U1010 ( .A(n1039), .B(n1043), .Z(n1041) );
  XNOR U1011 ( .A(n1000), .B(n1007), .Z(n1021) );
  NOR U1012 ( .A(n964), .B(n1044), .Z(n1007) );
  XOR U1013 ( .A(n1012), .B(n1011), .Z(n1000) );
  XNOR U1014 ( .A(n1045), .B(n1008), .Z(n1011) );
  XOR U1015 ( .A(n1046), .B(n1047), .Z(n1008) );
  AND U1016 ( .A(n1048), .B(n1049), .Z(n1047) );
  XOR U1017 ( .A(n1046), .B(n1050), .Z(n1048) );
  XNOR U1018 ( .A(n1051), .B(n1052), .Z(n1045) );
  NOR U1019 ( .A(n1053), .B(n1054), .Z(n1052) );
  XNOR U1020 ( .A(n1051), .B(n1055), .Z(n1053) );
  XOR U1021 ( .A(n1056), .B(n1057), .Z(n1012) );
  NOR U1022 ( .A(n1058), .B(n1059), .Z(n1057) );
  XNOR U1023 ( .A(n1056), .B(n1060), .Z(n1058) );
  XNOR U1024 ( .A(n945), .B(n1017), .Z(n1019) );
  XOR U1025 ( .A(n1061), .B(n1062), .Z(n945) );
  AND U1026 ( .A(n15), .B(n1063), .Z(n1062) );
  XOR U1027 ( .A(n1064), .B(n1061), .Z(n1063) );
  AND U1028 ( .A(n961), .B(n964), .Z(n1017) );
  XOR U1029 ( .A(n1065), .B(n1044), .Z(n964) );
  XNOR U1030 ( .A(p_input[256]), .B(p_input[32]), .Z(n1044) );
  XOR U1031 ( .A(n1032), .B(n1031), .Z(n1065) );
  XNOR U1032 ( .A(n1066), .B(n1038), .Z(n1031) );
  XNOR U1033 ( .A(n1027), .B(n1026), .Z(n1038) );
  XOR U1034 ( .A(n1067), .B(n1023), .Z(n1026) );
  XNOR U1035 ( .A(n952), .B(p_input[42]), .Z(n1023) );
  XNOR U1036 ( .A(p_input[267]), .B(p_input[43]), .Z(n1067) );
  XOR U1037 ( .A(p_input[268]), .B(p_input[44]), .Z(n1027) );
  XNOR U1038 ( .A(n1037), .B(n1028), .Z(n1066) );
  XNOR U1039 ( .A(n1068), .B(p_input[33]), .Z(n1028) );
  XOR U1040 ( .A(n1069), .B(n1043), .Z(n1037) );
  XNOR U1041 ( .A(p_input[271]), .B(p_input[47]), .Z(n1043) );
  XOR U1042 ( .A(n1034), .B(n1042), .Z(n1069) );
  XOR U1043 ( .A(n1070), .B(n1039), .Z(n1042) );
  XOR U1044 ( .A(p_input[269]), .B(p_input[45]), .Z(n1039) );
  XNOR U1045 ( .A(p_input[270]), .B(p_input[46]), .Z(n1070) );
  XNOR U1046 ( .A(n837), .B(p_input[41]), .Z(n1034) );
  XNOR U1047 ( .A(n1050), .B(n1049), .Z(n1032) );
  XNOR U1048 ( .A(n1071), .B(n1055), .Z(n1049) );
  XOR U1049 ( .A(p_input[264]), .B(p_input[40]), .Z(n1055) );
  XOR U1050 ( .A(n1046), .B(n1054), .Z(n1071) );
  XOR U1051 ( .A(n1072), .B(n1051), .Z(n1054) );
  XOR U1052 ( .A(p_input[262]), .B(p_input[38]), .Z(n1051) );
  XNOR U1053 ( .A(p_input[263]), .B(p_input[39]), .Z(n1072) );
  XNOR U1054 ( .A(n840), .B(p_input[34]), .Z(n1046) );
  XNOR U1055 ( .A(n1060), .B(n1059), .Z(n1050) );
  XOR U1056 ( .A(n1073), .B(n1056), .Z(n1059) );
  XOR U1057 ( .A(p_input[259]), .B(p_input[35]), .Z(n1056) );
  XNOR U1058 ( .A(p_input[260]), .B(p_input[36]), .Z(n1073) );
  XOR U1059 ( .A(p_input[261]), .B(p_input[37]), .Z(n1060) );
  XOR U1060 ( .A(n1074), .B(n1075), .Z(n961) );
  AND U1061 ( .A(n15), .B(n1076), .Z(n1075) );
  XNOR U1062 ( .A(n1077), .B(n1074), .Z(n1076) );
  XNOR U1063 ( .A(n1078), .B(n1079), .Z(n15) );
  AND U1064 ( .A(n1080), .B(n1081), .Z(n1079) );
  XOR U1065 ( .A(n974), .B(n1078), .Z(n1081) );
  AND U1066 ( .A(n1082), .B(n1083), .Z(n974) );
  XNOR U1067 ( .A(n971), .B(n1078), .Z(n1080) );
  XOR U1068 ( .A(n1084), .B(n1085), .Z(n971) );
  AND U1069 ( .A(n19), .B(n1086), .Z(n1085) );
  XOR U1070 ( .A(n1087), .B(n1084), .Z(n1086) );
  XOR U1071 ( .A(n1088), .B(n1089), .Z(n1078) );
  AND U1072 ( .A(n1090), .B(n1091), .Z(n1089) );
  XNOR U1073 ( .A(n1088), .B(n1082), .Z(n1091) );
  IV U1074 ( .A(n989), .Z(n1082) );
  XOR U1075 ( .A(n1092), .B(n1093), .Z(n989) );
  XOR U1076 ( .A(n1094), .B(n1083), .Z(n1093) );
  AND U1077 ( .A(n1016), .B(n1095), .Z(n1083) );
  AND U1078 ( .A(n1096), .B(n1097), .Z(n1094) );
  XOR U1079 ( .A(n1098), .B(n1092), .Z(n1096) );
  XNOR U1080 ( .A(n986), .B(n1088), .Z(n1090) );
  XOR U1081 ( .A(n1099), .B(n1100), .Z(n986) );
  AND U1082 ( .A(n19), .B(n1101), .Z(n1100) );
  XOR U1083 ( .A(n1102), .B(n1099), .Z(n1101) );
  XOR U1084 ( .A(n1103), .B(n1104), .Z(n1088) );
  AND U1085 ( .A(n1105), .B(n1106), .Z(n1104) );
  XNOR U1086 ( .A(n1103), .B(n1016), .Z(n1106) );
  XOR U1087 ( .A(n1107), .B(n1097), .Z(n1016) );
  XNOR U1088 ( .A(n1108), .B(n1092), .Z(n1097) );
  XOR U1089 ( .A(n1109), .B(n1110), .Z(n1092) );
  AND U1090 ( .A(n1111), .B(n1112), .Z(n1110) );
  XOR U1091 ( .A(n1113), .B(n1109), .Z(n1111) );
  XNOR U1092 ( .A(n1114), .B(n1115), .Z(n1108) );
  AND U1093 ( .A(n1116), .B(n1117), .Z(n1115) );
  XOR U1094 ( .A(n1114), .B(n1118), .Z(n1116) );
  XNOR U1095 ( .A(n1098), .B(n1095), .Z(n1107) );
  AND U1096 ( .A(n1119), .B(n1120), .Z(n1095) );
  XOR U1097 ( .A(n1121), .B(n1122), .Z(n1098) );
  AND U1098 ( .A(n1123), .B(n1124), .Z(n1122) );
  XOR U1099 ( .A(n1121), .B(n1125), .Z(n1123) );
  XNOR U1100 ( .A(n1013), .B(n1103), .Z(n1105) );
  XOR U1101 ( .A(n1126), .B(n1127), .Z(n1013) );
  AND U1102 ( .A(n19), .B(n1128), .Z(n1127) );
  XNOR U1103 ( .A(n1129), .B(n1126), .Z(n1128) );
  XOR U1104 ( .A(n1130), .B(n1131), .Z(n1103) );
  AND U1105 ( .A(n1132), .B(n1133), .Z(n1131) );
  XNOR U1106 ( .A(n1130), .B(n1119), .Z(n1133) );
  IV U1107 ( .A(n1064), .Z(n1119) );
  XNOR U1108 ( .A(n1134), .B(n1112), .Z(n1064) );
  XNOR U1109 ( .A(n1135), .B(n1118), .Z(n1112) );
  XOR U1110 ( .A(n1136), .B(n1137), .Z(n1118) );
  NOR U1111 ( .A(n1138), .B(n1139), .Z(n1137) );
  XNOR U1112 ( .A(n1136), .B(n1140), .Z(n1138) );
  XNOR U1113 ( .A(n1117), .B(n1109), .Z(n1135) );
  XOR U1114 ( .A(n1141), .B(n1142), .Z(n1109) );
  AND U1115 ( .A(n1143), .B(n1144), .Z(n1142) );
  XNOR U1116 ( .A(n1141), .B(n1145), .Z(n1143) );
  XNOR U1117 ( .A(n1146), .B(n1114), .Z(n1117) );
  XOR U1118 ( .A(n1147), .B(n1148), .Z(n1114) );
  AND U1119 ( .A(n1149), .B(n1150), .Z(n1148) );
  XOR U1120 ( .A(n1147), .B(n1151), .Z(n1149) );
  XNOR U1121 ( .A(n1152), .B(n1153), .Z(n1146) );
  NOR U1122 ( .A(n1154), .B(n1155), .Z(n1153) );
  XOR U1123 ( .A(n1152), .B(n1156), .Z(n1154) );
  XNOR U1124 ( .A(n1113), .B(n1120), .Z(n1134) );
  NOR U1125 ( .A(n1077), .B(n1157), .Z(n1120) );
  XOR U1126 ( .A(n1125), .B(n1124), .Z(n1113) );
  XNOR U1127 ( .A(n1158), .B(n1121), .Z(n1124) );
  XOR U1128 ( .A(n1159), .B(n1160), .Z(n1121) );
  AND U1129 ( .A(n1161), .B(n1162), .Z(n1160) );
  XOR U1130 ( .A(n1159), .B(n1163), .Z(n1161) );
  XNOR U1131 ( .A(n1164), .B(n1165), .Z(n1158) );
  NOR U1132 ( .A(n1166), .B(n1167), .Z(n1165) );
  XNOR U1133 ( .A(n1164), .B(n1168), .Z(n1166) );
  XOR U1134 ( .A(n1169), .B(n1170), .Z(n1125) );
  NOR U1135 ( .A(n1171), .B(n1172), .Z(n1170) );
  XNOR U1136 ( .A(n1169), .B(n1173), .Z(n1171) );
  XNOR U1137 ( .A(n1061), .B(n1130), .Z(n1132) );
  XOR U1138 ( .A(n1174), .B(n1175), .Z(n1061) );
  AND U1139 ( .A(n19), .B(n1176), .Z(n1175) );
  XOR U1140 ( .A(n1177), .B(n1174), .Z(n1176) );
  AND U1141 ( .A(n1074), .B(n1077), .Z(n1130) );
  XOR U1142 ( .A(n1178), .B(n1157), .Z(n1077) );
  XNOR U1143 ( .A(p_input[256]), .B(p_input[48]), .Z(n1157) );
  XOR U1144 ( .A(n1145), .B(n1144), .Z(n1178) );
  XNOR U1145 ( .A(n1179), .B(n1151), .Z(n1144) );
  XNOR U1146 ( .A(n1140), .B(n1139), .Z(n1151) );
  XOR U1147 ( .A(n1180), .B(n1136), .Z(n1139) );
  XNOR U1148 ( .A(n952), .B(p_input[58]), .Z(n1136) );
  XNOR U1149 ( .A(p_input[267]), .B(p_input[59]), .Z(n1180) );
  XOR U1150 ( .A(p_input[268]), .B(p_input[60]), .Z(n1140) );
  XNOR U1151 ( .A(n1150), .B(n1141), .Z(n1179) );
  XNOR U1152 ( .A(n1068), .B(p_input[49]), .Z(n1141) );
  XOR U1153 ( .A(n1181), .B(n1156), .Z(n1150) );
  XNOR U1154 ( .A(p_input[271]), .B(p_input[63]), .Z(n1156) );
  XOR U1155 ( .A(n1147), .B(n1155), .Z(n1181) );
  XOR U1156 ( .A(n1182), .B(n1152), .Z(n1155) );
  XOR U1157 ( .A(p_input[269]), .B(p_input[61]), .Z(n1152) );
  XNOR U1158 ( .A(p_input[270]), .B(p_input[62]), .Z(n1182) );
  XNOR U1159 ( .A(n837), .B(p_input[57]), .Z(n1147) );
  XNOR U1160 ( .A(n1163), .B(n1162), .Z(n1145) );
  XNOR U1161 ( .A(n1183), .B(n1168), .Z(n1162) );
  XOR U1162 ( .A(p_input[264]), .B(p_input[56]), .Z(n1168) );
  XOR U1163 ( .A(n1159), .B(n1167), .Z(n1183) );
  XOR U1164 ( .A(n1184), .B(n1164), .Z(n1167) );
  XOR U1165 ( .A(p_input[262]), .B(p_input[54]), .Z(n1164) );
  XNOR U1166 ( .A(p_input[263]), .B(p_input[55]), .Z(n1184) );
  XNOR U1167 ( .A(n840), .B(p_input[50]), .Z(n1159) );
  XNOR U1168 ( .A(n1173), .B(n1172), .Z(n1163) );
  XOR U1169 ( .A(n1185), .B(n1169), .Z(n1172) );
  XOR U1170 ( .A(p_input[259]), .B(p_input[51]), .Z(n1169) );
  XNOR U1171 ( .A(p_input[260]), .B(p_input[52]), .Z(n1185) );
  XOR U1172 ( .A(p_input[261]), .B(p_input[53]), .Z(n1173) );
  XOR U1173 ( .A(n1186), .B(n1187), .Z(n1074) );
  AND U1174 ( .A(n19), .B(n1188), .Z(n1187) );
  XNOR U1175 ( .A(n1189), .B(n1186), .Z(n1188) );
  XNOR U1176 ( .A(n1190), .B(n1191), .Z(n19) );
  AND U1177 ( .A(n1192), .B(n1193), .Z(n1191) );
  XOR U1178 ( .A(n1087), .B(n1190), .Z(n1193) );
  AND U1179 ( .A(n1194), .B(n1195), .Z(n1087) );
  XNOR U1180 ( .A(n1084), .B(n1190), .Z(n1192) );
  XOR U1181 ( .A(n1196), .B(n1197), .Z(n1084) );
  AND U1182 ( .A(n1198), .B(n23), .Z(n1197) );
  AND U1183 ( .A(n1196), .B(n1199), .Z(n1198) );
  XOR U1184 ( .A(n1200), .B(n1201), .Z(n1190) );
  AND U1185 ( .A(n1202), .B(n1203), .Z(n1201) );
  XNOR U1186 ( .A(n1200), .B(n1194), .Z(n1203) );
  IV U1187 ( .A(n1102), .Z(n1194) );
  XOR U1188 ( .A(n1204), .B(n1205), .Z(n1102) );
  XOR U1189 ( .A(n1206), .B(n1195), .Z(n1205) );
  AND U1190 ( .A(n1129), .B(n1207), .Z(n1195) );
  AND U1191 ( .A(n1208), .B(n1209), .Z(n1206) );
  XOR U1192 ( .A(n1210), .B(n1204), .Z(n1208) );
  XNOR U1193 ( .A(n1099), .B(n1200), .Z(n1202) );
  XOR U1194 ( .A(n1211), .B(n1212), .Z(n1099) );
  AND U1195 ( .A(n23), .B(n1213), .Z(n1212) );
  XOR U1196 ( .A(n1214), .B(n1211), .Z(n1213) );
  XOR U1197 ( .A(n1215), .B(n1216), .Z(n1200) );
  AND U1198 ( .A(n1217), .B(n1218), .Z(n1216) );
  XNOR U1199 ( .A(n1215), .B(n1129), .Z(n1218) );
  XOR U1200 ( .A(n1219), .B(n1209), .Z(n1129) );
  XNOR U1201 ( .A(n1220), .B(n1204), .Z(n1209) );
  XOR U1202 ( .A(n1221), .B(n1222), .Z(n1204) );
  AND U1203 ( .A(n1223), .B(n1224), .Z(n1222) );
  XOR U1204 ( .A(n1225), .B(n1221), .Z(n1223) );
  XNOR U1205 ( .A(n1226), .B(n1227), .Z(n1220) );
  AND U1206 ( .A(n1228), .B(n1229), .Z(n1227) );
  XOR U1207 ( .A(n1226), .B(n1230), .Z(n1228) );
  XNOR U1208 ( .A(n1210), .B(n1207), .Z(n1219) );
  AND U1209 ( .A(n1231), .B(n1232), .Z(n1207) );
  XOR U1210 ( .A(n1233), .B(n1234), .Z(n1210) );
  AND U1211 ( .A(n1235), .B(n1236), .Z(n1234) );
  XOR U1212 ( .A(n1233), .B(n1237), .Z(n1235) );
  XNOR U1213 ( .A(n1126), .B(n1215), .Z(n1217) );
  XOR U1214 ( .A(n1238), .B(n1239), .Z(n1126) );
  AND U1215 ( .A(n23), .B(n1240), .Z(n1239) );
  XNOR U1216 ( .A(n1241), .B(n1238), .Z(n1240) );
  XOR U1217 ( .A(n1242), .B(n1243), .Z(n1215) );
  AND U1218 ( .A(n1244), .B(n1245), .Z(n1243) );
  XNOR U1219 ( .A(n1242), .B(n1231), .Z(n1245) );
  IV U1220 ( .A(n1177), .Z(n1231) );
  XNOR U1221 ( .A(n1246), .B(n1224), .Z(n1177) );
  XNOR U1222 ( .A(n1247), .B(n1230), .Z(n1224) );
  XOR U1223 ( .A(n1248), .B(n1249), .Z(n1230) );
  NOR U1224 ( .A(n1250), .B(n1251), .Z(n1249) );
  XNOR U1225 ( .A(n1248), .B(n1252), .Z(n1250) );
  XNOR U1226 ( .A(n1229), .B(n1221), .Z(n1247) );
  XOR U1227 ( .A(n1253), .B(n1254), .Z(n1221) );
  AND U1228 ( .A(n1255), .B(n1256), .Z(n1254) );
  XNOR U1229 ( .A(n1253), .B(n1257), .Z(n1255) );
  XNOR U1230 ( .A(n1258), .B(n1226), .Z(n1229) );
  XOR U1231 ( .A(n1259), .B(n1260), .Z(n1226) );
  AND U1232 ( .A(n1261), .B(n1262), .Z(n1260) );
  XOR U1233 ( .A(n1259), .B(n1263), .Z(n1261) );
  XNOR U1234 ( .A(n1264), .B(n1265), .Z(n1258) );
  NOR U1235 ( .A(n1266), .B(n1267), .Z(n1265) );
  XOR U1236 ( .A(n1264), .B(n1268), .Z(n1266) );
  XNOR U1237 ( .A(n1225), .B(n1232), .Z(n1246) );
  NOR U1238 ( .A(n1189), .B(n1269), .Z(n1232) );
  XOR U1239 ( .A(n1237), .B(n1236), .Z(n1225) );
  XNOR U1240 ( .A(n1270), .B(n1233), .Z(n1236) );
  XOR U1241 ( .A(n1271), .B(n1272), .Z(n1233) );
  AND U1242 ( .A(n1273), .B(n1274), .Z(n1272) );
  XOR U1243 ( .A(n1271), .B(n1275), .Z(n1273) );
  XNOR U1244 ( .A(n1276), .B(n1277), .Z(n1270) );
  NOR U1245 ( .A(n1278), .B(n1279), .Z(n1277) );
  XNOR U1246 ( .A(n1276), .B(n1280), .Z(n1278) );
  XOR U1247 ( .A(n1281), .B(n1282), .Z(n1237) );
  NOR U1248 ( .A(n1283), .B(n1284), .Z(n1282) );
  XNOR U1249 ( .A(n1281), .B(n1285), .Z(n1283) );
  XNOR U1250 ( .A(n1174), .B(n1242), .Z(n1244) );
  XOR U1251 ( .A(n1286), .B(n1287), .Z(n1174) );
  AND U1252 ( .A(n23), .B(n1288), .Z(n1287) );
  XOR U1253 ( .A(n1289), .B(n1286), .Z(n1288) );
  AND U1254 ( .A(n1186), .B(n1189), .Z(n1242) );
  XOR U1255 ( .A(n1290), .B(n1269), .Z(n1189) );
  XNOR U1256 ( .A(p_input[256]), .B(p_input[64]), .Z(n1269) );
  XOR U1257 ( .A(n1257), .B(n1256), .Z(n1290) );
  XNOR U1258 ( .A(n1291), .B(n1263), .Z(n1256) );
  XNOR U1259 ( .A(n1252), .B(n1251), .Z(n1263) );
  XOR U1260 ( .A(n1292), .B(n1248), .Z(n1251) );
  XNOR U1261 ( .A(n952), .B(p_input[74]), .Z(n1248) );
  XNOR U1262 ( .A(p_input[267]), .B(p_input[75]), .Z(n1292) );
  XOR U1263 ( .A(p_input[268]), .B(p_input[76]), .Z(n1252) );
  XNOR U1264 ( .A(n1262), .B(n1253), .Z(n1291) );
  XNOR U1265 ( .A(n1068), .B(p_input[65]), .Z(n1253) );
  XOR U1266 ( .A(n1293), .B(n1268), .Z(n1262) );
  XNOR U1267 ( .A(p_input[271]), .B(p_input[79]), .Z(n1268) );
  XOR U1268 ( .A(n1259), .B(n1267), .Z(n1293) );
  XOR U1269 ( .A(n1294), .B(n1264), .Z(n1267) );
  XOR U1270 ( .A(p_input[269]), .B(p_input[77]), .Z(n1264) );
  XNOR U1271 ( .A(p_input[270]), .B(p_input[78]), .Z(n1294) );
  XNOR U1272 ( .A(n837), .B(p_input[73]), .Z(n1259) );
  XNOR U1273 ( .A(n1275), .B(n1274), .Z(n1257) );
  XNOR U1274 ( .A(n1295), .B(n1280), .Z(n1274) );
  XOR U1275 ( .A(p_input[264]), .B(p_input[72]), .Z(n1280) );
  XOR U1276 ( .A(n1271), .B(n1279), .Z(n1295) );
  XOR U1277 ( .A(n1296), .B(n1276), .Z(n1279) );
  XOR U1278 ( .A(p_input[262]), .B(p_input[70]), .Z(n1276) );
  XNOR U1279 ( .A(p_input[263]), .B(p_input[71]), .Z(n1296) );
  XNOR U1280 ( .A(n840), .B(p_input[66]), .Z(n1271) );
  XNOR U1281 ( .A(n1285), .B(n1284), .Z(n1275) );
  XOR U1282 ( .A(n1297), .B(n1281), .Z(n1284) );
  XOR U1283 ( .A(p_input[259]), .B(p_input[67]), .Z(n1281) );
  XNOR U1284 ( .A(p_input[260]), .B(p_input[68]), .Z(n1297) );
  XOR U1285 ( .A(p_input[261]), .B(p_input[69]), .Z(n1285) );
  XOR U1286 ( .A(n1298), .B(n1299), .Z(n1186) );
  AND U1287 ( .A(n23), .B(n1300), .Z(n1299) );
  XNOR U1288 ( .A(n1301), .B(n1298), .Z(n1300) );
  XNOR U1289 ( .A(n1302), .B(n1303), .Z(n23) );
  AND U1290 ( .A(n1304), .B(n1305), .Z(n1303) );
  XNOR U1291 ( .A(n1199), .B(n1302), .Z(n1305) );
  IV U1292 ( .A(n1306), .Z(n1199) );
  AND U1293 ( .A(n1307), .B(n1308), .Z(n1306) );
  XNOR U1294 ( .A(n1302), .B(n1196), .Z(n1304) );
  AND U1295 ( .A(n1309), .B(n1310), .Z(n1196) );
  XOR U1296 ( .A(n1311), .B(n1312), .Z(n1302) );
  AND U1297 ( .A(n1313), .B(n1314), .Z(n1312) );
  XNOR U1298 ( .A(n1311), .B(n1307), .Z(n1314) );
  IV U1299 ( .A(n1214), .Z(n1307) );
  XOR U1300 ( .A(n1315), .B(n1316), .Z(n1214) );
  XOR U1301 ( .A(n1317), .B(n1308), .Z(n1316) );
  AND U1302 ( .A(n1241), .B(n1318), .Z(n1308) );
  AND U1303 ( .A(n1319), .B(n1320), .Z(n1317) );
  XOR U1304 ( .A(n1321), .B(n1315), .Z(n1319) );
  XNOR U1305 ( .A(n1211), .B(n1311), .Z(n1313) );
  XOR U1306 ( .A(n1322), .B(n1323), .Z(n1211) );
  AND U1307 ( .A(n27), .B(n1324), .Z(n1323) );
  XOR U1308 ( .A(n1325), .B(n1322), .Z(n1324) );
  XOR U1309 ( .A(n1326), .B(n1327), .Z(n1311) );
  AND U1310 ( .A(n1328), .B(n1329), .Z(n1327) );
  XNOR U1311 ( .A(n1326), .B(n1241), .Z(n1329) );
  XOR U1312 ( .A(n1330), .B(n1320), .Z(n1241) );
  XNOR U1313 ( .A(n1331), .B(n1315), .Z(n1320) );
  XOR U1314 ( .A(n1332), .B(n1333), .Z(n1315) );
  AND U1315 ( .A(n1334), .B(n1335), .Z(n1333) );
  XOR U1316 ( .A(n1336), .B(n1332), .Z(n1334) );
  XNOR U1317 ( .A(n1337), .B(n1338), .Z(n1331) );
  AND U1318 ( .A(n1339), .B(n1340), .Z(n1338) );
  XOR U1319 ( .A(n1337), .B(n1341), .Z(n1339) );
  XNOR U1320 ( .A(n1321), .B(n1318), .Z(n1330) );
  AND U1321 ( .A(n1342), .B(n1343), .Z(n1318) );
  XOR U1322 ( .A(n1344), .B(n1345), .Z(n1321) );
  AND U1323 ( .A(n1346), .B(n1347), .Z(n1345) );
  XOR U1324 ( .A(n1344), .B(n1348), .Z(n1346) );
  XNOR U1325 ( .A(n1238), .B(n1326), .Z(n1328) );
  XOR U1326 ( .A(n1349), .B(n1350), .Z(n1238) );
  AND U1327 ( .A(n27), .B(n1351), .Z(n1350) );
  XNOR U1328 ( .A(n1352), .B(n1349), .Z(n1351) );
  XOR U1329 ( .A(n1353), .B(n1354), .Z(n1326) );
  AND U1330 ( .A(n1355), .B(n1356), .Z(n1354) );
  XNOR U1331 ( .A(n1353), .B(n1342), .Z(n1356) );
  IV U1332 ( .A(n1289), .Z(n1342) );
  XNOR U1333 ( .A(n1357), .B(n1335), .Z(n1289) );
  XNOR U1334 ( .A(n1358), .B(n1341), .Z(n1335) );
  XOR U1335 ( .A(n1359), .B(n1360), .Z(n1341) );
  NOR U1336 ( .A(n1361), .B(n1362), .Z(n1360) );
  XNOR U1337 ( .A(n1359), .B(n1363), .Z(n1361) );
  XNOR U1338 ( .A(n1340), .B(n1332), .Z(n1358) );
  XOR U1339 ( .A(n1364), .B(n1365), .Z(n1332) );
  AND U1340 ( .A(n1366), .B(n1367), .Z(n1365) );
  XNOR U1341 ( .A(n1364), .B(n1368), .Z(n1366) );
  XNOR U1342 ( .A(n1369), .B(n1337), .Z(n1340) );
  XOR U1343 ( .A(n1370), .B(n1371), .Z(n1337) );
  AND U1344 ( .A(n1372), .B(n1373), .Z(n1371) );
  XOR U1345 ( .A(n1370), .B(n1374), .Z(n1372) );
  XNOR U1346 ( .A(n1375), .B(n1376), .Z(n1369) );
  NOR U1347 ( .A(n1377), .B(n1378), .Z(n1376) );
  XOR U1348 ( .A(n1375), .B(n1379), .Z(n1377) );
  XNOR U1349 ( .A(n1336), .B(n1343), .Z(n1357) );
  NOR U1350 ( .A(n1301), .B(n1380), .Z(n1343) );
  XOR U1351 ( .A(n1348), .B(n1347), .Z(n1336) );
  XNOR U1352 ( .A(n1381), .B(n1344), .Z(n1347) );
  XOR U1353 ( .A(n1382), .B(n1383), .Z(n1344) );
  AND U1354 ( .A(n1384), .B(n1385), .Z(n1383) );
  XOR U1355 ( .A(n1382), .B(n1386), .Z(n1384) );
  XNOR U1356 ( .A(n1387), .B(n1388), .Z(n1381) );
  NOR U1357 ( .A(n1389), .B(n1390), .Z(n1388) );
  XNOR U1358 ( .A(n1387), .B(n1391), .Z(n1389) );
  XOR U1359 ( .A(n1392), .B(n1393), .Z(n1348) );
  NOR U1360 ( .A(n1394), .B(n1395), .Z(n1393) );
  XNOR U1361 ( .A(n1392), .B(n1396), .Z(n1394) );
  XNOR U1362 ( .A(n1286), .B(n1353), .Z(n1355) );
  XOR U1363 ( .A(n1397), .B(n1398), .Z(n1286) );
  AND U1364 ( .A(n27), .B(n1399), .Z(n1398) );
  XOR U1365 ( .A(n1400), .B(n1397), .Z(n1399) );
  AND U1366 ( .A(n1298), .B(n1301), .Z(n1353) );
  XOR U1367 ( .A(n1401), .B(n1380), .Z(n1301) );
  XNOR U1368 ( .A(p_input[256]), .B(p_input[80]), .Z(n1380) );
  XOR U1369 ( .A(n1368), .B(n1367), .Z(n1401) );
  XNOR U1370 ( .A(n1402), .B(n1374), .Z(n1367) );
  XNOR U1371 ( .A(n1363), .B(n1362), .Z(n1374) );
  XOR U1372 ( .A(n1403), .B(n1359), .Z(n1362) );
  XNOR U1373 ( .A(n952), .B(p_input[90]), .Z(n1359) );
  XNOR U1374 ( .A(p_input[267]), .B(p_input[91]), .Z(n1403) );
  XOR U1375 ( .A(p_input[268]), .B(p_input[92]), .Z(n1363) );
  XNOR U1376 ( .A(n1373), .B(n1364), .Z(n1402) );
  XNOR U1377 ( .A(n1068), .B(p_input[81]), .Z(n1364) );
  XOR U1378 ( .A(n1404), .B(n1379), .Z(n1373) );
  XNOR U1379 ( .A(p_input[271]), .B(p_input[95]), .Z(n1379) );
  XOR U1380 ( .A(n1370), .B(n1378), .Z(n1404) );
  XOR U1381 ( .A(n1405), .B(n1375), .Z(n1378) );
  XOR U1382 ( .A(p_input[269]), .B(p_input[93]), .Z(n1375) );
  XNOR U1383 ( .A(p_input[270]), .B(p_input[94]), .Z(n1405) );
  XNOR U1384 ( .A(n837), .B(p_input[89]), .Z(n1370) );
  XNOR U1385 ( .A(n1386), .B(n1385), .Z(n1368) );
  XNOR U1386 ( .A(n1406), .B(n1391), .Z(n1385) );
  XOR U1387 ( .A(p_input[264]), .B(p_input[88]), .Z(n1391) );
  XOR U1388 ( .A(n1382), .B(n1390), .Z(n1406) );
  XOR U1389 ( .A(n1407), .B(n1387), .Z(n1390) );
  XOR U1390 ( .A(p_input[262]), .B(p_input[86]), .Z(n1387) );
  XNOR U1391 ( .A(p_input[263]), .B(p_input[87]), .Z(n1407) );
  XNOR U1392 ( .A(n840), .B(p_input[82]), .Z(n1382) );
  XNOR U1393 ( .A(n1396), .B(n1395), .Z(n1386) );
  XOR U1394 ( .A(n1408), .B(n1392), .Z(n1395) );
  XOR U1395 ( .A(p_input[259]), .B(p_input[83]), .Z(n1392) );
  XNOR U1396 ( .A(p_input[260]), .B(p_input[84]), .Z(n1408) );
  XOR U1397 ( .A(p_input[261]), .B(p_input[85]), .Z(n1396) );
  XOR U1398 ( .A(n1409), .B(n1410), .Z(n1298) );
  AND U1399 ( .A(n27), .B(n1411), .Z(n1410) );
  XNOR U1400 ( .A(n1412), .B(n1409), .Z(n1411) );
  XNOR U1401 ( .A(n1413), .B(n1414), .Z(n27) );
  NOR U1402 ( .A(n1415), .B(n1416), .Z(n1414) );
  XOR U1403 ( .A(n1310), .B(n1413), .Z(n1416) );
  AND U1404 ( .A(n1417), .B(n1418), .Z(n1310) );
  NOR U1405 ( .A(n1413), .B(n1309), .Z(n1415) );
  AND U1406 ( .A(n1419), .B(n1420), .Z(n1309) );
  XOR U1407 ( .A(n1421), .B(n1422), .Z(n1413) );
  AND U1408 ( .A(n1423), .B(n1424), .Z(n1422) );
  XNOR U1409 ( .A(n1421), .B(n1419), .Z(n1424) );
  IV U1410 ( .A(n1325), .Z(n1419) );
  XOR U1411 ( .A(n1425), .B(n1426), .Z(n1325) );
  XOR U1412 ( .A(n1427), .B(n1420), .Z(n1426) );
  AND U1413 ( .A(n1352), .B(n1428), .Z(n1420) );
  AND U1414 ( .A(n1429), .B(n1430), .Z(n1427) );
  XOR U1415 ( .A(n1431), .B(n1425), .Z(n1429) );
  XNOR U1416 ( .A(n1322), .B(n1421), .Z(n1423) );
  XOR U1417 ( .A(n1432), .B(n1433), .Z(n1322) );
  AND U1418 ( .A(n31), .B(n1434), .Z(n1433) );
  XOR U1419 ( .A(n1435), .B(n1432), .Z(n1434) );
  XOR U1420 ( .A(n1436), .B(n1437), .Z(n1421) );
  AND U1421 ( .A(n1438), .B(n1439), .Z(n1437) );
  XNOR U1422 ( .A(n1436), .B(n1352), .Z(n1439) );
  XOR U1423 ( .A(n1440), .B(n1430), .Z(n1352) );
  XNOR U1424 ( .A(n1441), .B(n1425), .Z(n1430) );
  XOR U1425 ( .A(n1442), .B(n1443), .Z(n1425) );
  AND U1426 ( .A(n1444), .B(n1445), .Z(n1443) );
  XOR U1427 ( .A(n1446), .B(n1442), .Z(n1444) );
  XNOR U1428 ( .A(n1447), .B(n1448), .Z(n1441) );
  AND U1429 ( .A(n1449), .B(n1450), .Z(n1448) );
  XOR U1430 ( .A(n1447), .B(n1451), .Z(n1449) );
  XNOR U1431 ( .A(n1431), .B(n1428), .Z(n1440) );
  AND U1432 ( .A(n1452), .B(n1453), .Z(n1428) );
  XOR U1433 ( .A(n1454), .B(n1455), .Z(n1431) );
  AND U1434 ( .A(n1456), .B(n1457), .Z(n1455) );
  XOR U1435 ( .A(n1454), .B(n1458), .Z(n1456) );
  XNOR U1436 ( .A(n1349), .B(n1436), .Z(n1438) );
  XOR U1437 ( .A(n1459), .B(n1460), .Z(n1349) );
  AND U1438 ( .A(n31), .B(n1461), .Z(n1460) );
  XNOR U1439 ( .A(n1462), .B(n1459), .Z(n1461) );
  XOR U1440 ( .A(n1463), .B(n1464), .Z(n1436) );
  AND U1441 ( .A(n1465), .B(n1466), .Z(n1464) );
  XNOR U1442 ( .A(n1463), .B(n1452), .Z(n1466) );
  IV U1443 ( .A(n1400), .Z(n1452) );
  XNOR U1444 ( .A(n1467), .B(n1445), .Z(n1400) );
  XNOR U1445 ( .A(n1468), .B(n1451), .Z(n1445) );
  XNOR U1446 ( .A(n1469), .B(n1470), .Z(n1451) );
  NOR U1447 ( .A(n1471), .B(n1472), .Z(n1470) );
  XOR U1448 ( .A(n1469), .B(n1473), .Z(n1471) );
  XNOR U1449 ( .A(n1450), .B(n1442), .Z(n1468) );
  XOR U1450 ( .A(n1474), .B(n1475), .Z(n1442) );
  AND U1451 ( .A(n1476), .B(n1477), .Z(n1475) );
  XOR U1452 ( .A(n1474), .B(n1478), .Z(n1476) );
  XNOR U1453 ( .A(n1479), .B(n1447), .Z(n1450) );
  XOR U1454 ( .A(n1480), .B(n1481), .Z(n1447) );
  AND U1455 ( .A(n1482), .B(n1483), .Z(n1481) );
  XNOR U1456 ( .A(n1484), .B(n1485), .Z(n1482) );
  IV U1457 ( .A(n1480), .Z(n1484) );
  XNOR U1458 ( .A(n1486), .B(n1487), .Z(n1479) );
  NOR U1459 ( .A(n1488), .B(n1489), .Z(n1487) );
  XNOR U1460 ( .A(n1486), .B(n1490), .Z(n1488) );
  XNOR U1461 ( .A(n1446), .B(n1453), .Z(n1467) );
  NOR U1462 ( .A(n1412), .B(n1491), .Z(n1453) );
  XOR U1463 ( .A(n1458), .B(n1457), .Z(n1446) );
  XNOR U1464 ( .A(n1492), .B(n1454), .Z(n1457) );
  XOR U1465 ( .A(n1493), .B(n1494), .Z(n1454) );
  AND U1466 ( .A(n1495), .B(n1496), .Z(n1494) );
  XOR U1467 ( .A(n1493), .B(n1497), .Z(n1495) );
  XNOR U1468 ( .A(n1498), .B(n1499), .Z(n1492) );
  NOR U1469 ( .A(n1500), .B(n1501), .Z(n1499) );
  XNOR U1470 ( .A(n1498), .B(n1502), .Z(n1500) );
  XOR U1471 ( .A(n1503), .B(n1504), .Z(n1458) );
  NOR U1472 ( .A(n1505), .B(n1506), .Z(n1504) );
  XNOR U1473 ( .A(n1503), .B(n1507), .Z(n1505) );
  XNOR U1474 ( .A(n1397), .B(n1463), .Z(n1465) );
  XOR U1475 ( .A(n1508), .B(n1509), .Z(n1397) );
  AND U1476 ( .A(n31), .B(n1510), .Z(n1509) );
  XOR U1477 ( .A(n1511), .B(n1508), .Z(n1510) );
  AND U1478 ( .A(n1409), .B(n1412), .Z(n1463) );
  XOR U1479 ( .A(n1512), .B(n1491), .Z(n1412) );
  XNOR U1480 ( .A(p_input[256]), .B(p_input[96]), .Z(n1491) );
  XNOR U1481 ( .A(n1478), .B(n1477), .Z(n1512) );
  XNOR U1482 ( .A(n1513), .B(n1485), .Z(n1477) );
  XNOR U1483 ( .A(n1473), .B(n1472), .Z(n1485) );
  XNOR U1484 ( .A(n1514), .B(n1469), .Z(n1472) );
  XNOR U1485 ( .A(p_input[106]), .B(p_input[266]), .Z(n1469) );
  XOR U1486 ( .A(p_input[107]), .B(n831), .Z(n1514) );
  XOR U1487 ( .A(p_input[108]), .B(p_input[268]), .Z(n1473) );
  XNOR U1488 ( .A(n1483), .B(n1474), .Z(n1513) );
  XNOR U1489 ( .A(n1068), .B(p_input[97]), .Z(n1474) );
  XNOR U1490 ( .A(n1515), .B(n1490), .Z(n1483) );
  XNOR U1491 ( .A(p_input[111]), .B(n834), .Z(n1490) );
  XOR U1492 ( .A(n1480), .B(n1489), .Z(n1515) );
  XOR U1493 ( .A(n1516), .B(n1486), .Z(n1489) );
  XOR U1494 ( .A(p_input[109]), .B(p_input[269]), .Z(n1486) );
  XOR U1495 ( .A(p_input[110]), .B(n836), .Z(n1516) );
  XOR U1496 ( .A(p_input[105]), .B(p_input[265]), .Z(n1480) );
  XOR U1497 ( .A(n1497), .B(n1496), .Z(n1478) );
  XNOR U1498 ( .A(n1517), .B(n1502), .Z(n1496) );
  XOR U1499 ( .A(p_input[104]), .B(p_input[264]), .Z(n1502) );
  XOR U1500 ( .A(n1493), .B(n1501), .Z(n1517) );
  XOR U1501 ( .A(n1518), .B(n1498), .Z(n1501) );
  XOR U1502 ( .A(p_input[102]), .B(p_input[262]), .Z(n1498) );
  XOR U1503 ( .A(p_input[103]), .B(n958), .Z(n1518) );
  XNOR U1504 ( .A(n840), .B(p_input[98]), .Z(n1493) );
  XNOR U1505 ( .A(n1507), .B(n1506), .Z(n1497) );
  XOR U1506 ( .A(n1519), .B(n1503), .Z(n1506) );
  XOR U1507 ( .A(p_input[259]), .B(p_input[99]), .Z(n1503) );
  XOR U1508 ( .A(p_input[100]), .B(n960), .Z(n1519) );
  XOR U1509 ( .A(p_input[101]), .B(p_input[261]), .Z(n1507) );
  XOR U1510 ( .A(n1520), .B(n1521), .Z(n1409) );
  AND U1511 ( .A(n31), .B(n1522), .Z(n1521) );
  XNOR U1512 ( .A(n1523), .B(n1520), .Z(n1522) );
  XNOR U1513 ( .A(n1524), .B(n1525), .Z(n31) );
  NOR U1514 ( .A(n1526), .B(n1527), .Z(n1525) );
  XOR U1515 ( .A(n1418), .B(n1524), .Z(n1527) );
  AND U1516 ( .A(n1528), .B(n1529), .Z(n1418) );
  NOR U1517 ( .A(n1524), .B(n1417), .Z(n1526) );
  AND U1518 ( .A(n1530), .B(n1531), .Z(n1417) );
  XOR U1519 ( .A(n1532), .B(n1533), .Z(n1524) );
  AND U1520 ( .A(n1534), .B(n1535), .Z(n1533) );
  XNOR U1521 ( .A(n1532), .B(n1530), .Z(n1535) );
  IV U1522 ( .A(n1435), .Z(n1530) );
  XOR U1523 ( .A(n1536), .B(n1537), .Z(n1435) );
  XOR U1524 ( .A(n1538), .B(n1531), .Z(n1537) );
  AND U1525 ( .A(n1462), .B(n1539), .Z(n1531) );
  AND U1526 ( .A(n1540), .B(n1541), .Z(n1538) );
  XOR U1527 ( .A(n1542), .B(n1536), .Z(n1540) );
  XNOR U1528 ( .A(n1432), .B(n1532), .Z(n1534) );
  XOR U1529 ( .A(n1543), .B(n1544), .Z(n1432) );
  AND U1530 ( .A(n35), .B(n1545), .Z(n1544) );
  XOR U1531 ( .A(n1546), .B(n1543), .Z(n1545) );
  XOR U1532 ( .A(n1547), .B(n1548), .Z(n1532) );
  AND U1533 ( .A(n1549), .B(n1550), .Z(n1548) );
  XNOR U1534 ( .A(n1547), .B(n1462), .Z(n1550) );
  XOR U1535 ( .A(n1551), .B(n1541), .Z(n1462) );
  XNOR U1536 ( .A(n1552), .B(n1536), .Z(n1541) );
  XOR U1537 ( .A(n1553), .B(n1554), .Z(n1536) );
  AND U1538 ( .A(n1555), .B(n1556), .Z(n1554) );
  XOR U1539 ( .A(n1557), .B(n1553), .Z(n1555) );
  XNOR U1540 ( .A(n1558), .B(n1559), .Z(n1552) );
  AND U1541 ( .A(n1560), .B(n1561), .Z(n1559) );
  XOR U1542 ( .A(n1558), .B(n1562), .Z(n1560) );
  XNOR U1543 ( .A(n1542), .B(n1539), .Z(n1551) );
  AND U1544 ( .A(n1563), .B(n1564), .Z(n1539) );
  XOR U1545 ( .A(n1565), .B(n1566), .Z(n1542) );
  AND U1546 ( .A(n1567), .B(n1568), .Z(n1566) );
  XOR U1547 ( .A(n1565), .B(n1569), .Z(n1567) );
  XNOR U1548 ( .A(n1459), .B(n1547), .Z(n1549) );
  XOR U1549 ( .A(n1570), .B(n1571), .Z(n1459) );
  AND U1550 ( .A(n35), .B(n1572), .Z(n1571) );
  XNOR U1551 ( .A(n1573), .B(n1570), .Z(n1572) );
  XOR U1552 ( .A(n1574), .B(n1575), .Z(n1547) );
  AND U1553 ( .A(n1576), .B(n1577), .Z(n1575) );
  XNOR U1554 ( .A(n1574), .B(n1563), .Z(n1577) );
  IV U1555 ( .A(n1511), .Z(n1563) );
  XNOR U1556 ( .A(n1578), .B(n1556), .Z(n1511) );
  XNOR U1557 ( .A(n1579), .B(n1562), .Z(n1556) );
  XNOR U1558 ( .A(n1580), .B(n1581), .Z(n1562) );
  NOR U1559 ( .A(n1582), .B(n1583), .Z(n1581) );
  XOR U1560 ( .A(n1580), .B(n1584), .Z(n1582) );
  XNOR U1561 ( .A(n1561), .B(n1553), .Z(n1579) );
  XOR U1562 ( .A(n1585), .B(n1586), .Z(n1553) );
  AND U1563 ( .A(n1587), .B(n1588), .Z(n1586) );
  XOR U1564 ( .A(n1585), .B(n1589), .Z(n1587) );
  XNOR U1565 ( .A(n1590), .B(n1558), .Z(n1561) );
  XOR U1566 ( .A(n1591), .B(n1592), .Z(n1558) );
  AND U1567 ( .A(n1593), .B(n1594), .Z(n1592) );
  XNOR U1568 ( .A(n1595), .B(n1596), .Z(n1593) );
  IV U1569 ( .A(n1591), .Z(n1595) );
  XNOR U1570 ( .A(n1597), .B(n1598), .Z(n1590) );
  NOR U1571 ( .A(n1599), .B(n1600), .Z(n1598) );
  XNOR U1572 ( .A(n1597), .B(n1601), .Z(n1599) );
  XNOR U1573 ( .A(n1557), .B(n1564), .Z(n1578) );
  NOR U1574 ( .A(n1523), .B(n1602), .Z(n1564) );
  XOR U1575 ( .A(n1569), .B(n1568), .Z(n1557) );
  XNOR U1576 ( .A(n1603), .B(n1565), .Z(n1568) );
  XOR U1577 ( .A(n1604), .B(n1605), .Z(n1565) );
  AND U1578 ( .A(n1606), .B(n1607), .Z(n1605) );
  XNOR U1579 ( .A(n1608), .B(n1609), .Z(n1606) );
  IV U1580 ( .A(n1604), .Z(n1608) );
  XNOR U1581 ( .A(n1610), .B(n1611), .Z(n1603) );
  NOR U1582 ( .A(n1612), .B(n1613), .Z(n1611) );
  XNOR U1583 ( .A(n1610), .B(n1614), .Z(n1612) );
  XOR U1584 ( .A(n1615), .B(n1616), .Z(n1569) );
  NOR U1585 ( .A(n1617), .B(n1618), .Z(n1616) );
  XNOR U1586 ( .A(n1615), .B(n1619), .Z(n1617) );
  XNOR U1587 ( .A(n1508), .B(n1574), .Z(n1576) );
  XOR U1588 ( .A(n1620), .B(n1621), .Z(n1508) );
  AND U1589 ( .A(n35), .B(n1622), .Z(n1621) );
  XOR U1590 ( .A(n1623), .B(n1620), .Z(n1622) );
  AND U1591 ( .A(n1520), .B(n1523), .Z(n1574) );
  XOR U1592 ( .A(n1624), .B(n1602), .Z(n1523) );
  XNOR U1593 ( .A(p_input[112]), .B(p_input[256]), .Z(n1602) );
  XNOR U1594 ( .A(n1589), .B(n1588), .Z(n1624) );
  XNOR U1595 ( .A(n1625), .B(n1596), .Z(n1588) );
  XNOR U1596 ( .A(n1584), .B(n1583), .Z(n1596) );
  XNOR U1597 ( .A(n1626), .B(n1580), .Z(n1583) );
  XNOR U1598 ( .A(p_input[122]), .B(p_input[266]), .Z(n1580) );
  XOR U1599 ( .A(p_input[123]), .B(n831), .Z(n1626) );
  XOR U1600 ( .A(p_input[124]), .B(p_input[268]), .Z(n1584) );
  XOR U1601 ( .A(n1594), .B(n1627), .Z(n1625) );
  IV U1602 ( .A(n1585), .Z(n1627) );
  XOR U1603 ( .A(p_input[113]), .B(p_input[257]), .Z(n1585) );
  XNOR U1604 ( .A(n1628), .B(n1601), .Z(n1594) );
  XNOR U1605 ( .A(p_input[127]), .B(n834), .Z(n1601) );
  XOR U1606 ( .A(n1591), .B(n1600), .Z(n1628) );
  XOR U1607 ( .A(n1629), .B(n1597), .Z(n1600) );
  XOR U1608 ( .A(p_input[125]), .B(p_input[269]), .Z(n1597) );
  XOR U1609 ( .A(p_input[126]), .B(n836), .Z(n1629) );
  XOR U1610 ( .A(p_input[121]), .B(p_input[265]), .Z(n1591) );
  XOR U1611 ( .A(n1609), .B(n1607), .Z(n1589) );
  XNOR U1612 ( .A(n1630), .B(n1614), .Z(n1607) );
  XOR U1613 ( .A(p_input[120]), .B(p_input[264]), .Z(n1614) );
  XOR U1614 ( .A(n1604), .B(n1613), .Z(n1630) );
  XOR U1615 ( .A(n1631), .B(n1610), .Z(n1613) );
  XOR U1616 ( .A(p_input[118]), .B(p_input[262]), .Z(n1610) );
  XOR U1617 ( .A(p_input[119]), .B(n958), .Z(n1631) );
  XOR U1618 ( .A(p_input[114]), .B(p_input[258]), .Z(n1604) );
  XNOR U1619 ( .A(n1619), .B(n1618), .Z(n1609) );
  XOR U1620 ( .A(n1632), .B(n1615), .Z(n1618) );
  XOR U1621 ( .A(p_input[115]), .B(p_input[259]), .Z(n1615) );
  XOR U1622 ( .A(p_input[116]), .B(n960), .Z(n1632) );
  XOR U1623 ( .A(p_input[117]), .B(p_input[261]), .Z(n1619) );
  XOR U1624 ( .A(n1633), .B(n1634), .Z(n1520) );
  AND U1625 ( .A(n35), .B(n1635), .Z(n1634) );
  XNOR U1626 ( .A(n1636), .B(n1633), .Z(n1635) );
  XNOR U1627 ( .A(n1637), .B(n1638), .Z(n35) );
  NOR U1628 ( .A(n1639), .B(n1640), .Z(n1638) );
  XOR U1629 ( .A(n1529), .B(n1637), .Z(n1640) );
  AND U1630 ( .A(n1641), .B(n1642), .Z(n1529) );
  NOR U1631 ( .A(n1637), .B(n1528), .Z(n1639) );
  AND U1632 ( .A(n1643), .B(n1644), .Z(n1528) );
  XOR U1633 ( .A(n1645), .B(n1646), .Z(n1637) );
  AND U1634 ( .A(n1647), .B(n1648), .Z(n1646) );
  XNOR U1635 ( .A(n1645), .B(n1643), .Z(n1648) );
  IV U1636 ( .A(n1546), .Z(n1643) );
  XOR U1637 ( .A(n1649), .B(n1650), .Z(n1546) );
  XOR U1638 ( .A(n1651), .B(n1644), .Z(n1650) );
  AND U1639 ( .A(n1573), .B(n1652), .Z(n1644) );
  AND U1640 ( .A(n1653), .B(n1654), .Z(n1651) );
  XOR U1641 ( .A(n1655), .B(n1649), .Z(n1653) );
  XNOR U1642 ( .A(n1543), .B(n1645), .Z(n1647) );
  XOR U1643 ( .A(n1656), .B(n1657), .Z(n1543) );
  AND U1644 ( .A(n39), .B(n1658), .Z(n1657) );
  XOR U1645 ( .A(n1659), .B(n1656), .Z(n1658) );
  XOR U1646 ( .A(n1660), .B(n1661), .Z(n1645) );
  AND U1647 ( .A(n1662), .B(n1663), .Z(n1661) );
  XNOR U1648 ( .A(n1660), .B(n1573), .Z(n1663) );
  XOR U1649 ( .A(n1664), .B(n1654), .Z(n1573) );
  XNOR U1650 ( .A(n1665), .B(n1649), .Z(n1654) );
  XOR U1651 ( .A(n1666), .B(n1667), .Z(n1649) );
  AND U1652 ( .A(n1668), .B(n1669), .Z(n1667) );
  XOR U1653 ( .A(n1670), .B(n1666), .Z(n1668) );
  XNOR U1654 ( .A(n1671), .B(n1672), .Z(n1665) );
  AND U1655 ( .A(n1673), .B(n1674), .Z(n1672) );
  XOR U1656 ( .A(n1671), .B(n1675), .Z(n1673) );
  XNOR U1657 ( .A(n1655), .B(n1652), .Z(n1664) );
  AND U1658 ( .A(n1676), .B(n1677), .Z(n1652) );
  XOR U1659 ( .A(n1678), .B(n1679), .Z(n1655) );
  AND U1660 ( .A(n1680), .B(n1681), .Z(n1679) );
  XOR U1661 ( .A(n1678), .B(n1682), .Z(n1680) );
  XNOR U1662 ( .A(n1570), .B(n1660), .Z(n1662) );
  XOR U1663 ( .A(n1683), .B(n1684), .Z(n1570) );
  AND U1664 ( .A(n39), .B(n1685), .Z(n1684) );
  XNOR U1665 ( .A(n1686), .B(n1683), .Z(n1685) );
  XOR U1666 ( .A(n1687), .B(n1688), .Z(n1660) );
  AND U1667 ( .A(n1689), .B(n1690), .Z(n1688) );
  XNOR U1668 ( .A(n1687), .B(n1676), .Z(n1690) );
  IV U1669 ( .A(n1623), .Z(n1676) );
  XNOR U1670 ( .A(n1691), .B(n1669), .Z(n1623) );
  XNOR U1671 ( .A(n1692), .B(n1675), .Z(n1669) );
  XNOR U1672 ( .A(n1693), .B(n1694), .Z(n1675) );
  NOR U1673 ( .A(n1695), .B(n1696), .Z(n1694) );
  XOR U1674 ( .A(n1693), .B(n1697), .Z(n1695) );
  XNOR U1675 ( .A(n1674), .B(n1666), .Z(n1692) );
  XOR U1676 ( .A(n1698), .B(n1699), .Z(n1666) );
  AND U1677 ( .A(n1700), .B(n1701), .Z(n1699) );
  XOR U1678 ( .A(n1698), .B(n1702), .Z(n1700) );
  XNOR U1679 ( .A(n1703), .B(n1671), .Z(n1674) );
  XOR U1680 ( .A(n1704), .B(n1705), .Z(n1671) );
  AND U1681 ( .A(n1706), .B(n1707), .Z(n1705) );
  XNOR U1682 ( .A(n1708), .B(n1709), .Z(n1706) );
  IV U1683 ( .A(n1704), .Z(n1708) );
  XNOR U1684 ( .A(n1710), .B(n1711), .Z(n1703) );
  NOR U1685 ( .A(n1712), .B(n1713), .Z(n1711) );
  XNOR U1686 ( .A(n1710), .B(n1714), .Z(n1712) );
  XNOR U1687 ( .A(n1670), .B(n1677), .Z(n1691) );
  NOR U1688 ( .A(n1636), .B(n1715), .Z(n1677) );
  XOR U1689 ( .A(n1682), .B(n1681), .Z(n1670) );
  XNOR U1690 ( .A(n1716), .B(n1678), .Z(n1681) );
  XOR U1691 ( .A(n1717), .B(n1718), .Z(n1678) );
  AND U1692 ( .A(n1719), .B(n1720), .Z(n1718) );
  XNOR U1693 ( .A(n1721), .B(n1722), .Z(n1719) );
  IV U1694 ( .A(n1717), .Z(n1721) );
  XNOR U1695 ( .A(n1723), .B(n1724), .Z(n1716) );
  NOR U1696 ( .A(n1725), .B(n1726), .Z(n1724) );
  XNOR U1697 ( .A(n1723), .B(n1727), .Z(n1725) );
  XOR U1698 ( .A(n1728), .B(n1729), .Z(n1682) );
  NOR U1699 ( .A(n1730), .B(n1731), .Z(n1729) );
  XNOR U1700 ( .A(n1728), .B(n1732), .Z(n1730) );
  XNOR U1701 ( .A(n1620), .B(n1687), .Z(n1689) );
  XOR U1702 ( .A(n1733), .B(n1734), .Z(n1620) );
  AND U1703 ( .A(n39), .B(n1735), .Z(n1734) );
  XOR U1704 ( .A(n1736), .B(n1733), .Z(n1735) );
  AND U1705 ( .A(n1633), .B(n1636), .Z(n1687) );
  XOR U1706 ( .A(n1737), .B(n1715), .Z(n1636) );
  XNOR U1707 ( .A(p_input[128]), .B(p_input[256]), .Z(n1715) );
  XNOR U1708 ( .A(n1702), .B(n1701), .Z(n1737) );
  XNOR U1709 ( .A(n1738), .B(n1709), .Z(n1701) );
  XNOR U1710 ( .A(n1697), .B(n1696), .Z(n1709) );
  XNOR U1711 ( .A(n1739), .B(n1693), .Z(n1696) );
  XNOR U1712 ( .A(p_input[138]), .B(p_input[266]), .Z(n1693) );
  XOR U1713 ( .A(p_input[139]), .B(n831), .Z(n1739) );
  XOR U1714 ( .A(p_input[140]), .B(p_input[268]), .Z(n1697) );
  XOR U1715 ( .A(n1707), .B(n1740), .Z(n1738) );
  IV U1716 ( .A(n1698), .Z(n1740) );
  XOR U1717 ( .A(p_input[129]), .B(p_input[257]), .Z(n1698) );
  XNOR U1718 ( .A(n1741), .B(n1714), .Z(n1707) );
  XNOR U1719 ( .A(p_input[143]), .B(n834), .Z(n1714) );
  XOR U1720 ( .A(n1704), .B(n1713), .Z(n1741) );
  XOR U1721 ( .A(n1742), .B(n1710), .Z(n1713) );
  XOR U1722 ( .A(p_input[141]), .B(p_input[269]), .Z(n1710) );
  XOR U1723 ( .A(p_input[142]), .B(n836), .Z(n1742) );
  XOR U1724 ( .A(p_input[137]), .B(p_input[265]), .Z(n1704) );
  XOR U1725 ( .A(n1722), .B(n1720), .Z(n1702) );
  XNOR U1726 ( .A(n1743), .B(n1727), .Z(n1720) );
  XOR U1727 ( .A(p_input[136]), .B(p_input[264]), .Z(n1727) );
  XOR U1728 ( .A(n1717), .B(n1726), .Z(n1743) );
  XOR U1729 ( .A(n1744), .B(n1723), .Z(n1726) );
  XOR U1730 ( .A(p_input[134]), .B(p_input[262]), .Z(n1723) );
  XOR U1731 ( .A(p_input[135]), .B(n958), .Z(n1744) );
  XOR U1732 ( .A(p_input[130]), .B(p_input[258]), .Z(n1717) );
  XNOR U1733 ( .A(n1732), .B(n1731), .Z(n1722) );
  XOR U1734 ( .A(n1745), .B(n1728), .Z(n1731) );
  XOR U1735 ( .A(p_input[131]), .B(p_input[259]), .Z(n1728) );
  XOR U1736 ( .A(p_input[132]), .B(n960), .Z(n1745) );
  XOR U1737 ( .A(p_input[133]), .B(p_input[261]), .Z(n1732) );
  XOR U1738 ( .A(n1746), .B(n1747), .Z(n1633) );
  AND U1739 ( .A(n39), .B(n1748), .Z(n1747) );
  XNOR U1740 ( .A(n1749), .B(n1746), .Z(n1748) );
  XNOR U1741 ( .A(n1750), .B(n1751), .Z(n39) );
  NOR U1742 ( .A(n1752), .B(n1753), .Z(n1751) );
  XOR U1743 ( .A(n1642), .B(n1750), .Z(n1753) );
  AND U1744 ( .A(n1754), .B(n1755), .Z(n1642) );
  NOR U1745 ( .A(n1750), .B(n1641), .Z(n1752) );
  AND U1746 ( .A(n1756), .B(n1757), .Z(n1641) );
  XOR U1747 ( .A(n1758), .B(n1759), .Z(n1750) );
  AND U1748 ( .A(n1760), .B(n1761), .Z(n1759) );
  XNOR U1749 ( .A(n1758), .B(n1756), .Z(n1761) );
  IV U1750 ( .A(n1659), .Z(n1756) );
  XOR U1751 ( .A(n1762), .B(n1763), .Z(n1659) );
  XOR U1752 ( .A(n1764), .B(n1757), .Z(n1763) );
  AND U1753 ( .A(n1686), .B(n1765), .Z(n1757) );
  AND U1754 ( .A(n1766), .B(n1767), .Z(n1764) );
  XOR U1755 ( .A(n1768), .B(n1762), .Z(n1766) );
  XNOR U1756 ( .A(n1656), .B(n1758), .Z(n1760) );
  XOR U1757 ( .A(n1769), .B(n1770), .Z(n1656) );
  AND U1758 ( .A(n43), .B(n1771), .Z(n1770) );
  XOR U1759 ( .A(n1772), .B(n1769), .Z(n1771) );
  XOR U1760 ( .A(n1773), .B(n1774), .Z(n1758) );
  AND U1761 ( .A(n1775), .B(n1776), .Z(n1774) );
  XNOR U1762 ( .A(n1773), .B(n1686), .Z(n1776) );
  XOR U1763 ( .A(n1777), .B(n1767), .Z(n1686) );
  XNOR U1764 ( .A(n1778), .B(n1762), .Z(n1767) );
  XOR U1765 ( .A(n1779), .B(n1780), .Z(n1762) );
  AND U1766 ( .A(n1781), .B(n1782), .Z(n1780) );
  XOR U1767 ( .A(n1783), .B(n1779), .Z(n1781) );
  XNOR U1768 ( .A(n1784), .B(n1785), .Z(n1778) );
  AND U1769 ( .A(n1786), .B(n1787), .Z(n1785) );
  XOR U1770 ( .A(n1784), .B(n1788), .Z(n1786) );
  XNOR U1771 ( .A(n1768), .B(n1765), .Z(n1777) );
  AND U1772 ( .A(n1789), .B(n1790), .Z(n1765) );
  XOR U1773 ( .A(n1791), .B(n1792), .Z(n1768) );
  AND U1774 ( .A(n1793), .B(n1794), .Z(n1792) );
  XOR U1775 ( .A(n1791), .B(n1795), .Z(n1793) );
  XNOR U1776 ( .A(n1683), .B(n1773), .Z(n1775) );
  XOR U1777 ( .A(n1796), .B(n1797), .Z(n1683) );
  AND U1778 ( .A(n43), .B(n1798), .Z(n1797) );
  XNOR U1779 ( .A(n1799), .B(n1796), .Z(n1798) );
  XOR U1780 ( .A(n1800), .B(n1801), .Z(n1773) );
  AND U1781 ( .A(n1802), .B(n1803), .Z(n1801) );
  XNOR U1782 ( .A(n1800), .B(n1789), .Z(n1803) );
  IV U1783 ( .A(n1736), .Z(n1789) );
  XNOR U1784 ( .A(n1804), .B(n1782), .Z(n1736) );
  XNOR U1785 ( .A(n1805), .B(n1788), .Z(n1782) );
  XNOR U1786 ( .A(n1806), .B(n1807), .Z(n1788) );
  NOR U1787 ( .A(n1808), .B(n1809), .Z(n1807) );
  XOR U1788 ( .A(n1806), .B(n1810), .Z(n1808) );
  XNOR U1789 ( .A(n1787), .B(n1779), .Z(n1805) );
  XOR U1790 ( .A(n1811), .B(n1812), .Z(n1779) );
  AND U1791 ( .A(n1813), .B(n1814), .Z(n1812) );
  XOR U1792 ( .A(n1811), .B(n1815), .Z(n1813) );
  XNOR U1793 ( .A(n1816), .B(n1784), .Z(n1787) );
  XOR U1794 ( .A(n1817), .B(n1818), .Z(n1784) );
  AND U1795 ( .A(n1819), .B(n1820), .Z(n1818) );
  XNOR U1796 ( .A(n1821), .B(n1822), .Z(n1819) );
  IV U1797 ( .A(n1817), .Z(n1821) );
  XNOR U1798 ( .A(n1823), .B(n1824), .Z(n1816) );
  NOR U1799 ( .A(n1825), .B(n1826), .Z(n1824) );
  XNOR U1800 ( .A(n1823), .B(n1827), .Z(n1825) );
  XNOR U1801 ( .A(n1783), .B(n1790), .Z(n1804) );
  NOR U1802 ( .A(n1749), .B(n1828), .Z(n1790) );
  XOR U1803 ( .A(n1795), .B(n1794), .Z(n1783) );
  XNOR U1804 ( .A(n1829), .B(n1791), .Z(n1794) );
  XOR U1805 ( .A(n1830), .B(n1831), .Z(n1791) );
  AND U1806 ( .A(n1832), .B(n1833), .Z(n1831) );
  XNOR U1807 ( .A(n1834), .B(n1835), .Z(n1832) );
  IV U1808 ( .A(n1830), .Z(n1834) );
  XNOR U1809 ( .A(n1836), .B(n1837), .Z(n1829) );
  NOR U1810 ( .A(n1838), .B(n1839), .Z(n1837) );
  XNOR U1811 ( .A(n1836), .B(n1840), .Z(n1838) );
  XOR U1812 ( .A(n1841), .B(n1842), .Z(n1795) );
  NOR U1813 ( .A(n1843), .B(n1844), .Z(n1842) );
  XNOR U1814 ( .A(n1841), .B(n1845), .Z(n1843) );
  XNOR U1815 ( .A(n1733), .B(n1800), .Z(n1802) );
  XOR U1816 ( .A(n1846), .B(n1847), .Z(n1733) );
  AND U1817 ( .A(n43), .B(n1848), .Z(n1847) );
  XOR U1818 ( .A(n1849), .B(n1846), .Z(n1848) );
  AND U1819 ( .A(n1746), .B(n1749), .Z(n1800) );
  XOR U1820 ( .A(n1850), .B(n1828), .Z(n1749) );
  XNOR U1821 ( .A(p_input[144]), .B(p_input[256]), .Z(n1828) );
  XNOR U1822 ( .A(n1815), .B(n1814), .Z(n1850) );
  XNOR U1823 ( .A(n1851), .B(n1822), .Z(n1814) );
  XNOR U1824 ( .A(n1810), .B(n1809), .Z(n1822) );
  XNOR U1825 ( .A(n1852), .B(n1806), .Z(n1809) );
  XNOR U1826 ( .A(p_input[154]), .B(p_input[266]), .Z(n1806) );
  XOR U1827 ( .A(p_input[155]), .B(n831), .Z(n1852) );
  XOR U1828 ( .A(p_input[156]), .B(p_input[268]), .Z(n1810) );
  XOR U1829 ( .A(n1820), .B(n1853), .Z(n1851) );
  IV U1830 ( .A(n1811), .Z(n1853) );
  XOR U1831 ( .A(p_input[145]), .B(p_input[257]), .Z(n1811) );
  XNOR U1832 ( .A(n1854), .B(n1827), .Z(n1820) );
  XNOR U1833 ( .A(p_input[159]), .B(n834), .Z(n1827) );
  XOR U1834 ( .A(n1817), .B(n1826), .Z(n1854) );
  XOR U1835 ( .A(n1855), .B(n1823), .Z(n1826) );
  XOR U1836 ( .A(p_input[157]), .B(p_input[269]), .Z(n1823) );
  XOR U1837 ( .A(p_input[158]), .B(n836), .Z(n1855) );
  XOR U1838 ( .A(p_input[153]), .B(p_input[265]), .Z(n1817) );
  XOR U1839 ( .A(n1835), .B(n1833), .Z(n1815) );
  XNOR U1840 ( .A(n1856), .B(n1840), .Z(n1833) );
  XOR U1841 ( .A(p_input[152]), .B(p_input[264]), .Z(n1840) );
  XOR U1842 ( .A(n1830), .B(n1839), .Z(n1856) );
  XOR U1843 ( .A(n1857), .B(n1836), .Z(n1839) );
  XOR U1844 ( .A(p_input[150]), .B(p_input[262]), .Z(n1836) );
  XOR U1845 ( .A(p_input[151]), .B(n958), .Z(n1857) );
  XOR U1846 ( .A(p_input[146]), .B(p_input[258]), .Z(n1830) );
  XNOR U1847 ( .A(n1845), .B(n1844), .Z(n1835) );
  XOR U1848 ( .A(n1858), .B(n1841), .Z(n1844) );
  XOR U1849 ( .A(p_input[147]), .B(p_input[259]), .Z(n1841) );
  XOR U1850 ( .A(p_input[148]), .B(n960), .Z(n1858) );
  XOR U1851 ( .A(p_input[149]), .B(p_input[261]), .Z(n1845) );
  XOR U1852 ( .A(n1859), .B(n1860), .Z(n1746) );
  AND U1853 ( .A(n43), .B(n1861), .Z(n1860) );
  XNOR U1854 ( .A(n1862), .B(n1859), .Z(n1861) );
  XNOR U1855 ( .A(n1863), .B(n1864), .Z(n43) );
  NOR U1856 ( .A(n1865), .B(n1866), .Z(n1864) );
  XOR U1857 ( .A(n1755), .B(n1863), .Z(n1866) );
  AND U1858 ( .A(n1867), .B(n1868), .Z(n1755) );
  NOR U1859 ( .A(n1863), .B(n1754), .Z(n1865) );
  AND U1860 ( .A(n1869), .B(n1870), .Z(n1754) );
  XOR U1861 ( .A(n1871), .B(n1872), .Z(n1863) );
  AND U1862 ( .A(n1873), .B(n1874), .Z(n1872) );
  XNOR U1863 ( .A(n1871), .B(n1869), .Z(n1874) );
  IV U1864 ( .A(n1772), .Z(n1869) );
  XOR U1865 ( .A(n1875), .B(n1876), .Z(n1772) );
  XOR U1866 ( .A(n1877), .B(n1870), .Z(n1876) );
  AND U1867 ( .A(n1799), .B(n1878), .Z(n1870) );
  AND U1868 ( .A(n1879), .B(n1880), .Z(n1877) );
  XOR U1869 ( .A(n1881), .B(n1875), .Z(n1879) );
  XNOR U1870 ( .A(n1769), .B(n1871), .Z(n1873) );
  XOR U1871 ( .A(n1882), .B(n1883), .Z(n1769) );
  AND U1872 ( .A(n47), .B(n1884), .Z(n1883) );
  XOR U1873 ( .A(n1885), .B(n1882), .Z(n1884) );
  XOR U1874 ( .A(n1886), .B(n1887), .Z(n1871) );
  AND U1875 ( .A(n1888), .B(n1889), .Z(n1887) );
  XNOR U1876 ( .A(n1886), .B(n1799), .Z(n1889) );
  XOR U1877 ( .A(n1890), .B(n1880), .Z(n1799) );
  XNOR U1878 ( .A(n1891), .B(n1875), .Z(n1880) );
  XOR U1879 ( .A(n1892), .B(n1893), .Z(n1875) );
  AND U1880 ( .A(n1894), .B(n1895), .Z(n1893) );
  XOR U1881 ( .A(n1896), .B(n1892), .Z(n1894) );
  XNOR U1882 ( .A(n1897), .B(n1898), .Z(n1891) );
  AND U1883 ( .A(n1899), .B(n1900), .Z(n1898) );
  XOR U1884 ( .A(n1897), .B(n1901), .Z(n1899) );
  XNOR U1885 ( .A(n1881), .B(n1878), .Z(n1890) );
  AND U1886 ( .A(n1902), .B(n1903), .Z(n1878) );
  XOR U1887 ( .A(n1904), .B(n1905), .Z(n1881) );
  AND U1888 ( .A(n1906), .B(n1907), .Z(n1905) );
  XOR U1889 ( .A(n1904), .B(n1908), .Z(n1906) );
  XNOR U1890 ( .A(n1796), .B(n1886), .Z(n1888) );
  XOR U1891 ( .A(n1909), .B(n1910), .Z(n1796) );
  AND U1892 ( .A(n47), .B(n1911), .Z(n1910) );
  XNOR U1893 ( .A(n1912), .B(n1909), .Z(n1911) );
  XOR U1894 ( .A(n1913), .B(n1914), .Z(n1886) );
  AND U1895 ( .A(n1915), .B(n1916), .Z(n1914) );
  XNOR U1896 ( .A(n1913), .B(n1902), .Z(n1916) );
  IV U1897 ( .A(n1849), .Z(n1902) );
  XNOR U1898 ( .A(n1917), .B(n1895), .Z(n1849) );
  XNOR U1899 ( .A(n1918), .B(n1901), .Z(n1895) );
  XNOR U1900 ( .A(n1919), .B(n1920), .Z(n1901) );
  NOR U1901 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U1902 ( .A(n1919), .B(n1923), .Z(n1921) );
  XNOR U1903 ( .A(n1900), .B(n1892), .Z(n1918) );
  XOR U1904 ( .A(n1924), .B(n1925), .Z(n1892) );
  AND U1905 ( .A(n1926), .B(n1927), .Z(n1925) );
  XOR U1906 ( .A(n1924), .B(n1928), .Z(n1926) );
  XNOR U1907 ( .A(n1929), .B(n1897), .Z(n1900) );
  XOR U1908 ( .A(n1930), .B(n1931), .Z(n1897) );
  AND U1909 ( .A(n1932), .B(n1933), .Z(n1931) );
  XNOR U1910 ( .A(n1934), .B(n1935), .Z(n1932) );
  IV U1911 ( .A(n1930), .Z(n1934) );
  XNOR U1912 ( .A(n1936), .B(n1937), .Z(n1929) );
  NOR U1913 ( .A(n1938), .B(n1939), .Z(n1937) );
  XNOR U1914 ( .A(n1936), .B(n1940), .Z(n1938) );
  XNOR U1915 ( .A(n1896), .B(n1903), .Z(n1917) );
  NOR U1916 ( .A(n1862), .B(n1941), .Z(n1903) );
  XOR U1917 ( .A(n1908), .B(n1907), .Z(n1896) );
  XNOR U1918 ( .A(n1942), .B(n1904), .Z(n1907) );
  XOR U1919 ( .A(n1943), .B(n1944), .Z(n1904) );
  AND U1920 ( .A(n1945), .B(n1946), .Z(n1944) );
  XNOR U1921 ( .A(n1947), .B(n1948), .Z(n1945) );
  IV U1922 ( .A(n1943), .Z(n1947) );
  XNOR U1923 ( .A(n1949), .B(n1950), .Z(n1942) );
  NOR U1924 ( .A(n1951), .B(n1952), .Z(n1950) );
  XNOR U1925 ( .A(n1949), .B(n1953), .Z(n1951) );
  XOR U1926 ( .A(n1954), .B(n1955), .Z(n1908) );
  NOR U1927 ( .A(n1956), .B(n1957), .Z(n1955) );
  XNOR U1928 ( .A(n1954), .B(n1958), .Z(n1956) );
  XNOR U1929 ( .A(n1846), .B(n1913), .Z(n1915) );
  XOR U1930 ( .A(n1959), .B(n1960), .Z(n1846) );
  AND U1931 ( .A(n47), .B(n1961), .Z(n1960) );
  XOR U1932 ( .A(n1962), .B(n1959), .Z(n1961) );
  AND U1933 ( .A(n1859), .B(n1862), .Z(n1913) );
  XOR U1934 ( .A(n1963), .B(n1941), .Z(n1862) );
  XNOR U1935 ( .A(p_input[160]), .B(p_input[256]), .Z(n1941) );
  XNOR U1936 ( .A(n1928), .B(n1927), .Z(n1963) );
  XNOR U1937 ( .A(n1964), .B(n1935), .Z(n1927) );
  XNOR U1938 ( .A(n1923), .B(n1922), .Z(n1935) );
  XNOR U1939 ( .A(n1965), .B(n1919), .Z(n1922) );
  XNOR U1940 ( .A(p_input[170]), .B(p_input[266]), .Z(n1919) );
  XOR U1941 ( .A(p_input[171]), .B(n831), .Z(n1965) );
  XOR U1942 ( .A(p_input[172]), .B(p_input[268]), .Z(n1923) );
  XOR U1943 ( .A(n1933), .B(n1966), .Z(n1964) );
  IV U1944 ( .A(n1924), .Z(n1966) );
  XOR U1945 ( .A(p_input[161]), .B(p_input[257]), .Z(n1924) );
  XNOR U1946 ( .A(n1967), .B(n1940), .Z(n1933) );
  XNOR U1947 ( .A(p_input[175]), .B(n834), .Z(n1940) );
  XOR U1948 ( .A(n1930), .B(n1939), .Z(n1967) );
  XOR U1949 ( .A(n1968), .B(n1936), .Z(n1939) );
  XOR U1950 ( .A(p_input[173]), .B(p_input[269]), .Z(n1936) );
  XOR U1951 ( .A(p_input[174]), .B(n836), .Z(n1968) );
  XOR U1952 ( .A(p_input[169]), .B(p_input[265]), .Z(n1930) );
  XOR U1953 ( .A(n1948), .B(n1946), .Z(n1928) );
  XNOR U1954 ( .A(n1969), .B(n1953), .Z(n1946) );
  XOR U1955 ( .A(p_input[168]), .B(p_input[264]), .Z(n1953) );
  XOR U1956 ( .A(n1943), .B(n1952), .Z(n1969) );
  XOR U1957 ( .A(n1970), .B(n1949), .Z(n1952) );
  XOR U1958 ( .A(p_input[166]), .B(p_input[262]), .Z(n1949) );
  XOR U1959 ( .A(p_input[167]), .B(n958), .Z(n1970) );
  XOR U1960 ( .A(p_input[162]), .B(p_input[258]), .Z(n1943) );
  XNOR U1961 ( .A(n1958), .B(n1957), .Z(n1948) );
  XOR U1962 ( .A(n1971), .B(n1954), .Z(n1957) );
  XOR U1963 ( .A(p_input[163]), .B(p_input[259]), .Z(n1954) );
  XOR U1964 ( .A(p_input[164]), .B(n960), .Z(n1971) );
  XOR U1965 ( .A(p_input[165]), .B(p_input[261]), .Z(n1958) );
  XOR U1966 ( .A(n1972), .B(n1973), .Z(n1859) );
  AND U1967 ( .A(n47), .B(n1974), .Z(n1973) );
  XNOR U1968 ( .A(n1975), .B(n1972), .Z(n1974) );
  XNOR U1969 ( .A(n1976), .B(n1977), .Z(n47) );
  NOR U1970 ( .A(n1978), .B(n1979), .Z(n1977) );
  XOR U1971 ( .A(n1868), .B(n1976), .Z(n1979) );
  AND U1972 ( .A(n1980), .B(n1981), .Z(n1868) );
  NOR U1973 ( .A(n1976), .B(n1867), .Z(n1978) );
  AND U1974 ( .A(n1982), .B(n1983), .Z(n1867) );
  XOR U1975 ( .A(n1984), .B(n1985), .Z(n1976) );
  AND U1976 ( .A(n1986), .B(n1987), .Z(n1985) );
  XNOR U1977 ( .A(n1984), .B(n1982), .Z(n1987) );
  IV U1978 ( .A(n1885), .Z(n1982) );
  XOR U1979 ( .A(n1988), .B(n1989), .Z(n1885) );
  XOR U1980 ( .A(n1990), .B(n1983), .Z(n1989) );
  AND U1981 ( .A(n1912), .B(n1991), .Z(n1983) );
  AND U1982 ( .A(n1992), .B(n1993), .Z(n1990) );
  XOR U1983 ( .A(n1994), .B(n1988), .Z(n1992) );
  XNOR U1984 ( .A(n1882), .B(n1984), .Z(n1986) );
  XOR U1985 ( .A(n1995), .B(n1996), .Z(n1882) );
  AND U1986 ( .A(n51), .B(n1997), .Z(n1996) );
  XOR U1987 ( .A(n1998), .B(n1995), .Z(n1997) );
  XOR U1988 ( .A(n1999), .B(n2000), .Z(n1984) );
  AND U1989 ( .A(n2001), .B(n2002), .Z(n2000) );
  XNOR U1990 ( .A(n1999), .B(n1912), .Z(n2002) );
  XOR U1991 ( .A(n2003), .B(n1993), .Z(n1912) );
  XNOR U1992 ( .A(n2004), .B(n1988), .Z(n1993) );
  XOR U1993 ( .A(n2005), .B(n2006), .Z(n1988) );
  AND U1994 ( .A(n2007), .B(n2008), .Z(n2006) );
  XOR U1995 ( .A(n2009), .B(n2005), .Z(n2007) );
  XNOR U1996 ( .A(n2010), .B(n2011), .Z(n2004) );
  AND U1997 ( .A(n2012), .B(n2013), .Z(n2011) );
  XOR U1998 ( .A(n2010), .B(n2014), .Z(n2012) );
  XNOR U1999 ( .A(n1994), .B(n1991), .Z(n2003) );
  AND U2000 ( .A(n2015), .B(n2016), .Z(n1991) );
  XOR U2001 ( .A(n2017), .B(n2018), .Z(n1994) );
  AND U2002 ( .A(n2019), .B(n2020), .Z(n2018) );
  XOR U2003 ( .A(n2017), .B(n2021), .Z(n2019) );
  XNOR U2004 ( .A(n1909), .B(n1999), .Z(n2001) );
  XOR U2005 ( .A(n2022), .B(n2023), .Z(n1909) );
  AND U2006 ( .A(n51), .B(n2024), .Z(n2023) );
  XNOR U2007 ( .A(n2025), .B(n2022), .Z(n2024) );
  XOR U2008 ( .A(n2026), .B(n2027), .Z(n1999) );
  AND U2009 ( .A(n2028), .B(n2029), .Z(n2027) );
  XNOR U2010 ( .A(n2026), .B(n2015), .Z(n2029) );
  IV U2011 ( .A(n1962), .Z(n2015) );
  XNOR U2012 ( .A(n2030), .B(n2008), .Z(n1962) );
  XNOR U2013 ( .A(n2031), .B(n2014), .Z(n2008) );
  XNOR U2014 ( .A(n2032), .B(n2033), .Z(n2014) );
  NOR U2015 ( .A(n2034), .B(n2035), .Z(n2033) );
  XOR U2016 ( .A(n2032), .B(n2036), .Z(n2034) );
  XNOR U2017 ( .A(n2013), .B(n2005), .Z(n2031) );
  XOR U2018 ( .A(n2037), .B(n2038), .Z(n2005) );
  AND U2019 ( .A(n2039), .B(n2040), .Z(n2038) );
  XOR U2020 ( .A(n2037), .B(n2041), .Z(n2039) );
  XNOR U2021 ( .A(n2042), .B(n2010), .Z(n2013) );
  XOR U2022 ( .A(n2043), .B(n2044), .Z(n2010) );
  AND U2023 ( .A(n2045), .B(n2046), .Z(n2044) );
  XNOR U2024 ( .A(n2047), .B(n2048), .Z(n2045) );
  IV U2025 ( .A(n2043), .Z(n2047) );
  XNOR U2026 ( .A(n2049), .B(n2050), .Z(n2042) );
  NOR U2027 ( .A(n2051), .B(n2052), .Z(n2050) );
  XNOR U2028 ( .A(n2049), .B(n2053), .Z(n2051) );
  XNOR U2029 ( .A(n2009), .B(n2016), .Z(n2030) );
  NOR U2030 ( .A(n1975), .B(n2054), .Z(n2016) );
  XOR U2031 ( .A(n2021), .B(n2020), .Z(n2009) );
  XNOR U2032 ( .A(n2055), .B(n2017), .Z(n2020) );
  XOR U2033 ( .A(n2056), .B(n2057), .Z(n2017) );
  AND U2034 ( .A(n2058), .B(n2059), .Z(n2057) );
  XNOR U2035 ( .A(n2060), .B(n2061), .Z(n2058) );
  IV U2036 ( .A(n2056), .Z(n2060) );
  XNOR U2037 ( .A(n2062), .B(n2063), .Z(n2055) );
  NOR U2038 ( .A(n2064), .B(n2065), .Z(n2063) );
  XNOR U2039 ( .A(n2062), .B(n2066), .Z(n2064) );
  XOR U2040 ( .A(n2067), .B(n2068), .Z(n2021) );
  NOR U2041 ( .A(n2069), .B(n2070), .Z(n2068) );
  XNOR U2042 ( .A(n2067), .B(n2071), .Z(n2069) );
  XNOR U2043 ( .A(n1959), .B(n2026), .Z(n2028) );
  XOR U2044 ( .A(n2072), .B(n2073), .Z(n1959) );
  AND U2045 ( .A(n51), .B(n2074), .Z(n2073) );
  XOR U2046 ( .A(n2075), .B(n2072), .Z(n2074) );
  AND U2047 ( .A(n1972), .B(n1975), .Z(n2026) );
  XOR U2048 ( .A(n2076), .B(n2054), .Z(n1975) );
  XNOR U2049 ( .A(p_input[176]), .B(p_input[256]), .Z(n2054) );
  XNOR U2050 ( .A(n2041), .B(n2040), .Z(n2076) );
  XNOR U2051 ( .A(n2077), .B(n2048), .Z(n2040) );
  XNOR U2052 ( .A(n2036), .B(n2035), .Z(n2048) );
  XNOR U2053 ( .A(n2078), .B(n2032), .Z(n2035) );
  XNOR U2054 ( .A(p_input[186]), .B(p_input[266]), .Z(n2032) );
  XOR U2055 ( .A(p_input[187]), .B(n831), .Z(n2078) );
  XOR U2056 ( .A(p_input[188]), .B(p_input[268]), .Z(n2036) );
  XOR U2057 ( .A(n2046), .B(n2079), .Z(n2077) );
  IV U2058 ( .A(n2037), .Z(n2079) );
  XOR U2059 ( .A(p_input[177]), .B(p_input[257]), .Z(n2037) );
  XNOR U2060 ( .A(n2080), .B(n2053), .Z(n2046) );
  XNOR U2061 ( .A(p_input[191]), .B(n834), .Z(n2053) );
  XOR U2062 ( .A(n2043), .B(n2052), .Z(n2080) );
  XOR U2063 ( .A(n2081), .B(n2049), .Z(n2052) );
  XOR U2064 ( .A(p_input[189]), .B(p_input[269]), .Z(n2049) );
  XOR U2065 ( .A(p_input[190]), .B(n836), .Z(n2081) );
  XOR U2066 ( .A(p_input[185]), .B(p_input[265]), .Z(n2043) );
  XOR U2067 ( .A(n2061), .B(n2059), .Z(n2041) );
  XNOR U2068 ( .A(n2082), .B(n2066), .Z(n2059) );
  XOR U2069 ( .A(p_input[184]), .B(p_input[264]), .Z(n2066) );
  XOR U2070 ( .A(n2056), .B(n2065), .Z(n2082) );
  XOR U2071 ( .A(n2083), .B(n2062), .Z(n2065) );
  XOR U2072 ( .A(p_input[182]), .B(p_input[262]), .Z(n2062) );
  XOR U2073 ( .A(p_input[183]), .B(n958), .Z(n2083) );
  XOR U2074 ( .A(p_input[178]), .B(p_input[258]), .Z(n2056) );
  XNOR U2075 ( .A(n2071), .B(n2070), .Z(n2061) );
  XOR U2076 ( .A(n2084), .B(n2067), .Z(n2070) );
  XOR U2077 ( .A(p_input[179]), .B(p_input[259]), .Z(n2067) );
  XOR U2078 ( .A(p_input[180]), .B(n960), .Z(n2084) );
  XOR U2079 ( .A(p_input[181]), .B(p_input[261]), .Z(n2071) );
  XOR U2080 ( .A(n2085), .B(n2086), .Z(n1972) );
  AND U2081 ( .A(n51), .B(n2087), .Z(n2086) );
  XNOR U2082 ( .A(n2088), .B(n2085), .Z(n2087) );
  XNOR U2083 ( .A(n2089), .B(n2090), .Z(n51) );
  NOR U2084 ( .A(n2091), .B(n2092), .Z(n2090) );
  XOR U2085 ( .A(n1981), .B(n2089), .Z(n2092) );
  AND U2086 ( .A(n2093), .B(n2094), .Z(n1981) );
  NOR U2087 ( .A(n2089), .B(n1980), .Z(n2091) );
  AND U2088 ( .A(n2095), .B(n2096), .Z(n1980) );
  XOR U2089 ( .A(n2097), .B(n2098), .Z(n2089) );
  AND U2090 ( .A(n2099), .B(n2100), .Z(n2098) );
  XNOR U2091 ( .A(n2097), .B(n2095), .Z(n2100) );
  IV U2092 ( .A(n1998), .Z(n2095) );
  XOR U2093 ( .A(n2101), .B(n2102), .Z(n1998) );
  XOR U2094 ( .A(n2103), .B(n2096), .Z(n2102) );
  AND U2095 ( .A(n2025), .B(n2104), .Z(n2096) );
  AND U2096 ( .A(n2105), .B(n2106), .Z(n2103) );
  XOR U2097 ( .A(n2107), .B(n2101), .Z(n2105) );
  XNOR U2098 ( .A(n1995), .B(n2097), .Z(n2099) );
  XOR U2099 ( .A(n2108), .B(n2109), .Z(n1995) );
  AND U2100 ( .A(n55), .B(n2110), .Z(n2109) );
  XOR U2101 ( .A(n2111), .B(n2108), .Z(n2110) );
  XOR U2102 ( .A(n2112), .B(n2113), .Z(n2097) );
  AND U2103 ( .A(n2114), .B(n2115), .Z(n2113) );
  XNOR U2104 ( .A(n2112), .B(n2025), .Z(n2115) );
  XOR U2105 ( .A(n2116), .B(n2106), .Z(n2025) );
  XNOR U2106 ( .A(n2117), .B(n2101), .Z(n2106) );
  XOR U2107 ( .A(n2118), .B(n2119), .Z(n2101) );
  AND U2108 ( .A(n2120), .B(n2121), .Z(n2119) );
  XOR U2109 ( .A(n2122), .B(n2118), .Z(n2120) );
  XNOR U2110 ( .A(n2123), .B(n2124), .Z(n2117) );
  AND U2111 ( .A(n2125), .B(n2126), .Z(n2124) );
  XOR U2112 ( .A(n2123), .B(n2127), .Z(n2125) );
  XNOR U2113 ( .A(n2107), .B(n2104), .Z(n2116) );
  AND U2114 ( .A(n2128), .B(n2129), .Z(n2104) );
  XOR U2115 ( .A(n2130), .B(n2131), .Z(n2107) );
  AND U2116 ( .A(n2132), .B(n2133), .Z(n2131) );
  XOR U2117 ( .A(n2130), .B(n2134), .Z(n2132) );
  XNOR U2118 ( .A(n2022), .B(n2112), .Z(n2114) );
  XOR U2119 ( .A(n2135), .B(n2136), .Z(n2022) );
  AND U2120 ( .A(n55), .B(n2137), .Z(n2136) );
  XNOR U2121 ( .A(n2138), .B(n2135), .Z(n2137) );
  XOR U2122 ( .A(n2139), .B(n2140), .Z(n2112) );
  AND U2123 ( .A(n2141), .B(n2142), .Z(n2140) );
  XNOR U2124 ( .A(n2139), .B(n2128), .Z(n2142) );
  IV U2125 ( .A(n2075), .Z(n2128) );
  XNOR U2126 ( .A(n2143), .B(n2121), .Z(n2075) );
  XNOR U2127 ( .A(n2144), .B(n2127), .Z(n2121) );
  XNOR U2128 ( .A(n2145), .B(n2146), .Z(n2127) );
  NOR U2129 ( .A(n2147), .B(n2148), .Z(n2146) );
  XOR U2130 ( .A(n2145), .B(n2149), .Z(n2147) );
  XNOR U2131 ( .A(n2126), .B(n2118), .Z(n2144) );
  XOR U2132 ( .A(n2150), .B(n2151), .Z(n2118) );
  AND U2133 ( .A(n2152), .B(n2153), .Z(n2151) );
  XOR U2134 ( .A(n2150), .B(n2154), .Z(n2152) );
  XNOR U2135 ( .A(n2155), .B(n2123), .Z(n2126) );
  XOR U2136 ( .A(n2156), .B(n2157), .Z(n2123) );
  AND U2137 ( .A(n2158), .B(n2159), .Z(n2157) );
  XNOR U2138 ( .A(n2160), .B(n2161), .Z(n2158) );
  IV U2139 ( .A(n2156), .Z(n2160) );
  XNOR U2140 ( .A(n2162), .B(n2163), .Z(n2155) );
  NOR U2141 ( .A(n2164), .B(n2165), .Z(n2163) );
  XNOR U2142 ( .A(n2162), .B(n2166), .Z(n2164) );
  XNOR U2143 ( .A(n2122), .B(n2129), .Z(n2143) );
  NOR U2144 ( .A(n2088), .B(n2167), .Z(n2129) );
  XOR U2145 ( .A(n2134), .B(n2133), .Z(n2122) );
  XNOR U2146 ( .A(n2168), .B(n2130), .Z(n2133) );
  XOR U2147 ( .A(n2169), .B(n2170), .Z(n2130) );
  AND U2148 ( .A(n2171), .B(n2172), .Z(n2170) );
  XNOR U2149 ( .A(n2173), .B(n2174), .Z(n2171) );
  IV U2150 ( .A(n2169), .Z(n2173) );
  XNOR U2151 ( .A(n2175), .B(n2176), .Z(n2168) );
  NOR U2152 ( .A(n2177), .B(n2178), .Z(n2176) );
  XNOR U2153 ( .A(n2175), .B(n2179), .Z(n2177) );
  XOR U2154 ( .A(n2180), .B(n2181), .Z(n2134) );
  NOR U2155 ( .A(n2182), .B(n2183), .Z(n2181) );
  XNOR U2156 ( .A(n2180), .B(n2184), .Z(n2182) );
  XNOR U2157 ( .A(n2072), .B(n2139), .Z(n2141) );
  XOR U2158 ( .A(n2185), .B(n2186), .Z(n2072) );
  AND U2159 ( .A(n55), .B(n2187), .Z(n2186) );
  XOR U2160 ( .A(n2188), .B(n2185), .Z(n2187) );
  AND U2161 ( .A(n2085), .B(n2088), .Z(n2139) );
  XOR U2162 ( .A(n2189), .B(n2167), .Z(n2088) );
  XNOR U2163 ( .A(p_input[192]), .B(p_input[256]), .Z(n2167) );
  XNOR U2164 ( .A(n2154), .B(n2153), .Z(n2189) );
  XNOR U2165 ( .A(n2190), .B(n2161), .Z(n2153) );
  XNOR U2166 ( .A(n2149), .B(n2148), .Z(n2161) );
  XNOR U2167 ( .A(n2191), .B(n2145), .Z(n2148) );
  XNOR U2168 ( .A(p_input[202]), .B(p_input[266]), .Z(n2145) );
  XOR U2169 ( .A(p_input[203]), .B(n831), .Z(n2191) );
  XOR U2170 ( .A(p_input[204]), .B(p_input[268]), .Z(n2149) );
  XOR U2171 ( .A(n2159), .B(n2192), .Z(n2190) );
  IV U2172 ( .A(n2150), .Z(n2192) );
  XOR U2173 ( .A(p_input[193]), .B(p_input[257]), .Z(n2150) );
  XNOR U2174 ( .A(n2193), .B(n2166), .Z(n2159) );
  XNOR U2175 ( .A(p_input[207]), .B(n834), .Z(n2166) );
  XOR U2176 ( .A(n2156), .B(n2165), .Z(n2193) );
  XOR U2177 ( .A(n2194), .B(n2162), .Z(n2165) );
  XOR U2178 ( .A(p_input[205]), .B(p_input[269]), .Z(n2162) );
  XOR U2179 ( .A(p_input[206]), .B(n836), .Z(n2194) );
  XOR U2180 ( .A(p_input[201]), .B(p_input[265]), .Z(n2156) );
  XOR U2181 ( .A(n2174), .B(n2172), .Z(n2154) );
  XNOR U2182 ( .A(n2195), .B(n2179), .Z(n2172) );
  XOR U2183 ( .A(p_input[200]), .B(p_input[264]), .Z(n2179) );
  XOR U2184 ( .A(n2169), .B(n2178), .Z(n2195) );
  XOR U2185 ( .A(n2196), .B(n2175), .Z(n2178) );
  XOR U2186 ( .A(p_input[198]), .B(p_input[262]), .Z(n2175) );
  XOR U2187 ( .A(p_input[199]), .B(n958), .Z(n2196) );
  XOR U2188 ( .A(p_input[194]), .B(p_input[258]), .Z(n2169) );
  XNOR U2189 ( .A(n2184), .B(n2183), .Z(n2174) );
  XOR U2190 ( .A(n2197), .B(n2180), .Z(n2183) );
  XOR U2191 ( .A(p_input[195]), .B(p_input[259]), .Z(n2180) );
  XOR U2192 ( .A(p_input[196]), .B(n960), .Z(n2197) );
  XOR U2193 ( .A(p_input[197]), .B(p_input[261]), .Z(n2184) );
  XOR U2194 ( .A(n2198), .B(n2199), .Z(n2085) );
  AND U2195 ( .A(n55), .B(n2200), .Z(n2199) );
  XNOR U2196 ( .A(n2201), .B(n2198), .Z(n2200) );
  XNOR U2197 ( .A(n2202), .B(n2203), .Z(n55) );
  NOR U2198 ( .A(n2204), .B(n2205), .Z(n2203) );
  XOR U2199 ( .A(n2094), .B(n2202), .Z(n2205) );
  AND U2200 ( .A(n2206), .B(n2207), .Z(n2094) );
  NOR U2201 ( .A(n2202), .B(n2093), .Z(n2204) );
  AND U2202 ( .A(n2208), .B(n2209), .Z(n2093) );
  XOR U2203 ( .A(n2210), .B(n2211), .Z(n2202) );
  AND U2204 ( .A(n2212), .B(n2213), .Z(n2211) );
  XNOR U2205 ( .A(n2210), .B(n2208), .Z(n2213) );
  IV U2206 ( .A(n2111), .Z(n2208) );
  XOR U2207 ( .A(n2214), .B(n2215), .Z(n2111) );
  XOR U2208 ( .A(n2216), .B(n2209), .Z(n2215) );
  AND U2209 ( .A(n2138), .B(n2217), .Z(n2209) );
  AND U2210 ( .A(n2218), .B(n2219), .Z(n2216) );
  XOR U2211 ( .A(n2220), .B(n2214), .Z(n2218) );
  XNOR U2212 ( .A(n2108), .B(n2210), .Z(n2212) );
  XNOR U2213 ( .A(n2221), .B(n2222), .Z(n2108) );
  AND U2214 ( .A(n58), .B(n2223), .Z(n2222) );
  XNOR U2215 ( .A(n2224), .B(n2221), .Z(n2223) );
  XOR U2216 ( .A(n2225), .B(n2226), .Z(n2210) );
  AND U2217 ( .A(n2227), .B(n2228), .Z(n2226) );
  XNOR U2218 ( .A(n2225), .B(n2138), .Z(n2228) );
  XOR U2219 ( .A(n2229), .B(n2219), .Z(n2138) );
  XNOR U2220 ( .A(n2230), .B(n2214), .Z(n2219) );
  XOR U2221 ( .A(n2231), .B(n2232), .Z(n2214) );
  AND U2222 ( .A(n2233), .B(n2234), .Z(n2232) );
  XOR U2223 ( .A(n2235), .B(n2231), .Z(n2233) );
  XNOR U2224 ( .A(n2236), .B(n2237), .Z(n2230) );
  AND U2225 ( .A(n2238), .B(n2239), .Z(n2237) );
  XOR U2226 ( .A(n2236), .B(n2240), .Z(n2238) );
  XNOR U2227 ( .A(n2220), .B(n2217), .Z(n2229) );
  AND U2228 ( .A(n2241), .B(n2242), .Z(n2217) );
  XOR U2229 ( .A(n2243), .B(n2244), .Z(n2220) );
  AND U2230 ( .A(n2245), .B(n2246), .Z(n2244) );
  XOR U2231 ( .A(n2243), .B(n2247), .Z(n2245) );
  XNOR U2232 ( .A(n2135), .B(n2225), .Z(n2227) );
  XNOR U2233 ( .A(n2248), .B(n2249), .Z(n2135) );
  AND U2234 ( .A(n58), .B(n2250), .Z(n2249) );
  XOR U2235 ( .A(n2251), .B(n2248), .Z(n2250) );
  XOR U2236 ( .A(n2252), .B(n2253), .Z(n2225) );
  AND U2237 ( .A(n2254), .B(n2255), .Z(n2253) );
  XNOR U2238 ( .A(n2252), .B(n2241), .Z(n2255) );
  IV U2239 ( .A(n2188), .Z(n2241) );
  XNOR U2240 ( .A(n2256), .B(n2234), .Z(n2188) );
  XNOR U2241 ( .A(n2257), .B(n2240), .Z(n2234) );
  XNOR U2242 ( .A(n2258), .B(n2259), .Z(n2240) );
  NOR U2243 ( .A(n2260), .B(n2261), .Z(n2259) );
  XOR U2244 ( .A(n2258), .B(n2262), .Z(n2260) );
  XNOR U2245 ( .A(n2239), .B(n2231), .Z(n2257) );
  XOR U2246 ( .A(n2263), .B(n2264), .Z(n2231) );
  AND U2247 ( .A(n2265), .B(n2266), .Z(n2264) );
  XOR U2248 ( .A(n2263), .B(n2267), .Z(n2265) );
  XNOR U2249 ( .A(n2268), .B(n2236), .Z(n2239) );
  XOR U2250 ( .A(n2269), .B(n2270), .Z(n2236) );
  AND U2251 ( .A(n2271), .B(n2272), .Z(n2270) );
  XNOR U2252 ( .A(n2273), .B(n2274), .Z(n2271) );
  IV U2253 ( .A(n2269), .Z(n2273) );
  XNOR U2254 ( .A(n2275), .B(n2276), .Z(n2268) );
  NOR U2255 ( .A(n2277), .B(n2278), .Z(n2276) );
  XNOR U2256 ( .A(n2275), .B(n2279), .Z(n2277) );
  XNOR U2257 ( .A(n2235), .B(n2242), .Z(n2256) );
  NOR U2258 ( .A(n2201), .B(n2280), .Z(n2242) );
  XOR U2259 ( .A(n2247), .B(n2246), .Z(n2235) );
  XNOR U2260 ( .A(n2281), .B(n2243), .Z(n2246) );
  XOR U2261 ( .A(n2282), .B(n2283), .Z(n2243) );
  AND U2262 ( .A(n2284), .B(n2285), .Z(n2283) );
  XNOR U2263 ( .A(n2286), .B(n2287), .Z(n2284) );
  IV U2264 ( .A(n2282), .Z(n2286) );
  XNOR U2265 ( .A(n2288), .B(n2289), .Z(n2281) );
  NOR U2266 ( .A(n2290), .B(n2291), .Z(n2289) );
  XNOR U2267 ( .A(n2288), .B(n2292), .Z(n2290) );
  XOR U2268 ( .A(n2293), .B(n2294), .Z(n2247) );
  NOR U2269 ( .A(n2295), .B(n2296), .Z(n2294) );
  XNOR U2270 ( .A(n2293), .B(n2297), .Z(n2295) );
  XNOR U2271 ( .A(n2185), .B(n2252), .Z(n2254) );
  XNOR U2272 ( .A(n2298), .B(n2299), .Z(n2185) );
  AND U2273 ( .A(n58), .B(n2300), .Z(n2299) );
  XNOR U2274 ( .A(n2301), .B(n2298), .Z(n2300) );
  AND U2275 ( .A(n2198), .B(n2201), .Z(n2252) );
  XOR U2276 ( .A(n2302), .B(n2280), .Z(n2201) );
  XNOR U2277 ( .A(p_input[208]), .B(p_input[256]), .Z(n2280) );
  XNOR U2278 ( .A(n2267), .B(n2266), .Z(n2302) );
  XNOR U2279 ( .A(n2303), .B(n2274), .Z(n2266) );
  XNOR U2280 ( .A(n2262), .B(n2261), .Z(n2274) );
  XNOR U2281 ( .A(n2304), .B(n2258), .Z(n2261) );
  XNOR U2282 ( .A(p_input[218]), .B(p_input[266]), .Z(n2258) );
  XOR U2283 ( .A(p_input[219]), .B(n831), .Z(n2304) );
  XOR U2284 ( .A(p_input[220]), .B(p_input[268]), .Z(n2262) );
  XOR U2285 ( .A(n2272), .B(n2305), .Z(n2303) );
  IV U2286 ( .A(n2263), .Z(n2305) );
  XOR U2287 ( .A(p_input[209]), .B(p_input[257]), .Z(n2263) );
  XNOR U2288 ( .A(n2306), .B(n2279), .Z(n2272) );
  XNOR U2289 ( .A(p_input[223]), .B(n834), .Z(n2279) );
  XOR U2290 ( .A(n2269), .B(n2278), .Z(n2306) );
  XOR U2291 ( .A(n2307), .B(n2275), .Z(n2278) );
  XOR U2292 ( .A(p_input[221]), .B(p_input[269]), .Z(n2275) );
  XOR U2293 ( .A(p_input[222]), .B(n836), .Z(n2307) );
  XOR U2294 ( .A(p_input[217]), .B(p_input[265]), .Z(n2269) );
  XOR U2295 ( .A(n2287), .B(n2285), .Z(n2267) );
  XNOR U2296 ( .A(n2308), .B(n2292), .Z(n2285) );
  XOR U2297 ( .A(p_input[216]), .B(p_input[264]), .Z(n2292) );
  XOR U2298 ( .A(n2282), .B(n2291), .Z(n2308) );
  XOR U2299 ( .A(n2309), .B(n2288), .Z(n2291) );
  XOR U2300 ( .A(p_input[214]), .B(p_input[262]), .Z(n2288) );
  XOR U2301 ( .A(p_input[215]), .B(n958), .Z(n2309) );
  XOR U2302 ( .A(p_input[210]), .B(p_input[258]), .Z(n2282) );
  XNOR U2303 ( .A(n2297), .B(n2296), .Z(n2287) );
  XOR U2304 ( .A(n2310), .B(n2293), .Z(n2296) );
  XOR U2305 ( .A(p_input[211]), .B(p_input[259]), .Z(n2293) );
  XOR U2306 ( .A(p_input[212]), .B(n960), .Z(n2310) );
  XOR U2307 ( .A(p_input[213]), .B(p_input[261]), .Z(n2297) );
  XOR U2308 ( .A(n2311), .B(n2312), .Z(n2198) );
  AND U2309 ( .A(n58), .B(n2313), .Z(n2312) );
  XNOR U2310 ( .A(n2314), .B(n2311), .Z(n2313) );
  XNOR U2311 ( .A(n2315), .B(n2316), .Z(n58) );
  NOR U2312 ( .A(n2317), .B(n2318), .Z(n2316) );
  XOR U2313 ( .A(n2207), .B(n2315), .Z(n2318) );
  AND U2314 ( .A(n2221), .B(n2319), .Z(n2207) );
  NOR U2315 ( .A(n2315), .B(n2206), .Z(n2317) );
  AND U2316 ( .A(n2320), .B(n2321), .Z(n2206) );
  XOR U2317 ( .A(n2322), .B(n2323), .Z(n2315) );
  AND U2318 ( .A(n2324), .B(n2325), .Z(n2323) );
  XNOR U2319 ( .A(n2322), .B(n2320), .Z(n2325) );
  IV U2320 ( .A(n2224), .Z(n2320) );
  XOR U2321 ( .A(n2326), .B(n2327), .Z(n2224) );
  XOR U2322 ( .A(n2328), .B(n2321), .Z(n2327) );
  AND U2323 ( .A(n2251), .B(n2329), .Z(n2321) );
  AND U2324 ( .A(n2330), .B(n2331), .Z(n2328) );
  XOR U2325 ( .A(n2332), .B(n2326), .Z(n2330) );
  XNOR U2326 ( .A(n2333), .B(n2322), .Z(n2324) );
  IV U2327 ( .A(n2221), .Z(n2333) );
  XNOR U2328 ( .A(n2334), .B(n2335), .Z(n2221) );
  XOR U2329 ( .A(n2336), .B(n2319), .Z(n2335) );
  AND U2330 ( .A(n2248), .B(n2337), .Z(n2319) );
  AND U2331 ( .A(n2338), .B(n2339), .Z(n2336) );
  XNOR U2332 ( .A(n2334), .B(n2340), .Z(n2338) );
  XOR U2333 ( .A(n2341), .B(n2342), .Z(n2322) );
  AND U2334 ( .A(n2343), .B(n2344), .Z(n2342) );
  XNOR U2335 ( .A(n2341), .B(n2251), .Z(n2344) );
  XOR U2336 ( .A(n2345), .B(n2331), .Z(n2251) );
  XNOR U2337 ( .A(n2346), .B(n2326), .Z(n2331) );
  XOR U2338 ( .A(n2347), .B(n2348), .Z(n2326) );
  AND U2339 ( .A(n2349), .B(n2350), .Z(n2348) );
  XOR U2340 ( .A(n2351), .B(n2347), .Z(n2349) );
  XNOR U2341 ( .A(n2352), .B(n2353), .Z(n2346) );
  AND U2342 ( .A(n2354), .B(n2355), .Z(n2353) );
  XOR U2343 ( .A(n2352), .B(n2356), .Z(n2354) );
  XNOR U2344 ( .A(n2332), .B(n2329), .Z(n2345) );
  AND U2345 ( .A(n2357), .B(n2358), .Z(n2329) );
  XOR U2346 ( .A(n2359), .B(n2360), .Z(n2332) );
  AND U2347 ( .A(n2361), .B(n2362), .Z(n2360) );
  XOR U2348 ( .A(n2359), .B(n2363), .Z(n2361) );
  XOR U2349 ( .A(n2248), .B(n2341), .Z(n2343) );
  XNOR U2350 ( .A(n2364), .B(n2340), .Z(n2248) );
  XNOR U2351 ( .A(n2365), .B(n2366), .Z(n2340) );
  AND U2352 ( .A(n2367), .B(n2368), .Z(n2366) );
  XOR U2353 ( .A(n2365), .B(n2369), .Z(n2367) );
  XNOR U2354 ( .A(n2339), .B(n2337), .Z(n2364) );
  AND U2355 ( .A(n2298), .B(n2370), .Z(n2337) );
  XNOR U2356 ( .A(n2371), .B(n2334), .Z(n2339) );
  XOR U2357 ( .A(n2372), .B(n2373), .Z(n2334) );
  AND U2358 ( .A(n2374), .B(n2375), .Z(n2373) );
  XOR U2359 ( .A(n2372), .B(n2376), .Z(n2374) );
  XNOR U2360 ( .A(n2377), .B(n2378), .Z(n2371) );
  AND U2361 ( .A(n2379), .B(n2380), .Z(n2378) );
  XNOR U2362 ( .A(n2377), .B(n2381), .Z(n2379) );
  XOR U2363 ( .A(n2382), .B(n2383), .Z(n2341) );
  AND U2364 ( .A(n2384), .B(n2385), .Z(n2383) );
  XNOR U2365 ( .A(n2382), .B(n2357), .Z(n2385) );
  IV U2366 ( .A(n2301), .Z(n2357) );
  XNOR U2367 ( .A(n2386), .B(n2350), .Z(n2301) );
  XNOR U2368 ( .A(n2387), .B(n2356), .Z(n2350) );
  XNOR U2369 ( .A(n2388), .B(n2389), .Z(n2356) );
  NOR U2370 ( .A(n2390), .B(n2391), .Z(n2389) );
  XOR U2371 ( .A(n2388), .B(n2392), .Z(n2390) );
  XNOR U2372 ( .A(n2355), .B(n2347), .Z(n2387) );
  XOR U2373 ( .A(n2393), .B(n2394), .Z(n2347) );
  AND U2374 ( .A(n2395), .B(n2396), .Z(n2394) );
  XOR U2375 ( .A(n2393), .B(n2397), .Z(n2395) );
  XNOR U2376 ( .A(n2398), .B(n2352), .Z(n2355) );
  XOR U2377 ( .A(n2399), .B(n2400), .Z(n2352) );
  AND U2378 ( .A(n2401), .B(n2402), .Z(n2400) );
  XNOR U2379 ( .A(n2403), .B(n2404), .Z(n2401) );
  IV U2380 ( .A(n2399), .Z(n2403) );
  XNOR U2381 ( .A(n2405), .B(n2406), .Z(n2398) );
  NOR U2382 ( .A(n2407), .B(n2408), .Z(n2406) );
  XNOR U2383 ( .A(n2405), .B(n2409), .Z(n2407) );
  XNOR U2384 ( .A(n2351), .B(n2358), .Z(n2386) );
  NOR U2385 ( .A(n2314), .B(n2410), .Z(n2358) );
  XOR U2386 ( .A(n2363), .B(n2362), .Z(n2351) );
  XNOR U2387 ( .A(n2411), .B(n2359), .Z(n2362) );
  XOR U2388 ( .A(n2412), .B(n2413), .Z(n2359) );
  AND U2389 ( .A(n2414), .B(n2415), .Z(n2413) );
  XNOR U2390 ( .A(n2416), .B(n2417), .Z(n2414) );
  IV U2391 ( .A(n2412), .Z(n2416) );
  XNOR U2392 ( .A(n2418), .B(n2419), .Z(n2411) );
  NOR U2393 ( .A(n2420), .B(n2421), .Z(n2419) );
  XNOR U2394 ( .A(n2418), .B(n2422), .Z(n2420) );
  XOR U2395 ( .A(n2423), .B(n2424), .Z(n2363) );
  NOR U2396 ( .A(n2425), .B(n2426), .Z(n2424) );
  XNOR U2397 ( .A(n2423), .B(n2427), .Z(n2425) );
  XNOR U2398 ( .A(n2428), .B(n2382), .Z(n2384) );
  IV U2399 ( .A(n2298), .Z(n2428) );
  XOR U2400 ( .A(n2429), .B(n2376), .Z(n2298) );
  XOR U2401 ( .A(n2369), .B(n2368), .Z(n2376) );
  XNOR U2402 ( .A(n2430), .B(n2365), .Z(n2368) );
  XOR U2403 ( .A(n2431), .B(n2432), .Z(n2365) );
  AND U2404 ( .A(n2433), .B(n2434), .Z(n2432) );
  XOR U2405 ( .A(n2431), .B(n2435), .Z(n2433) );
  XNOR U2406 ( .A(n2436), .B(n2437), .Z(n2430) );
  NOR U2407 ( .A(n2438), .B(n2439), .Z(n2437) );
  XNOR U2408 ( .A(n2436), .B(n2440), .Z(n2438) );
  XOR U2409 ( .A(n2441), .B(n2442), .Z(n2369) );
  NOR U2410 ( .A(n2443), .B(n2444), .Z(n2442) );
  XNOR U2411 ( .A(n2441), .B(n2445), .Z(n2443) );
  XNOR U2412 ( .A(n2375), .B(n2370), .Z(n2429) );
  AND U2413 ( .A(n2311), .B(n2446), .Z(n2370) );
  XOR U2414 ( .A(n2447), .B(n2381), .Z(n2375) );
  XNOR U2415 ( .A(n2448), .B(n2449), .Z(n2381) );
  NOR U2416 ( .A(n2450), .B(n2451), .Z(n2449) );
  XNOR U2417 ( .A(n2448), .B(n2452), .Z(n2450) );
  XNOR U2418 ( .A(n2380), .B(n2372), .Z(n2447) );
  XOR U2419 ( .A(n2453), .B(n2454), .Z(n2372) );
  AND U2420 ( .A(n2455), .B(n2456), .Z(n2454) );
  XOR U2421 ( .A(n2453), .B(n2457), .Z(n2455) );
  XNOR U2422 ( .A(n2458), .B(n2377), .Z(n2380) );
  XOR U2423 ( .A(n2459), .B(n2460), .Z(n2377) );
  AND U2424 ( .A(n2461), .B(n2462), .Z(n2460) );
  XOR U2425 ( .A(n2459), .B(n2463), .Z(n2461) );
  XNOR U2426 ( .A(n2464), .B(n2465), .Z(n2458) );
  NOR U2427 ( .A(n2466), .B(n2467), .Z(n2465) );
  XOR U2428 ( .A(n2464), .B(n2468), .Z(n2466) );
  AND U2429 ( .A(n2311), .B(n2314), .Z(n2382) );
  XOR U2430 ( .A(n2469), .B(n2410), .Z(n2314) );
  XNOR U2431 ( .A(p_input[224]), .B(p_input[256]), .Z(n2410) );
  XNOR U2432 ( .A(n2397), .B(n2396), .Z(n2469) );
  XNOR U2433 ( .A(n2470), .B(n2404), .Z(n2396) );
  XNOR U2434 ( .A(n2392), .B(n2391), .Z(n2404) );
  XNOR U2435 ( .A(n2471), .B(n2388), .Z(n2391) );
  XNOR U2436 ( .A(p_input[234]), .B(p_input[266]), .Z(n2388) );
  XOR U2437 ( .A(p_input[235]), .B(n831), .Z(n2471) );
  XOR U2438 ( .A(p_input[236]), .B(p_input[268]), .Z(n2392) );
  XOR U2439 ( .A(n2402), .B(n2472), .Z(n2470) );
  IV U2440 ( .A(n2393), .Z(n2472) );
  XOR U2441 ( .A(p_input[225]), .B(p_input[257]), .Z(n2393) );
  XNOR U2442 ( .A(n2473), .B(n2409), .Z(n2402) );
  XNOR U2443 ( .A(p_input[239]), .B(n834), .Z(n2409) );
  IV U2444 ( .A(p_input[271]), .Z(n834) );
  XOR U2445 ( .A(n2399), .B(n2408), .Z(n2473) );
  XOR U2446 ( .A(n2474), .B(n2405), .Z(n2408) );
  XOR U2447 ( .A(p_input[237]), .B(p_input[269]), .Z(n2405) );
  XOR U2448 ( .A(p_input[238]), .B(n836), .Z(n2474) );
  XOR U2449 ( .A(p_input[233]), .B(p_input[265]), .Z(n2399) );
  XOR U2450 ( .A(n2417), .B(n2415), .Z(n2397) );
  XNOR U2451 ( .A(n2475), .B(n2422), .Z(n2415) );
  XOR U2452 ( .A(p_input[232]), .B(p_input[264]), .Z(n2422) );
  XOR U2453 ( .A(n2412), .B(n2421), .Z(n2475) );
  XOR U2454 ( .A(n2476), .B(n2418), .Z(n2421) );
  XOR U2455 ( .A(p_input[230]), .B(p_input[262]), .Z(n2418) );
  XOR U2456 ( .A(p_input[231]), .B(n958), .Z(n2476) );
  XOR U2457 ( .A(p_input[226]), .B(p_input[258]), .Z(n2412) );
  XNOR U2458 ( .A(n2427), .B(n2426), .Z(n2417) );
  XOR U2459 ( .A(n2477), .B(n2423), .Z(n2426) );
  XOR U2460 ( .A(p_input[227]), .B(p_input[259]), .Z(n2423) );
  XOR U2461 ( .A(p_input[228]), .B(n960), .Z(n2477) );
  XOR U2462 ( .A(p_input[229]), .B(p_input[261]), .Z(n2427) );
  XOR U2463 ( .A(n2478), .B(n2457), .Z(n2311) );
  XOR U2464 ( .A(n2435), .B(n2434), .Z(n2457) );
  XNOR U2465 ( .A(n2479), .B(n2440), .Z(n2434) );
  XOR U2466 ( .A(\knn_comb_/min_val_out[0][8] ), .B(p_input[264]), .Z(n2440)
         );
  XOR U2467 ( .A(n2431), .B(n2439), .Z(n2479) );
  XOR U2468 ( .A(n2480), .B(n2436), .Z(n2439) );
  XOR U2469 ( .A(\knn_comb_/min_val_out[0][6] ), .B(p_input[262]), .Z(n2436)
         );
  XOR U2470 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n958), .Z(n2480) );
  IV U2471 ( .A(p_input[263]), .Z(n958) );
  XNOR U2472 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n840), .Z(n2431) );
  IV U2473 ( .A(p_input[258]), .Z(n840) );
  XNOR U2474 ( .A(n2445), .B(n2444), .Z(n2435) );
  XOR U2475 ( .A(n2481), .B(n2441), .Z(n2444) );
  XOR U2476 ( .A(\knn_comb_/min_val_out[0][3] ), .B(p_input[259]), .Z(n2441)
         );
  XOR U2477 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n960), .Z(n2481) );
  IV U2478 ( .A(p_input[260]), .Z(n960) );
  XOR U2479 ( .A(\knn_comb_/min_val_out[0][5] ), .B(p_input[261]), .Z(n2445)
         );
  XNOR U2480 ( .A(n2456), .B(n2446), .Z(n2478) );
  XOR U2481 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[256]), .Z(n2446)
         );
  XNOR U2482 ( .A(n2482), .B(n2463), .Z(n2456) );
  XNOR U2483 ( .A(n2452), .B(n2451), .Z(n2463) );
  XOR U2484 ( .A(n2483), .B(n2448), .Z(n2451) );
  XNOR U2485 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n952), .Z(n2448) );
  IV U2486 ( .A(p_input[266]), .Z(n952) );
  XOR U2487 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n831), .Z(n2483) );
  IV U2488 ( .A(p_input[267]), .Z(n831) );
  XOR U2489 ( .A(\knn_comb_/min_val_out[0][12] ), .B(p_input[268]), .Z(n2452)
         );
  XNOR U2490 ( .A(n2462), .B(n2453), .Z(n2482) );
  XNOR U2491 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n1068), .Z(n2453) );
  IV U2492 ( .A(p_input[257]), .Z(n1068) );
  XOR U2493 ( .A(n2484), .B(n2468), .Z(n2462) );
  XNOR U2494 ( .A(\knn_comb_/min_val_out[0][15] ), .B(p_input[271]), .Z(n2468)
         );
  XOR U2495 ( .A(n2459), .B(n2467), .Z(n2484) );
  XOR U2496 ( .A(n2485), .B(n2464), .Z(n2467) );
  XOR U2497 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[269]), .Z(n2464)
         );
  XOR U2498 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n836), .Z(n2485) );
  IV U2499 ( .A(p_input[270]), .Z(n836) );
  XNOR U2500 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n837), .Z(n2459) );
  IV U2501 ( .A(p_input[265]), .Z(n837) );
endmodule

