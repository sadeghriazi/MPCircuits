
module knn_comb_BMR_W16_K1_N64 ( p_input, o );
  input [1039:0] p_input;
  output [15:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180;
  assign \knn_comb_/min_val_out[0][0]  = p_input[1008];
  assign \knn_comb_/min_val_out[0][1]  = p_input[1009];
  assign \knn_comb_/min_val_out[0][2]  = p_input[1010];
  assign \knn_comb_/min_val_out[0][3]  = p_input[1011];
  assign \knn_comb_/min_val_out[0][4]  = p_input[1012];
  assign \knn_comb_/min_val_out[0][5]  = p_input[1013];
  assign \knn_comb_/min_val_out[0][6]  = p_input[1014];
  assign \knn_comb_/min_val_out[0][7]  = p_input[1015];
  assign \knn_comb_/min_val_out[0][8]  = p_input[1016];
  assign \knn_comb_/min_val_out[0][9]  = p_input[1017];
  assign \knn_comb_/min_val_out[0][10]  = p_input[1018];
  assign \knn_comb_/min_val_out[0][11]  = p_input[1019];
  assign \knn_comb_/min_val_out[0][12]  = p_input[1020];
  assign \knn_comb_/min_val_out[0][13]  = p_input[1021];
  assign \knn_comb_/min_val_out[0][14]  = p_input[1022];
  assign \knn_comb_/min_val_out[0][15]  = p_input[1023];

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(n3), .B(n4), .Z(n1) );
  XNOR U3 ( .A(p_input[9]), .B(n2), .Z(n4) );
  XOR U4 ( .A(n5), .B(n6), .Z(n2) );
  AND U5 ( .A(n7), .B(n8), .Z(n6) );
  XNOR U6 ( .A(p_input[25]), .B(n5), .Z(n8) );
  XOR U7 ( .A(n9), .B(n10), .Z(n5) );
  AND U8 ( .A(n11), .B(n12), .Z(n10) );
  XNOR U9 ( .A(p_input[41]), .B(n9), .Z(n12) );
  XOR U10 ( .A(n13), .B(n14), .Z(n9) );
  AND U11 ( .A(n15), .B(n16), .Z(n14) );
  XNOR U12 ( .A(p_input[57]), .B(n13), .Z(n16) );
  XOR U13 ( .A(n17), .B(n18), .Z(n13) );
  AND U14 ( .A(n19), .B(n20), .Z(n18) );
  XNOR U15 ( .A(p_input[73]), .B(n17), .Z(n20) );
  XOR U16 ( .A(n21), .B(n22), .Z(n17) );
  AND U17 ( .A(n23), .B(n24), .Z(n22) );
  XNOR U18 ( .A(p_input[89]), .B(n21), .Z(n24) );
  XOR U19 ( .A(n25), .B(n26), .Z(n21) );
  AND U20 ( .A(n27), .B(n28), .Z(n26) );
  XNOR U21 ( .A(p_input[105]), .B(n25), .Z(n28) );
  XOR U22 ( .A(n29), .B(n30), .Z(n25) );
  AND U23 ( .A(n31), .B(n32), .Z(n30) );
  XNOR U24 ( .A(p_input[121]), .B(n29), .Z(n32) );
  XOR U25 ( .A(n33), .B(n34), .Z(n29) );
  AND U26 ( .A(n35), .B(n36), .Z(n34) );
  XNOR U27 ( .A(p_input[137]), .B(n33), .Z(n36) );
  XOR U28 ( .A(n37), .B(n38), .Z(n33) );
  AND U29 ( .A(n39), .B(n40), .Z(n38) );
  XNOR U30 ( .A(p_input[153]), .B(n37), .Z(n40) );
  XOR U31 ( .A(n41), .B(n42), .Z(n37) );
  AND U32 ( .A(n43), .B(n44), .Z(n42) );
  XNOR U33 ( .A(p_input[169]), .B(n41), .Z(n44) );
  XOR U34 ( .A(n45), .B(n46), .Z(n41) );
  AND U35 ( .A(n47), .B(n48), .Z(n46) );
  XNOR U36 ( .A(p_input[185]), .B(n45), .Z(n48) );
  XOR U37 ( .A(n49), .B(n50), .Z(n45) );
  AND U38 ( .A(n51), .B(n52), .Z(n50) );
  XNOR U39 ( .A(p_input[201]), .B(n49), .Z(n52) );
  XOR U40 ( .A(n53), .B(n54), .Z(n49) );
  AND U41 ( .A(n55), .B(n56), .Z(n54) );
  XNOR U42 ( .A(p_input[217]), .B(n53), .Z(n56) );
  XOR U43 ( .A(n57), .B(n58), .Z(n53) );
  AND U44 ( .A(n59), .B(n60), .Z(n58) );
  XNOR U45 ( .A(p_input[233]), .B(n57), .Z(n60) );
  XOR U46 ( .A(n61), .B(n62), .Z(n57) );
  AND U47 ( .A(n63), .B(n64), .Z(n62) );
  XNOR U48 ( .A(p_input[249]), .B(n61), .Z(n64) );
  XOR U49 ( .A(n65), .B(n66), .Z(n61) );
  AND U50 ( .A(n67), .B(n68), .Z(n66) );
  XNOR U51 ( .A(p_input[265]), .B(n65), .Z(n68) );
  XOR U52 ( .A(n69), .B(n70), .Z(n65) );
  AND U53 ( .A(n71), .B(n72), .Z(n70) );
  XNOR U54 ( .A(p_input[281]), .B(n69), .Z(n72) );
  XOR U55 ( .A(n73), .B(n74), .Z(n69) );
  AND U56 ( .A(n75), .B(n76), .Z(n74) );
  XNOR U57 ( .A(p_input[297]), .B(n73), .Z(n76) );
  XOR U58 ( .A(n77), .B(n78), .Z(n73) );
  AND U59 ( .A(n79), .B(n80), .Z(n78) );
  XNOR U60 ( .A(p_input[313]), .B(n77), .Z(n80) );
  XOR U61 ( .A(n81), .B(n82), .Z(n77) );
  AND U62 ( .A(n83), .B(n84), .Z(n82) );
  XNOR U63 ( .A(p_input[329]), .B(n81), .Z(n84) );
  XOR U64 ( .A(n85), .B(n86), .Z(n81) );
  AND U65 ( .A(n87), .B(n88), .Z(n86) );
  XNOR U66 ( .A(p_input[345]), .B(n85), .Z(n88) );
  XOR U67 ( .A(n89), .B(n90), .Z(n85) );
  AND U68 ( .A(n91), .B(n92), .Z(n90) );
  XNOR U69 ( .A(p_input[361]), .B(n89), .Z(n92) );
  XOR U70 ( .A(n93), .B(n94), .Z(n89) );
  AND U71 ( .A(n95), .B(n96), .Z(n94) );
  XNOR U72 ( .A(p_input[377]), .B(n93), .Z(n96) );
  XOR U73 ( .A(n97), .B(n98), .Z(n93) );
  AND U74 ( .A(n99), .B(n100), .Z(n98) );
  XNOR U75 ( .A(p_input[393]), .B(n97), .Z(n100) );
  XOR U76 ( .A(n101), .B(n102), .Z(n97) );
  AND U77 ( .A(n103), .B(n104), .Z(n102) );
  XNOR U78 ( .A(p_input[409]), .B(n101), .Z(n104) );
  XOR U79 ( .A(n105), .B(n106), .Z(n101) );
  AND U80 ( .A(n107), .B(n108), .Z(n106) );
  XNOR U81 ( .A(p_input[425]), .B(n105), .Z(n108) );
  XOR U82 ( .A(n109), .B(n110), .Z(n105) );
  AND U83 ( .A(n111), .B(n112), .Z(n110) );
  XNOR U84 ( .A(p_input[441]), .B(n109), .Z(n112) );
  XOR U85 ( .A(n113), .B(n114), .Z(n109) );
  AND U86 ( .A(n115), .B(n116), .Z(n114) );
  XNOR U87 ( .A(p_input[457]), .B(n113), .Z(n116) );
  XOR U88 ( .A(n117), .B(n118), .Z(n113) );
  AND U89 ( .A(n119), .B(n120), .Z(n118) );
  XNOR U90 ( .A(p_input[473]), .B(n117), .Z(n120) );
  XOR U91 ( .A(n121), .B(n122), .Z(n117) );
  AND U92 ( .A(n123), .B(n124), .Z(n122) );
  XNOR U93 ( .A(p_input[489]), .B(n121), .Z(n124) );
  XOR U94 ( .A(n125), .B(n126), .Z(n121) );
  AND U95 ( .A(n127), .B(n128), .Z(n126) );
  XNOR U96 ( .A(p_input[505]), .B(n125), .Z(n128) );
  XOR U97 ( .A(n129), .B(n130), .Z(n125) );
  AND U98 ( .A(n131), .B(n132), .Z(n130) );
  XNOR U99 ( .A(p_input[521]), .B(n129), .Z(n132) );
  XOR U100 ( .A(n133), .B(n134), .Z(n129) );
  AND U101 ( .A(n135), .B(n136), .Z(n134) );
  XNOR U102 ( .A(p_input[537]), .B(n133), .Z(n136) );
  XOR U103 ( .A(n137), .B(n138), .Z(n133) );
  AND U104 ( .A(n139), .B(n140), .Z(n138) );
  XNOR U105 ( .A(p_input[553]), .B(n137), .Z(n140) );
  XOR U106 ( .A(n141), .B(n142), .Z(n137) );
  AND U107 ( .A(n143), .B(n144), .Z(n142) );
  XNOR U108 ( .A(p_input[569]), .B(n141), .Z(n144) );
  XOR U109 ( .A(n145), .B(n146), .Z(n141) );
  AND U110 ( .A(n147), .B(n148), .Z(n146) );
  XNOR U111 ( .A(p_input[585]), .B(n145), .Z(n148) );
  XOR U112 ( .A(n149), .B(n150), .Z(n145) );
  AND U113 ( .A(n151), .B(n152), .Z(n150) );
  XNOR U114 ( .A(p_input[601]), .B(n149), .Z(n152) );
  XOR U115 ( .A(n153), .B(n154), .Z(n149) );
  AND U116 ( .A(n155), .B(n156), .Z(n154) );
  XNOR U117 ( .A(p_input[617]), .B(n153), .Z(n156) );
  XOR U118 ( .A(n157), .B(n158), .Z(n153) );
  AND U119 ( .A(n159), .B(n160), .Z(n158) );
  XNOR U120 ( .A(p_input[633]), .B(n157), .Z(n160) );
  XOR U121 ( .A(n161), .B(n162), .Z(n157) );
  AND U122 ( .A(n163), .B(n164), .Z(n162) );
  XNOR U123 ( .A(p_input[649]), .B(n161), .Z(n164) );
  XOR U124 ( .A(n165), .B(n166), .Z(n161) );
  AND U125 ( .A(n167), .B(n168), .Z(n166) );
  XNOR U126 ( .A(p_input[665]), .B(n165), .Z(n168) );
  XOR U127 ( .A(n169), .B(n170), .Z(n165) );
  AND U128 ( .A(n171), .B(n172), .Z(n170) );
  XNOR U129 ( .A(p_input[681]), .B(n169), .Z(n172) );
  XOR U130 ( .A(n173), .B(n174), .Z(n169) );
  AND U131 ( .A(n175), .B(n176), .Z(n174) );
  XNOR U132 ( .A(p_input[697]), .B(n173), .Z(n176) );
  XOR U133 ( .A(n177), .B(n178), .Z(n173) );
  AND U134 ( .A(n179), .B(n180), .Z(n178) );
  XNOR U135 ( .A(p_input[713]), .B(n177), .Z(n180) );
  XOR U136 ( .A(n181), .B(n182), .Z(n177) );
  AND U137 ( .A(n183), .B(n184), .Z(n182) );
  XNOR U138 ( .A(p_input[729]), .B(n181), .Z(n184) );
  XOR U139 ( .A(n185), .B(n186), .Z(n181) );
  AND U140 ( .A(n187), .B(n188), .Z(n186) );
  XNOR U141 ( .A(p_input[745]), .B(n185), .Z(n188) );
  XOR U142 ( .A(n189), .B(n190), .Z(n185) );
  AND U143 ( .A(n191), .B(n192), .Z(n190) );
  XNOR U144 ( .A(p_input[761]), .B(n189), .Z(n192) );
  XOR U145 ( .A(n193), .B(n194), .Z(n189) );
  AND U146 ( .A(n195), .B(n196), .Z(n194) );
  XNOR U147 ( .A(p_input[777]), .B(n193), .Z(n196) );
  XOR U148 ( .A(n197), .B(n198), .Z(n193) );
  AND U149 ( .A(n199), .B(n200), .Z(n198) );
  XNOR U150 ( .A(p_input[793]), .B(n197), .Z(n200) );
  XOR U151 ( .A(n201), .B(n202), .Z(n197) );
  AND U152 ( .A(n203), .B(n204), .Z(n202) );
  XNOR U153 ( .A(p_input[809]), .B(n201), .Z(n204) );
  XOR U154 ( .A(n205), .B(n206), .Z(n201) );
  AND U155 ( .A(n207), .B(n208), .Z(n206) );
  XNOR U156 ( .A(p_input[825]), .B(n205), .Z(n208) );
  XOR U157 ( .A(n209), .B(n210), .Z(n205) );
  AND U158 ( .A(n211), .B(n212), .Z(n210) );
  XNOR U159 ( .A(p_input[841]), .B(n209), .Z(n212) );
  XOR U160 ( .A(n213), .B(n214), .Z(n209) );
  AND U161 ( .A(n215), .B(n216), .Z(n214) );
  XNOR U162 ( .A(p_input[857]), .B(n213), .Z(n216) );
  XOR U163 ( .A(n217), .B(n218), .Z(n213) );
  AND U164 ( .A(n219), .B(n220), .Z(n218) );
  XNOR U165 ( .A(p_input[873]), .B(n217), .Z(n220) );
  XOR U166 ( .A(n221), .B(n222), .Z(n217) );
  AND U167 ( .A(n223), .B(n224), .Z(n222) );
  XNOR U168 ( .A(p_input[889]), .B(n221), .Z(n224) );
  XOR U169 ( .A(n225), .B(n226), .Z(n221) );
  AND U170 ( .A(n227), .B(n228), .Z(n226) );
  XNOR U171 ( .A(p_input[905]), .B(n225), .Z(n228) );
  XOR U172 ( .A(n229), .B(n230), .Z(n225) );
  AND U173 ( .A(n231), .B(n232), .Z(n230) );
  XNOR U174 ( .A(p_input[921]), .B(n229), .Z(n232) );
  XOR U175 ( .A(n233), .B(n234), .Z(n229) );
  AND U176 ( .A(n235), .B(n236), .Z(n234) );
  XNOR U177 ( .A(p_input[937]), .B(n233), .Z(n236) );
  XOR U178 ( .A(n237), .B(n238), .Z(n233) );
  AND U179 ( .A(n239), .B(n240), .Z(n238) );
  XNOR U180 ( .A(p_input[953]), .B(n237), .Z(n240) );
  XOR U181 ( .A(n241), .B(n242), .Z(n237) );
  AND U182 ( .A(n243), .B(n244), .Z(n242) );
  XNOR U183 ( .A(p_input[969]), .B(n241), .Z(n244) );
  XNOR U184 ( .A(n245), .B(n246), .Z(n241) );
  AND U185 ( .A(n247), .B(n248), .Z(n246) );
  XOR U186 ( .A(p_input[985]), .B(n245), .Z(n248) );
  XOR U187 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n249), .Z(n245) );
  AND U188 ( .A(n250), .B(n251), .Z(n249) );
  XOR U189 ( .A(p_input[1001]), .B(\knn_comb_/min_val_out[0][9] ), .Z(n251) );
  XNOR U190 ( .A(n252), .B(n253), .Z(o[8]) );
  AND U191 ( .A(n3), .B(n254), .Z(n252) );
  XNOR U192 ( .A(p_input[8]), .B(n253), .Z(n254) );
  XOR U193 ( .A(n255), .B(n256), .Z(n253) );
  AND U194 ( .A(n7), .B(n257), .Z(n256) );
  XNOR U195 ( .A(p_input[24]), .B(n255), .Z(n257) );
  XOR U196 ( .A(n258), .B(n259), .Z(n255) );
  AND U197 ( .A(n11), .B(n260), .Z(n259) );
  XNOR U198 ( .A(p_input[40]), .B(n258), .Z(n260) );
  XOR U199 ( .A(n261), .B(n262), .Z(n258) );
  AND U200 ( .A(n15), .B(n263), .Z(n262) );
  XNOR U201 ( .A(p_input[56]), .B(n261), .Z(n263) );
  XOR U202 ( .A(n264), .B(n265), .Z(n261) );
  AND U203 ( .A(n19), .B(n266), .Z(n265) );
  XNOR U204 ( .A(p_input[72]), .B(n264), .Z(n266) );
  XOR U205 ( .A(n267), .B(n268), .Z(n264) );
  AND U206 ( .A(n23), .B(n269), .Z(n268) );
  XNOR U207 ( .A(p_input[88]), .B(n267), .Z(n269) );
  XOR U208 ( .A(n270), .B(n271), .Z(n267) );
  AND U209 ( .A(n27), .B(n272), .Z(n271) );
  XNOR U210 ( .A(p_input[104]), .B(n270), .Z(n272) );
  XOR U211 ( .A(n273), .B(n274), .Z(n270) );
  AND U212 ( .A(n31), .B(n275), .Z(n274) );
  XNOR U213 ( .A(p_input[120]), .B(n273), .Z(n275) );
  XOR U214 ( .A(n276), .B(n277), .Z(n273) );
  AND U215 ( .A(n35), .B(n278), .Z(n277) );
  XNOR U216 ( .A(p_input[136]), .B(n276), .Z(n278) );
  XOR U217 ( .A(n279), .B(n280), .Z(n276) );
  AND U218 ( .A(n39), .B(n281), .Z(n280) );
  XNOR U219 ( .A(p_input[152]), .B(n279), .Z(n281) );
  XOR U220 ( .A(n282), .B(n283), .Z(n279) );
  AND U221 ( .A(n43), .B(n284), .Z(n283) );
  XNOR U222 ( .A(p_input[168]), .B(n282), .Z(n284) );
  XOR U223 ( .A(n285), .B(n286), .Z(n282) );
  AND U224 ( .A(n47), .B(n287), .Z(n286) );
  XNOR U225 ( .A(p_input[184]), .B(n285), .Z(n287) );
  XOR U226 ( .A(n288), .B(n289), .Z(n285) );
  AND U227 ( .A(n51), .B(n290), .Z(n289) );
  XNOR U228 ( .A(p_input[200]), .B(n288), .Z(n290) );
  XOR U229 ( .A(n291), .B(n292), .Z(n288) );
  AND U230 ( .A(n55), .B(n293), .Z(n292) );
  XNOR U231 ( .A(p_input[216]), .B(n291), .Z(n293) );
  XOR U232 ( .A(n294), .B(n295), .Z(n291) );
  AND U233 ( .A(n59), .B(n296), .Z(n295) );
  XNOR U234 ( .A(p_input[232]), .B(n294), .Z(n296) );
  XOR U235 ( .A(n297), .B(n298), .Z(n294) );
  AND U236 ( .A(n63), .B(n299), .Z(n298) );
  XNOR U237 ( .A(p_input[248]), .B(n297), .Z(n299) );
  XOR U238 ( .A(n300), .B(n301), .Z(n297) );
  AND U239 ( .A(n67), .B(n302), .Z(n301) );
  XNOR U240 ( .A(p_input[264]), .B(n300), .Z(n302) );
  XOR U241 ( .A(n303), .B(n304), .Z(n300) );
  AND U242 ( .A(n71), .B(n305), .Z(n304) );
  XNOR U243 ( .A(p_input[280]), .B(n303), .Z(n305) );
  XOR U244 ( .A(n306), .B(n307), .Z(n303) );
  AND U245 ( .A(n75), .B(n308), .Z(n307) );
  XNOR U246 ( .A(p_input[296]), .B(n306), .Z(n308) );
  XOR U247 ( .A(n309), .B(n310), .Z(n306) );
  AND U248 ( .A(n79), .B(n311), .Z(n310) );
  XNOR U249 ( .A(p_input[312]), .B(n309), .Z(n311) );
  XOR U250 ( .A(n312), .B(n313), .Z(n309) );
  AND U251 ( .A(n83), .B(n314), .Z(n313) );
  XNOR U252 ( .A(p_input[328]), .B(n312), .Z(n314) );
  XOR U253 ( .A(n315), .B(n316), .Z(n312) );
  AND U254 ( .A(n87), .B(n317), .Z(n316) );
  XNOR U255 ( .A(p_input[344]), .B(n315), .Z(n317) );
  XOR U256 ( .A(n318), .B(n319), .Z(n315) );
  AND U257 ( .A(n91), .B(n320), .Z(n319) );
  XNOR U258 ( .A(p_input[360]), .B(n318), .Z(n320) );
  XOR U259 ( .A(n321), .B(n322), .Z(n318) );
  AND U260 ( .A(n95), .B(n323), .Z(n322) );
  XNOR U261 ( .A(p_input[376]), .B(n321), .Z(n323) );
  XOR U262 ( .A(n324), .B(n325), .Z(n321) );
  AND U263 ( .A(n99), .B(n326), .Z(n325) );
  XNOR U264 ( .A(p_input[392]), .B(n324), .Z(n326) );
  XOR U265 ( .A(n327), .B(n328), .Z(n324) );
  AND U266 ( .A(n103), .B(n329), .Z(n328) );
  XNOR U267 ( .A(p_input[408]), .B(n327), .Z(n329) );
  XOR U268 ( .A(n330), .B(n331), .Z(n327) );
  AND U269 ( .A(n107), .B(n332), .Z(n331) );
  XNOR U270 ( .A(p_input[424]), .B(n330), .Z(n332) );
  XOR U271 ( .A(n333), .B(n334), .Z(n330) );
  AND U272 ( .A(n111), .B(n335), .Z(n334) );
  XNOR U273 ( .A(p_input[440]), .B(n333), .Z(n335) );
  XOR U274 ( .A(n336), .B(n337), .Z(n333) );
  AND U275 ( .A(n115), .B(n338), .Z(n337) );
  XNOR U276 ( .A(p_input[456]), .B(n336), .Z(n338) );
  XOR U277 ( .A(n339), .B(n340), .Z(n336) );
  AND U278 ( .A(n119), .B(n341), .Z(n340) );
  XNOR U279 ( .A(p_input[472]), .B(n339), .Z(n341) );
  XOR U280 ( .A(n342), .B(n343), .Z(n339) );
  AND U281 ( .A(n123), .B(n344), .Z(n343) );
  XNOR U282 ( .A(p_input[488]), .B(n342), .Z(n344) );
  XOR U283 ( .A(n345), .B(n346), .Z(n342) );
  AND U284 ( .A(n127), .B(n347), .Z(n346) );
  XNOR U285 ( .A(p_input[504]), .B(n345), .Z(n347) );
  XOR U286 ( .A(n348), .B(n349), .Z(n345) );
  AND U287 ( .A(n131), .B(n350), .Z(n349) );
  XNOR U288 ( .A(p_input[520]), .B(n348), .Z(n350) );
  XOR U289 ( .A(n351), .B(n352), .Z(n348) );
  AND U290 ( .A(n135), .B(n353), .Z(n352) );
  XNOR U291 ( .A(p_input[536]), .B(n351), .Z(n353) );
  XOR U292 ( .A(n354), .B(n355), .Z(n351) );
  AND U293 ( .A(n139), .B(n356), .Z(n355) );
  XNOR U294 ( .A(p_input[552]), .B(n354), .Z(n356) );
  XOR U295 ( .A(n357), .B(n358), .Z(n354) );
  AND U296 ( .A(n143), .B(n359), .Z(n358) );
  XNOR U297 ( .A(p_input[568]), .B(n357), .Z(n359) );
  XOR U298 ( .A(n360), .B(n361), .Z(n357) );
  AND U299 ( .A(n147), .B(n362), .Z(n361) );
  XNOR U300 ( .A(p_input[584]), .B(n360), .Z(n362) );
  XOR U301 ( .A(n363), .B(n364), .Z(n360) );
  AND U302 ( .A(n151), .B(n365), .Z(n364) );
  XNOR U303 ( .A(p_input[600]), .B(n363), .Z(n365) );
  XOR U304 ( .A(n366), .B(n367), .Z(n363) );
  AND U305 ( .A(n155), .B(n368), .Z(n367) );
  XNOR U306 ( .A(p_input[616]), .B(n366), .Z(n368) );
  XOR U307 ( .A(n369), .B(n370), .Z(n366) );
  AND U308 ( .A(n159), .B(n371), .Z(n370) );
  XNOR U309 ( .A(p_input[632]), .B(n369), .Z(n371) );
  XOR U310 ( .A(n372), .B(n373), .Z(n369) );
  AND U311 ( .A(n163), .B(n374), .Z(n373) );
  XNOR U312 ( .A(p_input[648]), .B(n372), .Z(n374) );
  XOR U313 ( .A(n375), .B(n376), .Z(n372) );
  AND U314 ( .A(n167), .B(n377), .Z(n376) );
  XNOR U315 ( .A(p_input[664]), .B(n375), .Z(n377) );
  XOR U316 ( .A(n378), .B(n379), .Z(n375) );
  AND U317 ( .A(n171), .B(n380), .Z(n379) );
  XNOR U318 ( .A(p_input[680]), .B(n378), .Z(n380) );
  XOR U319 ( .A(n381), .B(n382), .Z(n378) );
  AND U320 ( .A(n175), .B(n383), .Z(n382) );
  XNOR U321 ( .A(p_input[696]), .B(n381), .Z(n383) );
  XOR U322 ( .A(n384), .B(n385), .Z(n381) );
  AND U323 ( .A(n179), .B(n386), .Z(n385) );
  XNOR U324 ( .A(p_input[712]), .B(n384), .Z(n386) );
  XOR U325 ( .A(n387), .B(n388), .Z(n384) );
  AND U326 ( .A(n183), .B(n389), .Z(n388) );
  XNOR U327 ( .A(p_input[728]), .B(n387), .Z(n389) );
  XOR U328 ( .A(n390), .B(n391), .Z(n387) );
  AND U329 ( .A(n187), .B(n392), .Z(n391) );
  XNOR U330 ( .A(p_input[744]), .B(n390), .Z(n392) );
  XOR U331 ( .A(n393), .B(n394), .Z(n390) );
  AND U332 ( .A(n191), .B(n395), .Z(n394) );
  XNOR U333 ( .A(p_input[760]), .B(n393), .Z(n395) );
  XOR U334 ( .A(n396), .B(n397), .Z(n393) );
  AND U335 ( .A(n195), .B(n398), .Z(n397) );
  XNOR U336 ( .A(p_input[776]), .B(n396), .Z(n398) );
  XOR U337 ( .A(n399), .B(n400), .Z(n396) );
  AND U338 ( .A(n199), .B(n401), .Z(n400) );
  XNOR U339 ( .A(p_input[792]), .B(n399), .Z(n401) );
  XOR U340 ( .A(n402), .B(n403), .Z(n399) );
  AND U341 ( .A(n203), .B(n404), .Z(n403) );
  XNOR U342 ( .A(p_input[808]), .B(n402), .Z(n404) );
  XOR U343 ( .A(n405), .B(n406), .Z(n402) );
  AND U344 ( .A(n207), .B(n407), .Z(n406) );
  XNOR U345 ( .A(p_input[824]), .B(n405), .Z(n407) );
  XOR U346 ( .A(n408), .B(n409), .Z(n405) );
  AND U347 ( .A(n211), .B(n410), .Z(n409) );
  XNOR U348 ( .A(p_input[840]), .B(n408), .Z(n410) );
  XOR U349 ( .A(n411), .B(n412), .Z(n408) );
  AND U350 ( .A(n215), .B(n413), .Z(n412) );
  XNOR U351 ( .A(p_input[856]), .B(n411), .Z(n413) );
  XOR U352 ( .A(n414), .B(n415), .Z(n411) );
  AND U353 ( .A(n219), .B(n416), .Z(n415) );
  XNOR U354 ( .A(p_input[872]), .B(n414), .Z(n416) );
  XOR U355 ( .A(n417), .B(n418), .Z(n414) );
  AND U356 ( .A(n223), .B(n419), .Z(n418) );
  XNOR U357 ( .A(p_input[888]), .B(n417), .Z(n419) );
  XOR U358 ( .A(n420), .B(n421), .Z(n417) );
  AND U359 ( .A(n227), .B(n422), .Z(n421) );
  XNOR U360 ( .A(p_input[904]), .B(n420), .Z(n422) );
  XOR U361 ( .A(n423), .B(n424), .Z(n420) );
  AND U362 ( .A(n231), .B(n425), .Z(n424) );
  XNOR U363 ( .A(p_input[920]), .B(n423), .Z(n425) );
  XOR U364 ( .A(n426), .B(n427), .Z(n423) );
  AND U365 ( .A(n235), .B(n428), .Z(n427) );
  XNOR U366 ( .A(p_input[936]), .B(n426), .Z(n428) );
  XOR U367 ( .A(n429), .B(n430), .Z(n426) );
  AND U368 ( .A(n239), .B(n431), .Z(n430) );
  XNOR U369 ( .A(p_input[952]), .B(n429), .Z(n431) );
  XOR U370 ( .A(n432), .B(n433), .Z(n429) );
  AND U371 ( .A(n243), .B(n434), .Z(n433) );
  XNOR U372 ( .A(p_input[968]), .B(n432), .Z(n434) );
  XNOR U373 ( .A(n435), .B(n436), .Z(n432) );
  AND U374 ( .A(n247), .B(n437), .Z(n436) );
  XOR U375 ( .A(p_input[984]), .B(n435), .Z(n437) );
  XOR U376 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n438), .Z(n435) );
  AND U377 ( .A(n250), .B(n439), .Z(n438) );
  XOR U378 ( .A(p_input[1000]), .B(\knn_comb_/min_val_out[0][8] ), .Z(n439) );
  XNOR U379 ( .A(n440), .B(n441), .Z(o[7]) );
  AND U380 ( .A(n3), .B(n442), .Z(n440) );
  XNOR U381 ( .A(p_input[7]), .B(n441), .Z(n442) );
  XOR U382 ( .A(n443), .B(n444), .Z(n441) );
  AND U383 ( .A(n7), .B(n445), .Z(n444) );
  XNOR U384 ( .A(p_input[23]), .B(n443), .Z(n445) );
  XOR U385 ( .A(n446), .B(n447), .Z(n443) );
  AND U386 ( .A(n11), .B(n448), .Z(n447) );
  XNOR U387 ( .A(p_input[39]), .B(n446), .Z(n448) );
  XOR U388 ( .A(n449), .B(n450), .Z(n446) );
  AND U389 ( .A(n15), .B(n451), .Z(n450) );
  XNOR U390 ( .A(p_input[55]), .B(n449), .Z(n451) );
  XOR U391 ( .A(n452), .B(n453), .Z(n449) );
  AND U392 ( .A(n19), .B(n454), .Z(n453) );
  XNOR U393 ( .A(p_input[71]), .B(n452), .Z(n454) );
  XOR U394 ( .A(n455), .B(n456), .Z(n452) );
  AND U395 ( .A(n23), .B(n457), .Z(n456) );
  XNOR U396 ( .A(p_input[87]), .B(n455), .Z(n457) );
  XOR U397 ( .A(n458), .B(n459), .Z(n455) );
  AND U398 ( .A(n27), .B(n460), .Z(n459) );
  XNOR U399 ( .A(p_input[103]), .B(n458), .Z(n460) );
  XOR U400 ( .A(n461), .B(n462), .Z(n458) );
  AND U401 ( .A(n31), .B(n463), .Z(n462) );
  XNOR U402 ( .A(p_input[119]), .B(n461), .Z(n463) );
  XOR U403 ( .A(n464), .B(n465), .Z(n461) );
  AND U404 ( .A(n35), .B(n466), .Z(n465) );
  XNOR U405 ( .A(p_input[135]), .B(n464), .Z(n466) );
  XOR U406 ( .A(n467), .B(n468), .Z(n464) );
  AND U407 ( .A(n39), .B(n469), .Z(n468) );
  XNOR U408 ( .A(p_input[151]), .B(n467), .Z(n469) );
  XOR U409 ( .A(n470), .B(n471), .Z(n467) );
  AND U410 ( .A(n43), .B(n472), .Z(n471) );
  XNOR U411 ( .A(p_input[167]), .B(n470), .Z(n472) );
  XOR U412 ( .A(n473), .B(n474), .Z(n470) );
  AND U413 ( .A(n47), .B(n475), .Z(n474) );
  XNOR U414 ( .A(p_input[183]), .B(n473), .Z(n475) );
  XOR U415 ( .A(n476), .B(n477), .Z(n473) );
  AND U416 ( .A(n51), .B(n478), .Z(n477) );
  XNOR U417 ( .A(p_input[199]), .B(n476), .Z(n478) );
  XOR U418 ( .A(n479), .B(n480), .Z(n476) );
  AND U419 ( .A(n55), .B(n481), .Z(n480) );
  XNOR U420 ( .A(p_input[215]), .B(n479), .Z(n481) );
  XOR U421 ( .A(n482), .B(n483), .Z(n479) );
  AND U422 ( .A(n59), .B(n484), .Z(n483) );
  XNOR U423 ( .A(p_input[231]), .B(n482), .Z(n484) );
  XOR U424 ( .A(n485), .B(n486), .Z(n482) );
  AND U425 ( .A(n63), .B(n487), .Z(n486) );
  XNOR U426 ( .A(p_input[247]), .B(n485), .Z(n487) );
  XOR U427 ( .A(n488), .B(n489), .Z(n485) );
  AND U428 ( .A(n67), .B(n490), .Z(n489) );
  XNOR U429 ( .A(p_input[263]), .B(n488), .Z(n490) );
  XOR U430 ( .A(n491), .B(n492), .Z(n488) );
  AND U431 ( .A(n71), .B(n493), .Z(n492) );
  XNOR U432 ( .A(p_input[279]), .B(n491), .Z(n493) );
  XOR U433 ( .A(n494), .B(n495), .Z(n491) );
  AND U434 ( .A(n75), .B(n496), .Z(n495) );
  XNOR U435 ( .A(p_input[295]), .B(n494), .Z(n496) );
  XOR U436 ( .A(n497), .B(n498), .Z(n494) );
  AND U437 ( .A(n79), .B(n499), .Z(n498) );
  XNOR U438 ( .A(p_input[311]), .B(n497), .Z(n499) );
  XOR U439 ( .A(n500), .B(n501), .Z(n497) );
  AND U440 ( .A(n83), .B(n502), .Z(n501) );
  XNOR U441 ( .A(p_input[327]), .B(n500), .Z(n502) );
  XOR U442 ( .A(n503), .B(n504), .Z(n500) );
  AND U443 ( .A(n87), .B(n505), .Z(n504) );
  XNOR U444 ( .A(p_input[343]), .B(n503), .Z(n505) );
  XOR U445 ( .A(n506), .B(n507), .Z(n503) );
  AND U446 ( .A(n91), .B(n508), .Z(n507) );
  XNOR U447 ( .A(p_input[359]), .B(n506), .Z(n508) );
  XOR U448 ( .A(n509), .B(n510), .Z(n506) );
  AND U449 ( .A(n95), .B(n511), .Z(n510) );
  XNOR U450 ( .A(p_input[375]), .B(n509), .Z(n511) );
  XOR U451 ( .A(n512), .B(n513), .Z(n509) );
  AND U452 ( .A(n99), .B(n514), .Z(n513) );
  XNOR U453 ( .A(p_input[391]), .B(n512), .Z(n514) );
  XOR U454 ( .A(n515), .B(n516), .Z(n512) );
  AND U455 ( .A(n103), .B(n517), .Z(n516) );
  XNOR U456 ( .A(p_input[407]), .B(n515), .Z(n517) );
  XOR U457 ( .A(n518), .B(n519), .Z(n515) );
  AND U458 ( .A(n107), .B(n520), .Z(n519) );
  XNOR U459 ( .A(p_input[423]), .B(n518), .Z(n520) );
  XOR U460 ( .A(n521), .B(n522), .Z(n518) );
  AND U461 ( .A(n111), .B(n523), .Z(n522) );
  XNOR U462 ( .A(p_input[439]), .B(n521), .Z(n523) );
  XOR U463 ( .A(n524), .B(n525), .Z(n521) );
  AND U464 ( .A(n115), .B(n526), .Z(n525) );
  XNOR U465 ( .A(p_input[455]), .B(n524), .Z(n526) );
  XOR U466 ( .A(n527), .B(n528), .Z(n524) );
  AND U467 ( .A(n119), .B(n529), .Z(n528) );
  XNOR U468 ( .A(p_input[471]), .B(n527), .Z(n529) );
  XOR U469 ( .A(n530), .B(n531), .Z(n527) );
  AND U470 ( .A(n123), .B(n532), .Z(n531) );
  XNOR U471 ( .A(p_input[487]), .B(n530), .Z(n532) );
  XOR U472 ( .A(n533), .B(n534), .Z(n530) );
  AND U473 ( .A(n127), .B(n535), .Z(n534) );
  XNOR U474 ( .A(p_input[503]), .B(n533), .Z(n535) );
  XOR U475 ( .A(n536), .B(n537), .Z(n533) );
  AND U476 ( .A(n131), .B(n538), .Z(n537) );
  XNOR U477 ( .A(p_input[519]), .B(n536), .Z(n538) );
  XOR U478 ( .A(n539), .B(n540), .Z(n536) );
  AND U479 ( .A(n135), .B(n541), .Z(n540) );
  XNOR U480 ( .A(p_input[535]), .B(n539), .Z(n541) );
  XOR U481 ( .A(n542), .B(n543), .Z(n539) );
  AND U482 ( .A(n139), .B(n544), .Z(n543) );
  XNOR U483 ( .A(p_input[551]), .B(n542), .Z(n544) );
  XOR U484 ( .A(n545), .B(n546), .Z(n542) );
  AND U485 ( .A(n143), .B(n547), .Z(n546) );
  XNOR U486 ( .A(p_input[567]), .B(n545), .Z(n547) );
  XOR U487 ( .A(n548), .B(n549), .Z(n545) );
  AND U488 ( .A(n147), .B(n550), .Z(n549) );
  XNOR U489 ( .A(p_input[583]), .B(n548), .Z(n550) );
  XOR U490 ( .A(n551), .B(n552), .Z(n548) );
  AND U491 ( .A(n151), .B(n553), .Z(n552) );
  XNOR U492 ( .A(p_input[599]), .B(n551), .Z(n553) );
  XOR U493 ( .A(n554), .B(n555), .Z(n551) );
  AND U494 ( .A(n155), .B(n556), .Z(n555) );
  XNOR U495 ( .A(p_input[615]), .B(n554), .Z(n556) );
  XOR U496 ( .A(n557), .B(n558), .Z(n554) );
  AND U497 ( .A(n159), .B(n559), .Z(n558) );
  XNOR U498 ( .A(p_input[631]), .B(n557), .Z(n559) );
  XOR U499 ( .A(n560), .B(n561), .Z(n557) );
  AND U500 ( .A(n163), .B(n562), .Z(n561) );
  XNOR U501 ( .A(p_input[647]), .B(n560), .Z(n562) );
  XOR U502 ( .A(n563), .B(n564), .Z(n560) );
  AND U503 ( .A(n167), .B(n565), .Z(n564) );
  XNOR U504 ( .A(p_input[663]), .B(n563), .Z(n565) );
  XOR U505 ( .A(n566), .B(n567), .Z(n563) );
  AND U506 ( .A(n171), .B(n568), .Z(n567) );
  XNOR U507 ( .A(p_input[679]), .B(n566), .Z(n568) );
  XOR U508 ( .A(n569), .B(n570), .Z(n566) );
  AND U509 ( .A(n175), .B(n571), .Z(n570) );
  XNOR U510 ( .A(p_input[695]), .B(n569), .Z(n571) );
  XOR U511 ( .A(n572), .B(n573), .Z(n569) );
  AND U512 ( .A(n179), .B(n574), .Z(n573) );
  XNOR U513 ( .A(p_input[711]), .B(n572), .Z(n574) );
  XOR U514 ( .A(n575), .B(n576), .Z(n572) );
  AND U515 ( .A(n183), .B(n577), .Z(n576) );
  XNOR U516 ( .A(p_input[727]), .B(n575), .Z(n577) );
  XOR U517 ( .A(n578), .B(n579), .Z(n575) );
  AND U518 ( .A(n187), .B(n580), .Z(n579) );
  XNOR U519 ( .A(p_input[743]), .B(n578), .Z(n580) );
  XOR U520 ( .A(n581), .B(n582), .Z(n578) );
  AND U521 ( .A(n191), .B(n583), .Z(n582) );
  XNOR U522 ( .A(p_input[759]), .B(n581), .Z(n583) );
  XOR U523 ( .A(n584), .B(n585), .Z(n581) );
  AND U524 ( .A(n195), .B(n586), .Z(n585) );
  XNOR U525 ( .A(p_input[775]), .B(n584), .Z(n586) );
  XOR U526 ( .A(n587), .B(n588), .Z(n584) );
  AND U527 ( .A(n199), .B(n589), .Z(n588) );
  XNOR U528 ( .A(p_input[791]), .B(n587), .Z(n589) );
  XOR U529 ( .A(n590), .B(n591), .Z(n587) );
  AND U530 ( .A(n203), .B(n592), .Z(n591) );
  XNOR U531 ( .A(p_input[807]), .B(n590), .Z(n592) );
  XOR U532 ( .A(n593), .B(n594), .Z(n590) );
  AND U533 ( .A(n207), .B(n595), .Z(n594) );
  XNOR U534 ( .A(p_input[823]), .B(n593), .Z(n595) );
  XOR U535 ( .A(n596), .B(n597), .Z(n593) );
  AND U536 ( .A(n211), .B(n598), .Z(n597) );
  XNOR U537 ( .A(p_input[839]), .B(n596), .Z(n598) );
  XOR U538 ( .A(n599), .B(n600), .Z(n596) );
  AND U539 ( .A(n215), .B(n601), .Z(n600) );
  XNOR U540 ( .A(p_input[855]), .B(n599), .Z(n601) );
  XOR U541 ( .A(n602), .B(n603), .Z(n599) );
  AND U542 ( .A(n219), .B(n604), .Z(n603) );
  XNOR U543 ( .A(p_input[871]), .B(n602), .Z(n604) );
  XOR U544 ( .A(n605), .B(n606), .Z(n602) );
  AND U545 ( .A(n223), .B(n607), .Z(n606) );
  XNOR U546 ( .A(p_input[887]), .B(n605), .Z(n607) );
  XOR U547 ( .A(n608), .B(n609), .Z(n605) );
  AND U548 ( .A(n227), .B(n610), .Z(n609) );
  XNOR U549 ( .A(p_input[903]), .B(n608), .Z(n610) );
  XOR U550 ( .A(n611), .B(n612), .Z(n608) );
  AND U551 ( .A(n231), .B(n613), .Z(n612) );
  XNOR U552 ( .A(p_input[919]), .B(n611), .Z(n613) );
  XOR U553 ( .A(n614), .B(n615), .Z(n611) );
  AND U554 ( .A(n235), .B(n616), .Z(n615) );
  XNOR U555 ( .A(p_input[935]), .B(n614), .Z(n616) );
  XOR U556 ( .A(n617), .B(n618), .Z(n614) );
  AND U557 ( .A(n239), .B(n619), .Z(n618) );
  XNOR U558 ( .A(p_input[951]), .B(n617), .Z(n619) );
  XOR U559 ( .A(n620), .B(n621), .Z(n617) );
  AND U560 ( .A(n243), .B(n622), .Z(n621) );
  XNOR U561 ( .A(p_input[967]), .B(n620), .Z(n622) );
  XNOR U562 ( .A(n623), .B(n624), .Z(n620) );
  AND U563 ( .A(n247), .B(n625), .Z(n624) );
  XOR U564 ( .A(p_input[983]), .B(n623), .Z(n625) );
  XOR U565 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n626), .Z(n623) );
  AND U566 ( .A(n250), .B(n627), .Z(n626) );
  XOR U567 ( .A(p_input[999]), .B(\knn_comb_/min_val_out[0][7] ), .Z(n627) );
  XNOR U568 ( .A(n628), .B(n629), .Z(o[6]) );
  AND U569 ( .A(n3), .B(n630), .Z(n628) );
  XNOR U570 ( .A(p_input[6]), .B(n629), .Z(n630) );
  XOR U571 ( .A(n631), .B(n632), .Z(n629) );
  AND U572 ( .A(n7), .B(n633), .Z(n632) );
  XNOR U573 ( .A(p_input[22]), .B(n631), .Z(n633) );
  XOR U574 ( .A(n634), .B(n635), .Z(n631) );
  AND U575 ( .A(n11), .B(n636), .Z(n635) );
  XNOR U576 ( .A(p_input[38]), .B(n634), .Z(n636) );
  XOR U577 ( .A(n637), .B(n638), .Z(n634) );
  AND U578 ( .A(n15), .B(n639), .Z(n638) );
  XNOR U579 ( .A(p_input[54]), .B(n637), .Z(n639) );
  XOR U580 ( .A(n640), .B(n641), .Z(n637) );
  AND U581 ( .A(n19), .B(n642), .Z(n641) );
  XNOR U582 ( .A(p_input[70]), .B(n640), .Z(n642) );
  XOR U583 ( .A(n643), .B(n644), .Z(n640) );
  AND U584 ( .A(n23), .B(n645), .Z(n644) );
  XNOR U585 ( .A(p_input[86]), .B(n643), .Z(n645) );
  XOR U586 ( .A(n646), .B(n647), .Z(n643) );
  AND U587 ( .A(n27), .B(n648), .Z(n647) );
  XNOR U588 ( .A(p_input[102]), .B(n646), .Z(n648) );
  XOR U589 ( .A(n649), .B(n650), .Z(n646) );
  AND U590 ( .A(n31), .B(n651), .Z(n650) );
  XNOR U591 ( .A(p_input[118]), .B(n649), .Z(n651) );
  XOR U592 ( .A(n652), .B(n653), .Z(n649) );
  AND U593 ( .A(n35), .B(n654), .Z(n653) );
  XNOR U594 ( .A(p_input[134]), .B(n652), .Z(n654) );
  XOR U595 ( .A(n655), .B(n656), .Z(n652) );
  AND U596 ( .A(n39), .B(n657), .Z(n656) );
  XNOR U597 ( .A(p_input[150]), .B(n655), .Z(n657) );
  XOR U598 ( .A(n658), .B(n659), .Z(n655) );
  AND U599 ( .A(n43), .B(n660), .Z(n659) );
  XNOR U600 ( .A(p_input[166]), .B(n658), .Z(n660) );
  XOR U601 ( .A(n661), .B(n662), .Z(n658) );
  AND U602 ( .A(n47), .B(n663), .Z(n662) );
  XNOR U603 ( .A(p_input[182]), .B(n661), .Z(n663) );
  XOR U604 ( .A(n664), .B(n665), .Z(n661) );
  AND U605 ( .A(n51), .B(n666), .Z(n665) );
  XNOR U606 ( .A(p_input[198]), .B(n664), .Z(n666) );
  XOR U607 ( .A(n667), .B(n668), .Z(n664) );
  AND U608 ( .A(n55), .B(n669), .Z(n668) );
  XNOR U609 ( .A(p_input[214]), .B(n667), .Z(n669) );
  XOR U610 ( .A(n670), .B(n671), .Z(n667) );
  AND U611 ( .A(n59), .B(n672), .Z(n671) );
  XNOR U612 ( .A(p_input[230]), .B(n670), .Z(n672) );
  XOR U613 ( .A(n673), .B(n674), .Z(n670) );
  AND U614 ( .A(n63), .B(n675), .Z(n674) );
  XNOR U615 ( .A(p_input[246]), .B(n673), .Z(n675) );
  XOR U616 ( .A(n676), .B(n677), .Z(n673) );
  AND U617 ( .A(n67), .B(n678), .Z(n677) );
  XNOR U618 ( .A(p_input[262]), .B(n676), .Z(n678) );
  XOR U619 ( .A(n679), .B(n680), .Z(n676) );
  AND U620 ( .A(n71), .B(n681), .Z(n680) );
  XNOR U621 ( .A(p_input[278]), .B(n679), .Z(n681) );
  XOR U622 ( .A(n682), .B(n683), .Z(n679) );
  AND U623 ( .A(n75), .B(n684), .Z(n683) );
  XNOR U624 ( .A(p_input[294]), .B(n682), .Z(n684) );
  XOR U625 ( .A(n685), .B(n686), .Z(n682) );
  AND U626 ( .A(n79), .B(n687), .Z(n686) );
  XNOR U627 ( .A(p_input[310]), .B(n685), .Z(n687) );
  XOR U628 ( .A(n688), .B(n689), .Z(n685) );
  AND U629 ( .A(n83), .B(n690), .Z(n689) );
  XNOR U630 ( .A(p_input[326]), .B(n688), .Z(n690) );
  XOR U631 ( .A(n691), .B(n692), .Z(n688) );
  AND U632 ( .A(n87), .B(n693), .Z(n692) );
  XNOR U633 ( .A(p_input[342]), .B(n691), .Z(n693) );
  XOR U634 ( .A(n694), .B(n695), .Z(n691) );
  AND U635 ( .A(n91), .B(n696), .Z(n695) );
  XNOR U636 ( .A(p_input[358]), .B(n694), .Z(n696) );
  XOR U637 ( .A(n697), .B(n698), .Z(n694) );
  AND U638 ( .A(n95), .B(n699), .Z(n698) );
  XNOR U639 ( .A(p_input[374]), .B(n697), .Z(n699) );
  XOR U640 ( .A(n700), .B(n701), .Z(n697) );
  AND U641 ( .A(n99), .B(n702), .Z(n701) );
  XNOR U642 ( .A(p_input[390]), .B(n700), .Z(n702) );
  XOR U643 ( .A(n703), .B(n704), .Z(n700) );
  AND U644 ( .A(n103), .B(n705), .Z(n704) );
  XNOR U645 ( .A(p_input[406]), .B(n703), .Z(n705) );
  XOR U646 ( .A(n706), .B(n707), .Z(n703) );
  AND U647 ( .A(n107), .B(n708), .Z(n707) );
  XNOR U648 ( .A(p_input[422]), .B(n706), .Z(n708) );
  XOR U649 ( .A(n709), .B(n710), .Z(n706) );
  AND U650 ( .A(n111), .B(n711), .Z(n710) );
  XNOR U651 ( .A(p_input[438]), .B(n709), .Z(n711) );
  XOR U652 ( .A(n712), .B(n713), .Z(n709) );
  AND U653 ( .A(n115), .B(n714), .Z(n713) );
  XNOR U654 ( .A(p_input[454]), .B(n712), .Z(n714) );
  XOR U655 ( .A(n715), .B(n716), .Z(n712) );
  AND U656 ( .A(n119), .B(n717), .Z(n716) );
  XNOR U657 ( .A(p_input[470]), .B(n715), .Z(n717) );
  XOR U658 ( .A(n718), .B(n719), .Z(n715) );
  AND U659 ( .A(n123), .B(n720), .Z(n719) );
  XNOR U660 ( .A(p_input[486]), .B(n718), .Z(n720) );
  XOR U661 ( .A(n721), .B(n722), .Z(n718) );
  AND U662 ( .A(n127), .B(n723), .Z(n722) );
  XNOR U663 ( .A(p_input[502]), .B(n721), .Z(n723) );
  XOR U664 ( .A(n724), .B(n725), .Z(n721) );
  AND U665 ( .A(n131), .B(n726), .Z(n725) );
  XNOR U666 ( .A(p_input[518]), .B(n724), .Z(n726) );
  XOR U667 ( .A(n727), .B(n728), .Z(n724) );
  AND U668 ( .A(n135), .B(n729), .Z(n728) );
  XNOR U669 ( .A(p_input[534]), .B(n727), .Z(n729) );
  XOR U670 ( .A(n730), .B(n731), .Z(n727) );
  AND U671 ( .A(n139), .B(n732), .Z(n731) );
  XNOR U672 ( .A(p_input[550]), .B(n730), .Z(n732) );
  XOR U673 ( .A(n733), .B(n734), .Z(n730) );
  AND U674 ( .A(n143), .B(n735), .Z(n734) );
  XNOR U675 ( .A(p_input[566]), .B(n733), .Z(n735) );
  XOR U676 ( .A(n736), .B(n737), .Z(n733) );
  AND U677 ( .A(n147), .B(n738), .Z(n737) );
  XNOR U678 ( .A(p_input[582]), .B(n736), .Z(n738) );
  XOR U679 ( .A(n739), .B(n740), .Z(n736) );
  AND U680 ( .A(n151), .B(n741), .Z(n740) );
  XNOR U681 ( .A(p_input[598]), .B(n739), .Z(n741) );
  XOR U682 ( .A(n742), .B(n743), .Z(n739) );
  AND U683 ( .A(n155), .B(n744), .Z(n743) );
  XNOR U684 ( .A(p_input[614]), .B(n742), .Z(n744) );
  XOR U685 ( .A(n745), .B(n746), .Z(n742) );
  AND U686 ( .A(n159), .B(n747), .Z(n746) );
  XNOR U687 ( .A(p_input[630]), .B(n745), .Z(n747) );
  XOR U688 ( .A(n748), .B(n749), .Z(n745) );
  AND U689 ( .A(n163), .B(n750), .Z(n749) );
  XNOR U690 ( .A(p_input[646]), .B(n748), .Z(n750) );
  XOR U691 ( .A(n751), .B(n752), .Z(n748) );
  AND U692 ( .A(n167), .B(n753), .Z(n752) );
  XNOR U693 ( .A(p_input[662]), .B(n751), .Z(n753) );
  XOR U694 ( .A(n754), .B(n755), .Z(n751) );
  AND U695 ( .A(n171), .B(n756), .Z(n755) );
  XNOR U696 ( .A(p_input[678]), .B(n754), .Z(n756) );
  XOR U697 ( .A(n757), .B(n758), .Z(n754) );
  AND U698 ( .A(n175), .B(n759), .Z(n758) );
  XNOR U699 ( .A(p_input[694]), .B(n757), .Z(n759) );
  XOR U700 ( .A(n760), .B(n761), .Z(n757) );
  AND U701 ( .A(n179), .B(n762), .Z(n761) );
  XNOR U702 ( .A(p_input[710]), .B(n760), .Z(n762) );
  XOR U703 ( .A(n763), .B(n764), .Z(n760) );
  AND U704 ( .A(n183), .B(n765), .Z(n764) );
  XNOR U705 ( .A(p_input[726]), .B(n763), .Z(n765) );
  XOR U706 ( .A(n766), .B(n767), .Z(n763) );
  AND U707 ( .A(n187), .B(n768), .Z(n767) );
  XNOR U708 ( .A(p_input[742]), .B(n766), .Z(n768) );
  XOR U709 ( .A(n769), .B(n770), .Z(n766) );
  AND U710 ( .A(n191), .B(n771), .Z(n770) );
  XNOR U711 ( .A(p_input[758]), .B(n769), .Z(n771) );
  XOR U712 ( .A(n772), .B(n773), .Z(n769) );
  AND U713 ( .A(n195), .B(n774), .Z(n773) );
  XNOR U714 ( .A(p_input[774]), .B(n772), .Z(n774) );
  XOR U715 ( .A(n775), .B(n776), .Z(n772) );
  AND U716 ( .A(n199), .B(n777), .Z(n776) );
  XNOR U717 ( .A(p_input[790]), .B(n775), .Z(n777) );
  XOR U718 ( .A(n778), .B(n779), .Z(n775) );
  AND U719 ( .A(n203), .B(n780), .Z(n779) );
  XNOR U720 ( .A(p_input[806]), .B(n778), .Z(n780) );
  XOR U721 ( .A(n781), .B(n782), .Z(n778) );
  AND U722 ( .A(n207), .B(n783), .Z(n782) );
  XNOR U723 ( .A(p_input[822]), .B(n781), .Z(n783) );
  XOR U724 ( .A(n784), .B(n785), .Z(n781) );
  AND U725 ( .A(n211), .B(n786), .Z(n785) );
  XNOR U726 ( .A(p_input[838]), .B(n784), .Z(n786) );
  XOR U727 ( .A(n787), .B(n788), .Z(n784) );
  AND U728 ( .A(n215), .B(n789), .Z(n788) );
  XNOR U729 ( .A(p_input[854]), .B(n787), .Z(n789) );
  XOR U730 ( .A(n790), .B(n791), .Z(n787) );
  AND U731 ( .A(n219), .B(n792), .Z(n791) );
  XNOR U732 ( .A(p_input[870]), .B(n790), .Z(n792) );
  XOR U733 ( .A(n793), .B(n794), .Z(n790) );
  AND U734 ( .A(n223), .B(n795), .Z(n794) );
  XNOR U735 ( .A(p_input[886]), .B(n793), .Z(n795) );
  XOR U736 ( .A(n796), .B(n797), .Z(n793) );
  AND U737 ( .A(n227), .B(n798), .Z(n797) );
  XNOR U738 ( .A(p_input[902]), .B(n796), .Z(n798) );
  XOR U739 ( .A(n799), .B(n800), .Z(n796) );
  AND U740 ( .A(n231), .B(n801), .Z(n800) );
  XNOR U741 ( .A(p_input[918]), .B(n799), .Z(n801) );
  XOR U742 ( .A(n802), .B(n803), .Z(n799) );
  AND U743 ( .A(n235), .B(n804), .Z(n803) );
  XNOR U744 ( .A(p_input[934]), .B(n802), .Z(n804) );
  XOR U745 ( .A(n805), .B(n806), .Z(n802) );
  AND U746 ( .A(n239), .B(n807), .Z(n806) );
  XNOR U747 ( .A(p_input[950]), .B(n805), .Z(n807) );
  XOR U748 ( .A(n808), .B(n809), .Z(n805) );
  AND U749 ( .A(n243), .B(n810), .Z(n809) );
  XNOR U750 ( .A(p_input[966]), .B(n808), .Z(n810) );
  XNOR U751 ( .A(n811), .B(n812), .Z(n808) );
  AND U752 ( .A(n247), .B(n813), .Z(n812) );
  XOR U753 ( .A(p_input[982]), .B(n811), .Z(n813) );
  XOR U754 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n814), .Z(n811) );
  AND U755 ( .A(n250), .B(n815), .Z(n814) );
  XOR U756 ( .A(p_input[998]), .B(\knn_comb_/min_val_out[0][6] ), .Z(n815) );
  XNOR U757 ( .A(n816), .B(n817), .Z(o[5]) );
  AND U758 ( .A(n3), .B(n818), .Z(n816) );
  XNOR U759 ( .A(p_input[5]), .B(n817), .Z(n818) );
  XOR U760 ( .A(n819), .B(n820), .Z(n817) );
  AND U761 ( .A(n7), .B(n821), .Z(n820) );
  XNOR U762 ( .A(p_input[21]), .B(n819), .Z(n821) );
  XOR U763 ( .A(n822), .B(n823), .Z(n819) );
  AND U764 ( .A(n11), .B(n824), .Z(n823) );
  XNOR U765 ( .A(p_input[37]), .B(n822), .Z(n824) );
  XOR U766 ( .A(n825), .B(n826), .Z(n822) );
  AND U767 ( .A(n15), .B(n827), .Z(n826) );
  XNOR U768 ( .A(p_input[53]), .B(n825), .Z(n827) );
  XOR U769 ( .A(n828), .B(n829), .Z(n825) );
  AND U770 ( .A(n19), .B(n830), .Z(n829) );
  XNOR U771 ( .A(p_input[69]), .B(n828), .Z(n830) );
  XOR U772 ( .A(n831), .B(n832), .Z(n828) );
  AND U773 ( .A(n23), .B(n833), .Z(n832) );
  XNOR U774 ( .A(p_input[85]), .B(n831), .Z(n833) );
  XOR U775 ( .A(n834), .B(n835), .Z(n831) );
  AND U776 ( .A(n27), .B(n836), .Z(n835) );
  XNOR U777 ( .A(p_input[101]), .B(n834), .Z(n836) );
  XOR U778 ( .A(n837), .B(n838), .Z(n834) );
  AND U779 ( .A(n31), .B(n839), .Z(n838) );
  XNOR U780 ( .A(p_input[117]), .B(n837), .Z(n839) );
  XOR U781 ( .A(n840), .B(n841), .Z(n837) );
  AND U782 ( .A(n35), .B(n842), .Z(n841) );
  XNOR U783 ( .A(p_input[133]), .B(n840), .Z(n842) );
  XOR U784 ( .A(n843), .B(n844), .Z(n840) );
  AND U785 ( .A(n39), .B(n845), .Z(n844) );
  XNOR U786 ( .A(p_input[149]), .B(n843), .Z(n845) );
  XOR U787 ( .A(n846), .B(n847), .Z(n843) );
  AND U788 ( .A(n43), .B(n848), .Z(n847) );
  XNOR U789 ( .A(p_input[165]), .B(n846), .Z(n848) );
  XOR U790 ( .A(n849), .B(n850), .Z(n846) );
  AND U791 ( .A(n47), .B(n851), .Z(n850) );
  XNOR U792 ( .A(p_input[181]), .B(n849), .Z(n851) );
  XOR U793 ( .A(n852), .B(n853), .Z(n849) );
  AND U794 ( .A(n51), .B(n854), .Z(n853) );
  XNOR U795 ( .A(p_input[197]), .B(n852), .Z(n854) );
  XOR U796 ( .A(n855), .B(n856), .Z(n852) );
  AND U797 ( .A(n55), .B(n857), .Z(n856) );
  XNOR U798 ( .A(p_input[213]), .B(n855), .Z(n857) );
  XOR U799 ( .A(n858), .B(n859), .Z(n855) );
  AND U800 ( .A(n59), .B(n860), .Z(n859) );
  XNOR U801 ( .A(p_input[229]), .B(n858), .Z(n860) );
  XOR U802 ( .A(n861), .B(n862), .Z(n858) );
  AND U803 ( .A(n63), .B(n863), .Z(n862) );
  XNOR U804 ( .A(p_input[245]), .B(n861), .Z(n863) );
  XOR U805 ( .A(n864), .B(n865), .Z(n861) );
  AND U806 ( .A(n67), .B(n866), .Z(n865) );
  XNOR U807 ( .A(p_input[261]), .B(n864), .Z(n866) );
  XOR U808 ( .A(n867), .B(n868), .Z(n864) );
  AND U809 ( .A(n71), .B(n869), .Z(n868) );
  XNOR U810 ( .A(p_input[277]), .B(n867), .Z(n869) );
  XOR U811 ( .A(n870), .B(n871), .Z(n867) );
  AND U812 ( .A(n75), .B(n872), .Z(n871) );
  XNOR U813 ( .A(p_input[293]), .B(n870), .Z(n872) );
  XOR U814 ( .A(n873), .B(n874), .Z(n870) );
  AND U815 ( .A(n79), .B(n875), .Z(n874) );
  XNOR U816 ( .A(p_input[309]), .B(n873), .Z(n875) );
  XOR U817 ( .A(n876), .B(n877), .Z(n873) );
  AND U818 ( .A(n83), .B(n878), .Z(n877) );
  XNOR U819 ( .A(p_input[325]), .B(n876), .Z(n878) );
  XOR U820 ( .A(n879), .B(n880), .Z(n876) );
  AND U821 ( .A(n87), .B(n881), .Z(n880) );
  XNOR U822 ( .A(p_input[341]), .B(n879), .Z(n881) );
  XOR U823 ( .A(n882), .B(n883), .Z(n879) );
  AND U824 ( .A(n91), .B(n884), .Z(n883) );
  XNOR U825 ( .A(p_input[357]), .B(n882), .Z(n884) );
  XOR U826 ( .A(n885), .B(n886), .Z(n882) );
  AND U827 ( .A(n95), .B(n887), .Z(n886) );
  XNOR U828 ( .A(p_input[373]), .B(n885), .Z(n887) );
  XOR U829 ( .A(n888), .B(n889), .Z(n885) );
  AND U830 ( .A(n99), .B(n890), .Z(n889) );
  XNOR U831 ( .A(p_input[389]), .B(n888), .Z(n890) );
  XOR U832 ( .A(n891), .B(n892), .Z(n888) );
  AND U833 ( .A(n103), .B(n893), .Z(n892) );
  XNOR U834 ( .A(p_input[405]), .B(n891), .Z(n893) );
  XOR U835 ( .A(n894), .B(n895), .Z(n891) );
  AND U836 ( .A(n107), .B(n896), .Z(n895) );
  XNOR U837 ( .A(p_input[421]), .B(n894), .Z(n896) );
  XOR U838 ( .A(n897), .B(n898), .Z(n894) );
  AND U839 ( .A(n111), .B(n899), .Z(n898) );
  XNOR U840 ( .A(p_input[437]), .B(n897), .Z(n899) );
  XOR U841 ( .A(n900), .B(n901), .Z(n897) );
  AND U842 ( .A(n115), .B(n902), .Z(n901) );
  XNOR U843 ( .A(p_input[453]), .B(n900), .Z(n902) );
  XOR U844 ( .A(n903), .B(n904), .Z(n900) );
  AND U845 ( .A(n119), .B(n905), .Z(n904) );
  XNOR U846 ( .A(p_input[469]), .B(n903), .Z(n905) );
  XOR U847 ( .A(n906), .B(n907), .Z(n903) );
  AND U848 ( .A(n123), .B(n908), .Z(n907) );
  XNOR U849 ( .A(p_input[485]), .B(n906), .Z(n908) );
  XOR U850 ( .A(n909), .B(n910), .Z(n906) );
  AND U851 ( .A(n127), .B(n911), .Z(n910) );
  XNOR U852 ( .A(p_input[501]), .B(n909), .Z(n911) );
  XOR U853 ( .A(n912), .B(n913), .Z(n909) );
  AND U854 ( .A(n131), .B(n914), .Z(n913) );
  XNOR U855 ( .A(p_input[517]), .B(n912), .Z(n914) );
  XOR U856 ( .A(n915), .B(n916), .Z(n912) );
  AND U857 ( .A(n135), .B(n917), .Z(n916) );
  XNOR U858 ( .A(p_input[533]), .B(n915), .Z(n917) );
  XOR U859 ( .A(n918), .B(n919), .Z(n915) );
  AND U860 ( .A(n139), .B(n920), .Z(n919) );
  XNOR U861 ( .A(p_input[549]), .B(n918), .Z(n920) );
  XOR U862 ( .A(n921), .B(n922), .Z(n918) );
  AND U863 ( .A(n143), .B(n923), .Z(n922) );
  XNOR U864 ( .A(p_input[565]), .B(n921), .Z(n923) );
  XOR U865 ( .A(n924), .B(n925), .Z(n921) );
  AND U866 ( .A(n147), .B(n926), .Z(n925) );
  XNOR U867 ( .A(p_input[581]), .B(n924), .Z(n926) );
  XOR U868 ( .A(n927), .B(n928), .Z(n924) );
  AND U869 ( .A(n151), .B(n929), .Z(n928) );
  XNOR U870 ( .A(p_input[597]), .B(n927), .Z(n929) );
  XOR U871 ( .A(n930), .B(n931), .Z(n927) );
  AND U872 ( .A(n155), .B(n932), .Z(n931) );
  XNOR U873 ( .A(p_input[613]), .B(n930), .Z(n932) );
  XOR U874 ( .A(n933), .B(n934), .Z(n930) );
  AND U875 ( .A(n159), .B(n935), .Z(n934) );
  XNOR U876 ( .A(p_input[629]), .B(n933), .Z(n935) );
  XOR U877 ( .A(n936), .B(n937), .Z(n933) );
  AND U878 ( .A(n163), .B(n938), .Z(n937) );
  XNOR U879 ( .A(p_input[645]), .B(n936), .Z(n938) );
  XOR U880 ( .A(n939), .B(n940), .Z(n936) );
  AND U881 ( .A(n167), .B(n941), .Z(n940) );
  XNOR U882 ( .A(p_input[661]), .B(n939), .Z(n941) );
  XOR U883 ( .A(n942), .B(n943), .Z(n939) );
  AND U884 ( .A(n171), .B(n944), .Z(n943) );
  XNOR U885 ( .A(p_input[677]), .B(n942), .Z(n944) );
  XOR U886 ( .A(n945), .B(n946), .Z(n942) );
  AND U887 ( .A(n175), .B(n947), .Z(n946) );
  XNOR U888 ( .A(p_input[693]), .B(n945), .Z(n947) );
  XOR U889 ( .A(n948), .B(n949), .Z(n945) );
  AND U890 ( .A(n179), .B(n950), .Z(n949) );
  XNOR U891 ( .A(p_input[709]), .B(n948), .Z(n950) );
  XOR U892 ( .A(n951), .B(n952), .Z(n948) );
  AND U893 ( .A(n183), .B(n953), .Z(n952) );
  XNOR U894 ( .A(p_input[725]), .B(n951), .Z(n953) );
  XOR U895 ( .A(n954), .B(n955), .Z(n951) );
  AND U896 ( .A(n187), .B(n956), .Z(n955) );
  XNOR U897 ( .A(p_input[741]), .B(n954), .Z(n956) );
  XOR U898 ( .A(n957), .B(n958), .Z(n954) );
  AND U899 ( .A(n191), .B(n959), .Z(n958) );
  XNOR U900 ( .A(p_input[757]), .B(n957), .Z(n959) );
  XOR U901 ( .A(n960), .B(n961), .Z(n957) );
  AND U902 ( .A(n195), .B(n962), .Z(n961) );
  XNOR U903 ( .A(p_input[773]), .B(n960), .Z(n962) );
  XOR U904 ( .A(n963), .B(n964), .Z(n960) );
  AND U905 ( .A(n199), .B(n965), .Z(n964) );
  XNOR U906 ( .A(p_input[789]), .B(n963), .Z(n965) );
  XOR U907 ( .A(n966), .B(n967), .Z(n963) );
  AND U908 ( .A(n203), .B(n968), .Z(n967) );
  XNOR U909 ( .A(p_input[805]), .B(n966), .Z(n968) );
  XOR U910 ( .A(n969), .B(n970), .Z(n966) );
  AND U911 ( .A(n207), .B(n971), .Z(n970) );
  XNOR U912 ( .A(p_input[821]), .B(n969), .Z(n971) );
  XOR U913 ( .A(n972), .B(n973), .Z(n969) );
  AND U914 ( .A(n211), .B(n974), .Z(n973) );
  XNOR U915 ( .A(p_input[837]), .B(n972), .Z(n974) );
  XOR U916 ( .A(n975), .B(n976), .Z(n972) );
  AND U917 ( .A(n215), .B(n977), .Z(n976) );
  XNOR U918 ( .A(p_input[853]), .B(n975), .Z(n977) );
  XOR U919 ( .A(n978), .B(n979), .Z(n975) );
  AND U920 ( .A(n219), .B(n980), .Z(n979) );
  XNOR U921 ( .A(p_input[869]), .B(n978), .Z(n980) );
  XOR U922 ( .A(n981), .B(n982), .Z(n978) );
  AND U923 ( .A(n223), .B(n983), .Z(n982) );
  XNOR U924 ( .A(p_input[885]), .B(n981), .Z(n983) );
  XOR U925 ( .A(n984), .B(n985), .Z(n981) );
  AND U926 ( .A(n227), .B(n986), .Z(n985) );
  XNOR U927 ( .A(p_input[901]), .B(n984), .Z(n986) );
  XOR U928 ( .A(n987), .B(n988), .Z(n984) );
  AND U929 ( .A(n231), .B(n989), .Z(n988) );
  XNOR U930 ( .A(p_input[917]), .B(n987), .Z(n989) );
  XOR U931 ( .A(n990), .B(n991), .Z(n987) );
  AND U932 ( .A(n235), .B(n992), .Z(n991) );
  XNOR U933 ( .A(p_input[933]), .B(n990), .Z(n992) );
  XOR U934 ( .A(n993), .B(n994), .Z(n990) );
  AND U935 ( .A(n239), .B(n995), .Z(n994) );
  XNOR U936 ( .A(p_input[949]), .B(n993), .Z(n995) );
  XOR U937 ( .A(n996), .B(n997), .Z(n993) );
  AND U938 ( .A(n243), .B(n998), .Z(n997) );
  XNOR U939 ( .A(p_input[965]), .B(n996), .Z(n998) );
  XNOR U940 ( .A(n999), .B(n1000), .Z(n996) );
  AND U941 ( .A(n247), .B(n1001), .Z(n1000) );
  XOR U942 ( .A(p_input[981]), .B(n999), .Z(n1001) );
  XOR U943 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n1002), .Z(n999) );
  AND U944 ( .A(n250), .B(n1003), .Z(n1002) );
  XOR U945 ( .A(p_input[997]), .B(\knn_comb_/min_val_out[0][5] ), .Z(n1003) );
  XNOR U946 ( .A(n1004), .B(n1005), .Z(o[4]) );
  AND U947 ( .A(n3), .B(n1006), .Z(n1004) );
  XNOR U948 ( .A(p_input[4]), .B(n1005), .Z(n1006) );
  XOR U949 ( .A(n1007), .B(n1008), .Z(n1005) );
  AND U950 ( .A(n7), .B(n1009), .Z(n1008) );
  XNOR U951 ( .A(p_input[20]), .B(n1007), .Z(n1009) );
  XOR U952 ( .A(n1010), .B(n1011), .Z(n1007) );
  AND U953 ( .A(n11), .B(n1012), .Z(n1011) );
  XNOR U954 ( .A(p_input[36]), .B(n1010), .Z(n1012) );
  XOR U955 ( .A(n1013), .B(n1014), .Z(n1010) );
  AND U956 ( .A(n15), .B(n1015), .Z(n1014) );
  XNOR U957 ( .A(p_input[52]), .B(n1013), .Z(n1015) );
  XOR U958 ( .A(n1016), .B(n1017), .Z(n1013) );
  AND U959 ( .A(n19), .B(n1018), .Z(n1017) );
  XNOR U960 ( .A(p_input[68]), .B(n1016), .Z(n1018) );
  XOR U961 ( .A(n1019), .B(n1020), .Z(n1016) );
  AND U962 ( .A(n23), .B(n1021), .Z(n1020) );
  XNOR U963 ( .A(p_input[84]), .B(n1019), .Z(n1021) );
  XOR U964 ( .A(n1022), .B(n1023), .Z(n1019) );
  AND U965 ( .A(n27), .B(n1024), .Z(n1023) );
  XNOR U966 ( .A(p_input[100]), .B(n1022), .Z(n1024) );
  XOR U967 ( .A(n1025), .B(n1026), .Z(n1022) );
  AND U968 ( .A(n31), .B(n1027), .Z(n1026) );
  XNOR U969 ( .A(p_input[116]), .B(n1025), .Z(n1027) );
  XOR U970 ( .A(n1028), .B(n1029), .Z(n1025) );
  AND U971 ( .A(n35), .B(n1030), .Z(n1029) );
  XNOR U972 ( .A(p_input[132]), .B(n1028), .Z(n1030) );
  XOR U973 ( .A(n1031), .B(n1032), .Z(n1028) );
  AND U974 ( .A(n39), .B(n1033), .Z(n1032) );
  XNOR U975 ( .A(p_input[148]), .B(n1031), .Z(n1033) );
  XOR U976 ( .A(n1034), .B(n1035), .Z(n1031) );
  AND U977 ( .A(n43), .B(n1036), .Z(n1035) );
  XNOR U978 ( .A(p_input[164]), .B(n1034), .Z(n1036) );
  XOR U979 ( .A(n1037), .B(n1038), .Z(n1034) );
  AND U980 ( .A(n47), .B(n1039), .Z(n1038) );
  XNOR U981 ( .A(p_input[180]), .B(n1037), .Z(n1039) );
  XOR U982 ( .A(n1040), .B(n1041), .Z(n1037) );
  AND U983 ( .A(n51), .B(n1042), .Z(n1041) );
  XNOR U984 ( .A(p_input[196]), .B(n1040), .Z(n1042) );
  XOR U985 ( .A(n1043), .B(n1044), .Z(n1040) );
  AND U986 ( .A(n55), .B(n1045), .Z(n1044) );
  XNOR U987 ( .A(p_input[212]), .B(n1043), .Z(n1045) );
  XOR U988 ( .A(n1046), .B(n1047), .Z(n1043) );
  AND U989 ( .A(n59), .B(n1048), .Z(n1047) );
  XNOR U990 ( .A(p_input[228]), .B(n1046), .Z(n1048) );
  XOR U991 ( .A(n1049), .B(n1050), .Z(n1046) );
  AND U992 ( .A(n63), .B(n1051), .Z(n1050) );
  XNOR U993 ( .A(p_input[244]), .B(n1049), .Z(n1051) );
  XOR U994 ( .A(n1052), .B(n1053), .Z(n1049) );
  AND U995 ( .A(n67), .B(n1054), .Z(n1053) );
  XNOR U996 ( .A(p_input[260]), .B(n1052), .Z(n1054) );
  XOR U997 ( .A(n1055), .B(n1056), .Z(n1052) );
  AND U998 ( .A(n71), .B(n1057), .Z(n1056) );
  XNOR U999 ( .A(p_input[276]), .B(n1055), .Z(n1057) );
  XOR U1000 ( .A(n1058), .B(n1059), .Z(n1055) );
  AND U1001 ( .A(n75), .B(n1060), .Z(n1059) );
  XNOR U1002 ( .A(p_input[292]), .B(n1058), .Z(n1060) );
  XOR U1003 ( .A(n1061), .B(n1062), .Z(n1058) );
  AND U1004 ( .A(n79), .B(n1063), .Z(n1062) );
  XNOR U1005 ( .A(p_input[308]), .B(n1061), .Z(n1063) );
  XOR U1006 ( .A(n1064), .B(n1065), .Z(n1061) );
  AND U1007 ( .A(n83), .B(n1066), .Z(n1065) );
  XNOR U1008 ( .A(p_input[324]), .B(n1064), .Z(n1066) );
  XOR U1009 ( .A(n1067), .B(n1068), .Z(n1064) );
  AND U1010 ( .A(n87), .B(n1069), .Z(n1068) );
  XNOR U1011 ( .A(p_input[340]), .B(n1067), .Z(n1069) );
  XOR U1012 ( .A(n1070), .B(n1071), .Z(n1067) );
  AND U1013 ( .A(n91), .B(n1072), .Z(n1071) );
  XNOR U1014 ( .A(p_input[356]), .B(n1070), .Z(n1072) );
  XOR U1015 ( .A(n1073), .B(n1074), .Z(n1070) );
  AND U1016 ( .A(n95), .B(n1075), .Z(n1074) );
  XNOR U1017 ( .A(p_input[372]), .B(n1073), .Z(n1075) );
  XOR U1018 ( .A(n1076), .B(n1077), .Z(n1073) );
  AND U1019 ( .A(n99), .B(n1078), .Z(n1077) );
  XNOR U1020 ( .A(p_input[388]), .B(n1076), .Z(n1078) );
  XOR U1021 ( .A(n1079), .B(n1080), .Z(n1076) );
  AND U1022 ( .A(n103), .B(n1081), .Z(n1080) );
  XNOR U1023 ( .A(p_input[404]), .B(n1079), .Z(n1081) );
  XOR U1024 ( .A(n1082), .B(n1083), .Z(n1079) );
  AND U1025 ( .A(n107), .B(n1084), .Z(n1083) );
  XNOR U1026 ( .A(p_input[420]), .B(n1082), .Z(n1084) );
  XOR U1027 ( .A(n1085), .B(n1086), .Z(n1082) );
  AND U1028 ( .A(n111), .B(n1087), .Z(n1086) );
  XNOR U1029 ( .A(p_input[436]), .B(n1085), .Z(n1087) );
  XOR U1030 ( .A(n1088), .B(n1089), .Z(n1085) );
  AND U1031 ( .A(n115), .B(n1090), .Z(n1089) );
  XNOR U1032 ( .A(p_input[452]), .B(n1088), .Z(n1090) );
  XOR U1033 ( .A(n1091), .B(n1092), .Z(n1088) );
  AND U1034 ( .A(n119), .B(n1093), .Z(n1092) );
  XNOR U1035 ( .A(p_input[468]), .B(n1091), .Z(n1093) );
  XOR U1036 ( .A(n1094), .B(n1095), .Z(n1091) );
  AND U1037 ( .A(n123), .B(n1096), .Z(n1095) );
  XNOR U1038 ( .A(p_input[484]), .B(n1094), .Z(n1096) );
  XOR U1039 ( .A(n1097), .B(n1098), .Z(n1094) );
  AND U1040 ( .A(n127), .B(n1099), .Z(n1098) );
  XNOR U1041 ( .A(p_input[500]), .B(n1097), .Z(n1099) );
  XOR U1042 ( .A(n1100), .B(n1101), .Z(n1097) );
  AND U1043 ( .A(n131), .B(n1102), .Z(n1101) );
  XNOR U1044 ( .A(p_input[516]), .B(n1100), .Z(n1102) );
  XOR U1045 ( .A(n1103), .B(n1104), .Z(n1100) );
  AND U1046 ( .A(n135), .B(n1105), .Z(n1104) );
  XNOR U1047 ( .A(p_input[532]), .B(n1103), .Z(n1105) );
  XOR U1048 ( .A(n1106), .B(n1107), .Z(n1103) );
  AND U1049 ( .A(n139), .B(n1108), .Z(n1107) );
  XNOR U1050 ( .A(p_input[548]), .B(n1106), .Z(n1108) );
  XOR U1051 ( .A(n1109), .B(n1110), .Z(n1106) );
  AND U1052 ( .A(n143), .B(n1111), .Z(n1110) );
  XNOR U1053 ( .A(p_input[564]), .B(n1109), .Z(n1111) );
  XOR U1054 ( .A(n1112), .B(n1113), .Z(n1109) );
  AND U1055 ( .A(n147), .B(n1114), .Z(n1113) );
  XNOR U1056 ( .A(p_input[580]), .B(n1112), .Z(n1114) );
  XOR U1057 ( .A(n1115), .B(n1116), .Z(n1112) );
  AND U1058 ( .A(n151), .B(n1117), .Z(n1116) );
  XNOR U1059 ( .A(p_input[596]), .B(n1115), .Z(n1117) );
  XOR U1060 ( .A(n1118), .B(n1119), .Z(n1115) );
  AND U1061 ( .A(n155), .B(n1120), .Z(n1119) );
  XNOR U1062 ( .A(p_input[612]), .B(n1118), .Z(n1120) );
  XOR U1063 ( .A(n1121), .B(n1122), .Z(n1118) );
  AND U1064 ( .A(n159), .B(n1123), .Z(n1122) );
  XNOR U1065 ( .A(p_input[628]), .B(n1121), .Z(n1123) );
  XOR U1066 ( .A(n1124), .B(n1125), .Z(n1121) );
  AND U1067 ( .A(n163), .B(n1126), .Z(n1125) );
  XNOR U1068 ( .A(p_input[644]), .B(n1124), .Z(n1126) );
  XOR U1069 ( .A(n1127), .B(n1128), .Z(n1124) );
  AND U1070 ( .A(n167), .B(n1129), .Z(n1128) );
  XNOR U1071 ( .A(p_input[660]), .B(n1127), .Z(n1129) );
  XOR U1072 ( .A(n1130), .B(n1131), .Z(n1127) );
  AND U1073 ( .A(n171), .B(n1132), .Z(n1131) );
  XNOR U1074 ( .A(p_input[676]), .B(n1130), .Z(n1132) );
  XOR U1075 ( .A(n1133), .B(n1134), .Z(n1130) );
  AND U1076 ( .A(n175), .B(n1135), .Z(n1134) );
  XNOR U1077 ( .A(p_input[692]), .B(n1133), .Z(n1135) );
  XOR U1078 ( .A(n1136), .B(n1137), .Z(n1133) );
  AND U1079 ( .A(n179), .B(n1138), .Z(n1137) );
  XNOR U1080 ( .A(p_input[708]), .B(n1136), .Z(n1138) );
  XOR U1081 ( .A(n1139), .B(n1140), .Z(n1136) );
  AND U1082 ( .A(n183), .B(n1141), .Z(n1140) );
  XNOR U1083 ( .A(p_input[724]), .B(n1139), .Z(n1141) );
  XOR U1084 ( .A(n1142), .B(n1143), .Z(n1139) );
  AND U1085 ( .A(n187), .B(n1144), .Z(n1143) );
  XNOR U1086 ( .A(p_input[740]), .B(n1142), .Z(n1144) );
  XOR U1087 ( .A(n1145), .B(n1146), .Z(n1142) );
  AND U1088 ( .A(n191), .B(n1147), .Z(n1146) );
  XNOR U1089 ( .A(p_input[756]), .B(n1145), .Z(n1147) );
  XOR U1090 ( .A(n1148), .B(n1149), .Z(n1145) );
  AND U1091 ( .A(n195), .B(n1150), .Z(n1149) );
  XNOR U1092 ( .A(p_input[772]), .B(n1148), .Z(n1150) );
  XOR U1093 ( .A(n1151), .B(n1152), .Z(n1148) );
  AND U1094 ( .A(n199), .B(n1153), .Z(n1152) );
  XNOR U1095 ( .A(p_input[788]), .B(n1151), .Z(n1153) );
  XOR U1096 ( .A(n1154), .B(n1155), .Z(n1151) );
  AND U1097 ( .A(n203), .B(n1156), .Z(n1155) );
  XNOR U1098 ( .A(p_input[804]), .B(n1154), .Z(n1156) );
  XOR U1099 ( .A(n1157), .B(n1158), .Z(n1154) );
  AND U1100 ( .A(n207), .B(n1159), .Z(n1158) );
  XNOR U1101 ( .A(p_input[820]), .B(n1157), .Z(n1159) );
  XOR U1102 ( .A(n1160), .B(n1161), .Z(n1157) );
  AND U1103 ( .A(n211), .B(n1162), .Z(n1161) );
  XNOR U1104 ( .A(p_input[836]), .B(n1160), .Z(n1162) );
  XOR U1105 ( .A(n1163), .B(n1164), .Z(n1160) );
  AND U1106 ( .A(n215), .B(n1165), .Z(n1164) );
  XNOR U1107 ( .A(p_input[852]), .B(n1163), .Z(n1165) );
  XOR U1108 ( .A(n1166), .B(n1167), .Z(n1163) );
  AND U1109 ( .A(n219), .B(n1168), .Z(n1167) );
  XNOR U1110 ( .A(p_input[868]), .B(n1166), .Z(n1168) );
  XOR U1111 ( .A(n1169), .B(n1170), .Z(n1166) );
  AND U1112 ( .A(n223), .B(n1171), .Z(n1170) );
  XNOR U1113 ( .A(p_input[884]), .B(n1169), .Z(n1171) );
  XOR U1114 ( .A(n1172), .B(n1173), .Z(n1169) );
  AND U1115 ( .A(n227), .B(n1174), .Z(n1173) );
  XNOR U1116 ( .A(p_input[900]), .B(n1172), .Z(n1174) );
  XOR U1117 ( .A(n1175), .B(n1176), .Z(n1172) );
  AND U1118 ( .A(n231), .B(n1177), .Z(n1176) );
  XNOR U1119 ( .A(p_input[916]), .B(n1175), .Z(n1177) );
  XOR U1120 ( .A(n1178), .B(n1179), .Z(n1175) );
  AND U1121 ( .A(n235), .B(n1180), .Z(n1179) );
  XNOR U1122 ( .A(p_input[932]), .B(n1178), .Z(n1180) );
  XOR U1123 ( .A(n1181), .B(n1182), .Z(n1178) );
  AND U1124 ( .A(n239), .B(n1183), .Z(n1182) );
  XNOR U1125 ( .A(p_input[948]), .B(n1181), .Z(n1183) );
  XOR U1126 ( .A(n1184), .B(n1185), .Z(n1181) );
  AND U1127 ( .A(n243), .B(n1186), .Z(n1185) );
  XNOR U1128 ( .A(p_input[964]), .B(n1184), .Z(n1186) );
  XNOR U1129 ( .A(n1187), .B(n1188), .Z(n1184) );
  AND U1130 ( .A(n247), .B(n1189), .Z(n1188) );
  XOR U1131 ( .A(p_input[980]), .B(n1187), .Z(n1189) );
  XOR U1132 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n1190), .Z(n1187) );
  AND U1133 ( .A(n250), .B(n1191), .Z(n1190) );
  XOR U1134 ( .A(p_input[996]), .B(\knn_comb_/min_val_out[0][4] ), .Z(n1191)
         );
  XNOR U1135 ( .A(n1192), .B(n1193), .Z(o[3]) );
  AND U1136 ( .A(n3), .B(n1194), .Z(n1192) );
  XNOR U1137 ( .A(p_input[3]), .B(n1193), .Z(n1194) );
  XOR U1138 ( .A(n1195), .B(n1196), .Z(n1193) );
  AND U1139 ( .A(n7), .B(n1197), .Z(n1196) );
  XNOR U1140 ( .A(p_input[19]), .B(n1195), .Z(n1197) );
  XOR U1141 ( .A(n1198), .B(n1199), .Z(n1195) );
  AND U1142 ( .A(n11), .B(n1200), .Z(n1199) );
  XNOR U1143 ( .A(p_input[35]), .B(n1198), .Z(n1200) );
  XOR U1144 ( .A(n1201), .B(n1202), .Z(n1198) );
  AND U1145 ( .A(n15), .B(n1203), .Z(n1202) );
  XNOR U1146 ( .A(p_input[51]), .B(n1201), .Z(n1203) );
  XOR U1147 ( .A(n1204), .B(n1205), .Z(n1201) );
  AND U1148 ( .A(n19), .B(n1206), .Z(n1205) );
  XNOR U1149 ( .A(p_input[67]), .B(n1204), .Z(n1206) );
  XOR U1150 ( .A(n1207), .B(n1208), .Z(n1204) );
  AND U1151 ( .A(n23), .B(n1209), .Z(n1208) );
  XNOR U1152 ( .A(p_input[83]), .B(n1207), .Z(n1209) );
  XOR U1153 ( .A(n1210), .B(n1211), .Z(n1207) );
  AND U1154 ( .A(n27), .B(n1212), .Z(n1211) );
  XNOR U1155 ( .A(p_input[99]), .B(n1210), .Z(n1212) );
  XOR U1156 ( .A(n1213), .B(n1214), .Z(n1210) );
  AND U1157 ( .A(n31), .B(n1215), .Z(n1214) );
  XNOR U1158 ( .A(p_input[115]), .B(n1213), .Z(n1215) );
  XOR U1159 ( .A(n1216), .B(n1217), .Z(n1213) );
  AND U1160 ( .A(n35), .B(n1218), .Z(n1217) );
  XNOR U1161 ( .A(p_input[131]), .B(n1216), .Z(n1218) );
  XOR U1162 ( .A(n1219), .B(n1220), .Z(n1216) );
  AND U1163 ( .A(n39), .B(n1221), .Z(n1220) );
  XNOR U1164 ( .A(p_input[147]), .B(n1219), .Z(n1221) );
  XOR U1165 ( .A(n1222), .B(n1223), .Z(n1219) );
  AND U1166 ( .A(n43), .B(n1224), .Z(n1223) );
  XNOR U1167 ( .A(p_input[163]), .B(n1222), .Z(n1224) );
  XOR U1168 ( .A(n1225), .B(n1226), .Z(n1222) );
  AND U1169 ( .A(n47), .B(n1227), .Z(n1226) );
  XNOR U1170 ( .A(p_input[179]), .B(n1225), .Z(n1227) );
  XOR U1171 ( .A(n1228), .B(n1229), .Z(n1225) );
  AND U1172 ( .A(n51), .B(n1230), .Z(n1229) );
  XNOR U1173 ( .A(p_input[195]), .B(n1228), .Z(n1230) );
  XOR U1174 ( .A(n1231), .B(n1232), .Z(n1228) );
  AND U1175 ( .A(n55), .B(n1233), .Z(n1232) );
  XNOR U1176 ( .A(p_input[211]), .B(n1231), .Z(n1233) );
  XOR U1177 ( .A(n1234), .B(n1235), .Z(n1231) );
  AND U1178 ( .A(n59), .B(n1236), .Z(n1235) );
  XNOR U1179 ( .A(p_input[227]), .B(n1234), .Z(n1236) );
  XOR U1180 ( .A(n1237), .B(n1238), .Z(n1234) );
  AND U1181 ( .A(n63), .B(n1239), .Z(n1238) );
  XNOR U1182 ( .A(p_input[243]), .B(n1237), .Z(n1239) );
  XOR U1183 ( .A(n1240), .B(n1241), .Z(n1237) );
  AND U1184 ( .A(n67), .B(n1242), .Z(n1241) );
  XNOR U1185 ( .A(p_input[259]), .B(n1240), .Z(n1242) );
  XOR U1186 ( .A(n1243), .B(n1244), .Z(n1240) );
  AND U1187 ( .A(n71), .B(n1245), .Z(n1244) );
  XNOR U1188 ( .A(p_input[275]), .B(n1243), .Z(n1245) );
  XOR U1189 ( .A(n1246), .B(n1247), .Z(n1243) );
  AND U1190 ( .A(n75), .B(n1248), .Z(n1247) );
  XNOR U1191 ( .A(p_input[291]), .B(n1246), .Z(n1248) );
  XOR U1192 ( .A(n1249), .B(n1250), .Z(n1246) );
  AND U1193 ( .A(n79), .B(n1251), .Z(n1250) );
  XNOR U1194 ( .A(p_input[307]), .B(n1249), .Z(n1251) );
  XOR U1195 ( .A(n1252), .B(n1253), .Z(n1249) );
  AND U1196 ( .A(n83), .B(n1254), .Z(n1253) );
  XNOR U1197 ( .A(p_input[323]), .B(n1252), .Z(n1254) );
  XOR U1198 ( .A(n1255), .B(n1256), .Z(n1252) );
  AND U1199 ( .A(n87), .B(n1257), .Z(n1256) );
  XNOR U1200 ( .A(p_input[339]), .B(n1255), .Z(n1257) );
  XOR U1201 ( .A(n1258), .B(n1259), .Z(n1255) );
  AND U1202 ( .A(n91), .B(n1260), .Z(n1259) );
  XNOR U1203 ( .A(p_input[355]), .B(n1258), .Z(n1260) );
  XOR U1204 ( .A(n1261), .B(n1262), .Z(n1258) );
  AND U1205 ( .A(n95), .B(n1263), .Z(n1262) );
  XNOR U1206 ( .A(p_input[371]), .B(n1261), .Z(n1263) );
  XOR U1207 ( .A(n1264), .B(n1265), .Z(n1261) );
  AND U1208 ( .A(n99), .B(n1266), .Z(n1265) );
  XNOR U1209 ( .A(p_input[387]), .B(n1264), .Z(n1266) );
  XOR U1210 ( .A(n1267), .B(n1268), .Z(n1264) );
  AND U1211 ( .A(n103), .B(n1269), .Z(n1268) );
  XNOR U1212 ( .A(p_input[403]), .B(n1267), .Z(n1269) );
  XOR U1213 ( .A(n1270), .B(n1271), .Z(n1267) );
  AND U1214 ( .A(n107), .B(n1272), .Z(n1271) );
  XNOR U1215 ( .A(p_input[419]), .B(n1270), .Z(n1272) );
  XOR U1216 ( .A(n1273), .B(n1274), .Z(n1270) );
  AND U1217 ( .A(n111), .B(n1275), .Z(n1274) );
  XNOR U1218 ( .A(p_input[435]), .B(n1273), .Z(n1275) );
  XOR U1219 ( .A(n1276), .B(n1277), .Z(n1273) );
  AND U1220 ( .A(n115), .B(n1278), .Z(n1277) );
  XNOR U1221 ( .A(p_input[451]), .B(n1276), .Z(n1278) );
  XOR U1222 ( .A(n1279), .B(n1280), .Z(n1276) );
  AND U1223 ( .A(n119), .B(n1281), .Z(n1280) );
  XNOR U1224 ( .A(p_input[467]), .B(n1279), .Z(n1281) );
  XOR U1225 ( .A(n1282), .B(n1283), .Z(n1279) );
  AND U1226 ( .A(n123), .B(n1284), .Z(n1283) );
  XNOR U1227 ( .A(p_input[483]), .B(n1282), .Z(n1284) );
  XOR U1228 ( .A(n1285), .B(n1286), .Z(n1282) );
  AND U1229 ( .A(n127), .B(n1287), .Z(n1286) );
  XNOR U1230 ( .A(p_input[499]), .B(n1285), .Z(n1287) );
  XOR U1231 ( .A(n1288), .B(n1289), .Z(n1285) );
  AND U1232 ( .A(n131), .B(n1290), .Z(n1289) );
  XNOR U1233 ( .A(p_input[515]), .B(n1288), .Z(n1290) );
  XOR U1234 ( .A(n1291), .B(n1292), .Z(n1288) );
  AND U1235 ( .A(n135), .B(n1293), .Z(n1292) );
  XNOR U1236 ( .A(p_input[531]), .B(n1291), .Z(n1293) );
  XOR U1237 ( .A(n1294), .B(n1295), .Z(n1291) );
  AND U1238 ( .A(n139), .B(n1296), .Z(n1295) );
  XNOR U1239 ( .A(p_input[547]), .B(n1294), .Z(n1296) );
  XOR U1240 ( .A(n1297), .B(n1298), .Z(n1294) );
  AND U1241 ( .A(n143), .B(n1299), .Z(n1298) );
  XNOR U1242 ( .A(p_input[563]), .B(n1297), .Z(n1299) );
  XOR U1243 ( .A(n1300), .B(n1301), .Z(n1297) );
  AND U1244 ( .A(n147), .B(n1302), .Z(n1301) );
  XNOR U1245 ( .A(p_input[579]), .B(n1300), .Z(n1302) );
  XOR U1246 ( .A(n1303), .B(n1304), .Z(n1300) );
  AND U1247 ( .A(n151), .B(n1305), .Z(n1304) );
  XNOR U1248 ( .A(p_input[595]), .B(n1303), .Z(n1305) );
  XOR U1249 ( .A(n1306), .B(n1307), .Z(n1303) );
  AND U1250 ( .A(n155), .B(n1308), .Z(n1307) );
  XNOR U1251 ( .A(p_input[611]), .B(n1306), .Z(n1308) );
  XOR U1252 ( .A(n1309), .B(n1310), .Z(n1306) );
  AND U1253 ( .A(n159), .B(n1311), .Z(n1310) );
  XNOR U1254 ( .A(p_input[627]), .B(n1309), .Z(n1311) );
  XOR U1255 ( .A(n1312), .B(n1313), .Z(n1309) );
  AND U1256 ( .A(n163), .B(n1314), .Z(n1313) );
  XNOR U1257 ( .A(p_input[643]), .B(n1312), .Z(n1314) );
  XOR U1258 ( .A(n1315), .B(n1316), .Z(n1312) );
  AND U1259 ( .A(n167), .B(n1317), .Z(n1316) );
  XNOR U1260 ( .A(p_input[659]), .B(n1315), .Z(n1317) );
  XOR U1261 ( .A(n1318), .B(n1319), .Z(n1315) );
  AND U1262 ( .A(n171), .B(n1320), .Z(n1319) );
  XNOR U1263 ( .A(p_input[675]), .B(n1318), .Z(n1320) );
  XOR U1264 ( .A(n1321), .B(n1322), .Z(n1318) );
  AND U1265 ( .A(n175), .B(n1323), .Z(n1322) );
  XNOR U1266 ( .A(p_input[691]), .B(n1321), .Z(n1323) );
  XOR U1267 ( .A(n1324), .B(n1325), .Z(n1321) );
  AND U1268 ( .A(n179), .B(n1326), .Z(n1325) );
  XNOR U1269 ( .A(p_input[707]), .B(n1324), .Z(n1326) );
  XOR U1270 ( .A(n1327), .B(n1328), .Z(n1324) );
  AND U1271 ( .A(n183), .B(n1329), .Z(n1328) );
  XNOR U1272 ( .A(p_input[723]), .B(n1327), .Z(n1329) );
  XOR U1273 ( .A(n1330), .B(n1331), .Z(n1327) );
  AND U1274 ( .A(n187), .B(n1332), .Z(n1331) );
  XNOR U1275 ( .A(p_input[739]), .B(n1330), .Z(n1332) );
  XOR U1276 ( .A(n1333), .B(n1334), .Z(n1330) );
  AND U1277 ( .A(n191), .B(n1335), .Z(n1334) );
  XNOR U1278 ( .A(p_input[755]), .B(n1333), .Z(n1335) );
  XOR U1279 ( .A(n1336), .B(n1337), .Z(n1333) );
  AND U1280 ( .A(n195), .B(n1338), .Z(n1337) );
  XNOR U1281 ( .A(p_input[771]), .B(n1336), .Z(n1338) );
  XOR U1282 ( .A(n1339), .B(n1340), .Z(n1336) );
  AND U1283 ( .A(n199), .B(n1341), .Z(n1340) );
  XNOR U1284 ( .A(p_input[787]), .B(n1339), .Z(n1341) );
  XOR U1285 ( .A(n1342), .B(n1343), .Z(n1339) );
  AND U1286 ( .A(n203), .B(n1344), .Z(n1343) );
  XNOR U1287 ( .A(p_input[803]), .B(n1342), .Z(n1344) );
  XOR U1288 ( .A(n1345), .B(n1346), .Z(n1342) );
  AND U1289 ( .A(n207), .B(n1347), .Z(n1346) );
  XNOR U1290 ( .A(p_input[819]), .B(n1345), .Z(n1347) );
  XOR U1291 ( .A(n1348), .B(n1349), .Z(n1345) );
  AND U1292 ( .A(n211), .B(n1350), .Z(n1349) );
  XNOR U1293 ( .A(p_input[835]), .B(n1348), .Z(n1350) );
  XOR U1294 ( .A(n1351), .B(n1352), .Z(n1348) );
  AND U1295 ( .A(n215), .B(n1353), .Z(n1352) );
  XNOR U1296 ( .A(p_input[851]), .B(n1351), .Z(n1353) );
  XOR U1297 ( .A(n1354), .B(n1355), .Z(n1351) );
  AND U1298 ( .A(n219), .B(n1356), .Z(n1355) );
  XNOR U1299 ( .A(p_input[867]), .B(n1354), .Z(n1356) );
  XOR U1300 ( .A(n1357), .B(n1358), .Z(n1354) );
  AND U1301 ( .A(n223), .B(n1359), .Z(n1358) );
  XNOR U1302 ( .A(p_input[883]), .B(n1357), .Z(n1359) );
  XOR U1303 ( .A(n1360), .B(n1361), .Z(n1357) );
  AND U1304 ( .A(n227), .B(n1362), .Z(n1361) );
  XNOR U1305 ( .A(p_input[899]), .B(n1360), .Z(n1362) );
  XOR U1306 ( .A(n1363), .B(n1364), .Z(n1360) );
  AND U1307 ( .A(n231), .B(n1365), .Z(n1364) );
  XNOR U1308 ( .A(p_input[915]), .B(n1363), .Z(n1365) );
  XOR U1309 ( .A(n1366), .B(n1367), .Z(n1363) );
  AND U1310 ( .A(n235), .B(n1368), .Z(n1367) );
  XNOR U1311 ( .A(p_input[931]), .B(n1366), .Z(n1368) );
  XOR U1312 ( .A(n1369), .B(n1370), .Z(n1366) );
  AND U1313 ( .A(n239), .B(n1371), .Z(n1370) );
  XNOR U1314 ( .A(p_input[947]), .B(n1369), .Z(n1371) );
  XOR U1315 ( .A(n1372), .B(n1373), .Z(n1369) );
  AND U1316 ( .A(n243), .B(n1374), .Z(n1373) );
  XNOR U1317 ( .A(p_input[963]), .B(n1372), .Z(n1374) );
  XNOR U1318 ( .A(n1375), .B(n1376), .Z(n1372) );
  AND U1319 ( .A(n247), .B(n1377), .Z(n1376) );
  XOR U1320 ( .A(p_input[979]), .B(n1375), .Z(n1377) );
  XOR U1321 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n1378), .Z(n1375) );
  AND U1322 ( .A(n250), .B(n1379), .Z(n1378) );
  XOR U1323 ( .A(p_input[995]), .B(\knn_comb_/min_val_out[0][3] ), .Z(n1379)
         );
  XNOR U1324 ( .A(n1380), .B(n1381), .Z(o[2]) );
  AND U1325 ( .A(n3), .B(n1382), .Z(n1380) );
  XNOR U1326 ( .A(p_input[2]), .B(n1381), .Z(n1382) );
  XOR U1327 ( .A(n1383), .B(n1384), .Z(n1381) );
  AND U1328 ( .A(n7), .B(n1385), .Z(n1384) );
  XNOR U1329 ( .A(p_input[18]), .B(n1383), .Z(n1385) );
  XOR U1330 ( .A(n1386), .B(n1387), .Z(n1383) );
  AND U1331 ( .A(n11), .B(n1388), .Z(n1387) );
  XNOR U1332 ( .A(p_input[34]), .B(n1386), .Z(n1388) );
  XOR U1333 ( .A(n1389), .B(n1390), .Z(n1386) );
  AND U1334 ( .A(n15), .B(n1391), .Z(n1390) );
  XNOR U1335 ( .A(p_input[50]), .B(n1389), .Z(n1391) );
  XOR U1336 ( .A(n1392), .B(n1393), .Z(n1389) );
  AND U1337 ( .A(n19), .B(n1394), .Z(n1393) );
  XNOR U1338 ( .A(p_input[66]), .B(n1392), .Z(n1394) );
  XOR U1339 ( .A(n1395), .B(n1396), .Z(n1392) );
  AND U1340 ( .A(n23), .B(n1397), .Z(n1396) );
  XNOR U1341 ( .A(p_input[82]), .B(n1395), .Z(n1397) );
  XOR U1342 ( .A(n1398), .B(n1399), .Z(n1395) );
  AND U1343 ( .A(n27), .B(n1400), .Z(n1399) );
  XNOR U1344 ( .A(p_input[98]), .B(n1398), .Z(n1400) );
  XOR U1345 ( .A(n1401), .B(n1402), .Z(n1398) );
  AND U1346 ( .A(n31), .B(n1403), .Z(n1402) );
  XNOR U1347 ( .A(p_input[114]), .B(n1401), .Z(n1403) );
  XOR U1348 ( .A(n1404), .B(n1405), .Z(n1401) );
  AND U1349 ( .A(n35), .B(n1406), .Z(n1405) );
  XNOR U1350 ( .A(p_input[130]), .B(n1404), .Z(n1406) );
  XOR U1351 ( .A(n1407), .B(n1408), .Z(n1404) );
  AND U1352 ( .A(n39), .B(n1409), .Z(n1408) );
  XNOR U1353 ( .A(p_input[146]), .B(n1407), .Z(n1409) );
  XOR U1354 ( .A(n1410), .B(n1411), .Z(n1407) );
  AND U1355 ( .A(n43), .B(n1412), .Z(n1411) );
  XNOR U1356 ( .A(p_input[162]), .B(n1410), .Z(n1412) );
  XOR U1357 ( .A(n1413), .B(n1414), .Z(n1410) );
  AND U1358 ( .A(n47), .B(n1415), .Z(n1414) );
  XNOR U1359 ( .A(p_input[178]), .B(n1413), .Z(n1415) );
  XOR U1360 ( .A(n1416), .B(n1417), .Z(n1413) );
  AND U1361 ( .A(n51), .B(n1418), .Z(n1417) );
  XNOR U1362 ( .A(p_input[194]), .B(n1416), .Z(n1418) );
  XOR U1363 ( .A(n1419), .B(n1420), .Z(n1416) );
  AND U1364 ( .A(n55), .B(n1421), .Z(n1420) );
  XNOR U1365 ( .A(p_input[210]), .B(n1419), .Z(n1421) );
  XOR U1366 ( .A(n1422), .B(n1423), .Z(n1419) );
  AND U1367 ( .A(n59), .B(n1424), .Z(n1423) );
  XNOR U1368 ( .A(p_input[226]), .B(n1422), .Z(n1424) );
  XOR U1369 ( .A(n1425), .B(n1426), .Z(n1422) );
  AND U1370 ( .A(n63), .B(n1427), .Z(n1426) );
  XNOR U1371 ( .A(p_input[242]), .B(n1425), .Z(n1427) );
  XOR U1372 ( .A(n1428), .B(n1429), .Z(n1425) );
  AND U1373 ( .A(n67), .B(n1430), .Z(n1429) );
  XNOR U1374 ( .A(p_input[258]), .B(n1428), .Z(n1430) );
  XOR U1375 ( .A(n1431), .B(n1432), .Z(n1428) );
  AND U1376 ( .A(n71), .B(n1433), .Z(n1432) );
  XNOR U1377 ( .A(p_input[274]), .B(n1431), .Z(n1433) );
  XOR U1378 ( .A(n1434), .B(n1435), .Z(n1431) );
  AND U1379 ( .A(n75), .B(n1436), .Z(n1435) );
  XNOR U1380 ( .A(p_input[290]), .B(n1434), .Z(n1436) );
  XOR U1381 ( .A(n1437), .B(n1438), .Z(n1434) );
  AND U1382 ( .A(n79), .B(n1439), .Z(n1438) );
  XNOR U1383 ( .A(p_input[306]), .B(n1437), .Z(n1439) );
  XOR U1384 ( .A(n1440), .B(n1441), .Z(n1437) );
  AND U1385 ( .A(n83), .B(n1442), .Z(n1441) );
  XNOR U1386 ( .A(p_input[322]), .B(n1440), .Z(n1442) );
  XOR U1387 ( .A(n1443), .B(n1444), .Z(n1440) );
  AND U1388 ( .A(n87), .B(n1445), .Z(n1444) );
  XNOR U1389 ( .A(p_input[338]), .B(n1443), .Z(n1445) );
  XOR U1390 ( .A(n1446), .B(n1447), .Z(n1443) );
  AND U1391 ( .A(n91), .B(n1448), .Z(n1447) );
  XNOR U1392 ( .A(p_input[354]), .B(n1446), .Z(n1448) );
  XOR U1393 ( .A(n1449), .B(n1450), .Z(n1446) );
  AND U1394 ( .A(n95), .B(n1451), .Z(n1450) );
  XNOR U1395 ( .A(p_input[370]), .B(n1449), .Z(n1451) );
  XOR U1396 ( .A(n1452), .B(n1453), .Z(n1449) );
  AND U1397 ( .A(n99), .B(n1454), .Z(n1453) );
  XNOR U1398 ( .A(p_input[386]), .B(n1452), .Z(n1454) );
  XOR U1399 ( .A(n1455), .B(n1456), .Z(n1452) );
  AND U1400 ( .A(n103), .B(n1457), .Z(n1456) );
  XNOR U1401 ( .A(p_input[402]), .B(n1455), .Z(n1457) );
  XOR U1402 ( .A(n1458), .B(n1459), .Z(n1455) );
  AND U1403 ( .A(n107), .B(n1460), .Z(n1459) );
  XNOR U1404 ( .A(p_input[418]), .B(n1458), .Z(n1460) );
  XOR U1405 ( .A(n1461), .B(n1462), .Z(n1458) );
  AND U1406 ( .A(n111), .B(n1463), .Z(n1462) );
  XNOR U1407 ( .A(p_input[434]), .B(n1461), .Z(n1463) );
  XOR U1408 ( .A(n1464), .B(n1465), .Z(n1461) );
  AND U1409 ( .A(n115), .B(n1466), .Z(n1465) );
  XNOR U1410 ( .A(p_input[450]), .B(n1464), .Z(n1466) );
  XOR U1411 ( .A(n1467), .B(n1468), .Z(n1464) );
  AND U1412 ( .A(n119), .B(n1469), .Z(n1468) );
  XNOR U1413 ( .A(p_input[466]), .B(n1467), .Z(n1469) );
  XOR U1414 ( .A(n1470), .B(n1471), .Z(n1467) );
  AND U1415 ( .A(n123), .B(n1472), .Z(n1471) );
  XNOR U1416 ( .A(p_input[482]), .B(n1470), .Z(n1472) );
  XOR U1417 ( .A(n1473), .B(n1474), .Z(n1470) );
  AND U1418 ( .A(n127), .B(n1475), .Z(n1474) );
  XNOR U1419 ( .A(p_input[498]), .B(n1473), .Z(n1475) );
  XOR U1420 ( .A(n1476), .B(n1477), .Z(n1473) );
  AND U1421 ( .A(n131), .B(n1478), .Z(n1477) );
  XNOR U1422 ( .A(p_input[514]), .B(n1476), .Z(n1478) );
  XOR U1423 ( .A(n1479), .B(n1480), .Z(n1476) );
  AND U1424 ( .A(n135), .B(n1481), .Z(n1480) );
  XNOR U1425 ( .A(p_input[530]), .B(n1479), .Z(n1481) );
  XOR U1426 ( .A(n1482), .B(n1483), .Z(n1479) );
  AND U1427 ( .A(n139), .B(n1484), .Z(n1483) );
  XNOR U1428 ( .A(p_input[546]), .B(n1482), .Z(n1484) );
  XOR U1429 ( .A(n1485), .B(n1486), .Z(n1482) );
  AND U1430 ( .A(n143), .B(n1487), .Z(n1486) );
  XNOR U1431 ( .A(p_input[562]), .B(n1485), .Z(n1487) );
  XOR U1432 ( .A(n1488), .B(n1489), .Z(n1485) );
  AND U1433 ( .A(n147), .B(n1490), .Z(n1489) );
  XNOR U1434 ( .A(p_input[578]), .B(n1488), .Z(n1490) );
  XOR U1435 ( .A(n1491), .B(n1492), .Z(n1488) );
  AND U1436 ( .A(n151), .B(n1493), .Z(n1492) );
  XNOR U1437 ( .A(p_input[594]), .B(n1491), .Z(n1493) );
  XOR U1438 ( .A(n1494), .B(n1495), .Z(n1491) );
  AND U1439 ( .A(n155), .B(n1496), .Z(n1495) );
  XNOR U1440 ( .A(p_input[610]), .B(n1494), .Z(n1496) );
  XOR U1441 ( .A(n1497), .B(n1498), .Z(n1494) );
  AND U1442 ( .A(n159), .B(n1499), .Z(n1498) );
  XNOR U1443 ( .A(p_input[626]), .B(n1497), .Z(n1499) );
  XOR U1444 ( .A(n1500), .B(n1501), .Z(n1497) );
  AND U1445 ( .A(n163), .B(n1502), .Z(n1501) );
  XNOR U1446 ( .A(p_input[642]), .B(n1500), .Z(n1502) );
  XOR U1447 ( .A(n1503), .B(n1504), .Z(n1500) );
  AND U1448 ( .A(n167), .B(n1505), .Z(n1504) );
  XNOR U1449 ( .A(p_input[658]), .B(n1503), .Z(n1505) );
  XOR U1450 ( .A(n1506), .B(n1507), .Z(n1503) );
  AND U1451 ( .A(n171), .B(n1508), .Z(n1507) );
  XNOR U1452 ( .A(p_input[674]), .B(n1506), .Z(n1508) );
  XOR U1453 ( .A(n1509), .B(n1510), .Z(n1506) );
  AND U1454 ( .A(n175), .B(n1511), .Z(n1510) );
  XNOR U1455 ( .A(p_input[690]), .B(n1509), .Z(n1511) );
  XOR U1456 ( .A(n1512), .B(n1513), .Z(n1509) );
  AND U1457 ( .A(n179), .B(n1514), .Z(n1513) );
  XNOR U1458 ( .A(p_input[706]), .B(n1512), .Z(n1514) );
  XOR U1459 ( .A(n1515), .B(n1516), .Z(n1512) );
  AND U1460 ( .A(n183), .B(n1517), .Z(n1516) );
  XNOR U1461 ( .A(p_input[722]), .B(n1515), .Z(n1517) );
  XOR U1462 ( .A(n1518), .B(n1519), .Z(n1515) );
  AND U1463 ( .A(n187), .B(n1520), .Z(n1519) );
  XNOR U1464 ( .A(p_input[738]), .B(n1518), .Z(n1520) );
  XOR U1465 ( .A(n1521), .B(n1522), .Z(n1518) );
  AND U1466 ( .A(n191), .B(n1523), .Z(n1522) );
  XNOR U1467 ( .A(p_input[754]), .B(n1521), .Z(n1523) );
  XOR U1468 ( .A(n1524), .B(n1525), .Z(n1521) );
  AND U1469 ( .A(n195), .B(n1526), .Z(n1525) );
  XNOR U1470 ( .A(p_input[770]), .B(n1524), .Z(n1526) );
  XOR U1471 ( .A(n1527), .B(n1528), .Z(n1524) );
  AND U1472 ( .A(n199), .B(n1529), .Z(n1528) );
  XNOR U1473 ( .A(p_input[786]), .B(n1527), .Z(n1529) );
  XOR U1474 ( .A(n1530), .B(n1531), .Z(n1527) );
  AND U1475 ( .A(n203), .B(n1532), .Z(n1531) );
  XNOR U1476 ( .A(p_input[802]), .B(n1530), .Z(n1532) );
  XOR U1477 ( .A(n1533), .B(n1534), .Z(n1530) );
  AND U1478 ( .A(n207), .B(n1535), .Z(n1534) );
  XNOR U1479 ( .A(p_input[818]), .B(n1533), .Z(n1535) );
  XOR U1480 ( .A(n1536), .B(n1537), .Z(n1533) );
  AND U1481 ( .A(n211), .B(n1538), .Z(n1537) );
  XNOR U1482 ( .A(p_input[834]), .B(n1536), .Z(n1538) );
  XOR U1483 ( .A(n1539), .B(n1540), .Z(n1536) );
  AND U1484 ( .A(n215), .B(n1541), .Z(n1540) );
  XNOR U1485 ( .A(p_input[850]), .B(n1539), .Z(n1541) );
  XOR U1486 ( .A(n1542), .B(n1543), .Z(n1539) );
  AND U1487 ( .A(n219), .B(n1544), .Z(n1543) );
  XNOR U1488 ( .A(p_input[866]), .B(n1542), .Z(n1544) );
  XOR U1489 ( .A(n1545), .B(n1546), .Z(n1542) );
  AND U1490 ( .A(n223), .B(n1547), .Z(n1546) );
  XNOR U1491 ( .A(p_input[882]), .B(n1545), .Z(n1547) );
  XOR U1492 ( .A(n1548), .B(n1549), .Z(n1545) );
  AND U1493 ( .A(n227), .B(n1550), .Z(n1549) );
  XNOR U1494 ( .A(p_input[898]), .B(n1548), .Z(n1550) );
  XOR U1495 ( .A(n1551), .B(n1552), .Z(n1548) );
  AND U1496 ( .A(n231), .B(n1553), .Z(n1552) );
  XNOR U1497 ( .A(p_input[914]), .B(n1551), .Z(n1553) );
  XOR U1498 ( .A(n1554), .B(n1555), .Z(n1551) );
  AND U1499 ( .A(n235), .B(n1556), .Z(n1555) );
  XNOR U1500 ( .A(p_input[930]), .B(n1554), .Z(n1556) );
  XOR U1501 ( .A(n1557), .B(n1558), .Z(n1554) );
  AND U1502 ( .A(n239), .B(n1559), .Z(n1558) );
  XNOR U1503 ( .A(p_input[946]), .B(n1557), .Z(n1559) );
  XOR U1504 ( .A(n1560), .B(n1561), .Z(n1557) );
  AND U1505 ( .A(n243), .B(n1562), .Z(n1561) );
  XNOR U1506 ( .A(p_input[962]), .B(n1560), .Z(n1562) );
  XNOR U1507 ( .A(n1563), .B(n1564), .Z(n1560) );
  AND U1508 ( .A(n247), .B(n1565), .Z(n1564) );
  XOR U1509 ( .A(p_input[978]), .B(n1563), .Z(n1565) );
  XOR U1510 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n1566), .Z(n1563) );
  AND U1511 ( .A(n250), .B(n1567), .Z(n1566) );
  XOR U1512 ( .A(p_input[994]), .B(\knn_comb_/min_val_out[0][2] ), .Z(n1567)
         );
  XNOR U1513 ( .A(n1568), .B(n1569), .Z(o[1]) );
  AND U1514 ( .A(n3), .B(n1570), .Z(n1568) );
  XNOR U1515 ( .A(p_input[1]), .B(n1569), .Z(n1570) );
  XOR U1516 ( .A(n1571), .B(n1572), .Z(n1569) );
  AND U1517 ( .A(n7), .B(n1573), .Z(n1572) );
  XNOR U1518 ( .A(p_input[17]), .B(n1571), .Z(n1573) );
  XOR U1519 ( .A(n1574), .B(n1575), .Z(n1571) );
  AND U1520 ( .A(n11), .B(n1576), .Z(n1575) );
  XNOR U1521 ( .A(p_input[33]), .B(n1574), .Z(n1576) );
  XOR U1522 ( .A(n1577), .B(n1578), .Z(n1574) );
  AND U1523 ( .A(n15), .B(n1579), .Z(n1578) );
  XNOR U1524 ( .A(p_input[49]), .B(n1577), .Z(n1579) );
  XOR U1525 ( .A(n1580), .B(n1581), .Z(n1577) );
  AND U1526 ( .A(n19), .B(n1582), .Z(n1581) );
  XNOR U1527 ( .A(p_input[65]), .B(n1580), .Z(n1582) );
  XOR U1528 ( .A(n1583), .B(n1584), .Z(n1580) );
  AND U1529 ( .A(n23), .B(n1585), .Z(n1584) );
  XNOR U1530 ( .A(p_input[81]), .B(n1583), .Z(n1585) );
  XOR U1531 ( .A(n1586), .B(n1587), .Z(n1583) );
  AND U1532 ( .A(n27), .B(n1588), .Z(n1587) );
  XNOR U1533 ( .A(p_input[97]), .B(n1586), .Z(n1588) );
  XOR U1534 ( .A(n1589), .B(n1590), .Z(n1586) );
  AND U1535 ( .A(n31), .B(n1591), .Z(n1590) );
  XNOR U1536 ( .A(p_input[113]), .B(n1589), .Z(n1591) );
  XOR U1537 ( .A(n1592), .B(n1593), .Z(n1589) );
  AND U1538 ( .A(n35), .B(n1594), .Z(n1593) );
  XNOR U1539 ( .A(p_input[129]), .B(n1592), .Z(n1594) );
  XOR U1540 ( .A(n1595), .B(n1596), .Z(n1592) );
  AND U1541 ( .A(n39), .B(n1597), .Z(n1596) );
  XNOR U1542 ( .A(p_input[145]), .B(n1595), .Z(n1597) );
  XOR U1543 ( .A(n1598), .B(n1599), .Z(n1595) );
  AND U1544 ( .A(n43), .B(n1600), .Z(n1599) );
  XNOR U1545 ( .A(p_input[161]), .B(n1598), .Z(n1600) );
  XOR U1546 ( .A(n1601), .B(n1602), .Z(n1598) );
  AND U1547 ( .A(n47), .B(n1603), .Z(n1602) );
  XNOR U1548 ( .A(p_input[177]), .B(n1601), .Z(n1603) );
  XOR U1549 ( .A(n1604), .B(n1605), .Z(n1601) );
  AND U1550 ( .A(n51), .B(n1606), .Z(n1605) );
  XNOR U1551 ( .A(p_input[193]), .B(n1604), .Z(n1606) );
  XOR U1552 ( .A(n1607), .B(n1608), .Z(n1604) );
  AND U1553 ( .A(n55), .B(n1609), .Z(n1608) );
  XNOR U1554 ( .A(p_input[209]), .B(n1607), .Z(n1609) );
  XOR U1555 ( .A(n1610), .B(n1611), .Z(n1607) );
  AND U1556 ( .A(n59), .B(n1612), .Z(n1611) );
  XNOR U1557 ( .A(p_input[225]), .B(n1610), .Z(n1612) );
  XOR U1558 ( .A(n1613), .B(n1614), .Z(n1610) );
  AND U1559 ( .A(n63), .B(n1615), .Z(n1614) );
  XNOR U1560 ( .A(p_input[241]), .B(n1613), .Z(n1615) );
  XOR U1561 ( .A(n1616), .B(n1617), .Z(n1613) );
  AND U1562 ( .A(n67), .B(n1618), .Z(n1617) );
  XNOR U1563 ( .A(p_input[257]), .B(n1616), .Z(n1618) );
  XOR U1564 ( .A(n1619), .B(n1620), .Z(n1616) );
  AND U1565 ( .A(n71), .B(n1621), .Z(n1620) );
  XNOR U1566 ( .A(p_input[273]), .B(n1619), .Z(n1621) );
  XOR U1567 ( .A(n1622), .B(n1623), .Z(n1619) );
  AND U1568 ( .A(n75), .B(n1624), .Z(n1623) );
  XNOR U1569 ( .A(p_input[289]), .B(n1622), .Z(n1624) );
  XOR U1570 ( .A(n1625), .B(n1626), .Z(n1622) );
  AND U1571 ( .A(n79), .B(n1627), .Z(n1626) );
  XNOR U1572 ( .A(p_input[305]), .B(n1625), .Z(n1627) );
  XOR U1573 ( .A(n1628), .B(n1629), .Z(n1625) );
  AND U1574 ( .A(n83), .B(n1630), .Z(n1629) );
  XNOR U1575 ( .A(p_input[321]), .B(n1628), .Z(n1630) );
  XOR U1576 ( .A(n1631), .B(n1632), .Z(n1628) );
  AND U1577 ( .A(n87), .B(n1633), .Z(n1632) );
  XNOR U1578 ( .A(p_input[337]), .B(n1631), .Z(n1633) );
  XOR U1579 ( .A(n1634), .B(n1635), .Z(n1631) );
  AND U1580 ( .A(n91), .B(n1636), .Z(n1635) );
  XNOR U1581 ( .A(p_input[353]), .B(n1634), .Z(n1636) );
  XOR U1582 ( .A(n1637), .B(n1638), .Z(n1634) );
  AND U1583 ( .A(n95), .B(n1639), .Z(n1638) );
  XNOR U1584 ( .A(p_input[369]), .B(n1637), .Z(n1639) );
  XOR U1585 ( .A(n1640), .B(n1641), .Z(n1637) );
  AND U1586 ( .A(n99), .B(n1642), .Z(n1641) );
  XNOR U1587 ( .A(p_input[385]), .B(n1640), .Z(n1642) );
  XOR U1588 ( .A(n1643), .B(n1644), .Z(n1640) );
  AND U1589 ( .A(n103), .B(n1645), .Z(n1644) );
  XNOR U1590 ( .A(p_input[401]), .B(n1643), .Z(n1645) );
  XOR U1591 ( .A(n1646), .B(n1647), .Z(n1643) );
  AND U1592 ( .A(n107), .B(n1648), .Z(n1647) );
  XNOR U1593 ( .A(p_input[417]), .B(n1646), .Z(n1648) );
  XOR U1594 ( .A(n1649), .B(n1650), .Z(n1646) );
  AND U1595 ( .A(n111), .B(n1651), .Z(n1650) );
  XNOR U1596 ( .A(p_input[433]), .B(n1649), .Z(n1651) );
  XOR U1597 ( .A(n1652), .B(n1653), .Z(n1649) );
  AND U1598 ( .A(n115), .B(n1654), .Z(n1653) );
  XNOR U1599 ( .A(p_input[449]), .B(n1652), .Z(n1654) );
  XOR U1600 ( .A(n1655), .B(n1656), .Z(n1652) );
  AND U1601 ( .A(n119), .B(n1657), .Z(n1656) );
  XNOR U1602 ( .A(p_input[465]), .B(n1655), .Z(n1657) );
  XOR U1603 ( .A(n1658), .B(n1659), .Z(n1655) );
  AND U1604 ( .A(n123), .B(n1660), .Z(n1659) );
  XNOR U1605 ( .A(p_input[481]), .B(n1658), .Z(n1660) );
  XOR U1606 ( .A(n1661), .B(n1662), .Z(n1658) );
  AND U1607 ( .A(n127), .B(n1663), .Z(n1662) );
  XNOR U1608 ( .A(p_input[497]), .B(n1661), .Z(n1663) );
  XOR U1609 ( .A(n1664), .B(n1665), .Z(n1661) );
  AND U1610 ( .A(n131), .B(n1666), .Z(n1665) );
  XNOR U1611 ( .A(p_input[513]), .B(n1664), .Z(n1666) );
  XOR U1612 ( .A(n1667), .B(n1668), .Z(n1664) );
  AND U1613 ( .A(n135), .B(n1669), .Z(n1668) );
  XNOR U1614 ( .A(p_input[529]), .B(n1667), .Z(n1669) );
  XOR U1615 ( .A(n1670), .B(n1671), .Z(n1667) );
  AND U1616 ( .A(n139), .B(n1672), .Z(n1671) );
  XNOR U1617 ( .A(p_input[545]), .B(n1670), .Z(n1672) );
  XOR U1618 ( .A(n1673), .B(n1674), .Z(n1670) );
  AND U1619 ( .A(n143), .B(n1675), .Z(n1674) );
  XNOR U1620 ( .A(p_input[561]), .B(n1673), .Z(n1675) );
  XOR U1621 ( .A(n1676), .B(n1677), .Z(n1673) );
  AND U1622 ( .A(n147), .B(n1678), .Z(n1677) );
  XNOR U1623 ( .A(p_input[577]), .B(n1676), .Z(n1678) );
  XOR U1624 ( .A(n1679), .B(n1680), .Z(n1676) );
  AND U1625 ( .A(n151), .B(n1681), .Z(n1680) );
  XNOR U1626 ( .A(p_input[593]), .B(n1679), .Z(n1681) );
  XOR U1627 ( .A(n1682), .B(n1683), .Z(n1679) );
  AND U1628 ( .A(n155), .B(n1684), .Z(n1683) );
  XNOR U1629 ( .A(p_input[609]), .B(n1682), .Z(n1684) );
  XOR U1630 ( .A(n1685), .B(n1686), .Z(n1682) );
  AND U1631 ( .A(n159), .B(n1687), .Z(n1686) );
  XNOR U1632 ( .A(p_input[625]), .B(n1685), .Z(n1687) );
  XOR U1633 ( .A(n1688), .B(n1689), .Z(n1685) );
  AND U1634 ( .A(n163), .B(n1690), .Z(n1689) );
  XNOR U1635 ( .A(p_input[641]), .B(n1688), .Z(n1690) );
  XOR U1636 ( .A(n1691), .B(n1692), .Z(n1688) );
  AND U1637 ( .A(n167), .B(n1693), .Z(n1692) );
  XNOR U1638 ( .A(p_input[657]), .B(n1691), .Z(n1693) );
  XOR U1639 ( .A(n1694), .B(n1695), .Z(n1691) );
  AND U1640 ( .A(n171), .B(n1696), .Z(n1695) );
  XNOR U1641 ( .A(p_input[673]), .B(n1694), .Z(n1696) );
  XOR U1642 ( .A(n1697), .B(n1698), .Z(n1694) );
  AND U1643 ( .A(n175), .B(n1699), .Z(n1698) );
  XNOR U1644 ( .A(p_input[689]), .B(n1697), .Z(n1699) );
  XOR U1645 ( .A(n1700), .B(n1701), .Z(n1697) );
  AND U1646 ( .A(n179), .B(n1702), .Z(n1701) );
  XNOR U1647 ( .A(p_input[705]), .B(n1700), .Z(n1702) );
  XOR U1648 ( .A(n1703), .B(n1704), .Z(n1700) );
  AND U1649 ( .A(n183), .B(n1705), .Z(n1704) );
  XNOR U1650 ( .A(p_input[721]), .B(n1703), .Z(n1705) );
  XOR U1651 ( .A(n1706), .B(n1707), .Z(n1703) );
  AND U1652 ( .A(n187), .B(n1708), .Z(n1707) );
  XNOR U1653 ( .A(p_input[737]), .B(n1706), .Z(n1708) );
  XOR U1654 ( .A(n1709), .B(n1710), .Z(n1706) );
  AND U1655 ( .A(n191), .B(n1711), .Z(n1710) );
  XNOR U1656 ( .A(p_input[753]), .B(n1709), .Z(n1711) );
  XOR U1657 ( .A(n1712), .B(n1713), .Z(n1709) );
  AND U1658 ( .A(n195), .B(n1714), .Z(n1713) );
  XNOR U1659 ( .A(p_input[769]), .B(n1712), .Z(n1714) );
  XOR U1660 ( .A(n1715), .B(n1716), .Z(n1712) );
  AND U1661 ( .A(n199), .B(n1717), .Z(n1716) );
  XNOR U1662 ( .A(p_input[785]), .B(n1715), .Z(n1717) );
  XOR U1663 ( .A(n1718), .B(n1719), .Z(n1715) );
  AND U1664 ( .A(n203), .B(n1720), .Z(n1719) );
  XNOR U1665 ( .A(p_input[801]), .B(n1718), .Z(n1720) );
  XOR U1666 ( .A(n1721), .B(n1722), .Z(n1718) );
  AND U1667 ( .A(n207), .B(n1723), .Z(n1722) );
  XNOR U1668 ( .A(p_input[817]), .B(n1721), .Z(n1723) );
  XOR U1669 ( .A(n1724), .B(n1725), .Z(n1721) );
  AND U1670 ( .A(n211), .B(n1726), .Z(n1725) );
  XNOR U1671 ( .A(p_input[833]), .B(n1724), .Z(n1726) );
  XOR U1672 ( .A(n1727), .B(n1728), .Z(n1724) );
  AND U1673 ( .A(n215), .B(n1729), .Z(n1728) );
  XNOR U1674 ( .A(p_input[849]), .B(n1727), .Z(n1729) );
  XOR U1675 ( .A(n1730), .B(n1731), .Z(n1727) );
  AND U1676 ( .A(n219), .B(n1732), .Z(n1731) );
  XNOR U1677 ( .A(p_input[865]), .B(n1730), .Z(n1732) );
  XOR U1678 ( .A(n1733), .B(n1734), .Z(n1730) );
  AND U1679 ( .A(n223), .B(n1735), .Z(n1734) );
  XNOR U1680 ( .A(p_input[881]), .B(n1733), .Z(n1735) );
  XOR U1681 ( .A(n1736), .B(n1737), .Z(n1733) );
  AND U1682 ( .A(n227), .B(n1738), .Z(n1737) );
  XNOR U1683 ( .A(p_input[897]), .B(n1736), .Z(n1738) );
  XOR U1684 ( .A(n1739), .B(n1740), .Z(n1736) );
  AND U1685 ( .A(n231), .B(n1741), .Z(n1740) );
  XNOR U1686 ( .A(p_input[913]), .B(n1739), .Z(n1741) );
  XOR U1687 ( .A(n1742), .B(n1743), .Z(n1739) );
  AND U1688 ( .A(n235), .B(n1744), .Z(n1743) );
  XNOR U1689 ( .A(p_input[929]), .B(n1742), .Z(n1744) );
  XOR U1690 ( .A(n1745), .B(n1746), .Z(n1742) );
  AND U1691 ( .A(n239), .B(n1747), .Z(n1746) );
  XNOR U1692 ( .A(p_input[945]), .B(n1745), .Z(n1747) );
  XOR U1693 ( .A(n1748), .B(n1749), .Z(n1745) );
  AND U1694 ( .A(n243), .B(n1750), .Z(n1749) );
  XNOR U1695 ( .A(p_input[961]), .B(n1748), .Z(n1750) );
  XNOR U1696 ( .A(n1751), .B(n1752), .Z(n1748) );
  AND U1697 ( .A(n247), .B(n1753), .Z(n1752) );
  XOR U1698 ( .A(p_input[977]), .B(n1751), .Z(n1753) );
  XOR U1699 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n1754), .Z(n1751) );
  AND U1700 ( .A(n250), .B(n1755), .Z(n1754) );
  XOR U1701 ( .A(p_input[993]), .B(\knn_comb_/min_val_out[0][1] ), .Z(n1755)
         );
  XNOR U1702 ( .A(n1756), .B(n1757), .Z(o[15]) );
  AND U1703 ( .A(n3), .B(n1758), .Z(n1756) );
  XNOR U1704 ( .A(p_input[15]), .B(n1757), .Z(n1758) );
  XOR U1705 ( .A(n1759), .B(n1760), .Z(n1757) );
  AND U1706 ( .A(n7), .B(n1761), .Z(n1760) );
  XNOR U1707 ( .A(p_input[31]), .B(n1759), .Z(n1761) );
  XOR U1708 ( .A(n1762), .B(n1763), .Z(n1759) );
  AND U1709 ( .A(n11), .B(n1764), .Z(n1763) );
  XNOR U1710 ( .A(p_input[47]), .B(n1762), .Z(n1764) );
  XOR U1711 ( .A(n1765), .B(n1766), .Z(n1762) );
  AND U1712 ( .A(n15), .B(n1767), .Z(n1766) );
  XNOR U1713 ( .A(p_input[63]), .B(n1765), .Z(n1767) );
  XOR U1714 ( .A(n1768), .B(n1769), .Z(n1765) );
  AND U1715 ( .A(n19), .B(n1770), .Z(n1769) );
  XNOR U1716 ( .A(p_input[79]), .B(n1768), .Z(n1770) );
  XOR U1717 ( .A(n1771), .B(n1772), .Z(n1768) );
  AND U1718 ( .A(n23), .B(n1773), .Z(n1772) );
  XNOR U1719 ( .A(p_input[95]), .B(n1771), .Z(n1773) );
  XOR U1720 ( .A(n1774), .B(n1775), .Z(n1771) );
  AND U1721 ( .A(n27), .B(n1776), .Z(n1775) );
  XNOR U1722 ( .A(p_input[111]), .B(n1774), .Z(n1776) );
  XOR U1723 ( .A(n1777), .B(n1778), .Z(n1774) );
  AND U1724 ( .A(n31), .B(n1779), .Z(n1778) );
  XNOR U1725 ( .A(p_input[127]), .B(n1777), .Z(n1779) );
  XOR U1726 ( .A(n1780), .B(n1781), .Z(n1777) );
  AND U1727 ( .A(n35), .B(n1782), .Z(n1781) );
  XNOR U1728 ( .A(p_input[143]), .B(n1780), .Z(n1782) );
  XOR U1729 ( .A(n1783), .B(n1784), .Z(n1780) );
  AND U1730 ( .A(n39), .B(n1785), .Z(n1784) );
  XNOR U1731 ( .A(p_input[159]), .B(n1783), .Z(n1785) );
  XOR U1732 ( .A(n1786), .B(n1787), .Z(n1783) );
  AND U1733 ( .A(n43), .B(n1788), .Z(n1787) );
  XNOR U1734 ( .A(p_input[175]), .B(n1786), .Z(n1788) );
  XOR U1735 ( .A(n1789), .B(n1790), .Z(n1786) );
  AND U1736 ( .A(n47), .B(n1791), .Z(n1790) );
  XNOR U1737 ( .A(p_input[191]), .B(n1789), .Z(n1791) );
  XOR U1738 ( .A(n1792), .B(n1793), .Z(n1789) );
  AND U1739 ( .A(n51), .B(n1794), .Z(n1793) );
  XNOR U1740 ( .A(p_input[207]), .B(n1792), .Z(n1794) );
  XOR U1741 ( .A(n1795), .B(n1796), .Z(n1792) );
  AND U1742 ( .A(n55), .B(n1797), .Z(n1796) );
  XNOR U1743 ( .A(p_input[223]), .B(n1795), .Z(n1797) );
  XOR U1744 ( .A(n1798), .B(n1799), .Z(n1795) );
  AND U1745 ( .A(n59), .B(n1800), .Z(n1799) );
  XNOR U1746 ( .A(p_input[239]), .B(n1798), .Z(n1800) );
  XOR U1747 ( .A(n1801), .B(n1802), .Z(n1798) );
  AND U1748 ( .A(n63), .B(n1803), .Z(n1802) );
  XNOR U1749 ( .A(p_input[255]), .B(n1801), .Z(n1803) );
  XOR U1750 ( .A(n1804), .B(n1805), .Z(n1801) );
  AND U1751 ( .A(n67), .B(n1806), .Z(n1805) );
  XNOR U1752 ( .A(p_input[271]), .B(n1804), .Z(n1806) );
  XOR U1753 ( .A(n1807), .B(n1808), .Z(n1804) );
  AND U1754 ( .A(n71), .B(n1809), .Z(n1808) );
  XNOR U1755 ( .A(p_input[287]), .B(n1807), .Z(n1809) );
  XOR U1756 ( .A(n1810), .B(n1811), .Z(n1807) );
  AND U1757 ( .A(n75), .B(n1812), .Z(n1811) );
  XNOR U1758 ( .A(p_input[303]), .B(n1810), .Z(n1812) );
  XOR U1759 ( .A(n1813), .B(n1814), .Z(n1810) );
  AND U1760 ( .A(n79), .B(n1815), .Z(n1814) );
  XNOR U1761 ( .A(p_input[319]), .B(n1813), .Z(n1815) );
  XOR U1762 ( .A(n1816), .B(n1817), .Z(n1813) );
  AND U1763 ( .A(n83), .B(n1818), .Z(n1817) );
  XNOR U1764 ( .A(p_input[335]), .B(n1816), .Z(n1818) );
  XOR U1765 ( .A(n1819), .B(n1820), .Z(n1816) );
  AND U1766 ( .A(n87), .B(n1821), .Z(n1820) );
  XNOR U1767 ( .A(p_input[351]), .B(n1819), .Z(n1821) );
  XOR U1768 ( .A(n1822), .B(n1823), .Z(n1819) );
  AND U1769 ( .A(n91), .B(n1824), .Z(n1823) );
  XNOR U1770 ( .A(p_input[367]), .B(n1822), .Z(n1824) );
  XOR U1771 ( .A(n1825), .B(n1826), .Z(n1822) );
  AND U1772 ( .A(n95), .B(n1827), .Z(n1826) );
  XNOR U1773 ( .A(p_input[383]), .B(n1825), .Z(n1827) );
  XOR U1774 ( .A(n1828), .B(n1829), .Z(n1825) );
  AND U1775 ( .A(n99), .B(n1830), .Z(n1829) );
  XNOR U1776 ( .A(p_input[399]), .B(n1828), .Z(n1830) );
  XOR U1777 ( .A(n1831), .B(n1832), .Z(n1828) );
  AND U1778 ( .A(n103), .B(n1833), .Z(n1832) );
  XNOR U1779 ( .A(p_input[415]), .B(n1831), .Z(n1833) );
  XOR U1780 ( .A(n1834), .B(n1835), .Z(n1831) );
  AND U1781 ( .A(n107), .B(n1836), .Z(n1835) );
  XNOR U1782 ( .A(p_input[431]), .B(n1834), .Z(n1836) );
  XOR U1783 ( .A(n1837), .B(n1838), .Z(n1834) );
  AND U1784 ( .A(n111), .B(n1839), .Z(n1838) );
  XNOR U1785 ( .A(p_input[447]), .B(n1837), .Z(n1839) );
  XOR U1786 ( .A(n1840), .B(n1841), .Z(n1837) );
  AND U1787 ( .A(n115), .B(n1842), .Z(n1841) );
  XNOR U1788 ( .A(p_input[463]), .B(n1840), .Z(n1842) );
  XOR U1789 ( .A(n1843), .B(n1844), .Z(n1840) );
  AND U1790 ( .A(n119), .B(n1845), .Z(n1844) );
  XNOR U1791 ( .A(p_input[479]), .B(n1843), .Z(n1845) );
  XOR U1792 ( .A(n1846), .B(n1847), .Z(n1843) );
  AND U1793 ( .A(n123), .B(n1848), .Z(n1847) );
  XNOR U1794 ( .A(p_input[495]), .B(n1846), .Z(n1848) );
  XOR U1795 ( .A(n1849), .B(n1850), .Z(n1846) );
  AND U1796 ( .A(n127), .B(n1851), .Z(n1850) );
  XNOR U1797 ( .A(p_input[511]), .B(n1849), .Z(n1851) );
  XOR U1798 ( .A(n1852), .B(n1853), .Z(n1849) );
  AND U1799 ( .A(n131), .B(n1854), .Z(n1853) );
  XNOR U1800 ( .A(p_input[527]), .B(n1852), .Z(n1854) );
  XOR U1801 ( .A(n1855), .B(n1856), .Z(n1852) );
  AND U1802 ( .A(n135), .B(n1857), .Z(n1856) );
  XNOR U1803 ( .A(p_input[543]), .B(n1855), .Z(n1857) );
  XOR U1804 ( .A(n1858), .B(n1859), .Z(n1855) );
  AND U1805 ( .A(n139), .B(n1860), .Z(n1859) );
  XNOR U1806 ( .A(p_input[559]), .B(n1858), .Z(n1860) );
  XOR U1807 ( .A(n1861), .B(n1862), .Z(n1858) );
  AND U1808 ( .A(n143), .B(n1863), .Z(n1862) );
  XNOR U1809 ( .A(p_input[575]), .B(n1861), .Z(n1863) );
  XOR U1810 ( .A(n1864), .B(n1865), .Z(n1861) );
  AND U1811 ( .A(n147), .B(n1866), .Z(n1865) );
  XNOR U1812 ( .A(p_input[591]), .B(n1864), .Z(n1866) );
  XOR U1813 ( .A(n1867), .B(n1868), .Z(n1864) );
  AND U1814 ( .A(n151), .B(n1869), .Z(n1868) );
  XNOR U1815 ( .A(p_input[607]), .B(n1867), .Z(n1869) );
  XOR U1816 ( .A(n1870), .B(n1871), .Z(n1867) );
  AND U1817 ( .A(n155), .B(n1872), .Z(n1871) );
  XNOR U1818 ( .A(p_input[623]), .B(n1870), .Z(n1872) );
  XOR U1819 ( .A(n1873), .B(n1874), .Z(n1870) );
  AND U1820 ( .A(n159), .B(n1875), .Z(n1874) );
  XNOR U1821 ( .A(p_input[639]), .B(n1873), .Z(n1875) );
  XOR U1822 ( .A(n1876), .B(n1877), .Z(n1873) );
  AND U1823 ( .A(n163), .B(n1878), .Z(n1877) );
  XNOR U1824 ( .A(p_input[655]), .B(n1876), .Z(n1878) );
  XOR U1825 ( .A(n1879), .B(n1880), .Z(n1876) );
  AND U1826 ( .A(n167), .B(n1881), .Z(n1880) );
  XNOR U1827 ( .A(p_input[671]), .B(n1879), .Z(n1881) );
  XOR U1828 ( .A(n1882), .B(n1883), .Z(n1879) );
  AND U1829 ( .A(n171), .B(n1884), .Z(n1883) );
  XNOR U1830 ( .A(p_input[687]), .B(n1882), .Z(n1884) );
  XOR U1831 ( .A(n1885), .B(n1886), .Z(n1882) );
  AND U1832 ( .A(n175), .B(n1887), .Z(n1886) );
  XNOR U1833 ( .A(p_input[703]), .B(n1885), .Z(n1887) );
  XOR U1834 ( .A(n1888), .B(n1889), .Z(n1885) );
  AND U1835 ( .A(n179), .B(n1890), .Z(n1889) );
  XNOR U1836 ( .A(p_input[719]), .B(n1888), .Z(n1890) );
  XOR U1837 ( .A(n1891), .B(n1892), .Z(n1888) );
  AND U1838 ( .A(n183), .B(n1893), .Z(n1892) );
  XNOR U1839 ( .A(p_input[735]), .B(n1891), .Z(n1893) );
  XOR U1840 ( .A(n1894), .B(n1895), .Z(n1891) );
  AND U1841 ( .A(n187), .B(n1896), .Z(n1895) );
  XNOR U1842 ( .A(p_input[751]), .B(n1894), .Z(n1896) );
  XOR U1843 ( .A(n1897), .B(n1898), .Z(n1894) );
  AND U1844 ( .A(n191), .B(n1899), .Z(n1898) );
  XNOR U1845 ( .A(p_input[767]), .B(n1897), .Z(n1899) );
  XOR U1846 ( .A(n1900), .B(n1901), .Z(n1897) );
  AND U1847 ( .A(n195), .B(n1902), .Z(n1901) );
  XNOR U1848 ( .A(p_input[783]), .B(n1900), .Z(n1902) );
  XOR U1849 ( .A(n1903), .B(n1904), .Z(n1900) );
  AND U1850 ( .A(n199), .B(n1905), .Z(n1904) );
  XNOR U1851 ( .A(p_input[799]), .B(n1903), .Z(n1905) );
  XOR U1852 ( .A(n1906), .B(n1907), .Z(n1903) );
  AND U1853 ( .A(n203), .B(n1908), .Z(n1907) );
  XNOR U1854 ( .A(p_input[815]), .B(n1906), .Z(n1908) );
  XOR U1855 ( .A(n1909), .B(n1910), .Z(n1906) );
  AND U1856 ( .A(n207), .B(n1911), .Z(n1910) );
  XNOR U1857 ( .A(p_input[831]), .B(n1909), .Z(n1911) );
  XOR U1858 ( .A(n1912), .B(n1913), .Z(n1909) );
  AND U1859 ( .A(n211), .B(n1914), .Z(n1913) );
  XNOR U1860 ( .A(p_input[847]), .B(n1912), .Z(n1914) );
  XOR U1861 ( .A(n1915), .B(n1916), .Z(n1912) );
  AND U1862 ( .A(n215), .B(n1917), .Z(n1916) );
  XNOR U1863 ( .A(p_input[863]), .B(n1915), .Z(n1917) );
  XOR U1864 ( .A(n1918), .B(n1919), .Z(n1915) );
  AND U1865 ( .A(n219), .B(n1920), .Z(n1919) );
  XNOR U1866 ( .A(p_input[879]), .B(n1918), .Z(n1920) );
  XOR U1867 ( .A(n1921), .B(n1922), .Z(n1918) );
  AND U1868 ( .A(n223), .B(n1923), .Z(n1922) );
  XNOR U1869 ( .A(p_input[895]), .B(n1921), .Z(n1923) );
  XOR U1870 ( .A(n1924), .B(n1925), .Z(n1921) );
  AND U1871 ( .A(n227), .B(n1926), .Z(n1925) );
  XNOR U1872 ( .A(p_input[911]), .B(n1924), .Z(n1926) );
  XOR U1873 ( .A(n1927), .B(n1928), .Z(n1924) );
  AND U1874 ( .A(n231), .B(n1929), .Z(n1928) );
  XNOR U1875 ( .A(p_input[927]), .B(n1927), .Z(n1929) );
  XOR U1876 ( .A(n1930), .B(n1931), .Z(n1927) );
  AND U1877 ( .A(n235), .B(n1932), .Z(n1931) );
  XNOR U1878 ( .A(p_input[943]), .B(n1930), .Z(n1932) );
  XOR U1879 ( .A(n1933), .B(n1934), .Z(n1930) );
  AND U1880 ( .A(n239), .B(n1935), .Z(n1934) );
  XNOR U1881 ( .A(p_input[959]), .B(n1933), .Z(n1935) );
  XOR U1882 ( .A(n1936), .B(n1937), .Z(n1933) );
  AND U1883 ( .A(n243), .B(n1938), .Z(n1937) );
  XNOR U1884 ( .A(p_input[975]), .B(n1936), .Z(n1938) );
  XNOR U1885 ( .A(n1939), .B(n1940), .Z(n1936) );
  AND U1886 ( .A(n247), .B(n1941), .Z(n1940) );
  XOR U1887 ( .A(p_input[991]), .B(n1939), .Z(n1941) );
  XOR U1888 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n1942), .Z(n1939) );
  AND U1889 ( .A(n250), .B(n1943), .Z(n1942) );
  XOR U1890 ( .A(p_input[1007]), .B(\knn_comb_/min_val_out[0][15] ), .Z(n1943)
         );
  XNOR U1891 ( .A(n1944), .B(n1945), .Z(o[14]) );
  AND U1892 ( .A(n3), .B(n1946), .Z(n1944) );
  XNOR U1893 ( .A(p_input[14]), .B(n1945), .Z(n1946) );
  XOR U1894 ( .A(n1947), .B(n1948), .Z(n1945) );
  AND U1895 ( .A(n7), .B(n1949), .Z(n1948) );
  XNOR U1896 ( .A(p_input[30]), .B(n1947), .Z(n1949) );
  XOR U1897 ( .A(n1950), .B(n1951), .Z(n1947) );
  AND U1898 ( .A(n11), .B(n1952), .Z(n1951) );
  XNOR U1899 ( .A(p_input[46]), .B(n1950), .Z(n1952) );
  XOR U1900 ( .A(n1953), .B(n1954), .Z(n1950) );
  AND U1901 ( .A(n15), .B(n1955), .Z(n1954) );
  XNOR U1902 ( .A(p_input[62]), .B(n1953), .Z(n1955) );
  XOR U1903 ( .A(n1956), .B(n1957), .Z(n1953) );
  AND U1904 ( .A(n19), .B(n1958), .Z(n1957) );
  XNOR U1905 ( .A(p_input[78]), .B(n1956), .Z(n1958) );
  XOR U1906 ( .A(n1959), .B(n1960), .Z(n1956) );
  AND U1907 ( .A(n23), .B(n1961), .Z(n1960) );
  XNOR U1908 ( .A(p_input[94]), .B(n1959), .Z(n1961) );
  XOR U1909 ( .A(n1962), .B(n1963), .Z(n1959) );
  AND U1910 ( .A(n27), .B(n1964), .Z(n1963) );
  XNOR U1911 ( .A(p_input[110]), .B(n1962), .Z(n1964) );
  XOR U1912 ( .A(n1965), .B(n1966), .Z(n1962) );
  AND U1913 ( .A(n31), .B(n1967), .Z(n1966) );
  XNOR U1914 ( .A(p_input[126]), .B(n1965), .Z(n1967) );
  XOR U1915 ( .A(n1968), .B(n1969), .Z(n1965) );
  AND U1916 ( .A(n35), .B(n1970), .Z(n1969) );
  XNOR U1917 ( .A(p_input[142]), .B(n1968), .Z(n1970) );
  XOR U1918 ( .A(n1971), .B(n1972), .Z(n1968) );
  AND U1919 ( .A(n39), .B(n1973), .Z(n1972) );
  XNOR U1920 ( .A(p_input[158]), .B(n1971), .Z(n1973) );
  XOR U1921 ( .A(n1974), .B(n1975), .Z(n1971) );
  AND U1922 ( .A(n43), .B(n1976), .Z(n1975) );
  XNOR U1923 ( .A(p_input[174]), .B(n1974), .Z(n1976) );
  XOR U1924 ( .A(n1977), .B(n1978), .Z(n1974) );
  AND U1925 ( .A(n47), .B(n1979), .Z(n1978) );
  XNOR U1926 ( .A(p_input[190]), .B(n1977), .Z(n1979) );
  XOR U1927 ( .A(n1980), .B(n1981), .Z(n1977) );
  AND U1928 ( .A(n51), .B(n1982), .Z(n1981) );
  XNOR U1929 ( .A(p_input[206]), .B(n1980), .Z(n1982) );
  XOR U1930 ( .A(n1983), .B(n1984), .Z(n1980) );
  AND U1931 ( .A(n55), .B(n1985), .Z(n1984) );
  XNOR U1932 ( .A(p_input[222]), .B(n1983), .Z(n1985) );
  XOR U1933 ( .A(n1986), .B(n1987), .Z(n1983) );
  AND U1934 ( .A(n59), .B(n1988), .Z(n1987) );
  XNOR U1935 ( .A(p_input[238]), .B(n1986), .Z(n1988) );
  XOR U1936 ( .A(n1989), .B(n1990), .Z(n1986) );
  AND U1937 ( .A(n63), .B(n1991), .Z(n1990) );
  XNOR U1938 ( .A(p_input[254]), .B(n1989), .Z(n1991) );
  XOR U1939 ( .A(n1992), .B(n1993), .Z(n1989) );
  AND U1940 ( .A(n67), .B(n1994), .Z(n1993) );
  XNOR U1941 ( .A(p_input[270]), .B(n1992), .Z(n1994) );
  XOR U1942 ( .A(n1995), .B(n1996), .Z(n1992) );
  AND U1943 ( .A(n71), .B(n1997), .Z(n1996) );
  XNOR U1944 ( .A(p_input[286]), .B(n1995), .Z(n1997) );
  XOR U1945 ( .A(n1998), .B(n1999), .Z(n1995) );
  AND U1946 ( .A(n75), .B(n2000), .Z(n1999) );
  XNOR U1947 ( .A(p_input[302]), .B(n1998), .Z(n2000) );
  XOR U1948 ( .A(n2001), .B(n2002), .Z(n1998) );
  AND U1949 ( .A(n79), .B(n2003), .Z(n2002) );
  XNOR U1950 ( .A(p_input[318]), .B(n2001), .Z(n2003) );
  XOR U1951 ( .A(n2004), .B(n2005), .Z(n2001) );
  AND U1952 ( .A(n83), .B(n2006), .Z(n2005) );
  XNOR U1953 ( .A(p_input[334]), .B(n2004), .Z(n2006) );
  XOR U1954 ( .A(n2007), .B(n2008), .Z(n2004) );
  AND U1955 ( .A(n87), .B(n2009), .Z(n2008) );
  XNOR U1956 ( .A(p_input[350]), .B(n2007), .Z(n2009) );
  XOR U1957 ( .A(n2010), .B(n2011), .Z(n2007) );
  AND U1958 ( .A(n91), .B(n2012), .Z(n2011) );
  XNOR U1959 ( .A(p_input[366]), .B(n2010), .Z(n2012) );
  XOR U1960 ( .A(n2013), .B(n2014), .Z(n2010) );
  AND U1961 ( .A(n95), .B(n2015), .Z(n2014) );
  XNOR U1962 ( .A(p_input[382]), .B(n2013), .Z(n2015) );
  XOR U1963 ( .A(n2016), .B(n2017), .Z(n2013) );
  AND U1964 ( .A(n99), .B(n2018), .Z(n2017) );
  XNOR U1965 ( .A(p_input[398]), .B(n2016), .Z(n2018) );
  XOR U1966 ( .A(n2019), .B(n2020), .Z(n2016) );
  AND U1967 ( .A(n103), .B(n2021), .Z(n2020) );
  XNOR U1968 ( .A(p_input[414]), .B(n2019), .Z(n2021) );
  XOR U1969 ( .A(n2022), .B(n2023), .Z(n2019) );
  AND U1970 ( .A(n107), .B(n2024), .Z(n2023) );
  XNOR U1971 ( .A(p_input[430]), .B(n2022), .Z(n2024) );
  XOR U1972 ( .A(n2025), .B(n2026), .Z(n2022) );
  AND U1973 ( .A(n111), .B(n2027), .Z(n2026) );
  XNOR U1974 ( .A(p_input[446]), .B(n2025), .Z(n2027) );
  XOR U1975 ( .A(n2028), .B(n2029), .Z(n2025) );
  AND U1976 ( .A(n115), .B(n2030), .Z(n2029) );
  XNOR U1977 ( .A(p_input[462]), .B(n2028), .Z(n2030) );
  XOR U1978 ( .A(n2031), .B(n2032), .Z(n2028) );
  AND U1979 ( .A(n119), .B(n2033), .Z(n2032) );
  XNOR U1980 ( .A(p_input[478]), .B(n2031), .Z(n2033) );
  XOR U1981 ( .A(n2034), .B(n2035), .Z(n2031) );
  AND U1982 ( .A(n123), .B(n2036), .Z(n2035) );
  XNOR U1983 ( .A(p_input[494]), .B(n2034), .Z(n2036) );
  XOR U1984 ( .A(n2037), .B(n2038), .Z(n2034) );
  AND U1985 ( .A(n127), .B(n2039), .Z(n2038) );
  XNOR U1986 ( .A(p_input[510]), .B(n2037), .Z(n2039) );
  XOR U1987 ( .A(n2040), .B(n2041), .Z(n2037) );
  AND U1988 ( .A(n131), .B(n2042), .Z(n2041) );
  XNOR U1989 ( .A(p_input[526]), .B(n2040), .Z(n2042) );
  XOR U1990 ( .A(n2043), .B(n2044), .Z(n2040) );
  AND U1991 ( .A(n135), .B(n2045), .Z(n2044) );
  XNOR U1992 ( .A(p_input[542]), .B(n2043), .Z(n2045) );
  XOR U1993 ( .A(n2046), .B(n2047), .Z(n2043) );
  AND U1994 ( .A(n139), .B(n2048), .Z(n2047) );
  XNOR U1995 ( .A(p_input[558]), .B(n2046), .Z(n2048) );
  XOR U1996 ( .A(n2049), .B(n2050), .Z(n2046) );
  AND U1997 ( .A(n143), .B(n2051), .Z(n2050) );
  XNOR U1998 ( .A(p_input[574]), .B(n2049), .Z(n2051) );
  XOR U1999 ( .A(n2052), .B(n2053), .Z(n2049) );
  AND U2000 ( .A(n147), .B(n2054), .Z(n2053) );
  XNOR U2001 ( .A(p_input[590]), .B(n2052), .Z(n2054) );
  XOR U2002 ( .A(n2055), .B(n2056), .Z(n2052) );
  AND U2003 ( .A(n151), .B(n2057), .Z(n2056) );
  XNOR U2004 ( .A(p_input[606]), .B(n2055), .Z(n2057) );
  XOR U2005 ( .A(n2058), .B(n2059), .Z(n2055) );
  AND U2006 ( .A(n155), .B(n2060), .Z(n2059) );
  XNOR U2007 ( .A(p_input[622]), .B(n2058), .Z(n2060) );
  XOR U2008 ( .A(n2061), .B(n2062), .Z(n2058) );
  AND U2009 ( .A(n159), .B(n2063), .Z(n2062) );
  XNOR U2010 ( .A(p_input[638]), .B(n2061), .Z(n2063) );
  XOR U2011 ( .A(n2064), .B(n2065), .Z(n2061) );
  AND U2012 ( .A(n163), .B(n2066), .Z(n2065) );
  XNOR U2013 ( .A(p_input[654]), .B(n2064), .Z(n2066) );
  XOR U2014 ( .A(n2067), .B(n2068), .Z(n2064) );
  AND U2015 ( .A(n167), .B(n2069), .Z(n2068) );
  XNOR U2016 ( .A(p_input[670]), .B(n2067), .Z(n2069) );
  XOR U2017 ( .A(n2070), .B(n2071), .Z(n2067) );
  AND U2018 ( .A(n171), .B(n2072), .Z(n2071) );
  XNOR U2019 ( .A(p_input[686]), .B(n2070), .Z(n2072) );
  XOR U2020 ( .A(n2073), .B(n2074), .Z(n2070) );
  AND U2021 ( .A(n175), .B(n2075), .Z(n2074) );
  XNOR U2022 ( .A(p_input[702]), .B(n2073), .Z(n2075) );
  XOR U2023 ( .A(n2076), .B(n2077), .Z(n2073) );
  AND U2024 ( .A(n179), .B(n2078), .Z(n2077) );
  XNOR U2025 ( .A(p_input[718]), .B(n2076), .Z(n2078) );
  XOR U2026 ( .A(n2079), .B(n2080), .Z(n2076) );
  AND U2027 ( .A(n183), .B(n2081), .Z(n2080) );
  XNOR U2028 ( .A(p_input[734]), .B(n2079), .Z(n2081) );
  XOR U2029 ( .A(n2082), .B(n2083), .Z(n2079) );
  AND U2030 ( .A(n187), .B(n2084), .Z(n2083) );
  XNOR U2031 ( .A(p_input[750]), .B(n2082), .Z(n2084) );
  XOR U2032 ( .A(n2085), .B(n2086), .Z(n2082) );
  AND U2033 ( .A(n191), .B(n2087), .Z(n2086) );
  XNOR U2034 ( .A(p_input[766]), .B(n2085), .Z(n2087) );
  XOR U2035 ( .A(n2088), .B(n2089), .Z(n2085) );
  AND U2036 ( .A(n195), .B(n2090), .Z(n2089) );
  XNOR U2037 ( .A(p_input[782]), .B(n2088), .Z(n2090) );
  XOR U2038 ( .A(n2091), .B(n2092), .Z(n2088) );
  AND U2039 ( .A(n199), .B(n2093), .Z(n2092) );
  XNOR U2040 ( .A(p_input[798]), .B(n2091), .Z(n2093) );
  XOR U2041 ( .A(n2094), .B(n2095), .Z(n2091) );
  AND U2042 ( .A(n203), .B(n2096), .Z(n2095) );
  XNOR U2043 ( .A(p_input[814]), .B(n2094), .Z(n2096) );
  XOR U2044 ( .A(n2097), .B(n2098), .Z(n2094) );
  AND U2045 ( .A(n207), .B(n2099), .Z(n2098) );
  XNOR U2046 ( .A(p_input[830]), .B(n2097), .Z(n2099) );
  XOR U2047 ( .A(n2100), .B(n2101), .Z(n2097) );
  AND U2048 ( .A(n211), .B(n2102), .Z(n2101) );
  XNOR U2049 ( .A(p_input[846]), .B(n2100), .Z(n2102) );
  XOR U2050 ( .A(n2103), .B(n2104), .Z(n2100) );
  AND U2051 ( .A(n215), .B(n2105), .Z(n2104) );
  XNOR U2052 ( .A(p_input[862]), .B(n2103), .Z(n2105) );
  XOR U2053 ( .A(n2106), .B(n2107), .Z(n2103) );
  AND U2054 ( .A(n219), .B(n2108), .Z(n2107) );
  XNOR U2055 ( .A(p_input[878]), .B(n2106), .Z(n2108) );
  XOR U2056 ( .A(n2109), .B(n2110), .Z(n2106) );
  AND U2057 ( .A(n223), .B(n2111), .Z(n2110) );
  XNOR U2058 ( .A(p_input[894]), .B(n2109), .Z(n2111) );
  XOR U2059 ( .A(n2112), .B(n2113), .Z(n2109) );
  AND U2060 ( .A(n227), .B(n2114), .Z(n2113) );
  XNOR U2061 ( .A(p_input[910]), .B(n2112), .Z(n2114) );
  XOR U2062 ( .A(n2115), .B(n2116), .Z(n2112) );
  AND U2063 ( .A(n231), .B(n2117), .Z(n2116) );
  XNOR U2064 ( .A(p_input[926]), .B(n2115), .Z(n2117) );
  XOR U2065 ( .A(n2118), .B(n2119), .Z(n2115) );
  AND U2066 ( .A(n235), .B(n2120), .Z(n2119) );
  XNOR U2067 ( .A(p_input[942]), .B(n2118), .Z(n2120) );
  XOR U2068 ( .A(n2121), .B(n2122), .Z(n2118) );
  AND U2069 ( .A(n239), .B(n2123), .Z(n2122) );
  XNOR U2070 ( .A(p_input[958]), .B(n2121), .Z(n2123) );
  XOR U2071 ( .A(n2124), .B(n2125), .Z(n2121) );
  AND U2072 ( .A(n243), .B(n2126), .Z(n2125) );
  XNOR U2073 ( .A(p_input[974]), .B(n2124), .Z(n2126) );
  XNOR U2074 ( .A(n2127), .B(n2128), .Z(n2124) );
  AND U2075 ( .A(n247), .B(n2129), .Z(n2128) );
  XOR U2076 ( .A(p_input[990]), .B(n2127), .Z(n2129) );
  XOR U2077 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n2130), .Z(n2127) );
  AND U2078 ( .A(n250), .B(n2131), .Z(n2130) );
  XOR U2079 ( .A(p_input[1006]), .B(\knn_comb_/min_val_out[0][14] ), .Z(n2131)
         );
  XNOR U2080 ( .A(n2132), .B(n2133), .Z(o[13]) );
  AND U2081 ( .A(n3), .B(n2134), .Z(n2132) );
  XNOR U2082 ( .A(p_input[13]), .B(n2133), .Z(n2134) );
  XOR U2083 ( .A(n2135), .B(n2136), .Z(n2133) );
  AND U2084 ( .A(n7), .B(n2137), .Z(n2136) );
  XNOR U2085 ( .A(p_input[29]), .B(n2135), .Z(n2137) );
  XOR U2086 ( .A(n2138), .B(n2139), .Z(n2135) );
  AND U2087 ( .A(n11), .B(n2140), .Z(n2139) );
  XNOR U2088 ( .A(p_input[45]), .B(n2138), .Z(n2140) );
  XOR U2089 ( .A(n2141), .B(n2142), .Z(n2138) );
  AND U2090 ( .A(n15), .B(n2143), .Z(n2142) );
  XNOR U2091 ( .A(p_input[61]), .B(n2141), .Z(n2143) );
  XOR U2092 ( .A(n2144), .B(n2145), .Z(n2141) );
  AND U2093 ( .A(n19), .B(n2146), .Z(n2145) );
  XNOR U2094 ( .A(p_input[77]), .B(n2144), .Z(n2146) );
  XOR U2095 ( .A(n2147), .B(n2148), .Z(n2144) );
  AND U2096 ( .A(n23), .B(n2149), .Z(n2148) );
  XNOR U2097 ( .A(p_input[93]), .B(n2147), .Z(n2149) );
  XOR U2098 ( .A(n2150), .B(n2151), .Z(n2147) );
  AND U2099 ( .A(n27), .B(n2152), .Z(n2151) );
  XNOR U2100 ( .A(p_input[109]), .B(n2150), .Z(n2152) );
  XOR U2101 ( .A(n2153), .B(n2154), .Z(n2150) );
  AND U2102 ( .A(n31), .B(n2155), .Z(n2154) );
  XNOR U2103 ( .A(p_input[125]), .B(n2153), .Z(n2155) );
  XOR U2104 ( .A(n2156), .B(n2157), .Z(n2153) );
  AND U2105 ( .A(n35), .B(n2158), .Z(n2157) );
  XNOR U2106 ( .A(p_input[141]), .B(n2156), .Z(n2158) );
  XOR U2107 ( .A(n2159), .B(n2160), .Z(n2156) );
  AND U2108 ( .A(n39), .B(n2161), .Z(n2160) );
  XNOR U2109 ( .A(p_input[157]), .B(n2159), .Z(n2161) );
  XOR U2110 ( .A(n2162), .B(n2163), .Z(n2159) );
  AND U2111 ( .A(n43), .B(n2164), .Z(n2163) );
  XNOR U2112 ( .A(p_input[173]), .B(n2162), .Z(n2164) );
  XOR U2113 ( .A(n2165), .B(n2166), .Z(n2162) );
  AND U2114 ( .A(n47), .B(n2167), .Z(n2166) );
  XNOR U2115 ( .A(p_input[189]), .B(n2165), .Z(n2167) );
  XOR U2116 ( .A(n2168), .B(n2169), .Z(n2165) );
  AND U2117 ( .A(n51), .B(n2170), .Z(n2169) );
  XNOR U2118 ( .A(p_input[205]), .B(n2168), .Z(n2170) );
  XOR U2119 ( .A(n2171), .B(n2172), .Z(n2168) );
  AND U2120 ( .A(n55), .B(n2173), .Z(n2172) );
  XNOR U2121 ( .A(p_input[221]), .B(n2171), .Z(n2173) );
  XOR U2122 ( .A(n2174), .B(n2175), .Z(n2171) );
  AND U2123 ( .A(n59), .B(n2176), .Z(n2175) );
  XNOR U2124 ( .A(p_input[237]), .B(n2174), .Z(n2176) );
  XOR U2125 ( .A(n2177), .B(n2178), .Z(n2174) );
  AND U2126 ( .A(n63), .B(n2179), .Z(n2178) );
  XNOR U2127 ( .A(p_input[253]), .B(n2177), .Z(n2179) );
  XOR U2128 ( .A(n2180), .B(n2181), .Z(n2177) );
  AND U2129 ( .A(n67), .B(n2182), .Z(n2181) );
  XNOR U2130 ( .A(p_input[269]), .B(n2180), .Z(n2182) );
  XOR U2131 ( .A(n2183), .B(n2184), .Z(n2180) );
  AND U2132 ( .A(n71), .B(n2185), .Z(n2184) );
  XNOR U2133 ( .A(p_input[285]), .B(n2183), .Z(n2185) );
  XOR U2134 ( .A(n2186), .B(n2187), .Z(n2183) );
  AND U2135 ( .A(n75), .B(n2188), .Z(n2187) );
  XNOR U2136 ( .A(p_input[301]), .B(n2186), .Z(n2188) );
  XOR U2137 ( .A(n2189), .B(n2190), .Z(n2186) );
  AND U2138 ( .A(n79), .B(n2191), .Z(n2190) );
  XNOR U2139 ( .A(p_input[317]), .B(n2189), .Z(n2191) );
  XOR U2140 ( .A(n2192), .B(n2193), .Z(n2189) );
  AND U2141 ( .A(n83), .B(n2194), .Z(n2193) );
  XNOR U2142 ( .A(p_input[333]), .B(n2192), .Z(n2194) );
  XOR U2143 ( .A(n2195), .B(n2196), .Z(n2192) );
  AND U2144 ( .A(n87), .B(n2197), .Z(n2196) );
  XNOR U2145 ( .A(p_input[349]), .B(n2195), .Z(n2197) );
  XOR U2146 ( .A(n2198), .B(n2199), .Z(n2195) );
  AND U2147 ( .A(n91), .B(n2200), .Z(n2199) );
  XNOR U2148 ( .A(p_input[365]), .B(n2198), .Z(n2200) );
  XOR U2149 ( .A(n2201), .B(n2202), .Z(n2198) );
  AND U2150 ( .A(n95), .B(n2203), .Z(n2202) );
  XNOR U2151 ( .A(p_input[381]), .B(n2201), .Z(n2203) );
  XOR U2152 ( .A(n2204), .B(n2205), .Z(n2201) );
  AND U2153 ( .A(n99), .B(n2206), .Z(n2205) );
  XNOR U2154 ( .A(p_input[397]), .B(n2204), .Z(n2206) );
  XOR U2155 ( .A(n2207), .B(n2208), .Z(n2204) );
  AND U2156 ( .A(n103), .B(n2209), .Z(n2208) );
  XNOR U2157 ( .A(p_input[413]), .B(n2207), .Z(n2209) );
  XOR U2158 ( .A(n2210), .B(n2211), .Z(n2207) );
  AND U2159 ( .A(n107), .B(n2212), .Z(n2211) );
  XNOR U2160 ( .A(p_input[429]), .B(n2210), .Z(n2212) );
  XOR U2161 ( .A(n2213), .B(n2214), .Z(n2210) );
  AND U2162 ( .A(n111), .B(n2215), .Z(n2214) );
  XNOR U2163 ( .A(p_input[445]), .B(n2213), .Z(n2215) );
  XOR U2164 ( .A(n2216), .B(n2217), .Z(n2213) );
  AND U2165 ( .A(n115), .B(n2218), .Z(n2217) );
  XNOR U2166 ( .A(p_input[461]), .B(n2216), .Z(n2218) );
  XOR U2167 ( .A(n2219), .B(n2220), .Z(n2216) );
  AND U2168 ( .A(n119), .B(n2221), .Z(n2220) );
  XNOR U2169 ( .A(p_input[477]), .B(n2219), .Z(n2221) );
  XOR U2170 ( .A(n2222), .B(n2223), .Z(n2219) );
  AND U2171 ( .A(n123), .B(n2224), .Z(n2223) );
  XNOR U2172 ( .A(p_input[493]), .B(n2222), .Z(n2224) );
  XOR U2173 ( .A(n2225), .B(n2226), .Z(n2222) );
  AND U2174 ( .A(n127), .B(n2227), .Z(n2226) );
  XNOR U2175 ( .A(p_input[509]), .B(n2225), .Z(n2227) );
  XOR U2176 ( .A(n2228), .B(n2229), .Z(n2225) );
  AND U2177 ( .A(n131), .B(n2230), .Z(n2229) );
  XNOR U2178 ( .A(p_input[525]), .B(n2228), .Z(n2230) );
  XOR U2179 ( .A(n2231), .B(n2232), .Z(n2228) );
  AND U2180 ( .A(n135), .B(n2233), .Z(n2232) );
  XNOR U2181 ( .A(p_input[541]), .B(n2231), .Z(n2233) );
  XOR U2182 ( .A(n2234), .B(n2235), .Z(n2231) );
  AND U2183 ( .A(n139), .B(n2236), .Z(n2235) );
  XNOR U2184 ( .A(p_input[557]), .B(n2234), .Z(n2236) );
  XOR U2185 ( .A(n2237), .B(n2238), .Z(n2234) );
  AND U2186 ( .A(n143), .B(n2239), .Z(n2238) );
  XNOR U2187 ( .A(p_input[573]), .B(n2237), .Z(n2239) );
  XOR U2188 ( .A(n2240), .B(n2241), .Z(n2237) );
  AND U2189 ( .A(n147), .B(n2242), .Z(n2241) );
  XNOR U2190 ( .A(p_input[589]), .B(n2240), .Z(n2242) );
  XOR U2191 ( .A(n2243), .B(n2244), .Z(n2240) );
  AND U2192 ( .A(n151), .B(n2245), .Z(n2244) );
  XNOR U2193 ( .A(p_input[605]), .B(n2243), .Z(n2245) );
  XOR U2194 ( .A(n2246), .B(n2247), .Z(n2243) );
  AND U2195 ( .A(n155), .B(n2248), .Z(n2247) );
  XNOR U2196 ( .A(p_input[621]), .B(n2246), .Z(n2248) );
  XOR U2197 ( .A(n2249), .B(n2250), .Z(n2246) );
  AND U2198 ( .A(n159), .B(n2251), .Z(n2250) );
  XNOR U2199 ( .A(p_input[637]), .B(n2249), .Z(n2251) );
  XOR U2200 ( .A(n2252), .B(n2253), .Z(n2249) );
  AND U2201 ( .A(n163), .B(n2254), .Z(n2253) );
  XNOR U2202 ( .A(p_input[653]), .B(n2252), .Z(n2254) );
  XOR U2203 ( .A(n2255), .B(n2256), .Z(n2252) );
  AND U2204 ( .A(n167), .B(n2257), .Z(n2256) );
  XNOR U2205 ( .A(p_input[669]), .B(n2255), .Z(n2257) );
  XOR U2206 ( .A(n2258), .B(n2259), .Z(n2255) );
  AND U2207 ( .A(n171), .B(n2260), .Z(n2259) );
  XNOR U2208 ( .A(p_input[685]), .B(n2258), .Z(n2260) );
  XOR U2209 ( .A(n2261), .B(n2262), .Z(n2258) );
  AND U2210 ( .A(n175), .B(n2263), .Z(n2262) );
  XNOR U2211 ( .A(p_input[701]), .B(n2261), .Z(n2263) );
  XOR U2212 ( .A(n2264), .B(n2265), .Z(n2261) );
  AND U2213 ( .A(n179), .B(n2266), .Z(n2265) );
  XNOR U2214 ( .A(p_input[717]), .B(n2264), .Z(n2266) );
  XOR U2215 ( .A(n2267), .B(n2268), .Z(n2264) );
  AND U2216 ( .A(n183), .B(n2269), .Z(n2268) );
  XNOR U2217 ( .A(p_input[733]), .B(n2267), .Z(n2269) );
  XOR U2218 ( .A(n2270), .B(n2271), .Z(n2267) );
  AND U2219 ( .A(n187), .B(n2272), .Z(n2271) );
  XNOR U2220 ( .A(p_input[749]), .B(n2270), .Z(n2272) );
  XOR U2221 ( .A(n2273), .B(n2274), .Z(n2270) );
  AND U2222 ( .A(n191), .B(n2275), .Z(n2274) );
  XNOR U2223 ( .A(p_input[765]), .B(n2273), .Z(n2275) );
  XOR U2224 ( .A(n2276), .B(n2277), .Z(n2273) );
  AND U2225 ( .A(n195), .B(n2278), .Z(n2277) );
  XNOR U2226 ( .A(p_input[781]), .B(n2276), .Z(n2278) );
  XOR U2227 ( .A(n2279), .B(n2280), .Z(n2276) );
  AND U2228 ( .A(n199), .B(n2281), .Z(n2280) );
  XNOR U2229 ( .A(p_input[797]), .B(n2279), .Z(n2281) );
  XOR U2230 ( .A(n2282), .B(n2283), .Z(n2279) );
  AND U2231 ( .A(n203), .B(n2284), .Z(n2283) );
  XNOR U2232 ( .A(p_input[813]), .B(n2282), .Z(n2284) );
  XOR U2233 ( .A(n2285), .B(n2286), .Z(n2282) );
  AND U2234 ( .A(n207), .B(n2287), .Z(n2286) );
  XNOR U2235 ( .A(p_input[829]), .B(n2285), .Z(n2287) );
  XOR U2236 ( .A(n2288), .B(n2289), .Z(n2285) );
  AND U2237 ( .A(n211), .B(n2290), .Z(n2289) );
  XNOR U2238 ( .A(p_input[845]), .B(n2288), .Z(n2290) );
  XOR U2239 ( .A(n2291), .B(n2292), .Z(n2288) );
  AND U2240 ( .A(n215), .B(n2293), .Z(n2292) );
  XNOR U2241 ( .A(p_input[861]), .B(n2291), .Z(n2293) );
  XOR U2242 ( .A(n2294), .B(n2295), .Z(n2291) );
  AND U2243 ( .A(n219), .B(n2296), .Z(n2295) );
  XNOR U2244 ( .A(p_input[877]), .B(n2294), .Z(n2296) );
  XOR U2245 ( .A(n2297), .B(n2298), .Z(n2294) );
  AND U2246 ( .A(n223), .B(n2299), .Z(n2298) );
  XNOR U2247 ( .A(p_input[893]), .B(n2297), .Z(n2299) );
  XOR U2248 ( .A(n2300), .B(n2301), .Z(n2297) );
  AND U2249 ( .A(n227), .B(n2302), .Z(n2301) );
  XNOR U2250 ( .A(p_input[909]), .B(n2300), .Z(n2302) );
  XOR U2251 ( .A(n2303), .B(n2304), .Z(n2300) );
  AND U2252 ( .A(n231), .B(n2305), .Z(n2304) );
  XNOR U2253 ( .A(p_input[925]), .B(n2303), .Z(n2305) );
  XOR U2254 ( .A(n2306), .B(n2307), .Z(n2303) );
  AND U2255 ( .A(n235), .B(n2308), .Z(n2307) );
  XNOR U2256 ( .A(p_input[941]), .B(n2306), .Z(n2308) );
  XOR U2257 ( .A(n2309), .B(n2310), .Z(n2306) );
  AND U2258 ( .A(n239), .B(n2311), .Z(n2310) );
  XNOR U2259 ( .A(p_input[957]), .B(n2309), .Z(n2311) );
  XOR U2260 ( .A(n2312), .B(n2313), .Z(n2309) );
  AND U2261 ( .A(n243), .B(n2314), .Z(n2313) );
  XNOR U2262 ( .A(p_input[973]), .B(n2312), .Z(n2314) );
  XNOR U2263 ( .A(n2315), .B(n2316), .Z(n2312) );
  AND U2264 ( .A(n247), .B(n2317), .Z(n2316) );
  XOR U2265 ( .A(p_input[989]), .B(n2315), .Z(n2317) );
  XOR U2266 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n2318), .Z(n2315) );
  AND U2267 ( .A(n250), .B(n2319), .Z(n2318) );
  XOR U2268 ( .A(p_input[1005]), .B(\knn_comb_/min_val_out[0][13] ), .Z(n2319)
         );
  XNOR U2269 ( .A(n2320), .B(n2321), .Z(o[12]) );
  AND U2270 ( .A(n3), .B(n2322), .Z(n2320) );
  XNOR U2271 ( .A(p_input[12]), .B(n2321), .Z(n2322) );
  XOR U2272 ( .A(n2323), .B(n2324), .Z(n2321) );
  AND U2273 ( .A(n7), .B(n2325), .Z(n2324) );
  XNOR U2274 ( .A(p_input[28]), .B(n2323), .Z(n2325) );
  XOR U2275 ( .A(n2326), .B(n2327), .Z(n2323) );
  AND U2276 ( .A(n11), .B(n2328), .Z(n2327) );
  XNOR U2277 ( .A(p_input[44]), .B(n2326), .Z(n2328) );
  XOR U2278 ( .A(n2329), .B(n2330), .Z(n2326) );
  AND U2279 ( .A(n15), .B(n2331), .Z(n2330) );
  XNOR U2280 ( .A(p_input[60]), .B(n2329), .Z(n2331) );
  XOR U2281 ( .A(n2332), .B(n2333), .Z(n2329) );
  AND U2282 ( .A(n19), .B(n2334), .Z(n2333) );
  XNOR U2283 ( .A(p_input[76]), .B(n2332), .Z(n2334) );
  XOR U2284 ( .A(n2335), .B(n2336), .Z(n2332) );
  AND U2285 ( .A(n23), .B(n2337), .Z(n2336) );
  XNOR U2286 ( .A(p_input[92]), .B(n2335), .Z(n2337) );
  XOR U2287 ( .A(n2338), .B(n2339), .Z(n2335) );
  AND U2288 ( .A(n27), .B(n2340), .Z(n2339) );
  XNOR U2289 ( .A(p_input[108]), .B(n2338), .Z(n2340) );
  XOR U2290 ( .A(n2341), .B(n2342), .Z(n2338) );
  AND U2291 ( .A(n31), .B(n2343), .Z(n2342) );
  XNOR U2292 ( .A(p_input[124]), .B(n2341), .Z(n2343) );
  XOR U2293 ( .A(n2344), .B(n2345), .Z(n2341) );
  AND U2294 ( .A(n35), .B(n2346), .Z(n2345) );
  XNOR U2295 ( .A(p_input[140]), .B(n2344), .Z(n2346) );
  XOR U2296 ( .A(n2347), .B(n2348), .Z(n2344) );
  AND U2297 ( .A(n39), .B(n2349), .Z(n2348) );
  XNOR U2298 ( .A(p_input[156]), .B(n2347), .Z(n2349) );
  XOR U2299 ( .A(n2350), .B(n2351), .Z(n2347) );
  AND U2300 ( .A(n43), .B(n2352), .Z(n2351) );
  XNOR U2301 ( .A(p_input[172]), .B(n2350), .Z(n2352) );
  XOR U2302 ( .A(n2353), .B(n2354), .Z(n2350) );
  AND U2303 ( .A(n47), .B(n2355), .Z(n2354) );
  XNOR U2304 ( .A(p_input[188]), .B(n2353), .Z(n2355) );
  XOR U2305 ( .A(n2356), .B(n2357), .Z(n2353) );
  AND U2306 ( .A(n51), .B(n2358), .Z(n2357) );
  XNOR U2307 ( .A(p_input[204]), .B(n2356), .Z(n2358) );
  XOR U2308 ( .A(n2359), .B(n2360), .Z(n2356) );
  AND U2309 ( .A(n55), .B(n2361), .Z(n2360) );
  XNOR U2310 ( .A(p_input[220]), .B(n2359), .Z(n2361) );
  XOR U2311 ( .A(n2362), .B(n2363), .Z(n2359) );
  AND U2312 ( .A(n59), .B(n2364), .Z(n2363) );
  XNOR U2313 ( .A(p_input[236]), .B(n2362), .Z(n2364) );
  XOR U2314 ( .A(n2365), .B(n2366), .Z(n2362) );
  AND U2315 ( .A(n63), .B(n2367), .Z(n2366) );
  XNOR U2316 ( .A(p_input[252]), .B(n2365), .Z(n2367) );
  XOR U2317 ( .A(n2368), .B(n2369), .Z(n2365) );
  AND U2318 ( .A(n67), .B(n2370), .Z(n2369) );
  XNOR U2319 ( .A(p_input[268]), .B(n2368), .Z(n2370) );
  XOR U2320 ( .A(n2371), .B(n2372), .Z(n2368) );
  AND U2321 ( .A(n71), .B(n2373), .Z(n2372) );
  XNOR U2322 ( .A(p_input[284]), .B(n2371), .Z(n2373) );
  XOR U2323 ( .A(n2374), .B(n2375), .Z(n2371) );
  AND U2324 ( .A(n75), .B(n2376), .Z(n2375) );
  XNOR U2325 ( .A(p_input[300]), .B(n2374), .Z(n2376) );
  XOR U2326 ( .A(n2377), .B(n2378), .Z(n2374) );
  AND U2327 ( .A(n79), .B(n2379), .Z(n2378) );
  XNOR U2328 ( .A(p_input[316]), .B(n2377), .Z(n2379) );
  XOR U2329 ( .A(n2380), .B(n2381), .Z(n2377) );
  AND U2330 ( .A(n83), .B(n2382), .Z(n2381) );
  XNOR U2331 ( .A(p_input[332]), .B(n2380), .Z(n2382) );
  XOR U2332 ( .A(n2383), .B(n2384), .Z(n2380) );
  AND U2333 ( .A(n87), .B(n2385), .Z(n2384) );
  XNOR U2334 ( .A(p_input[348]), .B(n2383), .Z(n2385) );
  XOR U2335 ( .A(n2386), .B(n2387), .Z(n2383) );
  AND U2336 ( .A(n91), .B(n2388), .Z(n2387) );
  XNOR U2337 ( .A(p_input[364]), .B(n2386), .Z(n2388) );
  XOR U2338 ( .A(n2389), .B(n2390), .Z(n2386) );
  AND U2339 ( .A(n95), .B(n2391), .Z(n2390) );
  XNOR U2340 ( .A(p_input[380]), .B(n2389), .Z(n2391) );
  XOR U2341 ( .A(n2392), .B(n2393), .Z(n2389) );
  AND U2342 ( .A(n99), .B(n2394), .Z(n2393) );
  XNOR U2343 ( .A(p_input[396]), .B(n2392), .Z(n2394) );
  XOR U2344 ( .A(n2395), .B(n2396), .Z(n2392) );
  AND U2345 ( .A(n103), .B(n2397), .Z(n2396) );
  XNOR U2346 ( .A(p_input[412]), .B(n2395), .Z(n2397) );
  XOR U2347 ( .A(n2398), .B(n2399), .Z(n2395) );
  AND U2348 ( .A(n107), .B(n2400), .Z(n2399) );
  XNOR U2349 ( .A(p_input[428]), .B(n2398), .Z(n2400) );
  XOR U2350 ( .A(n2401), .B(n2402), .Z(n2398) );
  AND U2351 ( .A(n111), .B(n2403), .Z(n2402) );
  XNOR U2352 ( .A(p_input[444]), .B(n2401), .Z(n2403) );
  XOR U2353 ( .A(n2404), .B(n2405), .Z(n2401) );
  AND U2354 ( .A(n115), .B(n2406), .Z(n2405) );
  XNOR U2355 ( .A(p_input[460]), .B(n2404), .Z(n2406) );
  XOR U2356 ( .A(n2407), .B(n2408), .Z(n2404) );
  AND U2357 ( .A(n119), .B(n2409), .Z(n2408) );
  XNOR U2358 ( .A(p_input[476]), .B(n2407), .Z(n2409) );
  XOR U2359 ( .A(n2410), .B(n2411), .Z(n2407) );
  AND U2360 ( .A(n123), .B(n2412), .Z(n2411) );
  XNOR U2361 ( .A(p_input[492]), .B(n2410), .Z(n2412) );
  XOR U2362 ( .A(n2413), .B(n2414), .Z(n2410) );
  AND U2363 ( .A(n127), .B(n2415), .Z(n2414) );
  XNOR U2364 ( .A(p_input[508]), .B(n2413), .Z(n2415) );
  XOR U2365 ( .A(n2416), .B(n2417), .Z(n2413) );
  AND U2366 ( .A(n131), .B(n2418), .Z(n2417) );
  XNOR U2367 ( .A(p_input[524]), .B(n2416), .Z(n2418) );
  XOR U2368 ( .A(n2419), .B(n2420), .Z(n2416) );
  AND U2369 ( .A(n135), .B(n2421), .Z(n2420) );
  XNOR U2370 ( .A(p_input[540]), .B(n2419), .Z(n2421) );
  XOR U2371 ( .A(n2422), .B(n2423), .Z(n2419) );
  AND U2372 ( .A(n139), .B(n2424), .Z(n2423) );
  XNOR U2373 ( .A(p_input[556]), .B(n2422), .Z(n2424) );
  XOR U2374 ( .A(n2425), .B(n2426), .Z(n2422) );
  AND U2375 ( .A(n143), .B(n2427), .Z(n2426) );
  XNOR U2376 ( .A(p_input[572]), .B(n2425), .Z(n2427) );
  XOR U2377 ( .A(n2428), .B(n2429), .Z(n2425) );
  AND U2378 ( .A(n147), .B(n2430), .Z(n2429) );
  XNOR U2379 ( .A(p_input[588]), .B(n2428), .Z(n2430) );
  XOR U2380 ( .A(n2431), .B(n2432), .Z(n2428) );
  AND U2381 ( .A(n151), .B(n2433), .Z(n2432) );
  XNOR U2382 ( .A(p_input[604]), .B(n2431), .Z(n2433) );
  XOR U2383 ( .A(n2434), .B(n2435), .Z(n2431) );
  AND U2384 ( .A(n155), .B(n2436), .Z(n2435) );
  XNOR U2385 ( .A(p_input[620]), .B(n2434), .Z(n2436) );
  XOR U2386 ( .A(n2437), .B(n2438), .Z(n2434) );
  AND U2387 ( .A(n159), .B(n2439), .Z(n2438) );
  XNOR U2388 ( .A(p_input[636]), .B(n2437), .Z(n2439) );
  XOR U2389 ( .A(n2440), .B(n2441), .Z(n2437) );
  AND U2390 ( .A(n163), .B(n2442), .Z(n2441) );
  XNOR U2391 ( .A(p_input[652]), .B(n2440), .Z(n2442) );
  XOR U2392 ( .A(n2443), .B(n2444), .Z(n2440) );
  AND U2393 ( .A(n167), .B(n2445), .Z(n2444) );
  XNOR U2394 ( .A(p_input[668]), .B(n2443), .Z(n2445) );
  XOR U2395 ( .A(n2446), .B(n2447), .Z(n2443) );
  AND U2396 ( .A(n171), .B(n2448), .Z(n2447) );
  XNOR U2397 ( .A(p_input[684]), .B(n2446), .Z(n2448) );
  XOR U2398 ( .A(n2449), .B(n2450), .Z(n2446) );
  AND U2399 ( .A(n175), .B(n2451), .Z(n2450) );
  XNOR U2400 ( .A(p_input[700]), .B(n2449), .Z(n2451) );
  XOR U2401 ( .A(n2452), .B(n2453), .Z(n2449) );
  AND U2402 ( .A(n179), .B(n2454), .Z(n2453) );
  XNOR U2403 ( .A(p_input[716]), .B(n2452), .Z(n2454) );
  XOR U2404 ( .A(n2455), .B(n2456), .Z(n2452) );
  AND U2405 ( .A(n183), .B(n2457), .Z(n2456) );
  XNOR U2406 ( .A(p_input[732]), .B(n2455), .Z(n2457) );
  XOR U2407 ( .A(n2458), .B(n2459), .Z(n2455) );
  AND U2408 ( .A(n187), .B(n2460), .Z(n2459) );
  XNOR U2409 ( .A(p_input[748]), .B(n2458), .Z(n2460) );
  XOR U2410 ( .A(n2461), .B(n2462), .Z(n2458) );
  AND U2411 ( .A(n191), .B(n2463), .Z(n2462) );
  XNOR U2412 ( .A(p_input[764]), .B(n2461), .Z(n2463) );
  XOR U2413 ( .A(n2464), .B(n2465), .Z(n2461) );
  AND U2414 ( .A(n195), .B(n2466), .Z(n2465) );
  XNOR U2415 ( .A(p_input[780]), .B(n2464), .Z(n2466) );
  XOR U2416 ( .A(n2467), .B(n2468), .Z(n2464) );
  AND U2417 ( .A(n199), .B(n2469), .Z(n2468) );
  XNOR U2418 ( .A(p_input[796]), .B(n2467), .Z(n2469) );
  XOR U2419 ( .A(n2470), .B(n2471), .Z(n2467) );
  AND U2420 ( .A(n203), .B(n2472), .Z(n2471) );
  XNOR U2421 ( .A(p_input[812]), .B(n2470), .Z(n2472) );
  XOR U2422 ( .A(n2473), .B(n2474), .Z(n2470) );
  AND U2423 ( .A(n207), .B(n2475), .Z(n2474) );
  XNOR U2424 ( .A(p_input[828]), .B(n2473), .Z(n2475) );
  XOR U2425 ( .A(n2476), .B(n2477), .Z(n2473) );
  AND U2426 ( .A(n211), .B(n2478), .Z(n2477) );
  XNOR U2427 ( .A(p_input[844]), .B(n2476), .Z(n2478) );
  XOR U2428 ( .A(n2479), .B(n2480), .Z(n2476) );
  AND U2429 ( .A(n215), .B(n2481), .Z(n2480) );
  XNOR U2430 ( .A(p_input[860]), .B(n2479), .Z(n2481) );
  XOR U2431 ( .A(n2482), .B(n2483), .Z(n2479) );
  AND U2432 ( .A(n219), .B(n2484), .Z(n2483) );
  XNOR U2433 ( .A(p_input[876]), .B(n2482), .Z(n2484) );
  XOR U2434 ( .A(n2485), .B(n2486), .Z(n2482) );
  AND U2435 ( .A(n223), .B(n2487), .Z(n2486) );
  XNOR U2436 ( .A(p_input[892]), .B(n2485), .Z(n2487) );
  XOR U2437 ( .A(n2488), .B(n2489), .Z(n2485) );
  AND U2438 ( .A(n227), .B(n2490), .Z(n2489) );
  XNOR U2439 ( .A(p_input[908]), .B(n2488), .Z(n2490) );
  XOR U2440 ( .A(n2491), .B(n2492), .Z(n2488) );
  AND U2441 ( .A(n231), .B(n2493), .Z(n2492) );
  XNOR U2442 ( .A(p_input[924]), .B(n2491), .Z(n2493) );
  XOR U2443 ( .A(n2494), .B(n2495), .Z(n2491) );
  AND U2444 ( .A(n235), .B(n2496), .Z(n2495) );
  XNOR U2445 ( .A(p_input[940]), .B(n2494), .Z(n2496) );
  XOR U2446 ( .A(n2497), .B(n2498), .Z(n2494) );
  AND U2447 ( .A(n239), .B(n2499), .Z(n2498) );
  XNOR U2448 ( .A(p_input[956]), .B(n2497), .Z(n2499) );
  XOR U2449 ( .A(n2500), .B(n2501), .Z(n2497) );
  AND U2450 ( .A(n243), .B(n2502), .Z(n2501) );
  XNOR U2451 ( .A(p_input[972]), .B(n2500), .Z(n2502) );
  XNOR U2452 ( .A(n2503), .B(n2504), .Z(n2500) );
  AND U2453 ( .A(n247), .B(n2505), .Z(n2504) );
  XOR U2454 ( .A(p_input[988]), .B(n2503), .Z(n2505) );
  XOR U2455 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n2506), .Z(n2503) );
  AND U2456 ( .A(n250), .B(n2507), .Z(n2506) );
  XOR U2457 ( .A(p_input[1004]), .B(\knn_comb_/min_val_out[0][12] ), .Z(n2507)
         );
  XNOR U2458 ( .A(n2508), .B(n2509), .Z(o[11]) );
  AND U2459 ( .A(n3), .B(n2510), .Z(n2508) );
  XNOR U2460 ( .A(p_input[11]), .B(n2509), .Z(n2510) );
  XOR U2461 ( .A(n2511), .B(n2512), .Z(n2509) );
  AND U2462 ( .A(n7), .B(n2513), .Z(n2512) );
  XNOR U2463 ( .A(p_input[27]), .B(n2511), .Z(n2513) );
  XOR U2464 ( .A(n2514), .B(n2515), .Z(n2511) );
  AND U2465 ( .A(n11), .B(n2516), .Z(n2515) );
  XNOR U2466 ( .A(p_input[43]), .B(n2514), .Z(n2516) );
  XOR U2467 ( .A(n2517), .B(n2518), .Z(n2514) );
  AND U2468 ( .A(n15), .B(n2519), .Z(n2518) );
  XNOR U2469 ( .A(p_input[59]), .B(n2517), .Z(n2519) );
  XOR U2470 ( .A(n2520), .B(n2521), .Z(n2517) );
  AND U2471 ( .A(n19), .B(n2522), .Z(n2521) );
  XNOR U2472 ( .A(p_input[75]), .B(n2520), .Z(n2522) );
  XOR U2473 ( .A(n2523), .B(n2524), .Z(n2520) );
  AND U2474 ( .A(n23), .B(n2525), .Z(n2524) );
  XNOR U2475 ( .A(p_input[91]), .B(n2523), .Z(n2525) );
  XOR U2476 ( .A(n2526), .B(n2527), .Z(n2523) );
  AND U2477 ( .A(n27), .B(n2528), .Z(n2527) );
  XNOR U2478 ( .A(p_input[107]), .B(n2526), .Z(n2528) );
  XOR U2479 ( .A(n2529), .B(n2530), .Z(n2526) );
  AND U2480 ( .A(n31), .B(n2531), .Z(n2530) );
  XNOR U2481 ( .A(p_input[123]), .B(n2529), .Z(n2531) );
  XOR U2482 ( .A(n2532), .B(n2533), .Z(n2529) );
  AND U2483 ( .A(n35), .B(n2534), .Z(n2533) );
  XNOR U2484 ( .A(p_input[139]), .B(n2532), .Z(n2534) );
  XOR U2485 ( .A(n2535), .B(n2536), .Z(n2532) );
  AND U2486 ( .A(n39), .B(n2537), .Z(n2536) );
  XNOR U2487 ( .A(p_input[155]), .B(n2535), .Z(n2537) );
  XOR U2488 ( .A(n2538), .B(n2539), .Z(n2535) );
  AND U2489 ( .A(n43), .B(n2540), .Z(n2539) );
  XNOR U2490 ( .A(p_input[171]), .B(n2538), .Z(n2540) );
  XOR U2491 ( .A(n2541), .B(n2542), .Z(n2538) );
  AND U2492 ( .A(n47), .B(n2543), .Z(n2542) );
  XNOR U2493 ( .A(p_input[187]), .B(n2541), .Z(n2543) );
  XOR U2494 ( .A(n2544), .B(n2545), .Z(n2541) );
  AND U2495 ( .A(n51), .B(n2546), .Z(n2545) );
  XNOR U2496 ( .A(p_input[203]), .B(n2544), .Z(n2546) );
  XOR U2497 ( .A(n2547), .B(n2548), .Z(n2544) );
  AND U2498 ( .A(n55), .B(n2549), .Z(n2548) );
  XNOR U2499 ( .A(p_input[219]), .B(n2547), .Z(n2549) );
  XOR U2500 ( .A(n2550), .B(n2551), .Z(n2547) );
  AND U2501 ( .A(n59), .B(n2552), .Z(n2551) );
  XNOR U2502 ( .A(p_input[235]), .B(n2550), .Z(n2552) );
  XOR U2503 ( .A(n2553), .B(n2554), .Z(n2550) );
  AND U2504 ( .A(n63), .B(n2555), .Z(n2554) );
  XNOR U2505 ( .A(p_input[251]), .B(n2553), .Z(n2555) );
  XOR U2506 ( .A(n2556), .B(n2557), .Z(n2553) );
  AND U2507 ( .A(n67), .B(n2558), .Z(n2557) );
  XNOR U2508 ( .A(p_input[267]), .B(n2556), .Z(n2558) );
  XOR U2509 ( .A(n2559), .B(n2560), .Z(n2556) );
  AND U2510 ( .A(n71), .B(n2561), .Z(n2560) );
  XNOR U2511 ( .A(p_input[283]), .B(n2559), .Z(n2561) );
  XOR U2512 ( .A(n2562), .B(n2563), .Z(n2559) );
  AND U2513 ( .A(n75), .B(n2564), .Z(n2563) );
  XNOR U2514 ( .A(p_input[299]), .B(n2562), .Z(n2564) );
  XOR U2515 ( .A(n2565), .B(n2566), .Z(n2562) );
  AND U2516 ( .A(n79), .B(n2567), .Z(n2566) );
  XNOR U2517 ( .A(p_input[315]), .B(n2565), .Z(n2567) );
  XOR U2518 ( .A(n2568), .B(n2569), .Z(n2565) );
  AND U2519 ( .A(n83), .B(n2570), .Z(n2569) );
  XNOR U2520 ( .A(p_input[331]), .B(n2568), .Z(n2570) );
  XOR U2521 ( .A(n2571), .B(n2572), .Z(n2568) );
  AND U2522 ( .A(n87), .B(n2573), .Z(n2572) );
  XNOR U2523 ( .A(p_input[347]), .B(n2571), .Z(n2573) );
  XOR U2524 ( .A(n2574), .B(n2575), .Z(n2571) );
  AND U2525 ( .A(n91), .B(n2576), .Z(n2575) );
  XNOR U2526 ( .A(p_input[363]), .B(n2574), .Z(n2576) );
  XOR U2527 ( .A(n2577), .B(n2578), .Z(n2574) );
  AND U2528 ( .A(n95), .B(n2579), .Z(n2578) );
  XNOR U2529 ( .A(p_input[379]), .B(n2577), .Z(n2579) );
  XOR U2530 ( .A(n2580), .B(n2581), .Z(n2577) );
  AND U2531 ( .A(n99), .B(n2582), .Z(n2581) );
  XNOR U2532 ( .A(p_input[395]), .B(n2580), .Z(n2582) );
  XOR U2533 ( .A(n2583), .B(n2584), .Z(n2580) );
  AND U2534 ( .A(n103), .B(n2585), .Z(n2584) );
  XNOR U2535 ( .A(p_input[411]), .B(n2583), .Z(n2585) );
  XOR U2536 ( .A(n2586), .B(n2587), .Z(n2583) );
  AND U2537 ( .A(n107), .B(n2588), .Z(n2587) );
  XNOR U2538 ( .A(p_input[427]), .B(n2586), .Z(n2588) );
  XOR U2539 ( .A(n2589), .B(n2590), .Z(n2586) );
  AND U2540 ( .A(n111), .B(n2591), .Z(n2590) );
  XNOR U2541 ( .A(p_input[443]), .B(n2589), .Z(n2591) );
  XOR U2542 ( .A(n2592), .B(n2593), .Z(n2589) );
  AND U2543 ( .A(n115), .B(n2594), .Z(n2593) );
  XNOR U2544 ( .A(p_input[459]), .B(n2592), .Z(n2594) );
  XOR U2545 ( .A(n2595), .B(n2596), .Z(n2592) );
  AND U2546 ( .A(n119), .B(n2597), .Z(n2596) );
  XNOR U2547 ( .A(p_input[475]), .B(n2595), .Z(n2597) );
  XOR U2548 ( .A(n2598), .B(n2599), .Z(n2595) );
  AND U2549 ( .A(n123), .B(n2600), .Z(n2599) );
  XNOR U2550 ( .A(p_input[491]), .B(n2598), .Z(n2600) );
  XOR U2551 ( .A(n2601), .B(n2602), .Z(n2598) );
  AND U2552 ( .A(n127), .B(n2603), .Z(n2602) );
  XNOR U2553 ( .A(p_input[507]), .B(n2601), .Z(n2603) );
  XOR U2554 ( .A(n2604), .B(n2605), .Z(n2601) );
  AND U2555 ( .A(n131), .B(n2606), .Z(n2605) );
  XNOR U2556 ( .A(p_input[523]), .B(n2604), .Z(n2606) );
  XOR U2557 ( .A(n2607), .B(n2608), .Z(n2604) );
  AND U2558 ( .A(n135), .B(n2609), .Z(n2608) );
  XNOR U2559 ( .A(p_input[539]), .B(n2607), .Z(n2609) );
  XOR U2560 ( .A(n2610), .B(n2611), .Z(n2607) );
  AND U2561 ( .A(n139), .B(n2612), .Z(n2611) );
  XNOR U2562 ( .A(p_input[555]), .B(n2610), .Z(n2612) );
  XOR U2563 ( .A(n2613), .B(n2614), .Z(n2610) );
  AND U2564 ( .A(n143), .B(n2615), .Z(n2614) );
  XNOR U2565 ( .A(p_input[571]), .B(n2613), .Z(n2615) );
  XOR U2566 ( .A(n2616), .B(n2617), .Z(n2613) );
  AND U2567 ( .A(n147), .B(n2618), .Z(n2617) );
  XNOR U2568 ( .A(p_input[587]), .B(n2616), .Z(n2618) );
  XOR U2569 ( .A(n2619), .B(n2620), .Z(n2616) );
  AND U2570 ( .A(n151), .B(n2621), .Z(n2620) );
  XNOR U2571 ( .A(p_input[603]), .B(n2619), .Z(n2621) );
  XOR U2572 ( .A(n2622), .B(n2623), .Z(n2619) );
  AND U2573 ( .A(n155), .B(n2624), .Z(n2623) );
  XNOR U2574 ( .A(p_input[619]), .B(n2622), .Z(n2624) );
  XOR U2575 ( .A(n2625), .B(n2626), .Z(n2622) );
  AND U2576 ( .A(n159), .B(n2627), .Z(n2626) );
  XNOR U2577 ( .A(p_input[635]), .B(n2625), .Z(n2627) );
  XOR U2578 ( .A(n2628), .B(n2629), .Z(n2625) );
  AND U2579 ( .A(n163), .B(n2630), .Z(n2629) );
  XNOR U2580 ( .A(p_input[651]), .B(n2628), .Z(n2630) );
  XOR U2581 ( .A(n2631), .B(n2632), .Z(n2628) );
  AND U2582 ( .A(n167), .B(n2633), .Z(n2632) );
  XNOR U2583 ( .A(p_input[667]), .B(n2631), .Z(n2633) );
  XOR U2584 ( .A(n2634), .B(n2635), .Z(n2631) );
  AND U2585 ( .A(n171), .B(n2636), .Z(n2635) );
  XNOR U2586 ( .A(p_input[683]), .B(n2634), .Z(n2636) );
  XOR U2587 ( .A(n2637), .B(n2638), .Z(n2634) );
  AND U2588 ( .A(n175), .B(n2639), .Z(n2638) );
  XNOR U2589 ( .A(p_input[699]), .B(n2637), .Z(n2639) );
  XOR U2590 ( .A(n2640), .B(n2641), .Z(n2637) );
  AND U2591 ( .A(n179), .B(n2642), .Z(n2641) );
  XNOR U2592 ( .A(p_input[715]), .B(n2640), .Z(n2642) );
  XOR U2593 ( .A(n2643), .B(n2644), .Z(n2640) );
  AND U2594 ( .A(n183), .B(n2645), .Z(n2644) );
  XNOR U2595 ( .A(p_input[731]), .B(n2643), .Z(n2645) );
  XOR U2596 ( .A(n2646), .B(n2647), .Z(n2643) );
  AND U2597 ( .A(n187), .B(n2648), .Z(n2647) );
  XNOR U2598 ( .A(p_input[747]), .B(n2646), .Z(n2648) );
  XOR U2599 ( .A(n2649), .B(n2650), .Z(n2646) );
  AND U2600 ( .A(n191), .B(n2651), .Z(n2650) );
  XNOR U2601 ( .A(p_input[763]), .B(n2649), .Z(n2651) );
  XOR U2602 ( .A(n2652), .B(n2653), .Z(n2649) );
  AND U2603 ( .A(n195), .B(n2654), .Z(n2653) );
  XNOR U2604 ( .A(p_input[779]), .B(n2652), .Z(n2654) );
  XOR U2605 ( .A(n2655), .B(n2656), .Z(n2652) );
  AND U2606 ( .A(n199), .B(n2657), .Z(n2656) );
  XNOR U2607 ( .A(p_input[795]), .B(n2655), .Z(n2657) );
  XOR U2608 ( .A(n2658), .B(n2659), .Z(n2655) );
  AND U2609 ( .A(n203), .B(n2660), .Z(n2659) );
  XNOR U2610 ( .A(p_input[811]), .B(n2658), .Z(n2660) );
  XOR U2611 ( .A(n2661), .B(n2662), .Z(n2658) );
  AND U2612 ( .A(n207), .B(n2663), .Z(n2662) );
  XNOR U2613 ( .A(p_input[827]), .B(n2661), .Z(n2663) );
  XOR U2614 ( .A(n2664), .B(n2665), .Z(n2661) );
  AND U2615 ( .A(n211), .B(n2666), .Z(n2665) );
  XNOR U2616 ( .A(p_input[843]), .B(n2664), .Z(n2666) );
  XOR U2617 ( .A(n2667), .B(n2668), .Z(n2664) );
  AND U2618 ( .A(n215), .B(n2669), .Z(n2668) );
  XNOR U2619 ( .A(p_input[859]), .B(n2667), .Z(n2669) );
  XOR U2620 ( .A(n2670), .B(n2671), .Z(n2667) );
  AND U2621 ( .A(n219), .B(n2672), .Z(n2671) );
  XNOR U2622 ( .A(p_input[875]), .B(n2670), .Z(n2672) );
  XOR U2623 ( .A(n2673), .B(n2674), .Z(n2670) );
  AND U2624 ( .A(n223), .B(n2675), .Z(n2674) );
  XNOR U2625 ( .A(p_input[891]), .B(n2673), .Z(n2675) );
  XOR U2626 ( .A(n2676), .B(n2677), .Z(n2673) );
  AND U2627 ( .A(n227), .B(n2678), .Z(n2677) );
  XNOR U2628 ( .A(p_input[907]), .B(n2676), .Z(n2678) );
  XOR U2629 ( .A(n2679), .B(n2680), .Z(n2676) );
  AND U2630 ( .A(n231), .B(n2681), .Z(n2680) );
  XNOR U2631 ( .A(p_input[923]), .B(n2679), .Z(n2681) );
  XOR U2632 ( .A(n2682), .B(n2683), .Z(n2679) );
  AND U2633 ( .A(n235), .B(n2684), .Z(n2683) );
  XNOR U2634 ( .A(p_input[939]), .B(n2682), .Z(n2684) );
  XOR U2635 ( .A(n2685), .B(n2686), .Z(n2682) );
  AND U2636 ( .A(n239), .B(n2687), .Z(n2686) );
  XNOR U2637 ( .A(p_input[955]), .B(n2685), .Z(n2687) );
  XOR U2638 ( .A(n2688), .B(n2689), .Z(n2685) );
  AND U2639 ( .A(n243), .B(n2690), .Z(n2689) );
  XNOR U2640 ( .A(p_input[971]), .B(n2688), .Z(n2690) );
  XNOR U2641 ( .A(n2691), .B(n2692), .Z(n2688) );
  AND U2642 ( .A(n247), .B(n2693), .Z(n2692) );
  XOR U2643 ( .A(p_input[987]), .B(n2691), .Z(n2693) );
  XOR U2644 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n2694), .Z(n2691) );
  AND U2645 ( .A(n250), .B(n2695), .Z(n2694) );
  XOR U2646 ( .A(p_input[1003]), .B(\knn_comb_/min_val_out[0][11] ), .Z(n2695)
         );
  XNOR U2647 ( .A(n2696), .B(n2697), .Z(o[10]) );
  AND U2648 ( .A(n3), .B(n2698), .Z(n2696) );
  XNOR U2649 ( .A(p_input[10]), .B(n2697), .Z(n2698) );
  XOR U2650 ( .A(n2699), .B(n2700), .Z(n2697) );
  AND U2651 ( .A(n7), .B(n2701), .Z(n2700) );
  XNOR U2652 ( .A(p_input[26]), .B(n2699), .Z(n2701) );
  XOR U2653 ( .A(n2702), .B(n2703), .Z(n2699) );
  AND U2654 ( .A(n11), .B(n2704), .Z(n2703) );
  XNOR U2655 ( .A(p_input[42]), .B(n2702), .Z(n2704) );
  XOR U2656 ( .A(n2705), .B(n2706), .Z(n2702) );
  AND U2657 ( .A(n15), .B(n2707), .Z(n2706) );
  XNOR U2658 ( .A(p_input[58]), .B(n2705), .Z(n2707) );
  XOR U2659 ( .A(n2708), .B(n2709), .Z(n2705) );
  AND U2660 ( .A(n19), .B(n2710), .Z(n2709) );
  XNOR U2661 ( .A(p_input[74]), .B(n2708), .Z(n2710) );
  XOR U2662 ( .A(n2711), .B(n2712), .Z(n2708) );
  AND U2663 ( .A(n23), .B(n2713), .Z(n2712) );
  XNOR U2664 ( .A(p_input[90]), .B(n2711), .Z(n2713) );
  XOR U2665 ( .A(n2714), .B(n2715), .Z(n2711) );
  AND U2666 ( .A(n27), .B(n2716), .Z(n2715) );
  XNOR U2667 ( .A(p_input[106]), .B(n2714), .Z(n2716) );
  XOR U2668 ( .A(n2717), .B(n2718), .Z(n2714) );
  AND U2669 ( .A(n31), .B(n2719), .Z(n2718) );
  XNOR U2670 ( .A(p_input[122]), .B(n2717), .Z(n2719) );
  XOR U2671 ( .A(n2720), .B(n2721), .Z(n2717) );
  AND U2672 ( .A(n35), .B(n2722), .Z(n2721) );
  XNOR U2673 ( .A(p_input[138]), .B(n2720), .Z(n2722) );
  XOR U2674 ( .A(n2723), .B(n2724), .Z(n2720) );
  AND U2675 ( .A(n39), .B(n2725), .Z(n2724) );
  XNOR U2676 ( .A(p_input[154]), .B(n2723), .Z(n2725) );
  XOR U2677 ( .A(n2726), .B(n2727), .Z(n2723) );
  AND U2678 ( .A(n43), .B(n2728), .Z(n2727) );
  XNOR U2679 ( .A(p_input[170]), .B(n2726), .Z(n2728) );
  XOR U2680 ( .A(n2729), .B(n2730), .Z(n2726) );
  AND U2681 ( .A(n47), .B(n2731), .Z(n2730) );
  XNOR U2682 ( .A(p_input[186]), .B(n2729), .Z(n2731) );
  XOR U2683 ( .A(n2732), .B(n2733), .Z(n2729) );
  AND U2684 ( .A(n51), .B(n2734), .Z(n2733) );
  XNOR U2685 ( .A(p_input[202]), .B(n2732), .Z(n2734) );
  XOR U2686 ( .A(n2735), .B(n2736), .Z(n2732) );
  AND U2687 ( .A(n55), .B(n2737), .Z(n2736) );
  XNOR U2688 ( .A(p_input[218]), .B(n2735), .Z(n2737) );
  XOR U2689 ( .A(n2738), .B(n2739), .Z(n2735) );
  AND U2690 ( .A(n59), .B(n2740), .Z(n2739) );
  XNOR U2691 ( .A(p_input[234]), .B(n2738), .Z(n2740) );
  XOR U2692 ( .A(n2741), .B(n2742), .Z(n2738) );
  AND U2693 ( .A(n63), .B(n2743), .Z(n2742) );
  XNOR U2694 ( .A(p_input[250]), .B(n2741), .Z(n2743) );
  XOR U2695 ( .A(n2744), .B(n2745), .Z(n2741) );
  AND U2696 ( .A(n67), .B(n2746), .Z(n2745) );
  XNOR U2697 ( .A(p_input[266]), .B(n2744), .Z(n2746) );
  XOR U2698 ( .A(n2747), .B(n2748), .Z(n2744) );
  AND U2699 ( .A(n71), .B(n2749), .Z(n2748) );
  XNOR U2700 ( .A(p_input[282]), .B(n2747), .Z(n2749) );
  XOR U2701 ( .A(n2750), .B(n2751), .Z(n2747) );
  AND U2702 ( .A(n75), .B(n2752), .Z(n2751) );
  XNOR U2703 ( .A(p_input[298]), .B(n2750), .Z(n2752) );
  XOR U2704 ( .A(n2753), .B(n2754), .Z(n2750) );
  AND U2705 ( .A(n79), .B(n2755), .Z(n2754) );
  XNOR U2706 ( .A(p_input[314]), .B(n2753), .Z(n2755) );
  XOR U2707 ( .A(n2756), .B(n2757), .Z(n2753) );
  AND U2708 ( .A(n83), .B(n2758), .Z(n2757) );
  XNOR U2709 ( .A(p_input[330]), .B(n2756), .Z(n2758) );
  XOR U2710 ( .A(n2759), .B(n2760), .Z(n2756) );
  AND U2711 ( .A(n87), .B(n2761), .Z(n2760) );
  XNOR U2712 ( .A(p_input[346]), .B(n2759), .Z(n2761) );
  XOR U2713 ( .A(n2762), .B(n2763), .Z(n2759) );
  AND U2714 ( .A(n91), .B(n2764), .Z(n2763) );
  XNOR U2715 ( .A(p_input[362]), .B(n2762), .Z(n2764) );
  XOR U2716 ( .A(n2765), .B(n2766), .Z(n2762) );
  AND U2717 ( .A(n95), .B(n2767), .Z(n2766) );
  XNOR U2718 ( .A(p_input[378]), .B(n2765), .Z(n2767) );
  XOR U2719 ( .A(n2768), .B(n2769), .Z(n2765) );
  AND U2720 ( .A(n99), .B(n2770), .Z(n2769) );
  XNOR U2721 ( .A(p_input[394]), .B(n2768), .Z(n2770) );
  XOR U2722 ( .A(n2771), .B(n2772), .Z(n2768) );
  AND U2723 ( .A(n103), .B(n2773), .Z(n2772) );
  XNOR U2724 ( .A(p_input[410]), .B(n2771), .Z(n2773) );
  XOR U2725 ( .A(n2774), .B(n2775), .Z(n2771) );
  AND U2726 ( .A(n107), .B(n2776), .Z(n2775) );
  XNOR U2727 ( .A(p_input[426]), .B(n2774), .Z(n2776) );
  XOR U2728 ( .A(n2777), .B(n2778), .Z(n2774) );
  AND U2729 ( .A(n111), .B(n2779), .Z(n2778) );
  XNOR U2730 ( .A(p_input[442]), .B(n2777), .Z(n2779) );
  XOR U2731 ( .A(n2780), .B(n2781), .Z(n2777) );
  AND U2732 ( .A(n115), .B(n2782), .Z(n2781) );
  XNOR U2733 ( .A(p_input[458]), .B(n2780), .Z(n2782) );
  XOR U2734 ( .A(n2783), .B(n2784), .Z(n2780) );
  AND U2735 ( .A(n119), .B(n2785), .Z(n2784) );
  XNOR U2736 ( .A(p_input[474]), .B(n2783), .Z(n2785) );
  XOR U2737 ( .A(n2786), .B(n2787), .Z(n2783) );
  AND U2738 ( .A(n123), .B(n2788), .Z(n2787) );
  XNOR U2739 ( .A(p_input[490]), .B(n2786), .Z(n2788) );
  XOR U2740 ( .A(n2789), .B(n2790), .Z(n2786) );
  AND U2741 ( .A(n127), .B(n2791), .Z(n2790) );
  XNOR U2742 ( .A(p_input[506]), .B(n2789), .Z(n2791) );
  XOR U2743 ( .A(n2792), .B(n2793), .Z(n2789) );
  AND U2744 ( .A(n131), .B(n2794), .Z(n2793) );
  XNOR U2745 ( .A(p_input[522]), .B(n2792), .Z(n2794) );
  XOR U2746 ( .A(n2795), .B(n2796), .Z(n2792) );
  AND U2747 ( .A(n135), .B(n2797), .Z(n2796) );
  XNOR U2748 ( .A(p_input[538]), .B(n2795), .Z(n2797) );
  XOR U2749 ( .A(n2798), .B(n2799), .Z(n2795) );
  AND U2750 ( .A(n139), .B(n2800), .Z(n2799) );
  XNOR U2751 ( .A(p_input[554]), .B(n2798), .Z(n2800) );
  XOR U2752 ( .A(n2801), .B(n2802), .Z(n2798) );
  AND U2753 ( .A(n143), .B(n2803), .Z(n2802) );
  XNOR U2754 ( .A(p_input[570]), .B(n2801), .Z(n2803) );
  XOR U2755 ( .A(n2804), .B(n2805), .Z(n2801) );
  AND U2756 ( .A(n147), .B(n2806), .Z(n2805) );
  XNOR U2757 ( .A(p_input[586]), .B(n2804), .Z(n2806) );
  XOR U2758 ( .A(n2807), .B(n2808), .Z(n2804) );
  AND U2759 ( .A(n151), .B(n2809), .Z(n2808) );
  XNOR U2760 ( .A(p_input[602]), .B(n2807), .Z(n2809) );
  XOR U2761 ( .A(n2810), .B(n2811), .Z(n2807) );
  AND U2762 ( .A(n155), .B(n2812), .Z(n2811) );
  XNOR U2763 ( .A(p_input[618]), .B(n2810), .Z(n2812) );
  XOR U2764 ( .A(n2813), .B(n2814), .Z(n2810) );
  AND U2765 ( .A(n159), .B(n2815), .Z(n2814) );
  XNOR U2766 ( .A(p_input[634]), .B(n2813), .Z(n2815) );
  XOR U2767 ( .A(n2816), .B(n2817), .Z(n2813) );
  AND U2768 ( .A(n163), .B(n2818), .Z(n2817) );
  XNOR U2769 ( .A(p_input[650]), .B(n2816), .Z(n2818) );
  XOR U2770 ( .A(n2819), .B(n2820), .Z(n2816) );
  AND U2771 ( .A(n167), .B(n2821), .Z(n2820) );
  XNOR U2772 ( .A(p_input[666]), .B(n2819), .Z(n2821) );
  XOR U2773 ( .A(n2822), .B(n2823), .Z(n2819) );
  AND U2774 ( .A(n171), .B(n2824), .Z(n2823) );
  XNOR U2775 ( .A(p_input[682]), .B(n2822), .Z(n2824) );
  XOR U2776 ( .A(n2825), .B(n2826), .Z(n2822) );
  AND U2777 ( .A(n175), .B(n2827), .Z(n2826) );
  XNOR U2778 ( .A(p_input[698]), .B(n2825), .Z(n2827) );
  XOR U2779 ( .A(n2828), .B(n2829), .Z(n2825) );
  AND U2780 ( .A(n179), .B(n2830), .Z(n2829) );
  XNOR U2781 ( .A(p_input[714]), .B(n2828), .Z(n2830) );
  XOR U2782 ( .A(n2831), .B(n2832), .Z(n2828) );
  AND U2783 ( .A(n183), .B(n2833), .Z(n2832) );
  XNOR U2784 ( .A(p_input[730]), .B(n2831), .Z(n2833) );
  XOR U2785 ( .A(n2834), .B(n2835), .Z(n2831) );
  AND U2786 ( .A(n187), .B(n2836), .Z(n2835) );
  XNOR U2787 ( .A(p_input[746]), .B(n2834), .Z(n2836) );
  XOR U2788 ( .A(n2837), .B(n2838), .Z(n2834) );
  AND U2789 ( .A(n191), .B(n2839), .Z(n2838) );
  XNOR U2790 ( .A(p_input[762]), .B(n2837), .Z(n2839) );
  XOR U2791 ( .A(n2840), .B(n2841), .Z(n2837) );
  AND U2792 ( .A(n195), .B(n2842), .Z(n2841) );
  XNOR U2793 ( .A(p_input[778]), .B(n2840), .Z(n2842) );
  XOR U2794 ( .A(n2843), .B(n2844), .Z(n2840) );
  AND U2795 ( .A(n199), .B(n2845), .Z(n2844) );
  XNOR U2796 ( .A(p_input[794]), .B(n2843), .Z(n2845) );
  XOR U2797 ( .A(n2846), .B(n2847), .Z(n2843) );
  AND U2798 ( .A(n203), .B(n2848), .Z(n2847) );
  XNOR U2799 ( .A(p_input[810]), .B(n2846), .Z(n2848) );
  XOR U2800 ( .A(n2849), .B(n2850), .Z(n2846) );
  AND U2801 ( .A(n207), .B(n2851), .Z(n2850) );
  XNOR U2802 ( .A(p_input[826]), .B(n2849), .Z(n2851) );
  XOR U2803 ( .A(n2852), .B(n2853), .Z(n2849) );
  AND U2804 ( .A(n211), .B(n2854), .Z(n2853) );
  XNOR U2805 ( .A(p_input[842]), .B(n2852), .Z(n2854) );
  XOR U2806 ( .A(n2855), .B(n2856), .Z(n2852) );
  AND U2807 ( .A(n215), .B(n2857), .Z(n2856) );
  XNOR U2808 ( .A(p_input[858]), .B(n2855), .Z(n2857) );
  XOR U2809 ( .A(n2858), .B(n2859), .Z(n2855) );
  AND U2810 ( .A(n219), .B(n2860), .Z(n2859) );
  XNOR U2811 ( .A(p_input[874]), .B(n2858), .Z(n2860) );
  XOR U2812 ( .A(n2861), .B(n2862), .Z(n2858) );
  AND U2813 ( .A(n223), .B(n2863), .Z(n2862) );
  XNOR U2814 ( .A(p_input[890]), .B(n2861), .Z(n2863) );
  XOR U2815 ( .A(n2864), .B(n2865), .Z(n2861) );
  AND U2816 ( .A(n227), .B(n2866), .Z(n2865) );
  XNOR U2817 ( .A(p_input[906]), .B(n2864), .Z(n2866) );
  XOR U2818 ( .A(n2867), .B(n2868), .Z(n2864) );
  AND U2819 ( .A(n231), .B(n2869), .Z(n2868) );
  XNOR U2820 ( .A(p_input[922]), .B(n2867), .Z(n2869) );
  XOR U2821 ( .A(n2870), .B(n2871), .Z(n2867) );
  AND U2822 ( .A(n235), .B(n2872), .Z(n2871) );
  XNOR U2823 ( .A(p_input[938]), .B(n2870), .Z(n2872) );
  XOR U2824 ( .A(n2873), .B(n2874), .Z(n2870) );
  AND U2825 ( .A(n239), .B(n2875), .Z(n2874) );
  XNOR U2826 ( .A(p_input[954]), .B(n2873), .Z(n2875) );
  XOR U2827 ( .A(n2876), .B(n2877), .Z(n2873) );
  AND U2828 ( .A(n243), .B(n2878), .Z(n2877) );
  XNOR U2829 ( .A(p_input[970]), .B(n2876), .Z(n2878) );
  XNOR U2830 ( .A(n2879), .B(n2880), .Z(n2876) );
  AND U2831 ( .A(n247), .B(n2881), .Z(n2880) );
  XOR U2832 ( .A(p_input[986]), .B(n2879), .Z(n2881) );
  XOR U2833 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n2882), .Z(n2879) );
  AND U2834 ( .A(n250), .B(n2883), .Z(n2882) );
  XOR U2835 ( .A(p_input[1002]), .B(\knn_comb_/min_val_out[0][10] ), .Z(n2883)
         );
  XNOR U2836 ( .A(n2884), .B(n2885), .Z(o[0]) );
  AND U2837 ( .A(n3), .B(n2886), .Z(n2884) );
  XNOR U2838 ( .A(p_input[0]), .B(n2885), .Z(n2886) );
  XOR U2839 ( .A(n2887), .B(n2888), .Z(n2885) );
  AND U2840 ( .A(n7), .B(n2889), .Z(n2888) );
  XNOR U2841 ( .A(p_input[16]), .B(n2887), .Z(n2889) );
  XOR U2842 ( .A(n2890), .B(n2891), .Z(n2887) );
  AND U2843 ( .A(n11), .B(n2892), .Z(n2891) );
  XNOR U2844 ( .A(p_input[32]), .B(n2890), .Z(n2892) );
  XOR U2845 ( .A(n2893), .B(n2894), .Z(n2890) );
  AND U2846 ( .A(n15), .B(n2895), .Z(n2894) );
  XNOR U2847 ( .A(p_input[48]), .B(n2893), .Z(n2895) );
  XOR U2848 ( .A(n2896), .B(n2897), .Z(n2893) );
  AND U2849 ( .A(n19), .B(n2898), .Z(n2897) );
  XNOR U2850 ( .A(p_input[64]), .B(n2896), .Z(n2898) );
  XOR U2851 ( .A(n2899), .B(n2900), .Z(n2896) );
  AND U2852 ( .A(n23), .B(n2901), .Z(n2900) );
  XNOR U2853 ( .A(p_input[80]), .B(n2899), .Z(n2901) );
  XOR U2854 ( .A(n2902), .B(n2903), .Z(n2899) );
  AND U2855 ( .A(n27), .B(n2904), .Z(n2903) );
  XNOR U2856 ( .A(p_input[96]), .B(n2902), .Z(n2904) );
  XOR U2857 ( .A(n2905), .B(n2906), .Z(n2902) );
  AND U2858 ( .A(n31), .B(n2907), .Z(n2906) );
  XNOR U2859 ( .A(p_input[112]), .B(n2905), .Z(n2907) );
  XOR U2860 ( .A(n2908), .B(n2909), .Z(n2905) );
  AND U2861 ( .A(n35), .B(n2910), .Z(n2909) );
  XNOR U2862 ( .A(p_input[128]), .B(n2908), .Z(n2910) );
  XOR U2863 ( .A(n2911), .B(n2912), .Z(n2908) );
  AND U2864 ( .A(n39), .B(n2913), .Z(n2912) );
  XNOR U2865 ( .A(p_input[144]), .B(n2911), .Z(n2913) );
  XOR U2866 ( .A(n2914), .B(n2915), .Z(n2911) );
  AND U2867 ( .A(n43), .B(n2916), .Z(n2915) );
  XNOR U2868 ( .A(p_input[160]), .B(n2914), .Z(n2916) );
  XOR U2869 ( .A(n2917), .B(n2918), .Z(n2914) );
  AND U2870 ( .A(n47), .B(n2919), .Z(n2918) );
  XNOR U2871 ( .A(p_input[176]), .B(n2917), .Z(n2919) );
  XOR U2872 ( .A(n2920), .B(n2921), .Z(n2917) );
  AND U2873 ( .A(n51), .B(n2922), .Z(n2921) );
  XNOR U2874 ( .A(p_input[192]), .B(n2920), .Z(n2922) );
  XOR U2875 ( .A(n2923), .B(n2924), .Z(n2920) );
  AND U2876 ( .A(n55), .B(n2925), .Z(n2924) );
  XNOR U2877 ( .A(p_input[208]), .B(n2923), .Z(n2925) );
  XOR U2878 ( .A(n2926), .B(n2927), .Z(n2923) );
  AND U2879 ( .A(n59), .B(n2928), .Z(n2927) );
  XNOR U2880 ( .A(p_input[224]), .B(n2926), .Z(n2928) );
  XOR U2881 ( .A(n2929), .B(n2930), .Z(n2926) );
  AND U2882 ( .A(n63), .B(n2931), .Z(n2930) );
  XNOR U2883 ( .A(p_input[240]), .B(n2929), .Z(n2931) );
  XOR U2884 ( .A(n2932), .B(n2933), .Z(n2929) );
  AND U2885 ( .A(n67), .B(n2934), .Z(n2933) );
  XNOR U2886 ( .A(p_input[256]), .B(n2932), .Z(n2934) );
  XOR U2887 ( .A(n2935), .B(n2936), .Z(n2932) );
  AND U2888 ( .A(n71), .B(n2937), .Z(n2936) );
  XNOR U2889 ( .A(p_input[272]), .B(n2935), .Z(n2937) );
  XOR U2890 ( .A(n2938), .B(n2939), .Z(n2935) );
  AND U2891 ( .A(n75), .B(n2940), .Z(n2939) );
  XNOR U2892 ( .A(p_input[288]), .B(n2938), .Z(n2940) );
  XOR U2893 ( .A(n2941), .B(n2942), .Z(n2938) );
  AND U2894 ( .A(n79), .B(n2943), .Z(n2942) );
  XNOR U2895 ( .A(p_input[304]), .B(n2941), .Z(n2943) );
  XOR U2896 ( .A(n2944), .B(n2945), .Z(n2941) );
  AND U2897 ( .A(n83), .B(n2946), .Z(n2945) );
  XNOR U2898 ( .A(p_input[320]), .B(n2944), .Z(n2946) );
  XOR U2899 ( .A(n2947), .B(n2948), .Z(n2944) );
  AND U2900 ( .A(n87), .B(n2949), .Z(n2948) );
  XNOR U2901 ( .A(p_input[336]), .B(n2947), .Z(n2949) );
  XOR U2902 ( .A(n2950), .B(n2951), .Z(n2947) );
  AND U2903 ( .A(n91), .B(n2952), .Z(n2951) );
  XNOR U2904 ( .A(p_input[352]), .B(n2950), .Z(n2952) );
  XOR U2905 ( .A(n2953), .B(n2954), .Z(n2950) );
  AND U2906 ( .A(n95), .B(n2955), .Z(n2954) );
  XNOR U2907 ( .A(p_input[368]), .B(n2953), .Z(n2955) );
  XOR U2908 ( .A(n2956), .B(n2957), .Z(n2953) );
  AND U2909 ( .A(n99), .B(n2958), .Z(n2957) );
  XNOR U2910 ( .A(p_input[384]), .B(n2956), .Z(n2958) );
  XOR U2911 ( .A(n2959), .B(n2960), .Z(n2956) );
  AND U2912 ( .A(n103), .B(n2961), .Z(n2960) );
  XNOR U2913 ( .A(p_input[400]), .B(n2959), .Z(n2961) );
  XOR U2914 ( .A(n2962), .B(n2963), .Z(n2959) );
  AND U2915 ( .A(n107), .B(n2964), .Z(n2963) );
  XNOR U2916 ( .A(p_input[416]), .B(n2962), .Z(n2964) );
  XOR U2917 ( .A(n2965), .B(n2966), .Z(n2962) );
  AND U2918 ( .A(n111), .B(n2967), .Z(n2966) );
  XNOR U2919 ( .A(p_input[432]), .B(n2965), .Z(n2967) );
  XOR U2920 ( .A(n2968), .B(n2969), .Z(n2965) );
  AND U2921 ( .A(n115), .B(n2970), .Z(n2969) );
  XNOR U2922 ( .A(p_input[448]), .B(n2968), .Z(n2970) );
  XOR U2923 ( .A(n2971), .B(n2972), .Z(n2968) );
  AND U2924 ( .A(n119), .B(n2973), .Z(n2972) );
  XNOR U2925 ( .A(p_input[464]), .B(n2971), .Z(n2973) );
  XOR U2926 ( .A(n2974), .B(n2975), .Z(n2971) );
  AND U2927 ( .A(n123), .B(n2976), .Z(n2975) );
  XNOR U2928 ( .A(p_input[480]), .B(n2974), .Z(n2976) );
  XOR U2929 ( .A(n2977), .B(n2978), .Z(n2974) );
  AND U2930 ( .A(n127), .B(n2979), .Z(n2978) );
  XNOR U2931 ( .A(p_input[496]), .B(n2977), .Z(n2979) );
  XOR U2932 ( .A(n2980), .B(n2981), .Z(n2977) );
  AND U2933 ( .A(n131), .B(n2982), .Z(n2981) );
  XNOR U2934 ( .A(p_input[512]), .B(n2980), .Z(n2982) );
  XOR U2935 ( .A(n2983), .B(n2984), .Z(n2980) );
  AND U2936 ( .A(n135), .B(n2985), .Z(n2984) );
  XNOR U2937 ( .A(p_input[528]), .B(n2983), .Z(n2985) );
  XOR U2938 ( .A(n2986), .B(n2987), .Z(n2983) );
  AND U2939 ( .A(n139), .B(n2988), .Z(n2987) );
  XNOR U2940 ( .A(p_input[544]), .B(n2986), .Z(n2988) );
  XOR U2941 ( .A(n2989), .B(n2990), .Z(n2986) );
  AND U2942 ( .A(n143), .B(n2991), .Z(n2990) );
  XNOR U2943 ( .A(p_input[560]), .B(n2989), .Z(n2991) );
  XOR U2944 ( .A(n2992), .B(n2993), .Z(n2989) );
  AND U2945 ( .A(n147), .B(n2994), .Z(n2993) );
  XNOR U2946 ( .A(p_input[576]), .B(n2992), .Z(n2994) );
  XOR U2947 ( .A(n2995), .B(n2996), .Z(n2992) );
  AND U2948 ( .A(n151), .B(n2997), .Z(n2996) );
  XNOR U2949 ( .A(p_input[592]), .B(n2995), .Z(n2997) );
  XOR U2950 ( .A(n2998), .B(n2999), .Z(n2995) );
  AND U2951 ( .A(n155), .B(n3000), .Z(n2999) );
  XNOR U2952 ( .A(p_input[608]), .B(n2998), .Z(n3000) );
  XOR U2953 ( .A(n3001), .B(n3002), .Z(n2998) );
  AND U2954 ( .A(n159), .B(n3003), .Z(n3002) );
  XNOR U2955 ( .A(p_input[624]), .B(n3001), .Z(n3003) );
  XOR U2956 ( .A(n3004), .B(n3005), .Z(n3001) );
  AND U2957 ( .A(n163), .B(n3006), .Z(n3005) );
  XNOR U2958 ( .A(p_input[640]), .B(n3004), .Z(n3006) );
  XOR U2959 ( .A(n3007), .B(n3008), .Z(n3004) );
  AND U2960 ( .A(n167), .B(n3009), .Z(n3008) );
  XNOR U2961 ( .A(p_input[656]), .B(n3007), .Z(n3009) );
  XOR U2962 ( .A(n3010), .B(n3011), .Z(n3007) );
  AND U2963 ( .A(n171), .B(n3012), .Z(n3011) );
  XNOR U2964 ( .A(p_input[672]), .B(n3010), .Z(n3012) );
  XOR U2965 ( .A(n3013), .B(n3014), .Z(n3010) );
  AND U2966 ( .A(n175), .B(n3015), .Z(n3014) );
  XNOR U2967 ( .A(p_input[688]), .B(n3013), .Z(n3015) );
  XOR U2968 ( .A(n3016), .B(n3017), .Z(n3013) );
  AND U2969 ( .A(n179), .B(n3018), .Z(n3017) );
  XNOR U2970 ( .A(p_input[704]), .B(n3016), .Z(n3018) );
  XOR U2971 ( .A(n3019), .B(n3020), .Z(n3016) );
  AND U2972 ( .A(n183), .B(n3021), .Z(n3020) );
  XNOR U2973 ( .A(p_input[720]), .B(n3019), .Z(n3021) );
  XOR U2974 ( .A(n3022), .B(n3023), .Z(n3019) );
  AND U2975 ( .A(n187), .B(n3024), .Z(n3023) );
  XNOR U2976 ( .A(p_input[736]), .B(n3022), .Z(n3024) );
  XOR U2977 ( .A(n3025), .B(n3026), .Z(n3022) );
  AND U2978 ( .A(n191), .B(n3027), .Z(n3026) );
  XNOR U2979 ( .A(p_input[752]), .B(n3025), .Z(n3027) );
  XOR U2980 ( .A(n3028), .B(n3029), .Z(n3025) );
  AND U2981 ( .A(n195), .B(n3030), .Z(n3029) );
  XNOR U2982 ( .A(p_input[768]), .B(n3028), .Z(n3030) );
  XOR U2983 ( .A(n3031), .B(n3032), .Z(n3028) );
  AND U2984 ( .A(n199), .B(n3033), .Z(n3032) );
  XNOR U2985 ( .A(p_input[784]), .B(n3031), .Z(n3033) );
  XOR U2986 ( .A(n3034), .B(n3035), .Z(n3031) );
  AND U2987 ( .A(n203), .B(n3036), .Z(n3035) );
  XNOR U2988 ( .A(p_input[800]), .B(n3034), .Z(n3036) );
  XOR U2989 ( .A(n3037), .B(n3038), .Z(n3034) );
  AND U2990 ( .A(n207), .B(n3039), .Z(n3038) );
  XNOR U2991 ( .A(p_input[816]), .B(n3037), .Z(n3039) );
  XOR U2992 ( .A(n3040), .B(n3041), .Z(n3037) );
  AND U2993 ( .A(n211), .B(n3042), .Z(n3041) );
  XNOR U2994 ( .A(p_input[832]), .B(n3040), .Z(n3042) );
  XOR U2995 ( .A(n3043), .B(n3044), .Z(n3040) );
  AND U2996 ( .A(n215), .B(n3045), .Z(n3044) );
  XNOR U2997 ( .A(p_input[848]), .B(n3043), .Z(n3045) );
  XOR U2998 ( .A(n3046), .B(n3047), .Z(n3043) );
  AND U2999 ( .A(n219), .B(n3048), .Z(n3047) );
  XNOR U3000 ( .A(p_input[864]), .B(n3046), .Z(n3048) );
  XOR U3001 ( .A(n3049), .B(n3050), .Z(n3046) );
  AND U3002 ( .A(n223), .B(n3051), .Z(n3050) );
  XNOR U3003 ( .A(p_input[880]), .B(n3049), .Z(n3051) );
  XOR U3004 ( .A(n3052), .B(n3053), .Z(n3049) );
  AND U3005 ( .A(n227), .B(n3054), .Z(n3053) );
  XNOR U3006 ( .A(p_input[896]), .B(n3052), .Z(n3054) );
  XOR U3007 ( .A(n3055), .B(n3056), .Z(n3052) );
  AND U3008 ( .A(n231), .B(n3057), .Z(n3056) );
  XNOR U3009 ( .A(p_input[912]), .B(n3055), .Z(n3057) );
  XOR U3010 ( .A(n3058), .B(n3059), .Z(n3055) );
  AND U3011 ( .A(n235), .B(n3060), .Z(n3059) );
  XNOR U3012 ( .A(p_input[928]), .B(n3058), .Z(n3060) );
  XOR U3013 ( .A(n3061), .B(n3062), .Z(n3058) );
  AND U3014 ( .A(n239), .B(n3063), .Z(n3062) );
  XNOR U3015 ( .A(p_input[944]), .B(n3061), .Z(n3063) );
  XOR U3016 ( .A(n3064), .B(n3065), .Z(n3061) );
  AND U3017 ( .A(n243), .B(n3066), .Z(n3065) );
  XNOR U3018 ( .A(p_input[960]), .B(n3064), .Z(n3066) );
  XNOR U3019 ( .A(n3067), .B(n3068), .Z(n3064) );
  AND U3020 ( .A(n247), .B(n3069), .Z(n3068) );
  XOR U3021 ( .A(p_input[976]), .B(n3067), .Z(n3069) );
  XOR U3022 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n3070), .Z(n3067) );
  AND U3023 ( .A(n250), .B(n3071), .Z(n3070) );
  XOR U3024 ( .A(p_input[992]), .B(\knn_comb_/min_val_out[0][0] ), .Z(n3071)
         );
  XNOR U3025 ( .A(n3072), .B(n3073), .Z(n3) );
  AND U3026 ( .A(n3074), .B(n3075), .Z(n3073) );
  XOR U3027 ( .A(n3076), .B(n3072), .Z(n3075) );
  AND U3028 ( .A(n3077), .B(n3078), .Z(n3076) );
  XOR U3029 ( .A(n3079), .B(n3072), .Z(n3074) );
  XNOR U3030 ( .A(n3080), .B(n3081), .Z(n3079) );
  AND U3031 ( .A(n7), .B(n3082), .Z(n3081) );
  XOR U3032 ( .A(n3083), .B(n3080), .Z(n3082) );
  XOR U3033 ( .A(n3084), .B(n3085), .Z(n3072) );
  AND U3034 ( .A(n3086), .B(n3087), .Z(n3085) );
  XNOR U3035 ( .A(n3084), .B(n3077), .Z(n3087) );
  XNOR U3036 ( .A(n3088), .B(n3089), .Z(n3077) );
  XOR U3037 ( .A(n3090), .B(n3078), .Z(n3089) );
  AND U3038 ( .A(n3091), .B(n3092), .Z(n3078) );
  AND U3039 ( .A(n3093), .B(n3094), .Z(n3090) );
  XOR U3040 ( .A(n3095), .B(n3088), .Z(n3093) );
  XOR U3041 ( .A(n3096), .B(n3084), .Z(n3086) );
  XNOR U3042 ( .A(n3097), .B(n3098), .Z(n3096) );
  AND U3043 ( .A(n7), .B(n3099), .Z(n3098) );
  XOR U3044 ( .A(n3100), .B(n3097), .Z(n3099) );
  XOR U3045 ( .A(n3101), .B(n3102), .Z(n3084) );
  AND U3046 ( .A(n3103), .B(n3104), .Z(n3102) );
  XNOR U3047 ( .A(n3101), .B(n3091), .Z(n3104) );
  XOR U3048 ( .A(n3105), .B(n3094), .Z(n3091) );
  XNOR U3049 ( .A(n3106), .B(n3088), .Z(n3094) );
  XOR U3050 ( .A(n3107), .B(n3108), .Z(n3088) );
  AND U3051 ( .A(n3109), .B(n3110), .Z(n3108) );
  XOR U3052 ( .A(n3111), .B(n3107), .Z(n3109) );
  XNOR U3053 ( .A(n3112), .B(n3113), .Z(n3106) );
  AND U3054 ( .A(n3114), .B(n3115), .Z(n3113) );
  XOR U3055 ( .A(n3112), .B(n3116), .Z(n3114) );
  XNOR U3056 ( .A(n3095), .B(n3092), .Z(n3105) );
  AND U3057 ( .A(n3117), .B(n3118), .Z(n3092) );
  XOR U3058 ( .A(n3119), .B(n3120), .Z(n3095) );
  AND U3059 ( .A(n3121), .B(n3122), .Z(n3120) );
  XOR U3060 ( .A(n3119), .B(n3123), .Z(n3121) );
  XOR U3061 ( .A(n3124), .B(n3101), .Z(n3103) );
  XNOR U3062 ( .A(n3125), .B(n3126), .Z(n3124) );
  AND U3063 ( .A(n7), .B(n3127), .Z(n3126) );
  XNOR U3064 ( .A(n3128), .B(n3125), .Z(n3127) );
  XOR U3065 ( .A(n3129), .B(n3130), .Z(n3101) );
  AND U3066 ( .A(n3131), .B(n3132), .Z(n3130) );
  XNOR U3067 ( .A(n3129), .B(n3117), .Z(n3132) );
  XOR U3068 ( .A(n3133), .B(n3110), .Z(n3117) );
  XNOR U3069 ( .A(n3134), .B(n3116), .Z(n3110) );
  XOR U3070 ( .A(n3135), .B(n3136), .Z(n3116) );
  NOR U3071 ( .A(n3137), .B(n3138), .Z(n3136) );
  XNOR U3072 ( .A(n3135), .B(n3139), .Z(n3137) );
  XNOR U3073 ( .A(n3115), .B(n3107), .Z(n3134) );
  XOR U3074 ( .A(n3140), .B(n3141), .Z(n3107) );
  AND U3075 ( .A(n3142), .B(n3143), .Z(n3141) );
  XNOR U3076 ( .A(n3140), .B(n3144), .Z(n3142) );
  XNOR U3077 ( .A(n3145), .B(n3112), .Z(n3115) );
  XOR U3078 ( .A(n3146), .B(n3147), .Z(n3112) );
  AND U3079 ( .A(n3148), .B(n3149), .Z(n3147) );
  XOR U3080 ( .A(n3146), .B(n3150), .Z(n3148) );
  XNOR U3081 ( .A(n3151), .B(n3152), .Z(n3145) );
  NOR U3082 ( .A(n3153), .B(n3154), .Z(n3152) );
  XOR U3083 ( .A(n3151), .B(n3155), .Z(n3153) );
  XNOR U3084 ( .A(n3111), .B(n3118), .Z(n3133) );
  NOR U3085 ( .A(n3156), .B(n3157), .Z(n3118) );
  XOR U3086 ( .A(n3123), .B(n3122), .Z(n3111) );
  XNOR U3087 ( .A(n3158), .B(n3119), .Z(n3122) );
  XOR U3088 ( .A(n3159), .B(n3160), .Z(n3119) );
  AND U3089 ( .A(n3161), .B(n3162), .Z(n3160) );
  XNOR U3090 ( .A(n3163), .B(n3164), .Z(n3161) );
  XNOR U3091 ( .A(n3165), .B(n3166), .Z(n3158) );
  NOR U3092 ( .A(n3167), .B(n3168), .Z(n3166) );
  XNOR U3093 ( .A(n3165), .B(n3169), .Z(n3167) );
  XOR U3094 ( .A(n3170), .B(n3171), .Z(n3123) );
  NOR U3095 ( .A(n3172), .B(n3173), .Z(n3171) );
  XNOR U3096 ( .A(n3170), .B(n3174), .Z(n3172) );
  XNOR U3097 ( .A(n3175), .B(n3176), .Z(n3131) );
  XOR U3098 ( .A(n3129), .B(n3177), .Z(n3176) );
  AND U3099 ( .A(n7), .B(n3178), .Z(n3177) );
  XOR U3100 ( .A(n3179), .B(n3175), .Z(n3178) );
  AND U3101 ( .A(n3180), .B(n3156), .Z(n3129) );
  XOR U3102 ( .A(n3181), .B(n3157), .Z(n3156) );
  XNOR U3103 ( .A(p_input[0]), .B(p_input[1024]), .Z(n3157) );
  XOR U3104 ( .A(n3144), .B(n3143), .Z(n3181) );
  XNOR U3105 ( .A(n3182), .B(n3150), .Z(n3143) );
  XNOR U3106 ( .A(n3139), .B(n3138), .Z(n3150) );
  XOR U3107 ( .A(n3183), .B(n3135), .Z(n3138) );
  XOR U3108 ( .A(p_input[1034]), .B(p_input[10]), .Z(n3135) );
  XNOR U3109 ( .A(p_input[1035]), .B(p_input[11]), .Z(n3183) );
  XOR U3110 ( .A(p_input[1036]), .B(p_input[12]), .Z(n3139) );
  XOR U3111 ( .A(n3149), .B(n3184), .Z(n3182) );
  IV U3112 ( .A(n3140), .Z(n3184) );
  XOR U3113 ( .A(p_input[1025]), .B(p_input[1]), .Z(n3140) );
  XOR U3114 ( .A(n3185), .B(n3155), .Z(n3149) );
  XNOR U3115 ( .A(p_input[1039]), .B(p_input[15]), .Z(n3155) );
  XOR U3116 ( .A(n3146), .B(n3154), .Z(n3185) );
  XOR U3117 ( .A(n3186), .B(n3151), .Z(n3154) );
  XOR U3118 ( .A(p_input[1037]), .B(p_input[13]), .Z(n3151) );
  XNOR U3119 ( .A(p_input[1038]), .B(p_input[14]), .Z(n3186) );
  XOR U3120 ( .A(p_input[1033]), .B(p_input[9]), .Z(n3146) );
  XNOR U3121 ( .A(n3164), .B(n3162), .Z(n3144) );
  XNOR U3122 ( .A(n3187), .B(n3169), .Z(n3162) );
  XOR U3123 ( .A(p_input[1032]), .B(p_input[8]), .Z(n3169) );
  XOR U3124 ( .A(n3159), .B(n3168), .Z(n3187) );
  XOR U3125 ( .A(n3188), .B(n3165), .Z(n3168) );
  XOR U3126 ( .A(p_input[1030]), .B(p_input[6]), .Z(n3165) );
  XNOR U3127 ( .A(p_input[1031]), .B(p_input[7]), .Z(n3188) );
  IV U3128 ( .A(n3163), .Z(n3159) );
  XNOR U3129 ( .A(p_input[1026]), .B(p_input[2]), .Z(n3163) );
  XNOR U3130 ( .A(n3174), .B(n3173), .Z(n3164) );
  XOR U3131 ( .A(n3189), .B(n3170), .Z(n3173) );
  XOR U3132 ( .A(p_input[1027]), .B(p_input[3]), .Z(n3170) );
  XNOR U3133 ( .A(p_input[1028]), .B(p_input[4]), .Z(n3189) );
  XOR U3134 ( .A(p_input[1029]), .B(p_input[5]), .Z(n3174) );
  XNOR U3135 ( .A(n3190), .B(n3191), .Z(n3180) );
  AND U3136 ( .A(n7), .B(n3192), .Z(n3191) );
  XNOR U3137 ( .A(n3193), .B(n3194), .Z(n3192) );
  XNOR U3138 ( .A(n3195), .B(n3196), .Z(n7) );
  AND U3139 ( .A(n3197), .B(n3198), .Z(n3196) );
  XOR U3140 ( .A(n3083), .B(n3195), .Z(n3198) );
  AND U3141 ( .A(n3199), .B(n3200), .Z(n3083) );
  XNOR U3142 ( .A(n3080), .B(n3195), .Z(n3197) );
  XOR U3143 ( .A(n3201), .B(n3202), .Z(n3080) );
  AND U3144 ( .A(n11), .B(n3203), .Z(n3202) );
  XOR U3145 ( .A(n3204), .B(n3201), .Z(n3203) );
  XOR U3146 ( .A(n3205), .B(n3206), .Z(n3195) );
  AND U3147 ( .A(n3207), .B(n3208), .Z(n3206) );
  XNOR U3148 ( .A(n3205), .B(n3199), .Z(n3208) );
  IV U3149 ( .A(n3100), .Z(n3199) );
  XOR U3150 ( .A(n3209), .B(n3210), .Z(n3100) );
  XOR U3151 ( .A(n3211), .B(n3200), .Z(n3210) );
  AND U3152 ( .A(n3128), .B(n3212), .Z(n3200) );
  AND U3153 ( .A(n3213), .B(n3214), .Z(n3211) );
  XOR U3154 ( .A(n3215), .B(n3209), .Z(n3213) );
  XNOR U3155 ( .A(n3097), .B(n3205), .Z(n3207) );
  XOR U3156 ( .A(n3216), .B(n3217), .Z(n3097) );
  AND U3157 ( .A(n11), .B(n3218), .Z(n3217) );
  XOR U3158 ( .A(n3219), .B(n3216), .Z(n3218) );
  XOR U3159 ( .A(n3220), .B(n3221), .Z(n3205) );
  AND U3160 ( .A(n3222), .B(n3223), .Z(n3221) );
  XNOR U3161 ( .A(n3220), .B(n3128), .Z(n3223) );
  XOR U3162 ( .A(n3224), .B(n3214), .Z(n3128) );
  XNOR U3163 ( .A(n3225), .B(n3209), .Z(n3214) );
  XOR U3164 ( .A(n3226), .B(n3227), .Z(n3209) );
  AND U3165 ( .A(n3228), .B(n3229), .Z(n3227) );
  XOR U3166 ( .A(n3230), .B(n3226), .Z(n3228) );
  XNOR U3167 ( .A(n3231), .B(n3232), .Z(n3225) );
  AND U3168 ( .A(n3233), .B(n3234), .Z(n3232) );
  XOR U3169 ( .A(n3231), .B(n3235), .Z(n3233) );
  XNOR U3170 ( .A(n3215), .B(n3212), .Z(n3224) );
  AND U3171 ( .A(n3236), .B(n3237), .Z(n3212) );
  XOR U3172 ( .A(n3238), .B(n3239), .Z(n3215) );
  AND U3173 ( .A(n3240), .B(n3241), .Z(n3239) );
  XOR U3174 ( .A(n3238), .B(n3242), .Z(n3240) );
  XNOR U3175 ( .A(n3125), .B(n3220), .Z(n3222) );
  XOR U3176 ( .A(n3243), .B(n3244), .Z(n3125) );
  AND U3177 ( .A(n11), .B(n3245), .Z(n3244) );
  XNOR U3178 ( .A(n3246), .B(n3243), .Z(n3245) );
  XOR U3179 ( .A(n3247), .B(n3248), .Z(n3220) );
  AND U3180 ( .A(n3249), .B(n3250), .Z(n3248) );
  XNOR U3181 ( .A(n3247), .B(n3236), .Z(n3250) );
  IV U3182 ( .A(n3179), .Z(n3236) );
  XNOR U3183 ( .A(n3251), .B(n3229), .Z(n3179) );
  XNOR U3184 ( .A(n3252), .B(n3235), .Z(n3229) );
  XOR U3185 ( .A(n3253), .B(n3254), .Z(n3235) );
  NOR U3186 ( .A(n3255), .B(n3256), .Z(n3254) );
  XNOR U3187 ( .A(n3253), .B(n3257), .Z(n3255) );
  XNOR U3188 ( .A(n3234), .B(n3226), .Z(n3252) );
  XOR U3189 ( .A(n3258), .B(n3259), .Z(n3226) );
  AND U3190 ( .A(n3260), .B(n3261), .Z(n3259) );
  XNOR U3191 ( .A(n3258), .B(n3262), .Z(n3260) );
  XNOR U3192 ( .A(n3263), .B(n3231), .Z(n3234) );
  XOR U3193 ( .A(n3264), .B(n3265), .Z(n3231) );
  AND U3194 ( .A(n3266), .B(n3267), .Z(n3265) );
  XOR U3195 ( .A(n3264), .B(n3268), .Z(n3266) );
  XNOR U3196 ( .A(n3269), .B(n3270), .Z(n3263) );
  NOR U3197 ( .A(n3271), .B(n3272), .Z(n3270) );
  XOR U3198 ( .A(n3269), .B(n3273), .Z(n3271) );
  XNOR U3199 ( .A(n3230), .B(n3237), .Z(n3251) );
  NOR U3200 ( .A(n3193), .B(n3274), .Z(n3237) );
  XOR U3201 ( .A(n3242), .B(n3241), .Z(n3230) );
  XNOR U3202 ( .A(n3275), .B(n3238), .Z(n3241) );
  XOR U3203 ( .A(n3276), .B(n3277), .Z(n3238) );
  AND U3204 ( .A(n3278), .B(n3279), .Z(n3277) );
  XOR U3205 ( .A(n3276), .B(n3280), .Z(n3278) );
  XNOR U3206 ( .A(n3281), .B(n3282), .Z(n3275) );
  NOR U3207 ( .A(n3283), .B(n3284), .Z(n3282) );
  XNOR U3208 ( .A(n3281), .B(n3285), .Z(n3283) );
  XOR U3209 ( .A(n3286), .B(n3287), .Z(n3242) );
  NOR U3210 ( .A(n3288), .B(n3289), .Z(n3287) );
  XNOR U3211 ( .A(n3286), .B(n3290), .Z(n3288) );
  XNOR U3212 ( .A(n3175), .B(n3247), .Z(n3249) );
  XOR U3213 ( .A(n3291), .B(n3292), .Z(n3175) );
  AND U3214 ( .A(n11), .B(n3293), .Z(n3292) );
  XOR U3215 ( .A(n3294), .B(n3291), .Z(n3293) );
  AND U3216 ( .A(n3194), .B(n3193), .Z(n3247) );
  XOR U3217 ( .A(n3295), .B(n3274), .Z(n3193) );
  XNOR U3218 ( .A(p_input[1024]), .B(p_input[16]), .Z(n3274) );
  XOR U3219 ( .A(n3262), .B(n3261), .Z(n3295) );
  XNOR U3220 ( .A(n3296), .B(n3268), .Z(n3261) );
  XNOR U3221 ( .A(n3257), .B(n3256), .Z(n3268) );
  XOR U3222 ( .A(n3297), .B(n3253), .Z(n3256) );
  XOR U3223 ( .A(p_input[1034]), .B(p_input[26]), .Z(n3253) );
  XNOR U3224 ( .A(p_input[1035]), .B(p_input[27]), .Z(n3297) );
  XOR U3225 ( .A(p_input[1036]), .B(p_input[28]), .Z(n3257) );
  XNOR U3226 ( .A(n3267), .B(n3258), .Z(n3296) );
  XNOR U3227 ( .A(n3298), .B(p_input[17]), .Z(n3258) );
  XOR U3228 ( .A(n3299), .B(n3273), .Z(n3267) );
  XNOR U3229 ( .A(p_input[1039]), .B(p_input[31]), .Z(n3273) );
  XOR U3230 ( .A(n3264), .B(n3272), .Z(n3299) );
  XOR U3231 ( .A(n3300), .B(n3269), .Z(n3272) );
  XOR U3232 ( .A(p_input[1037]), .B(p_input[29]), .Z(n3269) );
  XNOR U3233 ( .A(p_input[1038]), .B(p_input[30]), .Z(n3300) );
  XOR U3234 ( .A(p_input[1033]), .B(p_input[25]), .Z(n3264) );
  XNOR U3235 ( .A(n3280), .B(n3279), .Z(n3262) );
  XNOR U3236 ( .A(n3301), .B(n3285), .Z(n3279) );
  XOR U3237 ( .A(p_input[1032]), .B(p_input[24]), .Z(n3285) );
  XOR U3238 ( .A(n3276), .B(n3284), .Z(n3301) );
  XOR U3239 ( .A(n3302), .B(n3281), .Z(n3284) );
  XOR U3240 ( .A(p_input[1030]), .B(p_input[22]), .Z(n3281) );
  XNOR U3241 ( .A(p_input[1031]), .B(p_input[23]), .Z(n3302) );
  XOR U3242 ( .A(p_input[1026]), .B(p_input[18]), .Z(n3276) );
  XNOR U3243 ( .A(n3290), .B(n3289), .Z(n3280) );
  XOR U3244 ( .A(n3303), .B(n3286), .Z(n3289) );
  XOR U3245 ( .A(p_input[1027]), .B(p_input[19]), .Z(n3286) );
  XNOR U3246 ( .A(p_input[1028]), .B(p_input[20]), .Z(n3303) );
  XOR U3247 ( .A(p_input[1029]), .B(p_input[21]), .Z(n3290) );
  IV U3248 ( .A(n3190), .Z(n3194) );
  XNOR U3249 ( .A(n3304), .B(n3305), .Z(n3190) );
  AND U3250 ( .A(n11), .B(n3306), .Z(n3305) );
  XNOR U3251 ( .A(n3307), .B(n3304), .Z(n3306) );
  XNOR U3252 ( .A(n3308), .B(n3309), .Z(n11) );
  AND U3253 ( .A(n3310), .B(n3311), .Z(n3309) );
  XOR U3254 ( .A(n3204), .B(n3308), .Z(n3311) );
  AND U3255 ( .A(n3312), .B(n3313), .Z(n3204) );
  XNOR U3256 ( .A(n3201), .B(n3308), .Z(n3310) );
  XOR U3257 ( .A(n3314), .B(n3315), .Z(n3201) );
  AND U3258 ( .A(n15), .B(n3316), .Z(n3315) );
  XOR U3259 ( .A(n3317), .B(n3314), .Z(n3316) );
  XOR U3260 ( .A(n3318), .B(n3319), .Z(n3308) );
  AND U3261 ( .A(n3320), .B(n3321), .Z(n3319) );
  XNOR U3262 ( .A(n3318), .B(n3312), .Z(n3321) );
  IV U3263 ( .A(n3219), .Z(n3312) );
  XOR U3264 ( .A(n3322), .B(n3323), .Z(n3219) );
  XOR U3265 ( .A(n3324), .B(n3313), .Z(n3323) );
  AND U3266 ( .A(n3246), .B(n3325), .Z(n3313) );
  AND U3267 ( .A(n3326), .B(n3327), .Z(n3324) );
  XOR U3268 ( .A(n3328), .B(n3322), .Z(n3326) );
  XNOR U3269 ( .A(n3216), .B(n3318), .Z(n3320) );
  XOR U3270 ( .A(n3329), .B(n3330), .Z(n3216) );
  AND U3271 ( .A(n15), .B(n3331), .Z(n3330) );
  XOR U3272 ( .A(n3332), .B(n3329), .Z(n3331) );
  XOR U3273 ( .A(n3333), .B(n3334), .Z(n3318) );
  AND U3274 ( .A(n3335), .B(n3336), .Z(n3334) );
  XNOR U3275 ( .A(n3333), .B(n3246), .Z(n3336) );
  XOR U3276 ( .A(n3337), .B(n3327), .Z(n3246) );
  XNOR U3277 ( .A(n3338), .B(n3322), .Z(n3327) );
  XOR U3278 ( .A(n3339), .B(n3340), .Z(n3322) );
  AND U3279 ( .A(n3341), .B(n3342), .Z(n3340) );
  XOR U3280 ( .A(n3343), .B(n3339), .Z(n3341) );
  XNOR U3281 ( .A(n3344), .B(n3345), .Z(n3338) );
  AND U3282 ( .A(n3346), .B(n3347), .Z(n3345) );
  XOR U3283 ( .A(n3344), .B(n3348), .Z(n3346) );
  XNOR U3284 ( .A(n3328), .B(n3325), .Z(n3337) );
  AND U3285 ( .A(n3349), .B(n3350), .Z(n3325) );
  XOR U3286 ( .A(n3351), .B(n3352), .Z(n3328) );
  AND U3287 ( .A(n3353), .B(n3354), .Z(n3352) );
  XOR U3288 ( .A(n3351), .B(n3355), .Z(n3353) );
  XNOR U3289 ( .A(n3243), .B(n3333), .Z(n3335) );
  XOR U3290 ( .A(n3356), .B(n3357), .Z(n3243) );
  AND U3291 ( .A(n15), .B(n3358), .Z(n3357) );
  XNOR U3292 ( .A(n3359), .B(n3356), .Z(n3358) );
  XOR U3293 ( .A(n3360), .B(n3361), .Z(n3333) );
  AND U3294 ( .A(n3362), .B(n3363), .Z(n3361) );
  XNOR U3295 ( .A(n3360), .B(n3349), .Z(n3363) );
  IV U3296 ( .A(n3294), .Z(n3349) );
  XNOR U3297 ( .A(n3364), .B(n3342), .Z(n3294) );
  XNOR U3298 ( .A(n3365), .B(n3348), .Z(n3342) );
  XOR U3299 ( .A(n3366), .B(n3367), .Z(n3348) );
  NOR U3300 ( .A(n3368), .B(n3369), .Z(n3367) );
  XNOR U3301 ( .A(n3366), .B(n3370), .Z(n3368) );
  XNOR U3302 ( .A(n3347), .B(n3339), .Z(n3365) );
  XOR U3303 ( .A(n3371), .B(n3372), .Z(n3339) );
  AND U3304 ( .A(n3373), .B(n3374), .Z(n3372) );
  XNOR U3305 ( .A(n3371), .B(n3375), .Z(n3373) );
  XNOR U3306 ( .A(n3376), .B(n3344), .Z(n3347) );
  XOR U3307 ( .A(n3377), .B(n3378), .Z(n3344) );
  AND U3308 ( .A(n3379), .B(n3380), .Z(n3378) );
  XOR U3309 ( .A(n3377), .B(n3381), .Z(n3379) );
  XNOR U3310 ( .A(n3382), .B(n3383), .Z(n3376) );
  NOR U3311 ( .A(n3384), .B(n3385), .Z(n3383) );
  XOR U3312 ( .A(n3382), .B(n3386), .Z(n3384) );
  XNOR U3313 ( .A(n3343), .B(n3350), .Z(n3364) );
  NOR U3314 ( .A(n3307), .B(n3387), .Z(n3350) );
  XOR U3315 ( .A(n3355), .B(n3354), .Z(n3343) );
  XNOR U3316 ( .A(n3388), .B(n3351), .Z(n3354) );
  XOR U3317 ( .A(n3389), .B(n3390), .Z(n3351) );
  AND U3318 ( .A(n3391), .B(n3392), .Z(n3390) );
  XOR U3319 ( .A(n3389), .B(n3393), .Z(n3391) );
  XNOR U3320 ( .A(n3394), .B(n3395), .Z(n3388) );
  NOR U3321 ( .A(n3396), .B(n3397), .Z(n3395) );
  XNOR U3322 ( .A(n3394), .B(n3398), .Z(n3396) );
  XOR U3323 ( .A(n3399), .B(n3400), .Z(n3355) );
  NOR U3324 ( .A(n3401), .B(n3402), .Z(n3400) );
  XNOR U3325 ( .A(n3399), .B(n3403), .Z(n3401) );
  XNOR U3326 ( .A(n3291), .B(n3360), .Z(n3362) );
  XOR U3327 ( .A(n3404), .B(n3405), .Z(n3291) );
  AND U3328 ( .A(n15), .B(n3406), .Z(n3405) );
  XOR U3329 ( .A(n3407), .B(n3404), .Z(n3406) );
  AND U3330 ( .A(n3304), .B(n3307), .Z(n3360) );
  XOR U3331 ( .A(n3408), .B(n3387), .Z(n3307) );
  XNOR U3332 ( .A(p_input[1024]), .B(p_input[32]), .Z(n3387) );
  XOR U3333 ( .A(n3375), .B(n3374), .Z(n3408) );
  XNOR U3334 ( .A(n3409), .B(n3381), .Z(n3374) );
  XNOR U3335 ( .A(n3370), .B(n3369), .Z(n3381) );
  XOR U3336 ( .A(n3410), .B(n3366), .Z(n3369) );
  XOR U3337 ( .A(p_input[1034]), .B(p_input[42]), .Z(n3366) );
  XNOR U3338 ( .A(p_input[1035]), .B(p_input[43]), .Z(n3410) );
  XOR U3339 ( .A(p_input[1036]), .B(p_input[44]), .Z(n3370) );
  XNOR U3340 ( .A(n3380), .B(n3371), .Z(n3409) );
  XNOR U3341 ( .A(n3298), .B(p_input[33]), .Z(n3371) );
  XOR U3342 ( .A(n3411), .B(n3386), .Z(n3380) );
  XNOR U3343 ( .A(p_input[1039]), .B(p_input[47]), .Z(n3386) );
  XOR U3344 ( .A(n3377), .B(n3385), .Z(n3411) );
  XOR U3345 ( .A(n3412), .B(n3382), .Z(n3385) );
  XOR U3346 ( .A(p_input[1037]), .B(p_input[45]), .Z(n3382) );
  XNOR U3347 ( .A(p_input[1038]), .B(p_input[46]), .Z(n3412) );
  XOR U3348 ( .A(p_input[1033]), .B(p_input[41]), .Z(n3377) );
  XNOR U3349 ( .A(n3393), .B(n3392), .Z(n3375) );
  XNOR U3350 ( .A(n3413), .B(n3398), .Z(n3392) );
  XOR U3351 ( .A(p_input[1032]), .B(p_input[40]), .Z(n3398) );
  XOR U3352 ( .A(n3389), .B(n3397), .Z(n3413) );
  XOR U3353 ( .A(n3414), .B(n3394), .Z(n3397) );
  XOR U3354 ( .A(p_input[1030]), .B(p_input[38]), .Z(n3394) );
  XNOR U3355 ( .A(p_input[1031]), .B(p_input[39]), .Z(n3414) );
  XOR U3356 ( .A(p_input[1026]), .B(p_input[34]), .Z(n3389) );
  XNOR U3357 ( .A(n3403), .B(n3402), .Z(n3393) );
  XOR U3358 ( .A(n3415), .B(n3399), .Z(n3402) );
  XOR U3359 ( .A(p_input[1027]), .B(p_input[35]), .Z(n3399) );
  XNOR U3360 ( .A(p_input[1028]), .B(p_input[36]), .Z(n3415) );
  XOR U3361 ( .A(p_input[1029]), .B(p_input[37]), .Z(n3403) );
  XOR U3362 ( .A(n3416), .B(n3417), .Z(n3304) );
  AND U3363 ( .A(n15), .B(n3418), .Z(n3417) );
  XNOR U3364 ( .A(n3419), .B(n3416), .Z(n3418) );
  XNOR U3365 ( .A(n3420), .B(n3421), .Z(n15) );
  AND U3366 ( .A(n3422), .B(n3423), .Z(n3421) );
  XOR U3367 ( .A(n3317), .B(n3420), .Z(n3423) );
  AND U3368 ( .A(n3424), .B(n3425), .Z(n3317) );
  XNOR U3369 ( .A(n3314), .B(n3420), .Z(n3422) );
  XOR U3370 ( .A(n3426), .B(n3427), .Z(n3314) );
  AND U3371 ( .A(n19), .B(n3428), .Z(n3427) );
  XOR U3372 ( .A(n3429), .B(n3426), .Z(n3428) );
  XOR U3373 ( .A(n3430), .B(n3431), .Z(n3420) );
  AND U3374 ( .A(n3432), .B(n3433), .Z(n3431) );
  XNOR U3375 ( .A(n3430), .B(n3424), .Z(n3433) );
  IV U3376 ( .A(n3332), .Z(n3424) );
  XOR U3377 ( .A(n3434), .B(n3435), .Z(n3332) );
  XOR U3378 ( .A(n3436), .B(n3425), .Z(n3435) );
  AND U3379 ( .A(n3359), .B(n3437), .Z(n3425) );
  AND U3380 ( .A(n3438), .B(n3439), .Z(n3436) );
  XOR U3381 ( .A(n3440), .B(n3434), .Z(n3438) );
  XNOR U3382 ( .A(n3329), .B(n3430), .Z(n3432) );
  XOR U3383 ( .A(n3441), .B(n3442), .Z(n3329) );
  AND U3384 ( .A(n19), .B(n3443), .Z(n3442) );
  XOR U3385 ( .A(n3444), .B(n3441), .Z(n3443) );
  XOR U3386 ( .A(n3445), .B(n3446), .Z(n3430) );
  AND U3387 ( .A(n3447), .B(n3448), .Z(n3446) );
  XNOR U3388 ( .A(n3445), .B(n3359), .Z(n3448) );
  XOR U3389 ( .A(n3449), .B(n3439), .Z(n3359) );
  XNOR U3390 ( .A(n3450), .B(n3434), .Z(n3439) );
  XOR U3391 ( .A(n3451), .B(n3452), .Z(n3434) );
  AND U3392 ( .A(n3453), .B(n3454), .Z(n3452) );
  XOR U3393 ( .A(n3455), .B(n3451), .Z(n3453) );
  XNOR U3394 ( .A(n3456), .B(n3457), .Z(n3450) );
  AND U3395 ( .A(n3458), .B(n3459), .Z(n3457) );
  XOR U3396 ( .A(n3456), .B(n3460), .Z(n3458) );
  XNOR U3397 ( .A(n3440), .B(n3437), .Z(n3449) );
  AND U3398 ( .A(n3461), .B(n3462), .Z(n3437) );
  XOR U3399 ( .A(n3463), .B(n3464), .Z(n3440) );
  AND U3400 ( .A(n3465), .B(n3466), .Z(n3464) );
  XOR U3401 ( .A(n3463), .B(n3467), .Z(n3465) );
  XNOR U3402 ( .A(n3356), .B(n3445), .Z(n3447) );
  XOR U3403 ( .A(n3468), .B(n3469), .Z(n3356) );
  AND U3404 ( .A(n19), .B(n3470), .Z(n3469) );
  XNOR U3405 ( .A(n3471), .B(n3468), .Z(n3470) );
  XOR U3406 ( .A(n3472), .B(n3473), .Z(n3445) );
  AND U3407 ( .A(n3474), .B(n3475), .Z(n3473) );
  XNOR U3408 ( .A(n3472), .B(n3461), .Z(n3475) );
  IV U3409 ( .A(n3407), .Z(n3461) );
  XNOR U3410 ( .A(n3476), .B(n3454), .Z(n3407) );
  XNOR U3411 ( .A(n3477), .B(n3460), .Z(n3454) );
  XOR U3412 ( .A(n3478), .B(n3479), .Z(n3460) );
  NOR U3413 ( .A(n3480), .B(n3481), .Z(n3479) );
  XNOR U3414 ( .A(n3478), .B(n3482), .Z(n3480) );
  XNOR U3415 ( .A(n3459), .B(n3451), .Z(n3477) );
  XOR U3416 ( .A(n3483), .B(n3484), .Z(n3451) );
  AND U3417 ( .A(n3485), .B(n3486), .Z(n3484) );
  XNOR U3418 ( .A(n3483), .B(n3487), .Z(n3485) );
  XNOR U3419 ( .A(n3488), .B(n3456), .Z(n3459) );
  XOR U3420 ( .A(n3489), .B(n3490), .Z(n3456) );
  AND U3421 ( .A(n3491), .B(n3492), .Z(n3490) );
  XOR U3422 ( .A(n3489), .B(n3493), .Z(n3491) );
  XNOR U3423 ( .A(n3494), .B(n3495), .Z(n3488) );
  NOR U3424 ( .A(n3496), .B(n3497), .Z(n3495) );
  XOR U3425 ( .A(n3494), .B(n3498), .Z(n3496) );
  XNOR U3426 ( .A(n3455), .B(n3462), .Z(n3476) );
  NOR U3427 ( .A(n3419), .B(n3499), .Z(n3462) );
  XOR U3428 ( .A(n3467), .B(n3466), .Z(n3455) );
  XNOR U3429 ( .A(n3500), .B(n3463), .Z(n3466) );
  XOR U3430 ( .A(n3501), .B(n3502), .Z(n3463) );
  AND U3431 ( .A(n3503), .B(n3504), .Z(n3502) );
  XOR U3432 ( .A(n3501), .B(n3505), .Z(n3503) );
  XNOR U3433 ( .A(n3506), .B(n3507), .Z(n3500) );
  NOR U3434 ( .A(n3508), .B(n3509), .Z(n3507) );
  XNOR U3435 ( .A(n3506), .B(n3510), .Z(n3508) );
  XOR U3436 ( .A(n3511), .B(n3512), .Z(n3467) );
  NOR U3437 ( .A(n3513), .B(n3514), .Z(n3512) );
  XNOR U3438 ( .A(n3511), .B(n3515), .Z(n3513) );
  XNOR U3439 ( .A(n3404), .B(n3472), .Z(n3474) );
  XOR U3440 ( .A(n3516), .B(n3517), .Z(n3404) );
  AND U3441 ( .A(n19), .B(n3518), .Z(n3517) );
  XOR U3442 ( .A(n3519), .B(n3516), .Z(n3518) );
  AND U3443 ( .A(n3416), .B(n3419), .Z(n3472) );
  XOR U3444 ( .A(n3520), .B(n3499), .Z(n3419) );
  XNOR U3445 ( .A(p_input[1024]), .B(p_input[48]), .Z(n3499) );
  XOR U3446 ( .A(n3487), .B(n3486), .Z(n3520) );
  XNOR U3447 ( .A(n3521), .B(n3493), .Z(n3486) );
  XNOR U3448 ( .A(n3482), .B(n3481), .Z(n3493) );
  XOR U3449 ( .A(n3522), .B(n3478), .Z(n3481) );
  XOR U3450 ( .A(p_input[1034]), .B(p_input[58]), .Z(n3478) );
  XNOR U3451 ( .A(p_input[1035]), .B(p_input[59]), .Z(n3522) );
  XOR U3452 ( .A(p_input[1036]), .B(p_input[60]), .Z(n3482) );
  XNOR U3453 ( .A(n3492), .B(n3483), .Z(n3521) );
  XNOR U3454 ( .A(n3298), .B(p_input[49]), .Z(n3483) );
  XOR U3455 ( .A(n3523), .B(n3498), .Z(n3492) );
  XNOR U3456 ( .A(p_input[1039]), .B(p_input[63]), .Z(n3498) );
  XOR U3457 ( .A(n3489), .B(n3497), .Z(n3523) );
  XOR U3458 ( .A(n3524), .B(n3494), .Z(n3497) );
  XOR U3459 ( .A(p_input[1037]), .B(p_input[61]), .Z(n3494) );
  XNOR U3460 ( .A(p_input[1038]), .B(p_input[62]), .Z(n3524) );
  XOR U3461 ( .A(p_input[1033]), .B(p_input[57]), .Z(n3489) );
  XNOR U3462 ( .A(n3505), .B(n3504), .Z(n3487) );
  XNOR U3463 ( .A(n3525), .B(n3510), .Z(n3504) );
  XOR U3464 ( .A(p_input[1032]), .B(p_input[56]), .Z(n3510) );
  XOR U3465 ( .A(n3501), .B(n3509), .Z(n3525) );
  XOR U3466 ( .A(n3526), .B(n3506), .Z(n3509) );
  XOR U3467 ( .A(p_input[1030]), .B(p_input[54]), .Z(n3506) );
  XNOR U3468 ( .A(p_input[1031]), .B(p_input[55]), .Z(n3526) );
  XOR U3469 ( .A(p_input[1026]), .B(p_input[50]), .Z(n3501) );
  XNOR U3470 ( .A(n3515), .B(n3514), .Z(n3505) );
  XOR U3471 ( .A(n3527), .B(n3511), .Z(n3514) );
  XOR U3472 ( .A(p_input[1027]), .B(p_input[51]), .Z(n3511) );
  XNOR U3473 ( .A(p_input[1028]), .B(p_input[52]), .Z(n3527) );
  XOR U3474 ( .A(p_input[1029]), .B(p_input[53]), .Z(n3515) );
  XOR U3475 ( .A(n3528), .B(n3529), .Z(n3416) );
  AND U3476 ( .A(n19), .B(n3530), .Z(n3529) );
  XNOR U3477 ( .A(n3531), .B(n3528), .Z(n3530) );
  XNOR U3478 ( .A(n3532), .B(n3533), .Z(n19) );
  AND U3479 ( .A(n3534), .B(n3535), .Z(n3533) );
  XOR U3480 ( .A(n3429), .B(n3532), .Z(n3535) );
  AND U3481 ( .A(n3536), .B(n3537), .Z(n3429) );
  XNOR U3482 ( .A(n3426), .B(n3532), .Z(n3534) );
  XOR U3483 ( .A(n3538), .B(n3539), .Z(n3426) );
  AND U3484 ( .A(n23), .B(n3540), .Z(n3539) );
  XOR U3485 ( .A(n3541), .B(n3538), .Z(n3540) );
  XOR U3486 ( .A(n3542), .B(n3543), .Z(n3532) );
  AND U3487 ( .A(n3544), .B(n3545), .Z(n3543) );
  XNOR U3488 ( .A(n3542), .B(n3536), .Z(n3545) );
  IV U3489 ( .A(n3444), .Z(n3536) );
  XOR U3490 ( .A(n3546), .B(n3547), .Z(n3444) );
  XOR U3491 ( .A(n3548), .B(n3537), .Z(n3547) );
  AND U3492 ( .A(n3471), .B(n3549), .Z(n3537) );
  AND U3493 ( .A(n3550), .B(n3551), .Z(n3548) );
  XOR U3494 ( .A(n3552), .B(n3546), .Z(n3550) );
  XNOR U3495 ( .A(n3441), .B(n3542), .Z(n3544) );
  XOR U3496 ( .A(n3553), .B(n3554), .Z(n3441) );
  AND U3497 ( .A(n23), .B(n3555), .Z(n3554) );
  XOR U3498 ( .A(n3556), .B(n3553), .Z(n3555) );
  XOR U3499 ( .A(n3557), .B(n3558), .Z(n3542) );
  AND U3500 ( .A(n3559), .B(n3560), .Z(n3558) );
  XNOR U3501 ( .A(n3557), .B(n3471), .Z(n3560) );
  XOR U3502 ( .A(n3561), .B(n3551), .Z(n3471) );
  XNOR U3503 ( .A(n3562), .B(n3546), .Z(n3551) );
  XOR U3504 ( .A(n3563), .B(n3564), .Z(n3546) );
  AND U3505 ( .A(n3565), .B(n3566), .Z(n3564) );
  XOR U3506 ( .A(n3567), .B(n3563), .Z(n3565) );
  XNOR U3507 ( .A(n3568), .B(n3569), .Z(n3562) );
  AND U3508 ( .A(n3570), .B(n3571), .Z(n3569) );
  XOR U3509 ( .A(n3568), .B(n3572), .Z(n3570) );
  XNOR U3510 ( .A(n3552), .B(n3549), .Z(n3561) );
  AND U3511 ( .A(n3573), .B(n3574), .Z(n3549) );
  XOR U3512 ( .A(n3575), .B(n3576), .Z(n3552) );
  AND U3513 ( .A(n3577), .B(n3578), .Z(n3576) );
  XOR U3514 ( .A(n3575), .B(n3579), .Z(n3577) );
  XNOR U3515 ( .A(n3468), .B(n3557), .Z(n3559) );
  XOR U3516 ( .A(n3580), .B(n3581), .Z(n3468) );
  AND U3517 ( .A(n23), .B(n3582), .Z(n3581) );
  XNOR U3518 ( .A(n3583), .B(n3580), .Z(n3582) );
  XOR U3519 ( .A(n3584), .B(n3585), .Z(n3557) );
  AND U3520 ( .A(n3586), .B(n3587), .Z(n3585) );
  XNOR U3521 ( .A(n3584), .B(n3573), .Z(n3587) );
  IV U3522 ( .A(n3519), .Z(n3573) );
  XNOR U3523 ( .A(n3588), .B(n3566), .Z(n3519) );
  XNOR U3524 ( .A(n3589), .B(n3572), .Z(n3566) );
  XOR U3525 ( .A(n3590), .B(n3591), .Z(n3572) );
  NOR U3526 ( .A(n3592), .B(n3593), .Z(n3591) );
  XNOR U3527 ( .A(n3590), .B(n3594), .Z(n3592) );
  XNOR U3528 ( .A(n3571), .B(n3563), .Z(n3589) );
  XOR U3529 ( .A(n3595), .B(n3596), .Z(n3563) );
  AND U3530 ( .A(n3597), .B(n3598), .Z(n3596) );
  XNOR U3531 ( .A(n3595), .B(n3599), .Z(n3597) );
  XNOR U3532 ( .A(n3600), .B(n3568), .Z(n3571) );
  XOR U3533 ( .A(n3601), .B(n3602), .Z(n3568) );
  AND U3534 ( .A(n3603), .B(n3604), .Z(n3602) );
  XOR U3535 ( .A(n3601), .B(n3605), .Z(n3603) );
  XNOR U3536 ( .A(n3606), .B(n3607), .Z(n3600) );
  NOR U3537 ( .A(n3608), .B(n3609), .Z(n3607) );
  XOR U3538 ( .A(n3606), .B(n3610), .Z(n3608) );
  XNOR U3539 ( .A(n3567), .B(n3574), .Z(n3588) );
  NOR U3540 ( .A(n3531), .B(n3611), .Z(n3574) );
  XOR U3541 ( .A(n3579), .B(n3578), .Z(n3567) );
  XNOR U3542 ( .A(n3612), .B(n3575), .Z(n3578) );
  XOR U3543 ( .A(n3613), .B(n3614), .Z(n3575) );
  AND U3544 ( .A(n3615), .B(n3616), .Z(n3614) );
  XOR U3545 ( .A(n3613), .B(n3617), .Z(n3615) );
  XNOR U3546 ( .A(n3618), .B(n3619), .Z(n3612) );
  NOR U3547 ( .A(n3620), .B(n3621), .Z(n3619) );
  XNOR U3548 ( .A(n3618), .B(n3622), .Z(n3620) );
  XOR U3549 ( .A(n3623), .B(n3624), .Z(n3579) );
  NOR U3550 ( .A(n3625), .B(n3626), .Z(n3624) );
  XNOR U3551 ( .A(n3623), .B(n3627), .Z(n3625) );
  XNOR U3552 ( .A(n3516), .B(n3584), .Z(n3586) );
  XOR U3553 ( .A(n3628), .B(n3629), .Z(n3516) );
  AND U3554 ( .A(n23), .B(n3630), .Z(n3629) );
  XOR U3555 ( .A(n3631), .B(n3628), .Z(n3630) );
  AND U3556 ( .A(n3528), .B(n3531), .Z(n3584) );
  XOR U3557 ( .A(n3632), .B(n3611), .Z(n3531) );
  XNOR U3558 ( .A(p_input[1024]), .B(p_input[64]), .Z(n3611) );
  XOR U3559 ( .A(n3599), .B(n3598), .Z(n3632) );
  XNOR U3560 ( .A(n3633), .B(n3605), .Z(n3598) );
  XNOR U3561 ( .A(n3594), .B(n3593), .Z(n3605) );
  XOR U3562 ( .A(n3634), .B(n3590), .Z(n3593) );
  XOR U3563 ( .A(p_input[1034]), .B(p_input[74]), .Z(n3590) );
  XNOR U3564 ( .A(p_input[1035]), .B(p_input[75]), .Z(n3634) );
  XOR U3565 ( .A(p_input[1036]), .B(p_input[76]), .Z(n3594) );
  XNOR U3566 ( .A(n3604), .B(n3595), .Z(n3633) );
  XNOR U3567 ( .A(n3298), .B(p_input[65]), .Z(n3595) );
  XOR U3568 ( .A(n3635), .B(n3610), .Z(n3604) );
  XNOR U3569 ( .A(p_input[1039]), .B(p_input[79]), .Z(n3610) );
  XOR U3570 ( .A(n3601), .B(n3609), .Z(n3635) );
  XOR U3571 ( .A(n3636), .B(n3606), .Z(n3609) );
  XOR U3572 ( .A(p_input[1037]), .B(p_input[77]), .Z(n3606) );
  XNOR U3573 ( .A(p_input[1038]), .B(p_input[78]), .Z(n3636) );
  XOR U3574 ( .A(p_input[1033]), .B(p_input[73]), .Z(n3601) );
  XNOR U3575 ( .A(n3617), .B(n3616), .Z(n3599) );
  XNOR U3576 ( .A(n3637), .B(n3622), .Z(n3616) );
  XOR U3577 ( .A(p_input[1032]), .B(p_input[72]), .Z(n3622) );
  XOR U3578 ( .A(n3613), .B(n3621), .Z(n3637) );
  XOR U3579 ( .A(n3638), .B(n3618), .Z(n3621) );
  XOR U3580 ( .A(p_input[1030]), .B(p_input[70]), .Z(n3618) );
  XNOR U3581 ( .A(p_input[1031]), .B(p_input[71]), .Z(n3638) );
  XOR U3582 ( .A(p_input[1026]), .B(p_input[66]), .Z(n3613) );
  XNOR U3583 ( .A(n3627), .B(n3626), .Z(n3617) );
  XOR U3584 ( .A(n3639), .B(n3623), .Z(n3626) );
  XOR U3585 ( .A(p_input[1027]), .B(p_input[67]), .Z(n3623) );
  XNOR U3586 ( .A(p_input[1028]), .B(p_input[68]), .Z(n3639) );
  XOR U3587 ( .A(p_input[1029]), .B(p_input[69]), .Z(n3627) );
  XOR U3588 ( .A(n3640), .B(n3641), .Z(n3528) );
  AND U3589 ( .A(n23), .B(n3642), .Z(n3641) );
  XNOR U3590 ( .A(n3643), .B(n3640), .Z(n3642) );
  XNOR U3591 ( .A(n3644), .B(n3645), .Z(n23) );
  AND U3592 ( .A(n3646), .B(n3647), .Z(n3645) );
  XOR U3593 ( .A(n3541), .B(n3644), .Z(n3647) );
  AND U3594 ( .A(n3648), .B(n3649), .Z(n3541) );
  XNOR U3595 ( .A(n3538), .B(n3644), .Z(n3646) );
  XOR U3596 ( .A(n3650), .B(n3651), .Z(n3538) );
  AND U3597 ( .A(n27), .B(n3652), .Z(n3651) );
  XOR U3598 ( .A(n3653), .B(n3650), .Z(n3652) );
  XOR U3599 ( .A(n3654), .B(n3655), .Z(n3644) );
  AND U3600 ( .A(n3656), .B(n3657), .Z(n3655) );
  XNOR U3601 ( .A(n3654), .B(n3648), .Z(n3657) );
  IV U3602 ( .A(n3556), .Z(n3648) );
  XOR U3603 ( .A(n3658), .B(n3659), .Z(n3556) );
  XOR U3604 ( .A(n3660), .B(n3649), .Z(n3659) );
  AND U3605 ( .A(n3583), .B(n3661), .Z(n3649) );
  AND U3606 ( .A(n3662), .B(n3663), .Z(n3660) );
  XOR U3607 ( .A(n3664), .B(n3658), .Z(n3662) );
  XNOR U3608 ( .A(n3553), .B(n3654), .Z(n3656) );
  XOR U3609 ( .A(n3665), .B(n3666), .Z(n3553) );
  AND U3610 ( .A(n27), .B(n3667), .Z(n3666) );
  XOR U3611 ( .A(n3668), .B(n3665), .Z(n3667) );
  XOR U3612 ( .A(n3669), .B(n3670), .Z(n3654) );
  AND U3613 ( .A(n3671), .B(n3672), .Z(n3670) );
  XNOR U3614 ( .A(n3669), .B(n3583), .Z(n3672) );
  XOR U3615 ( .A(n3673), .B(n3663), .Z(n3583) );
  XNOR U3616 ( .A(n3674), .B(n3658), .Z(n3663) );
  XOR U3617 ( .A(n3675), .B(n3676), .Z(n3658) );
  AND U3618 ( .A(n3677), .B(n3678), .Z(n3676) );
  XOR U3619 ( .A(n3679), .B(n3675), .Z(n3677) );
  XNOR U3620 ( .A(n3680), .B(n3681), .Z(n3674) );
  AND U3621 ( .A(n3682), .B(n3683), .Z(n3681) );
  XOR U3622 ( .A(n3680), .B(n3684), .Z(n3682) );
  XNOR U3623 ( .A(n3664), .B(n3661), .Z(n3673) );
  AND U3624 ( .A(n3685), .B(n3686), .Z(n3661) );
  XOR U3625 ( .A(n3687), .B(n3688), .Z(n3664) );
  AND U3626 ( .A(n3689), .B(n3690), .Z(n3688) );
  XOR U3627 ( .A(n3687), .B(n3691), .Z(n3689) );
  XNOR U3628 ( .A(n3580), .B(n3669), .Z(n3671) );
  XOR U3629 ( .A(n3692), .B(n3693), .Z(n3580) );
  AND U3630 ( .A(n27), .B(n3694), .Z(n3693) );
  XNOR U3631 ( .A(n3695), .B(n3692), .Z(n3694) );
  XOR U3632 ( .A(n3696), .B(n3697), .Z(n3669) );
  AND U3633 ( .A(n3698), .B(n3699), .Z(n3697) );
  XNOR U3634 ( .A(n3696), .B(n3685), .Z(n3699) );
  IV U3635 ( .A(n3631), .Z(n3685) );
  XNOR U3636 ( .A(n3700), .B(n3678), .Z(n3631) );
  XNOR U3637 ( .A(n3701), .B(n3684), .Z(n3678) );
  XOR U3638 ( .A(n3702), .B(n3703), .Z(n3684) );
  NOR U3639 ( .A(n3704), .B(n3705), .Z(n3703) );
  XNOR U3640 ( .A(n3702), .B(n3706), .Z(n3704) );
  XNOR U3641 ( .A(n3683), .B(n3675), .Z(n3701) );
  XOR U3642 ( .A(n3707), .B(n3708), .Z(n3675) );
  AND U3643 ( .A(n3709), .B(n3710), .Z(n3708) );
  XNOR U3644 ( .A(n3707), .B(n3711), .Z(n3709) );
  XNOR U3645 ( .A(n3712), .B(n3680), .Z(n3683) );
  XOR U3646 ( .A(n3713), .B(n3714), .Z(n3680) );
  AND U3647 ( .A(n3715), .B(n3716), .Z(n3714) );
  XOR U3648 ( .A(n3713), .B(n3717), .Z(n3715) );
  XNOR U3649 ( .A(n3718), .B(n3719), .Z(n3712) );
  NOR U3650 ( .A(n3720), .B(n3721), .Z(n3719) );
  XOR U3651 ( .A(n3718), .B(n3722), .Z(n3720) );
  XNOR U3652 ( .A(n3679), .B(n3686), .Z(n3700) );
  NOR U3653 ( .A(n3643), .B(n3723), .Z(n3686) );
  XOR U3654 ( .A(n3691), .B(n3690), .Z(n3679) );
  XNOR U3655 ( .A(n3724), .B(n3687), .Z(n3690) );
  XOR U3656 ( .A(n3725), .B(n3726), .Z(n3687) );
  AND U3657 ( .A(n3727), .B(n3728), .Z(n3726) );
  XOR U3658 ( .A(n3725), .B(n3729), .Z(n3727) );
  XNOR U3659 ( .A(n3730), .B(n3731), .Z(n3724) );
  NOR U3660 ( .A(n3732), .B(n3733), .Z(n3731) );
  XNOR U3661 ( .A(n3730), .B(n3734), .Z(n3732) );
  XOR U3662 ( .A(n3735), .B(n3736), .Z(n3691) );
  NOR U3663 ( .A(n3737), .B(n3738), .Z(n3736) );
  XNOR U3664 ( .A(n3735), .B(n3739), .Z(n3737) );
  XNOR U3665 ( .A(n3628), .B(n3696), .Z(n3698) );
  XOR U3666 ( .A(n3740), .B(n3741), .Z(n3628) );
  AND U3667 ( .A(n27), .B(n3742), .Z(n3741) );
  XOR U3668 ( .A(n3743), .B(n3740), .Z(n3742) );
  AND U3669 ( .A(n3640), .B(n3643), .Z(n3696) );
  XOR U3670 ( .A(n3744), .B(n3723), .Z(n3643) );
  XNOR U3671 ( .A(p_input[1024]), .B(p_input[80]), .Z(n3723) );
  XOR U3672 ( .A(n3711), .B(n3710), .Z(n3744) );
  XNOR U3673 ( .A(n3745), .B(n3717), .Z(n3710) );
  XNOR U3674 ( .A(n3706), .B(n3705), .Z(n3717) );
  XOR U3675 ( .A(n3746), .B(n3702), .Z(n3705) );
  XOR U3676 ( .A(p_input[1034]), .B(p_input[90]), .Z(n3702) );
  XNOR U3677 ( .A(p_input[1035]), .B(p_input[91]), .Z(n3746) );
  XOR U3678 ( .A(p_input[1036]), .B(p_input[92]), .Z(n3706) );
  XNOR U3679 ( .A(n3716), .B(n3707), .Z(n3745) );
  XNOR U3680 ( .A(n3298), .B(p_input[81]), .Z(n3707) );
  XOR U3681 ( .A(n3747), .B(n3722), .Z(n3716) );
  XNOR U3682 ( .A(p_input[1039]), .B(p_input[95]), .Z(n3722) );
  XOR U3683 ( .A(n3713), .B(n3721), .Z(n3747) );
  XOR U3684 ( .A(n3748), .B(n3718), .Z(n3721) );
  XOR U3685 ( .A(p_input[1037]), .B(p_input[93]), .Z(n3718) );
  XNOR U3686 ( .A(p_input[1038]), .B(p_input[94]), .Z(n3748) );
  XOR U3687 ( .A(p_input[1033]), .B(p_input[89]), .Z(n3713) );
  XNOR U3688 ( .A(n3729), .B(n3728), .Z(n3711) );
  XNOR U3689 ( .A(n3749), .B(n3734), .Z(n3728) );
  XOR U3690 ( .A(p_input[1032]), .B(p_input[88]), .Z(n3734) );
  XOR U3691 ( .A(n3725), .B(n3733), .Z(n3749) );
  XOR U3692 ( .A(n3750), .B(n3730), .Z(n3733) );
  XOR U3693 ( .A(p_input[1030]), .B(p_input[86]), .Z(n3730) );
  XNOR U3694 ( .A(p_input[1031]), .B(p_input[87]), .Z(n3750) );
  XOR U3695 ( .A(p_input[1026]), .B(p_input[82]), .Z(n3725) );
  XNOR U3696 ( .A(n3739), .B(n3738), .Z(n3729) );
  XOR U3697 ( .A(n3751), .B(n3735), .Z(n3738) );
  XOR U3698 ( .A(p_input[1027]), .B(p_input[83]), .Z(n3735) );
  XNOR U3699 ( .A(p_input[1028]), .B(p_input[84]), .Z(n3751) );
  XOR U3700 ( .A(p_input[1029]), .B(p_input[85]), .Z(n3739) );
  XOR U3701 ( .A(n3752), .B(n3753), .Z(n3640) );
  AND U3702 ( .A(n27), .B(n3754), .Z(n3753) );
  XNOR U3703 ( .A(n3755), .B(n3752), .Z(n3754) );
  XNOR U3704 ( .A(n3756), .B(n3757), .Z(n27) );
  AND U3705 ( .A(n3758), .B(n3759), .Z(n3757) );
  XOR U3706 ( .A(n3653), .B(n3756), .Z(n3759) );
  AND U3707 ( .A(n3760), .B(n3761), .Z(n3653) );
  XNOR U3708 ( .A(n3650), .B(n3756), .Z(n3758) );
  XOR U3709 ( .A(n3762), .B(n3763), .Z(n3650) );
  AND U3710 ( .A(n31), .B(n3764), .Z(n3763) );
  XOR U3711 ( .A(n3765), .B(n3762), .Z(n3764) );
  XOR U3712 ( .A(n3766), .B(n3767), .Z(n3756) );
  AND U3713 ( .A(n3768), .B(n3769), .Z(n3767) );
  XNOR U3714 ( .A(n3766), .B(n3760), .Z(n3769) );
  IV U3715 ( .A(n3668), .Z(n3760) );
  XOR U3716 ( .A(n3770), .B(n3771), .Z(n3668) );
  XOR U3717 ( .A(n3772), .B(n3761), .Z(n3771) );
  AND U3718 ( .A(n3695), .B(n3773), .Z(n3761) );
  AND U3719 ( .A(n3774), .B(n3775), .Z(n3772) );
  XOR U3720 ( .A(n3776), .B(n3770), .Z(n3774) );
  XNOR U3721 ( .A(n3665), .B(n3766), .Z(n3768) );
  XOR U3722 ( .A(n3777), .B(n3778), .Z(n3665) );
  AND U3723 ( .A(n31), .B(n3779), .Z(n3778) );
  XOR U3724 ( .A(n3780), .B(n3777), .Z(n3779) );
  XOR U3725 ( .A(n3781), .B(n3782), .Z(n3766) );
  AND U3726 ( .A(n3783), .B(n3784), .Z(n3782) );
  XNOR U3727 ( .A(n3781), .B(n3695), .Z(n3784) );
  XOR U3728 ( .A(n3785), .B(n3775), .Z(n3695) );
  XNOR U3729 ( .A(n3786), .B(n3770), .Z(n3775) );
  XOR U3730 ( .A(n3787), .B(n3788), .Z(n3770) );
  AND U3731 ( .A(n3789), .B(n3790), .Z(n3788) );
  XOR U3732 ( .A(n3791), .B(n3787), .Z(n3789) );
  XNOR U3733 ( .A(n3792), .B(n3793), .Z(n3786) );
  AND U3734 ( .A(n3794), .B(n3795), .Z(n3793) );
  XOR U3735 ( .A(n3792), .B(n3796), .Z(n3794) );
  XNOR U3736 ( .A(n3776), .B(n3773), .Z(n3785) );
  AND U3737 ( .A(n3797), .B(n3798), .Z(n3773) );
  XOR U3738 ( .A(n3799), .B(n3800), .Z(n3776) );
  AND U3739 ( .A(n3801), .B(n3802), .Z(n3800) );
  XOR U3740 ( .A(n3799), .B(n3803), .Z(n3801) );
  XNOR U3741 ( .A(n3692), .B(n3781), .Z(n3783) );
  XOR U3742 ( .A(n3804), .B(n3805), .Z(n3692) );
  AND U3743 ( .A(n31), .B(n3806), .Z(n3805) );
  XNOR U3744 ( .A(n3807), .B(n3804), .Z(n3806) );
  XOR U3745 ( .A(n3808), .B(n3809), .Z(n3781) );
  AND U3746 ( .A(n3810), .B(n3811), .Z(n3809) );
  XNOR U3747 ( .A(n3808), .B(n3797), .Z(n3811) );
  IV U3748 ( .A(n3743), .Z(n3797) );
  XNOR U3749 ( .A(n3812), .B(n3790), .Z(n3743) );
  XNOR U3750 ( .A(n3813), .B(n3796), .Z(n3790) );
  XOR U3751 ( .A(n3814), .B(n3815), .Z(n3796) );
  NOR U3752 ( .A(n3816), .B(n3817), .Z(n3815) );
  XNOR U3753 ( .A(n3814), .B(n3818), .Z(n3816) );
  XNOR U3754 ( .A(n3795), .B(n3787), .Z(n3813) );
  XOR U3755 ( .A(n3819), .B(n3820), .Z(n3787) );
  AND U3756 ( .A(n3821), .B(n3822), .Z(n3820) );
  XNOR U3757 ( .A(n3819), .B(n3823), .Z(n3821) );
  XNOR U3758 ( .A(n3824), .B(n3792), .Z(n3795) );
  XOR U3759 ( .A(n3825), .B(n3826), .Z(n3792) );
  AND U3760 ( .A(n3827), .B(n3828), .Z(n3826) );
  XOR U3761 ( .A(n3825), .B(n3829), .Z(n3827) );
  XNOR U3762 ( .A(n3830), .B(n3831), .Z(n3824) );
  NOR U3763 ( .A(n3832), .B(n3833), .Z(n3831) );
  XOR U3764 ( .A(n3830), .B(n3834), .Z(n3832) );
  XNOR U3765 ( .A(n3791), .B(n3798), .Z(n3812) );
  NOR U3766 ( .A(n3755), .B(n3835), .Z(n3798) );
  XOR U3767 ( .A(n3803), .B(n3802), .Z(n3791) );
  XNOR U3768 ( .A(n3836), .B(n3799), .Z(n3802) );
  XOR U3769 ( .A(n3837), .B(n3838), .Z(n3799) );
  AND U3770 ( .A(n3839), .B(n3840), .Z(n3838) );
  XOR U3771 ( .A(n3837), .B(n3841), .Z(n3839) );
  XNOR U3772 ( .A(n3842), .B(n3843), .Z(n3836) );
  NOR U3773 ( .A(n3844), .B(n3845), .Z(n3843) );
  XNOR U3774 ( .A(n3842), .B(n3846), .Z(n3844) );
  XOR U3775 ( .A(n3847), .B(n3848), .Z(n3803) );
  NOR U3776 ( .A(n3849), .B(n3850), .Z(n3848) );
  XNOR U3777 ( .A(n3847), .B(n3851), .Z(n3849) );
  XNOR U3778 ( .A(n3740), .B(n3808), .Z(n3810) );
  XOR U3779 ( .A(n3852), .B(n3853), .Z(n3740) );
  AND U3780 ( .A(n31), .B(n3854), .Z(n3853) );
  XOR U3781 ( .A(n3855), .B(n3852), .Z(n3854) );
  AND U3782 ( .A(n3752), .B(n3755), .Z(n3808) );
  XOR U3783 ( .A(n3856), .B(n3835), .Z(n3755) );
  XNOR U3784 ( .A(p_input[1024]), .B(p_input[96]), .Z(n3835) );
  XOR U3785 ( .A(n3823), .B(n3822), .Z(n3856) );
  XNOR U3786 ( .A(n3857), .B(n3829), .Z(n3822) );
  XNOR U3787 ( .A(n3818), .B(n3817), .Z(n3829) );
  XOR U3788 ( .A(n3858), .B(n3814), .Z(n3817) );
  XOR U3789 ( .A(p_input[1034]), .B(p_input[106]), .Z(n3814) );
  XNOR U3790 ( .A(p_input[1035]), .B(p_input[107]), .Z(n3858) );
  XOR U3791 ( .A(p_input[1036]), .B(p_input[108]), .Z(n3818) );
  XNOR U3792 ( .A(n3828), .B(n3819), .Z(n3857) );
  XNOR U3793 ( .A(n3298), .B(p_input[97]), .Z(n3819) );
  XOR U3794 ( .A(n3859), .B(n3834), .Z(n3828) );
  XNOR U3795 ( .A(p_input[1039]), .B(p_input[111]), .Z(n3834) );
  XOR U3796 ( .A(n3825), .B(n3833), .Z(n3859) );
  XOR U3797 ( .A(n3860), .B(n3830), .Z(n3833) );
  XOR U3798 ( .A(p_input[1037]), .B(p_input[109]), .Z(n3830) );
  XNOR U3799 ( .A(p_input[1038]), .B(p_input[110]), .Z(n3860) );
  XOR U3800 ( .A(p_input[1033]), .B(p_input[105]), .Z(n3825) );
  XNOR U3801 ( .A(n3841), .B(n3840), .Z(n3823) );
  XNOR U3802 ( .A(n3861), .B(n3846), .Z(n3840) );
  XOR U3803 ( .A(p_input[1032]), .B(p_input[104]), .Z(n3846) );
  XOR U3804 ( .A(n3837), .B(n3845), .Z(n3861) );
  XOR U3805 ( .A(n3862), .B(n3842), .Z(n3845) );
  XOR U3806 ( .A(p_input[102]), .B(p_input[1030]), .Z(n3842) );
  XNOR U3807 ( .A(p_input[1031]), .B(p_input[103]), .Z(n3862) );
  XOR U3808 ( .A(p_input[1026]), .B(p_input[98]), .Z(n3837) );
  XNOR U3809 ( .A(n3851), .B(n3850), .Z(n3841) );
  XOR U3810 ( .A(n3863), .B(n3847), .Z(n3850) );
  XOR U3811 ( .A(p_input[1027]), .B(p_input[99]), .Z(n3847) );
  XOR U3812 ( .A(p_input[100]), .B(n3864), .Z(n3863) );
  XOR U3813 ( .A(p_input[101]), .B(p_input[1029]), .Z(n3851) );
  XOR U3814 ( .A(n3865), .B(n3866), .Z(n3752) );
  AND U3815 ( .A(n31), .B(n3867), .Z(n3866) );
  XNOR U3816 ( .A(n3868), .B(n3865), .Z(n3867) );
  XNOR U3817 ( .A(n3869), .B(n3870), .Z(n31) );
  AND U3818 ( .A(n3871), .B(n3872), .Z(n3870) );
  XOR U3819 ( .A(n3765), .B(n3869), .Z(n3872) );
  AND U3820 ( .A(n3873), .B(n3874), .Z(n3765) );
  XNOR U3821 ( .A(n3762), .B(n3869), .Z(n3871) );
  XOR U3822 ( .A(n3875), .B(n3876), .Z(n3762) );
  AND U3823 ( .A(n35), .B(n3877), .Z(n3876) );
  XOR U3824 ( .A(n3878), .B(n3875), .Z(n3877) );
  XOR U3825 ( .A(n3879), .B(n3880), .Z(n3869) );
  AND U3826 ( .A(n3881), .B(n3882), .Z(n3880) );
  XNOR U3827 ( .A(n3879), .B(n3873), .Z(n3882) );
  IV U3828 ( .A(n3780), .Z(n3873) );
  XOR U3829 ( .A(n3883), .B(n3884), .Z(n3780) );
  XOR U3830 ( .A(n3885), .B(n3874), .Z(n3884) );
  AND U3831 ( .A(n3807), .B(n3886), .Z(n3874) );
  AND U3832 ( .A(n3887), .B(n3888), .Z(n3885) );
  XOR U3833 ( .A(n3889), .B(n3883), .Z(n3887) );
  XNOR U3834 ( .A(n3777), .B(n3879), .Z(n3881) );
  XOR U3835 ( .A(n3890), .B(n3891), .Z(n3777) );
  AND U3836 ( .A(n35), .B(n3892), .Z(n3891) );
  XOR U3837 ( .A(n3893), .B(n3890), .Z(n3892) );
  XOR U3838 ( .A(n3894), .B(n3895), .Z(n3879) );
  AND U3839 ( .A(n3896), .B(n3897), .Z(n3895) );
  XNOR U3840 ( .A(n3894), .B(n3807), .Z(n3897) );
  XOR U3841 ( .A(n3898), .B(n3888), .Z(n3807) );
  XNOR U3842 ( .A(n3899), .B(n3883), .Z(n3888) );
  XOR U3843 ( .A(n3900), .B(n3901), .Z(n3883) );
  AND U3844 ( .A(n3902), .B(n3903), .Z(n3901) );
  XOR U3845 ( .A(n3904), .B(n3900), .Z(n3902) );
  XNOR U3846 ( .A(n3905), .B(n3906), .Z(n3899) );
  AND U3847 ( .A(n3907), .B(n3908), .Z(n3906) );
  XOR U3848 ( .A(n3905), .B(n3909), .Z(n3907) );
  XNOR U3849 ( .A(n3889), .B(n3886), .Z(n3898) );
  AND U3850 ( .A(n3910), .B(n3911), .Z(n3886) );
  XOR U3851 ( .A(n3912), .B(n3913), .Z(n3889) );
  AND U3852 ( .A(n3914), .B(n3915), .Z(n3913) );
  XOR U3853 ( .A(n3912), .B(n3916), .Z(n3914) );
  XNOR U3854 ( .A(n3804), .B(n3894), .Z(n3896) );
  XOR U3855 ( .A(n3917), .B(n3918), .Z(n3804) );
  AND U3856 ( .A(n35), .B(n3919), .Z(n3918) );
  XNOR U3857 ( .A(n3920), .B(n3917), .Z(n3919) );
  XOR U3858 ( .A(n3921), .B(n3922), .Z(n3894) );
  AND U3859 ( .A(n3923), .B(n3924), .Z(n3922) );
  XNOR U3860 ( .A(n3921), .B(n3910), .Z(n3924) );
  IV U3861 ( .A(n3855), .Z(n3910) );
  XNOR U3862 ( .A(n3925), .B(n3903), .Z(n3855) );
  XNOR U3863 ( .A(n3926), .B(n3909), .Z(n3903) );
  XOR U3864 ( .A(n3927), .B(n3928), .Z(n3909) );
  NOR U3865 ( .A(n3929), .B(n3930), .Z(n3928) );
  XNOR U3866 ( .A(n3927), .B(n3931), .Z(n3929) );
  XNOR U3867 ( .A(n3908), .B(n3900), .Z(n3926) );
  XOR U3868 ( .A(n3932), .B(n3933), .Z(n3900) );
  AND U3869 ( .A(n3934), .B(n3935), .Z(n3933) );
  XNOR U3870 ( .A(n3932), .B(n3936), .Z(n3934) );
  XNOR U3871 ( .A(n3937), .B(n3905), .Z(n3908) );
  XOR U3872 ( .A(n3938), .B(n3939), .Z(n3905) );
  AND U3873 ( .A(n3940), .B(n3941), .Z(n3939) );
  XOR U3874 ( .A(n3938), .B(n3942), .Z(n3940) );
  XNOR U3875 ( .A(n3943), .B(n3944), .Z(n3937) );
  NOR U3876 ( .A(n3945), .B(n3946), .Z(n3944) );
  XOR U3877 ( .A(n3943), .B(n3947), .Z(n3945) );
  XNOR U3878 ( .A(n3904), .B(n3911), .Z(n3925) );
  NOR U3879 ( .A(n3868), .B(n3948), .Z(n3911) );
  XOR U3880 ( .A(n3916), .B(n3915), .Z(n3904) );
  XNOR U3881 ( .A(n3949), .B(n3912), .Z(n3915) );
  XOR U3882 ( .A(n3950), .B(n3951), .Z(n3912) );
  AND U3883 ( .A(n3952), .B(n3953), .Z(n3951) );
  XOR U3884 ( .A(n3950), .B(n3954), .Z(n3952) );
  XNOR U3885 ( .A(n3955), .B(n3956), .Z(n3949) );
  NOR U3886 ( .A(n3957), .B(n3958), .Z(n3956) );
  XNOR U3887 ( .A(n3955), .B(n3959), .Z(n3957) );
  XOR U3888 ( .A(n3960), .B(n3961), .Z(n3916) );
  NOR U3889 ( .A(n3962), .B(n3963), .Z(n3961) );
  XNOR U3890 ( .A(n3960), .B(n3964), .Z(n3962) );
  XNOR U3891 ( .A(n3852), .B(n3921), .Z(n3923) );
  XOR U3892 ( .A(n3965), .B(n3966), .Z(n3852) );
  AND U3893 ( .A(n35), .B(n3967), .Z(n3966) );
  XOR U3894 ( .A(n3968), .B(n3965), .Z(n3967) );
  AND U3895 ( .A(n3865), .B(n3868), .Z(n3921) );
  XOR U3896 ( .A(n3969), .B(n3948), .Z(n3868) );
  XNOR U3897 ( .A(p_input[1024]), .B(p_input[112]), .Z(n3948) );
  XOR U3898 ( .A(n3936), .B(n3935), .Z(n3969) );
  XNOR U3899 ( .A(n3970), .B(n3942), .Z(n3935) );
  XNOR U3900 ( .A(n3931), .B(n3930), .Z(n3942) );
  XOR U3901 ( .A(n3971), .B(n3927), .Z(n3930) );
  XOR U3902 ( .A(p_input[1034]), .B(p_input[122]), .Z(n3927) );
  XNOR U3903 ( .A(p_input[1035]), .B(p_input[123]), .Z(n3971) );
  XOR U3904 ( .A(p_input[1036]), .B(p_input[124]), .Z(n3931) );
  XNOR U3905 ( .A(n3941), .B(n3932), .Z(n3970) );
  XNOR U3906 ( .A(n3298), .B(p_input[113]), .Z(n3932) );
  XOR U3907 ( .A(n3972), .B(n3947), .Z(n3941) );
  XNOR U3908 ( .A(p_input[1039]), .B(p_input[127]), .Z(n3947) );
  XOR U3909 ( .A(n3938), .B(n3946), .Z(n3972) );
  XOR U3910 ( .A(n3973), .B(n3943), .Z(n3946) );
  XOR U3911 ( .A(p_input[1037]), .B(p_input[125]), .Z(n3943) );
  XNOR U3912 ( .A(p_input[1038]), .B(p_input[126]), .Z(n3973) );
  XOR U3913 ( .A(p_input[1033]), .B(p_input[121]), .Z(n3938) );
  XNOR U3914 ( .A(n3954), .B(n3953), .Z(n3936) );
  XNOR U3915 ( .A(n3974), .B(n3959), .Z(n3953) );
  XOR U3916 ( .A(p_input[1032]), .B(p_input[120]), .Z(n3959) );
  XOR U3917 ( .A(n3950), .B(n3958), .Z(n3974) );
  XOR U3918 ( .A(n3975), .B(n3955), .Z(n3958) );
  XOR U3919 ( .A(p_input[1030]), .B(p_input[118]), .Z(n3955) );
  XNOR U3920 ( .A(p_input[1031]), .B(p_input[119]), .Z(n3975) );
  XOR U3921 ( .A(p_input[1026]), .B(p_input[114]), .Z(n3950) );
  XNOR U3922 ( .A(n3964), .B(n3963), .Z(n3954) );
  XOR U3923 ( .A(n3976), .B(n3960), .Z(n3963) );
  XOR U3924 ( .A(p_input[1027]), .B(p_input[115]), .Z(n3960) );
  XNOR U3925 ( .A(p_input[1028]), .B(p_input[116]), .Z(n3976) );
  XOR U3926 ( .A(p_input[1029]), .B(p_input[117]), .Z(n3964) );
  XOR U3927 ( .A(n3977), .B(n3978), .Z(n3865) );
  AND U3928 ( .A(n35), .B(n3979), .Z(n3978) );
  XNOR U3929 ( .A(n3980), .B(n3977), .Z(n3979) );
  XNOR U3930 ( .A(n3981), .B(n3982), .Z(n35) );
  AND U3931 ( .A(n3983), .B(n3984), .Z(n3982) );
  XOR U3932 ( .A(n3878), .B(n3981), .Z(n3984) );
  AND U3933 ( .A(n3985), .B(n3986), .Z(n3878) );
  XNOR U3934 ( .A(n3875), .B(n3981), .Z(n3983) );
  XOR U3935 ( .A(n3987), .B(n3988), .Z(n3875) );
  AND U3936 ( .A(n39), .B(n3989), .Z(n3988) );
  XOR U3937 ( .A(n3990), .B(n3987), .Z(n3989) );
  XOR U3938 ( .A(n3991), .B(n3992), .Z(n3981) );
  AND U3939 ( .A(n3993), .B(n3994), .Z(n3992) );
  XNOR U3940 ( .A(n3991), .B(n3985), .Z(n3994) );
  IV U3941 ( .A(n3893), .Z(n3985) );
  XOR U3942 ( .A(n3995), .B(n3996), .Z(n3893) );
  XOR U3943 ( .A(n3997), .B(n3986), .Z(n3996) );
  AND U3944 ( .A(n3920), .B(n3998), .Z(n3986) );
  AND U3945 ( .A(n3999), .B(n4000), .Z(n3997) );
  XOR U3946 ( .A(n4001), .B(n3995), .Z(n3999) );
  XNOR U3947 ( .A(n3890), .B(n3991), .Z(n3993) );
  XOR U3948 ( .A(n4002), .B(n4003), .Z(n3890) );
  AND U3949 ( .A(n39), .B(n4004), .Z(n4003) );
  XOR U3950 ( .A(n4005), .B(n4002), .Z(n4004) );
  XOR U3951 ( .A(n4006), .B(n4007), .Z(n3991) );
  AND U3952 ( .A(n4008), .B(n4009), .Z(n4007) );
  XNOR U3953 ( .A(n4006), .B(n3920), .Z(n4009) );
  XOR U3954 ( .A(n4010), .B(n4000), .Z(n3920) );
  XNOR U3955 ( .A(n4011), .B(n3995), .Z(n4000) );
  XOR U3956 ( .A(n4012), .B(n4013), .Z(n3995) );
  AND U3957 ( .A(n4014), .B(n4015), .Z(n4013) );
  XOR U3958 ( .A(n4016), .B(n4012), .Z(n4014) );
  XNOR U3959 ( .A(n4017), .B(n4018), .Z(n4011) );
  AND U3960 ( .A(n4019), .B(n4020), .Z(n4018) );
  XOR U3961 ( .A(n4017), .B(n4021), .Z(n4019) );
  XNOR U3962 ( .A(n4001), .B(n3998), .Z(n4010) );
  AND U3963 ( .A(n4022), .B(n4023), .Z(n3998) );
  XOR U3964 ( .A(n4024), .B(n4025), .Z(n4001) );
  AND U3965 ( .A(n4026), .B(n4027), .Z(n4025) );
  XOR U3966 ( .A(n4024), .B(n4028), .Z(n4026) );
  XNOR U3967 ( .A(n3917), .B(n4006), .Z(n4008) );
  XOR U3968 ( .A(n4029), .B(n4030), .Z(n3917) );
  AND U3969 ( .A(n39), .B(n4031), .Z(n4030) );
  XNOR U3970 ( .A(n4032), .B(n4029), .Z(n4031) );
  XOR U3971 ( .A(n4033), .B(n4034), .Z(n4006) );
  AND U3972 ( .A(n4035), .B(n4036), .Z(n4034) );
  XNOR U3973 ( .A(n4033), .B(n4022), .Z(n4036) );
  IV U3974 ( .A(n3968), .Z(n4022) );
  XNOR U3975 ( .A(n4037), .B(n4015), .Z(n3968) );
  XNOR U3976 ( .A(n4038), .B(n4021), .Z(n4015) );
  XOR U3977 ( .A(n4039), .B(n4040), .Z(n4021) );
  NOR U3978 ( .A(n4041), .B(n4042), .Z(n4040) );
  XNOR U3979 ( .A(n4039), .B(n4043), .Z(n4041) );
  XNOR U3980 ( .A(n4020), .B(n4012), .Z(n4038) );
  XOR U3981 ( .A(n4044), .B(n4045), .Z(n4012) );
  AND U3982 ( .A(n4046), .B(n4047), .Z(n4045) );
  XNOR U3983 ( .A(n4044), .B(n4048), .Z(n4046) );
  XNOR U3984 ( .A(n4049), .B(n4017), .Z(n4020) );
  XOR U3985 ( .A(n4050), .B(n4051), .Z(n4017) );
  AND U3986 ( .A(n4052), .B(n4053), .Z(n4051) );
  XOR U3987 ( .A(n4050), .B(n4054), .Z(n4052) );
  XNOR U3988 ( .A(n4055), .B(n4056), .Z(n4049) );
  NOR U3989 ( .A(n4057), .B(n4058), .Z(n4056) );
  XOR U3990 ( .A(n4055), .B(n4059), .Z(n4057) );
  XNOR U3991 ( .A(n4016), .B(n4023), .Z(n4037) );
  NOR U3992 ( .A(n3980), .B(n4060), .Z(n4023) );
  XOR U3993 ( .A(n4028), .B(n4027), .Z(n4016) );
  XNOR U3994 ( .A(n4061), .B(n4024), .Z(n4027) );
  XOR U3995 ( .A(n4062), .B(n4063), .Z(n4024) );
  AND U3996 ( .A(n4064), .B(n4065), .Z(n4063) );
  XOR U3997 ( .A(n4062), .B(n4066), .Z(n4064) );
  XNOR U3998 ( .A(n4067), .B(n4068), .Z(n4061) );
  NOR U3999 ( .A(n4069), .B(n4070), .Z(n4068) );
  XNOR U4000 ( .A(n4067), .B(n4071), .Z(n4069) );
  XOR U4001 ( .A(n4072), .B(n4073), .Z(n4028) );
  NOR U4002 ( .A(n4074), .B(n4075), .Z(n4073) );
  XNOR U4003 ( .A(n4072), .B(n4076), .Z(n4074) );
  XNOR U4004 ( .A(n3965), .B(n4033), .Z(n4035) );
  XOR U4005 ( .A(n4077), .B(n4078), .Z(n3965) );
  AND U4006 ( .A(n39), .B(n4079), .Z(n4078) );
  XOR U4007 ( .A(n4080), .B(n4077), .Z(n4079) );
  AND U4008 ( .A(n3977), .B(n3980), .Z(n4033) );
  XOR U4009 ( .A(n4081), .B(n4060), .Z(n3980) );
  XNOR U4010 ( .A(p_input[1024]), .B(p_input[128]), .Z(n4060) );
  XOR U4011 ( .A(n4048), .B(n4047), .Z(n4081) );
  XNOR U4012 ( .A(n4082), .B(n4054), .Z(n4047) );
  XNOR U4013 ( .A(n4043), .B(n4042), .Z(n4054) );
  XOR U4014 ( .A(n4083), .B(n4039), .Z(n4042) );
  XOR U4015 ( .A(p_input[1034]), .B(p_input[138]), .Z(n4039) );
  XNOR U4016 ( .A(p_input[1035]), .B(p_input[139]), .Z(n4083) );
  XOR U4017 ( .A(p_input[1036]), .B(p_input[140]), .Z(n4043) );
  XNOR U4018 ( .A(n4053), .B(n4044), .Z(n4082) );
  XNOR U4019 ( .A(n3298), .B(p_input[129]), .Z(n4044) );
  XOR U4020 ( .A(n4084), .B(n4059), .Z(n4053) );
  XNOR U4021 ( .A(p_input[1039]), .B(p_input[143]), .Z(n4059) );
  XOR U4022 ( .A(n4050), .B(n4058), .Z(n4084) );
  XOR U4023 ( .A(n4085), .B(n4055), .Z(n4058) );
  XOR U4024 ( .A(p_input[1037]), .B(p_input[141]), .Z(n4055) );
  XNOR U4025 ( .A(p_input[1038]), .B(p_input[142]), .Z(n4085) );
  XOR U4026 ( .A(p_input[1033]), .B(p_input[137]), .Z(n4050) );
  XNOR U4027 ( .A(n4066), .B(n4065), .Z(n4048) );
  XNOR U4028 ( .A(n4086), .B(n4071), .Z(n4065) );
  XOR U4029 ( .A(p_input[1032]), .B(p_input[136]), .Z(n4071) );
  XOR U4030 ( .A(n4062), .B(n4070), .Z(n4086) );
  XOR U4031 ( .A(n4087), .B(n4067), .Z(n4070) );
  XOR U4032 ( .A(p_input[1030]), .B(p_input[134]), .Z(n4067) );
  XNOR U4033 ( .A(p_input[1031]), .B(p_input[135]), .Z(n4087) );
  XOR U4034 ( .A(p_input[1026]), .B(p_input[130]), .Z(n4062) );
  XNOR U4035 ( .A(n4076), .B(n4075), .Z(n4066) );
  XOR U4036 ( .A(n4088), .B(n4072), .Z(n4075) );
  XOR U4037 ( .A(p_input[1027]), .B(p_input[131]), .Z(n4072) );
  XNOR U4038 ( .A(p_input[1028]), .B(p_input[132]), .Z(n4088) );
  XOR U4039 ( .A(p_input[1029]), .B(p_input[133]), .Z(n4076) );
  XOR U4040 ( .A(n4089), .B(n4090), .Z(n3977) );
  AND U4041 ( .A(n39), .B(n4091), .Z(n4090) );
  XNOR U4042 ( .A(n4092), .B(n4089), .Z(n4091) );
  XNOR U4043 ( .A(n4093), .B(n4094), .Z(n39) );
  AND U4044 ( .A(n4095), .B(n4096), .Z(n4094) );
  XOR U4045 ( .A(n3990), .B(n4093), .Z(n4096) );
  AND U4046 ( .A(n4097), .B(n4098), .Z(n3990) );
  XNOR U4047 ( .A(n3987), .B(n4093), .Z(n4095) );
  XOR U4048 ( .A(n4099), .B(n4100), .Z(n3987) );
  AND U4049 ( .A(n43), .B(n4101), .Z(n4100) );
  XOR U4050 ( .A(n4102), .B(n4099), .Z(n4101) );
  XOR U4051 ( .A(n4103), .B(n4104), .Z(n4093) );
  AND U4052 ( .A(n4105), .B(n4106), .Z(n4104) );
  XNOR U4053 ( .A(n4103), .B(n4097), .Z(n4106) );
  IV U4054 ( .A(n4005), .Z(n4097) );
  XOR U4055 ( .A(n4107), .B(n4108), .Z(n4005) );
  XOR U4056 ( .A(n4109), .B(n4098), .Z(n4108) );
  AND U4057 ( .A(n4032), .B(n4110), .Z(n4098) );
  AND U4058 ( .A(n4111), .B(n4112), .Z(n4109) );
  XOR U4059 ( .A(n4113), .B(n4107), .Z(n4111) );
  XNOR U4060 ( .A(n4002), .B(n4103), .Z(n4105) );
  XOR U4061 ( .A(n4114), .B(n4115), .Z(n4002) );
  AND U4062 ( .A(n43), .B(n4116), .Z(n4115) );
  XOR U4063 ( .A(n4117), .B(n4114), .Z(n4116) );
  XOR U4064 ( .A(n4118), .B(n4119), .Z(n4103) );
  AND U4065 ( .A(n4120), .B(n4121), .Z(n4119) );
  XNOR U4066 ( .A(n4118), .B(n4032), .Z(n4121) );
  XOR U4067 ( .A(n4122), .B(n4112), .Z(n4032) );
  XNOR U4068 ( .A(n4123), .B(n4107), .Z(n4112) );
  XOR U4069 ( .A(n4124), .B(n4125), .Z(n4107) );
  AND U4070 ( .A(n4126), .B(n4127), .Z(n4125) );
  XOR U4071 ( .A(n4128), .B(n4124), .Z(n4126) );
  XNOR U4072 ( .A(n4129), .B(n4130), .Z(n4123) );
  AND U4073 ( .A(n4131), .B(n4132), .Z(n4130) );
  XOR U4074 ( .A(n4129), .B(n4133), .Z(n4131) );
  XNOR U4075 ( .A(n4113), .B(n4110), .Z(n4122) );
  AND U4076 ( .A(n4134), .B(n4135), .Z(n4110) );
  XOR U4077 ( .A(n4136), .B(n4137), .Z(n4113) );
  AND U4078 ( .A(n4138), .B(n4139), .Z(n4137) );
  XOR U4079 ( .A(n4136), .B(n4140), .Z(n4138) );
  XNOR U4080 ( .A(n4029), .B(n4118), .Z(n4120) );
  XOR U4081 ( .A(n4141), .B(n4142), .Z(n4029) );
  AND U4082 ( .A(n43), .B(n4143), .Z(n4142) );
  XNOR U4083 ( .A(n4144), .B(n4141), .Z(n4143) );
  XOR U4084 ( .A(n4145), .B(n4146), .Z(n4118) );
  AND U4085 ( .A(n4147), .B(n4148), .Z(n4146) );
  XNOR U4086 ( .A(n4145), .B(n4134), .Z(n4148) );
  IV U4087 ( .A(n4080), .Z(n4134) );
  XNOR U4088 ( .A(n4149), .B(n4127), .Z(n4080) );
  XNOR U4089 ( .A(n4150), .B(n4133), .Z(n4127) );
  XOR U4090 ( .A(n4151), .B(n4152), .Z(n4133) );
  NOR U4091 ( .A(n4153), .B(n4154), .Z(n4152) );
  XNOR U4092 ( .A(n4151), .B(n4155), .Z(n4153) );
  XNOR U4093 ( .A(n4132), .B(n4124), .Z(n4150) );
  XOR U4094 ( .A(n4156), .B(n4157), .Z(n4124) );
  AND U4095 ( .A(n4158), .B(n4159), .Z(n4157) );
  XNOR U4096 ( .A(n4156), .B(n4160), .Z(n4158) );
  XNOR U4097 ( .A(n4161), .B(n4129), .Z(n4132) );
  XOR U4098 ( .A(n4162), .B(n4163), .Z(n4129) );
  AND U4099 ( .A(n4164), .B(n4165), .Z(n4163) );
  XOR U4100 ( .A(n4162), .B(n4166), .Z(n4164) );
  XNOR U4101 ( .A(n4167), .B(n4168), .Z(n4161) );
  NOR U4102 ( .A(n4169), .B(n4170), .Z(n4168) );
  XOR U4103 ( .A(n4167), .B(n4171), .Z(n4169) );
  XNOR U4104 ( .A(n4128), .B(n4135), .Z(n4149) );
  NOR U4105 ( .A(n4092), .B(n4172), .Z(n4135) );
  XOR U4106 ( .A(n4140), .B(n4139), .Z(n4128) );
  XNOR U4107 ( .A(n4173), .B(n4136), .Z(n4139) );
  XOR U4108 ( .A(n4174), .B(n4175), .Z(n4136) );
  AND U4109 ( .A(n4176), .B(n4177), .Z(n4175) );
  XOR U4110 ( .A(n4174), .B(n4178), .Z(n4176) );
  XNOR U4111 ( .A(n4179), .B(n4180), .Z(n4173) );
  NOR U4112 ( .A(n4181), .B(n4182), .Z(n4180) );
  XNOR U4113 ( .A(n4179), .B(n4183), .Z(n4181) );
  XOR U4114 ( .A(n4184), .B(n4185), .Z(n4140) );
  NOR U4115 ( .A(n4186), .B(n4187), .Z(n4185) );
  XNOR U4116 ( .A(n4184), .B(n4188), .Z(n4186) );
  XNOR U4117 ( .A(n4077), .B(n4145), .Z(n4147) );
  XOR U4118 ( .A(n4189), .B(n4190), .Z(n4077) );
  AND U4119 ( .A(n43), .B(n4191), .Z(n4190) );
  XOR U4120 ( .A(n4192), .B(n4189), .Z(n4191) );
  AND U4121 ( .A(n4089), .B(n4092), .Z(n4145) );
  XOR U4122 ( .A(n4193), .B(n4172), .Z(n4092) );
  XNOR U4123 ( .A(p_input[1024]), .B(p_input[144]), .Z(n4172) );
  XOR U4124 ( .A(n4160), .B(n4159), .Z(n4193) );
  XNOR U4125 ( .A(n4194), .B(n4166), .Z(n4159) );
  XNOR U4126 ( .A(n4155), .B(n4154), .Z(n4166) );
  XOR U4127 ( .A(n4195), .B(n4151), .Z(n4154) );
  XOR U4128 ( .A(p_input[1034]), .B(p_input[154]), .Z(n4151) );
  XNOR U4129 ( .A(p_input[1035]), .B(p_input[155]), .Z(n4195) );
  XOR U4130 ( .A(p_input[1036]), .B(p_input[156]), .Z(n4155) );
  XNOR U4131 ( .A(n4165), .B(n4156), .Z(n4194) );
  XNOR U4132 ( .A(n3298), .B(p_input[145]), .Z(n4156) );
  XOR U4133 ( .A(n4196), .B(n4171), .Z(n4165) );
  XNOR U4134 ( .A(p_input[1039]), .B(p_input[159]), .Z(n4171) );
  XOR U4135 ( .A(n4162), .B(n4170), .Z(n4196) );
  XOR U4136 ( .A(n4197), .B(n4167), .Z(n4170) );
  XOR U4137 ( .A(p_input[1037]), .B(p_input[157]), .Z(n4167) );
  XNOR U4138 ( .A(p_input[1038]), .B(p_input[158]), .Z(n4197) );
  XOR U4139 ( .A(p_input[1033]), .B(p_input[153]), .Z(n4162) );
  XNOR U4140 ( .A(n4178), .B(n4177), .Z(n4160) );
  XNOR U4141 ( .A(n4198), .B(n4183), .Z(n4177) );
  XOR U4142 ( .A(p_input[1032]), .B(p_input[152]), .Z(n4183) );
  XOR U4143 ( .A(n4174), .B(n4182), .Z(n4198) );
  XOR U4144 ( .A(n4199), .B(n4179), .Z(n4182) );
  XOR U4145 ( .A(p_input[1030]), .B(p_input[150]), .Z(n4179) );
  XNOR U4146 ( .A(p_input[1031]), .B(p_input[151]), .Z(n4199) );
  XOR U4147 ( .A(p_input[1026]), .B(p_input[146]), .Z(n4174) );
  XNOR U4148 ( .A(n4188), .B(n4187), .Z(n4178) );
  XOR U4149 ( .A(n4200), .B(n4184), .Z(n4187) );
  XOR U4150 ( .A(p_input[1027]), .B(p_input[147]), .Z(n4184) );
  XNOR U4151 ( .A(p_input[1028]), .B(p_input[148]), .Z(n4200) );
  XOR U4152 ( .A(p_input[1029]), .B(p_input[149]), .Z(n4188) );
  XOR U4153 ( .A(n4201), .B(n4202), .Z(n4089) );
  AND U4154 ( .A(n43), .B(n4203), .Z(n4202) );
  XNOR U4155 ( .A(n4204), .B(n4201), .Z(n4203) );
  XNOR U4156 ( .A(n4205), .B(n4206), .Z(n43) );
  AND U4157 ( .A(n4207), .B(n4208), .Z(n4206) );
  XOR U4158 ( .A(n4102), .B(n4205), .Z(n4208) );
  AND U4159 ( .A(n4209), .B(n4210), .Z(n4102) );
  XNOR U4160 ( .A(n4099), .B(n4205), .Z(n4207) );
  XOR U4161 ( .A(n4211), .B(n4212), .Z(n4099) );
  AND U4162 ( .A(n47), .B(n4213), .Z(n4212) );
  XOR U4163 ( .A(n4214), .B(n4211), .Z(n4213) );
  XOR U4164 ( .A(n4215), .B(n4216), .Z(n4205) );
  AND U4165 ( .A(n4217), .B(n4218), .Z(n4216) );
  XNOR U4166 ( .A(n4215), .B(n4209), .Z(n4218) );
  IV U4167 ( .A(n4117), .Z(n4209) );
  XOR U4168 ( .A(n4219), .B(n4220), .Z(n4117) );
  XOR U4169 ( .A(n4221), .B(n4210), .Z(n4220) );
  AND U4170 ( .A(n4144), .B(n4222), .Z(n4210) );
  AND U4171 ( .A(n4223), .B(n4224), .Z(n4221) );
  XOR U4172 ( .A(n4225), .B(n4219), .Z(n4223) );
  XNOR U4173 ( .A(n4114), .B(n4215), .Z(n4217) );
  XOR U4174 ( .A(n4226), .B(n4227), .Z(n4114) );
  AND U4175 ( .A(n47), .B(n4228), .Z(n4227) );
  XOR U4176 ( .A(n4229), .B(n4226), .Z(n4228) );
  XOR U4177 ( .A(n4230), .B(n4231), .Z(n4215) );
  AND U4178 ( .A(n4232), .B(n4233), .Z(n4231) );
  XNOR U4179 ( .A(n4230), .B(n4144), .Z(n4233) );
  XOR U4180 ( .A(n4234), .B(n4224), .Z(n4144) );
  XNOR U4181 ( .A(n4235), .B(n4219), .Z(n4224) );
  XOR U4182 ( .A(n4236), .B(n4237), .Z(n4219) );
  AND U4183 ( .A(n4238), .B(n4239), .Z(n4237) );
  XOR U4184 ( .A(n4240), .B(n4236), .Z(n4238) );
  XNOR U4185 ( .A(n4241), .B(n4242), .Z(n4235) );
  AND U4186 ( .A(n4243), .B(n4244), .Z(n4242) );
  XOR U4187 ( .A(n4241), .B(n4245), .Z(n4243) );
  XNOR U4188 ( .A(n4225), .B(n4222), .Z(n4234) );
  AND U4189 ( .A(n4246), .B(n4247), .Z(n4222) );
  XOR U4190 ( .A(n4248), .B(n4249), .Z(n4225) );
  AND U4191 ( .A(n4250), .B(n4251), .Z(n4249) );
  XOR U4192 ( .A(n4248), .B(n4252), .Z(n4250) );
  XNOR U4193 ( .A(n4141), .B(n4230), .Z(n4232) );
  XOR U4194 ( .A(n4253), .B(n4254), .Z(n4141) );
  AND U4195 ( .A(n47), .B(n4255), .Z(n4254) );
  XNOR U4196 ( .A(n4256), .B(n4253), .Z(n4255) );
  XOR U4197 ( .A(n4257), .B(n4258), .Z(n4230) );
  AND U4198 ( .A(n4259), .B(n4260), .Z(n4258) );
  XNOR U4199 ( .A(n4257), .B(n4246), .Z(n4260) );
  IV U4200 ( .A(n4192), .Z(n4246) );
  XNOR U4201 ( .A(n4261), .B(n4239), .Z(n4192) );
  XNOR U4202 ( .A(n4262), .B(n4245), .Z(n4239) );
  XOR U4203 ( .A(n4263), .B(n4264), .Z(n4245) );
  NOR U4204 ( .A(n4265), .B(n4266), .Z(n4264) );
  XNOR U4205 ( .A(n4263), .B(n4267), .Z(n4265) );
  XNOR U4206 ( .A(n4244), .B(n4236), .Z(n4262) );
  XOR U4207 ( .A(n4268), .B(n4269), .Z(n4236) );
  AND U4208 ( .A(n4270), .B(n4271), .Z(n4269) );
  XNOR U4209 ( .A(n4268), .B(n4272), .Z(n4270) );
  XNOR U4210 ( .A(n4273), .B(n4241), .Z(n4244) );
  XOR U4211 ( .A(n4274), .B(n4275), .Z(n4241) );
  AND U4212 ( .A(n4276), .B(n4277), .Z(n4275) );
  XOR U4213 ( .A(n4274), .B(n4278), .Z(n4276) );
  XNOR U4214 ( .A(n4279), .B(n4280), .Z(n4273) );
  NOR U4215 ( .A(n4281), .B(n4282), .Z(n4280) );
  XOR U4216 ( .A(n4279), .B(n4283), .Z(n4281) );
  XNOR U4217 ( .A(n4240), .B(n4247), .Z(n4261) );
  NOR U4218 ( .A(n4204), .B(n4284), .Z(n4247) );
  XOR U4219 ( .A(n4252), .B(n4251), .Z(n4240) );
  XNOR U4220 ( .A(n4285), .B(n4248), .Z(n4251) );
  XOR U4221 ( .A(n4286), .B(n4287), .Z(n4248) );
  AND U4222 ( .A(n4288), .B(n4289), .Z(n4287) );
  XOR U4223 ( .A(n4286), .B(n4290), .Z(n4288) );
  XNOR U4224 ( .A(n4291), .B(n4292), .Z(n4285) );
  NOR U4225 ( .A(n4293), .B(n4294), .Z(n4292) );
  XNOR U4226 ( .A(n4291), .B(n4295), .Z(n4293) );
  XOR U4227 ( .A(n4296), .B(n4297), .Z(n4252) );
  NOR U4228 ( .A(n4298), .B(n4299), .Z(n4297) );
  XNOR U4229 ( .A(n4296), .B(n4300), .Z(n4298) );
  XNOR U4230 ( .A(n4189), .B(n4257), .Z(n4259) );
  XOR U4231 ( .A(n4301), .B(n4302), .Z(n4189) );
  AND U4232 ( .A(n47), .B(n4303), .Z(n4302) );
  XOR U4233 ( .A(n4304), .B(n4301), .Z(n4303) );
  AND U4234 ( .A(n4201), .B(n4204), .Z(n4257) );
  XOR U4235 ( .A(n4305), .B(n4284), .Z(n4204) );
  XNOR U4236 ( .A(p_input[1024]), .B(p_input[160]), .Z(n4284) );
  XOR U4237 ( .A(n4272), .B(n4271), .Z(n4305) );
  XNOR U4238 ( .A(n4306), .B(n4278), .Z(n4271) );
  XNOR U4239 ( .A(n4267), .B(n4266), .Z(n4278) );
  XOR U4240 ( .A(n4307), .B(n4263), .Z(n4266) );
  XOR U4241 ( .A(p_input[1034]), .B(p_input[170]), .Z(n4263) );
  XNOR U4242 ( .A(p_input[1035]), .B(p_input[171]), .Z(n4307) );
  XOR U4243 ( .A(p_input[1036]), .B(p_input[172]), .Z(n4267) );
  XNOR U4244 ( .A(n4277), .B(n4268), .Z(n4306) );
  XNOR U4245 ( .A(n3298), .B(p_input[161]), .Z(n4268) );
  XOR U4246 ( .A(n4308), .B(n4283), .Z(n4277) );
  XNOR U4247 ( .A(p_input[1039]), .B(p_input[175]), .Z(n4283) );
  XOR U4248 ( .A(n4274), .B(n4282), .Z(n4308) );
  XOR U4249 ( .A(n4309), .B(n4279), .Z(n4282) );
  XOR U4250 ( .A(p_input[1037]), .B(p_input[173]), .Z(n4279) );
  XNOR U4251 ( .A(p_input[1038]), .B(p_input[174]), .Z(n4309) );
  XOR U4252 ( .A(p_input[1033]), .B(p_input[169]), .Z(n4274) );
  XNOR U4253 ( .A(n4290), .B(n4289), .Z(n4272) );
  XNOR U4254 ( .A(n4310), .B(n4295), .Z(n4289) );
  XOR U4255 ( .A(p_input[1032]), .B(p_input[168]), .Z(n4295) );
  XOR U4256 ( .A(n4286), .B(n4294), .Z(n4310) );
  XOR U4257 ( .A(n4311), .B(n4291), .Z(n4294) );
  XOR U4258 ( .A(p_input[1030]), .B(p_input[166]), .Z(n4291) );
  XNOR U4259 ( .A(p_input[1031]), .B(p_input[167]), .Z(n4311) );
  XOR U4260 ( .A(p_input[1026]), .B(p_input[162]), .Z(n4286) );
  XNOR U4261 ( .A(n4300), .B(n4299), .Z(n4290) );
  XOR U4262 ( .A(n4312), .B(n4296), .Z(n4299) );
  XOR U4263 ( .A(p_input[1027]), .B(p_input[163]), .Z(n4296) );
  XNOR U4264 ( .A(p_input[1028]), .B(p_input[164]), .Z(n4312) );
  XOR U4265 ( .A(p_input[1029]), .B(p_input[165]), .Z(n4300) );
  XOR U4266 ( .A(n4313), .B(n4314), .Z(n4201) );
  AND U4267 ( .A(n47), .B(n4315), .Z(n4314) );
  XNOR U4268 ( .A(n4316), .B(n4313), .Z(n4315) );
  XNOR U4269 ( .A(n4317), .B(n4318), .Z(n47) );
  AND U4270 ( .A(n4319), .B(n4320), .Z(n4318) );
  XOR U4271 ( .A(n4214), .B(n4317), .Z(n4320) );
  AND U4272 ( .A(n4321), .B(n4322), .Z(n4214) );
  XNOR U4273 ( .A(n4211), .B(n4317), .Z(n4319) );
  XOR U4274 ( .A(n4323), .B(n4324), .Z(n4211) );
  AND U4275 ( .A(n51), .B(n4325), .Z(n4324) );
  XOR U4276 ( .A(n4326), .B(n4323), .Z(n4325) );
  XOR U4277 ( .A(n4327), .B(n4328), .Z(n4317) );
  AND U4278 ( .A(n4329), .B(n4330), .Z(n4328) );
  XNOR U4279 ( .A(n4327), .B(n4321), .Z(n4330) );
  IV U4280 ( .A(n4229), .Z(n4321) );
  XOR U4281 ( .A(n4331), .B(n4332), .Z(n4229) );
  XOR U4282 ( .A(n4333), .B(n4322), .Z(n4332) );
  AND U4283 ( .A(n4256), .B(n4334), .Z(n4322) );
  AND U4284 ( .A(n4335), .B(n4336), .Z(n4333) );
  XOR U4285 ( .A(n4337), .B(n4331), .Z(n4335) );
  XNOR U4286 ( .A(n4226), .B(n4327), .Z(n4329) );
  XOR U4287 ( .A(n4338), .B(n4339), .Z(n4226) );
  AND U4288 ( .A(n51), .B(n4340), .Z(n4339) );
  XOR U4289 ( .A(n4341), .B(n4338), .Z(n4340) );
  XOR U4290 ( .A(n4342), .B(n4343), .Z(n4327) );
  AND U4291 ( .A(n4344), .B(n4345), .Z(n4343) );
  XNOR U4292 ( .A(n4342), .B(n4256), .Z(n4345) );
  XOR U4293 ( .A(n4346), .B(n4336), .Z(n4256) );
  XNOR U4294 ( .A(n4347), .B(n4331), .Z(n4336) );
  XOR U4295 ( .A(n4348), .B(n4349), .Z(n4331) );
  AND U4296 ( .A(n4350), .B(n4351), .Z(n4349) );
  XOR U4297 ( .A(n4352), .B(n4348), .Z(n4350) );
  XNOR U4298 ( .A(n4353), .B(n4354), .Z(n4347) );
  AND U4299 ( .A(n4355), .B(n4356), .Z(n4354) );
  XOR U4300 ( .A(n4353), .B(n4357), .Z(n4355) );
  XNOR U4301 ( .A(n4337), .B(n4334), .Z(n4346) );
  AND U4302 ( .A(n4358), .B(n4359), .Z(n4334) );
  XOR U4303 ( .A(n4360), .B(n4361), .Z(n4337) );
  AND U4304 ( .A(n4362), .B(n4363), .Z(n4361) );
  XOR U4305 ( .A(n4360), .B(n4364), .Z(n4362) );
  XNOR U4306 ( .A(n4253), .B(n4342), .Z(n4344) );
  XOR U4307 ( .A(n4365), .B(n4366), .Z(n4253) );
  AND U4308 ( .A(n51), .B(n4367), .Z(n4366) );
  XNOR U4309 ( .A(n4368), .B(n4365), .Z(n4367) );
  XOR U4310 ( .A(n4369), .B(n4370), .Z(n4342) );
  AND U4311 ( .A(n4371), .B(n4372), .Z(n4370) );
  XNOR U4312 ( .A(n4369), .B(n4358), .Z(n4372) );
  IV U4313 ( .A(n4304), .Z(n4358) );
  XNOR U4314 ( .A(n4373), .B(n4351), .Z(n4304) );
  XNOR U4315 ( .A(n4374), .B(n4357), .Z(n4351) );
  XOR U4316 ( .A(n4375), .B(n4376), .Z(n4357) );
  NOR U4317 ( .A(n4377), .B(n4378), .Z(n4376) );
  XNOR U4318 ( .A(n4375), .B(n4379), .Z(n4377) );
  XNOR U4319 ( .A(n4356), .B(n4348), .Z(n4374) );
  XOR U4320 ( .A(n4380), .B(n4381), .Z(n4348) );
  AND U4321 ( .A(n4382), .B(n4383), .Z(n4381) );
  XNOR U4322 ( .A(n4380), .B(n4384), .Z(n4382) );
  XNOR U4323 ( .A(n4385), .B(n4353), .Z(n4356) );
  XOR U4324 ( .A(n4386), .B(n4387), .Z(n4353) );
  AND U4325 ( .A(n4388), .B(n4389), .Z(n4387) );
  XOR U4326 ( .A(n4386), .B(n4390), .Z(n4388) );
  XNOR U4327 ( .A(n4391), .B(n4392), .Z(n4385) );
  NOR U4328 ( .A(n4393), .B(n4394), .Z(n4392) );
  XOR U4329 ( .A(n4391), .B(n4395), .Z(n4393) );
  XNOR U4330 ( .A(n4352), .B(n4359), .Z(n4373) );
  NOR U4331 ( .A(n4316), .B(n4396), .Z(n4359) );
  XOR U4332 ( .A(n4364), .B(n4363), .Z(n4352) );
  XNOR U4333 ( .A(n4397), .B(n4360), .Z(n4363) );
  XOR U4334 ( .A(n4398), .B(n4399), .Z(n4360) );
  AND U4335 ( .A(n4400), .B(n4401), .Z(n4399) );
  XOR U4336 ( .A(n4398), .B(n4402), .Z(n4400) );
  XNOR U4337 ( .A(n4403), .B(n4404), .Z(n4397) );
  NOR U4338 ( .A(n4405), .B(n4406), .Z(n4404) );
  XNOR U4339 ( .A(n4403), .B(n4407), .Z(n4405) );
  XOR U4340 ( .A(n4408), .B(n4409), .Z(n4364) );
  NOR U4341 ( .A(n4410), .B(n4411), .Z(n4409) );
  XNOR U4342 ( .A(n4408), .B(n4412), .Z(n4410) );
  XNOR U4343 ( .A(n4301), .B(n4369), .Z(n4371) );
  XOR U4344 ( .A(n4413), .B(n4414), .Z(n4301) );
  AND U4345 ( .A(n51), .B(n4415), .Z(n4414) );
  XOR U4346 ( .A(n4416), .B(n4413), .Z(n4415) );
  AND U4347 ( .A(n4313), .B(n4316), .Z(n4369) );
  XOR U4348 ( .A(n4417), .B(n4396), .Z(n4316) );
  XNOR U4349 ( .A(p_input[1024]), .B(p_input[176]), .Z(n4396) );
  XOR U4350 ( .A(n4384), .B(n4383), .Z(n4417) );
  XNOR U4351 ( .A(n4418), .B(n4390), .Z(n4383) );
  XNOR U4352 ( .A(n4379), .B(n4378), .Z(n4390) );
  XOR U4353 ( .A(n4419), .B(n4375), .Z(n4378) );
  XOR U4354 ( .A(p_input[1034]), .B(p_input[186]), .Z(n4375) );
  XNOR U4355 ( .A(p_input[1035]), .B(p_input[187]), .Z(n4419) );
  XOR U4356 ( .A(p_input[1036]), .B(p_input[188]), .Z(n4379) );
  XNOR U4357 ( .A(n4389), .B(n4380), .Z(n4418) );
  XNOR U4358 ( .A(n3298), .B(p_input[177]), .Z(n4380) );
  XOR U4359 ( .A(n4420), .B(n4395), .Z(n4389) );
  XNOR U4360 ( .A(p_input[1039]), .B(p_input[191]), .Z(n4395) );
  XOR U4361 ( .A(n4386), .B(n4394), .Z(n4420) );
  XOR U4362 ( .A(n4421), .B(n4391), .Z(n4394) );
  XOR U4363 ( .A(p_input[1037]), .B(p_input[189]), .Z(n4391) );
  XNOR U4364 ( .A(p_input[1038]), .B(p_input[190]), .Z(n4421) );
  XOR U4365 ( .A(p_input[1033]), .B(p_input[185]), .Z(n4386) );
  XNOR U4366 ( .A(n4402), .B(n4401), .Z(n4384) );
  XNOR U4367 ( .A(n4422), .B(n4407), .Z(n4401) );
  XOR U4368 ( .A(p_input[1032]), .B(p_input[184]), .Z(n4407) );
  XOR U4369 ( .A(n4398), .B(n4406), .Z(n4422) );
  XOR U4370 ( .A(n4423), .B(n4403), .Z(n4406) );
  XOR U4371 ( .A(p_input[1030]), .B(p_input[182]), .Z(n4403) );
  XNOR U4372 ( .A(p_input[1031]), .B(p_input[183]), .Z(n4423) );
  XOR U4373 ( .A(p_input[1026]), .B(p_input[178]), .Z(n4398) );
  XNOR U4374 ( .A(n4412), .B(n4411), .Z(n4402) );
  XOR U4375 ( .A(n4424), .B(n4408), .Z(n4411) );
  XOR U4376 ( .A(p_input[1027]), .B(p_input[179]), .Z(n4408) );
  XNOR U4377 ( .A(p_input[1028]), .B(p_input[180]), .Z(n4424) );
  XOR U4378 ( .A(p_input[1029]), .B(p_input[181]), .Z(n4412) );
  XOR U4379 ( .A(n4425), .B(n4426), .Z(n4313) );
  AND U4380 ( .A(n51), .B(n4427), .Z(n4426) );
  XNOR U4381 ( .A(n4428), .B(n4425), .Z(n4427) );
  XNOR U4382 ( .A(n4429), .B(n4430), .Z(n51) );
  AND U4383 ( .A(n4431), .B(n4432), .Z(n4430) );
  XOR U4384 ( .A(n4326), .B(n4429), .Z(n4432) );
  AND U4385 ( .A(n4433), .B(n4434), .Z(n4326) );
  XNOR U4386 ( .A(n4323), .B(n4429), .Z(n4431) );
  XOR U4387 ( .A(n4435), .B(n4436), .Z(n4323) );
  AND U4388 ( .A(n55), .B(n4437), .Z(n4436) );
  XOR U4389 ( .A(n4438), .B(n4435), .Z(n4437) );
  XOR U4390 ( .A(n4439), .B(n4440), .Z(n4429) );
  AND U4391 ( .A(n4441), .B(n4442), .Z(n4440) );
  XNOR U4392 ( .A(n4439), .B(n4433), .Z(n4442) );
  IV U4393 ( .A(n4341), .Z(n4433) );
  XOR U4394 ( .A(n4443), .B(n4444), .Z(n4341) );
  XOR U4395 ( .A(n4445), .B(n4434), .Z(n4444) );
  AND U4396 ( .A(n4368), .B(n4446), .Z(n4434) );
  AND U4397 ( .A(n4447), .B(n4448), .Z(n4445) );
  XOR U4398 ( .A(n4449), .B(n4443), .Z(n4447) );
  XNOR U4399 ( .A(n4338), .B(n4439), .Z(n4441) );
  XOR U4400 ( .A(n4450), .B(n4451), .Z(n4338) );
  AND U4401 ( .A(n55), .B(n4452), .Z(n4451) );
  XOR U4402 ( .A(n4453), .B(n4450), .Z(n4452) );
  XOR U4403 ( .A(n4454), .B(n4455), .Z(n4439) );
  AND U4404 ( .A(n4456), .B(n4457), .Z(n4455) );
  XNOR U4405 ( .A(n4454), .B(n4368), .Z(n4457) );
  XOR U4406 ( .A(n4458), .B(n4448), .Z(n4368) );
  XNOR U4407 ( .A(n4459), .B(n4443), .Z(n4448) );
  XOR U4408 ( .A(n4460), .B(n4461), .Z(n4443) );
  AND U4409 ( .A(n4462), .B(n4463), .Z(n4461) );
  XOR U4410 ( .A(n4464), .B(n4460), .Z(n4462) );
  XNOR U4411 ( .A(n4465), .B(n4466), .Z(n4459) );
  AND U4412 ( .A(n4467), .B(n4468), .Z(n4466) );
  XOR U4413 ( .A(n4465), .B(n4469), .Z(n4467) );
  XNOR U4414 ( .A(n4449), .B(n4446), .Z(n4458) );
  AND U4415 ( .A(n4470), .B(n4471), .Z(n4446) );
  XOR U4416 ( .A(n4472), .B(n4473), .Z(n4449) );
  AND U4417 ( .A(n4474), .B(n4475), .Z(n4473) );
  XOR U4418 ( .A(n4472), .B(n4476), .Z(n4474) );
  XNOR U4419 ( .A(n4365), .B(n4454), .Z(n4456) );
  XOR U4420 ( .A(n4477), .B(n4478), .Z(n4365) );
  AND U4421 ( .A(n55), .B(n4479), .Z(n4478) );
  XNOR U4422 ( .A(n4480), .B(n4477), .Z(n4479) );
  XOR U4423 ( .A(n4481), .B(n4482), .Z(n4454) );
  AND U4424 ( .A(n4483), .B(n4484), .Z(n4482) );
  XNOR U4425 ( .A(n4481), .B(n4470), .Z(n4484) );
  IV U4426 ( .A(n4416), .Z(n4470) );
  XNOR U4427 ( .A(n4485), .B(n4463), .Z(n4416) );
  XNOR U4428 ( .A(n4486), .B(n4469), .Z(n4463) );
  XOR U4429 ( .A(n4487), .B(n4488), .Z(n4469) );
  NOR U4430 ( .A(n4489), .B(n4490), .Z(n4488) );
  XNOR U4431 ( .A(n4487), .B(n4491), .Z(n4489) );
  XNOR U4432 ( .A(n4468), .B(n4460), .Z(n4486) );
  XOR U4433 ( .A(n4492), .B(n4493), .Z(n4460) );
  AND U4434 ( .A(n4494), .B(n4495), .Z(n4493) );
  XNOR U4435 ( .A(n4492), .B(n4496), .Z(n4494) );
  XNOR U4436 ( .A(n4497), .B(n4465), .Z(n4468) );
  XOR U4437 ( .A(n4498), .B(n4499), .Z(n4465) );
  AND U4438 ( .A(n4500), .B(n4501), .Z(n4499) );
  XOR U4439 ( .A(n4498), .B(n4502), .Z(n4500) );
  XNOR U4440 ( .A(n4503), .B(n4504), .Z(n4497) );
  NOR U4441 ( .A(n4505), .B(n4506), .Z(n4504) );
  XOR U4442 ( .A(n4503), .B(n4507), .Z(n4505) );
  XNOR U4443 ( .A(n4464), .B(n4471), .Z(n4485) );
  NOR U4444 ( .A(n4428), .B(n4508), .Z(n4471) );
  XOR U4445 ( .A(n4476), .B(n4475), .Z(n4464) );
  XNOR U4446 ( .A(n4509), .B(n4472), .Z(n4475) );
  XOR U4447 ( .A(n4510), .B(n4511), .Z(n4472) );
  AND U4448 ( .A(n4512), .B(n4513), .Z(n4511) );
  XOR U4449 ( .A(n4510), .B(n4514), .Z(n4512) );
  XNOR U4450 ( .A(n4515), .B(n4516), .Z(n4509) );
  NOR U4451 ( .A(n4517), .B(n4518), .Z(n4516) );
  XNOR U4452 ( .A(n4515), .B(n4519), .Z(n4517) );
  XOR U4453 ( .A(n4520), .B(n4521), .Z(n4476) );
  NOR U4454 ( .A(n4522), .B(n4523), .Z(n4521) );
  XNOR U4455 ( .A(n4520), .B(n4524), .Z(n4522) );
  XNOR U4456 ( .A(n4413), .B(n4481), .Z(n4483) );
  XOR U4457 ( .A(n4525), .B(n4526), .Z(n4413) );
  AND U4458 ( .A(n55), .B(n4527), .Z(n4526) );
  XOR U4459 ( .A(n4528), .B(n4525), .Z(n4527) );
  AND U4460 ( .A(n4425), .B(n4428), .Z(n4481) );
  XOR U4461 ( .A(n4529), .B(n4508), .Z(n4428) );
  XNOR U4462 ( .A(p_input[1024]), .B(p_input[192]), .Z(n4508) );
  XOR U4463 ( .A(n4496), .B(n4495), .Z(n4529) );
  XNOR U4464 ( .A(n4530), .B(n4502), .Z(n4495) );
  XNOR U4465 ( .A(n4491), .B(n4490), .Z(n4502) );
  XOR U4466 ( .A(n4531), .B(n4487), .Z(n4490) );
  XOR U4467 ( .A(p_input[1034]), .B(p_input[202]), .Z(n4487) );
  XNOR U4468 ( .A(p_input[1035]), .B(p_input[203]), .Z(n4531) );
  XOR U4469 ( .A(p_input[1036]), .B(p_input[204]), .Z(n4491) );
  XNOR U4470 ( .A(n4501), .B(n4492), .Z(n4530) );
  XNOR U4471 ( .A(n3298), .B(p_input[193]), .Z(n4492) );
  XOR U4472 ( .A(n4532), .B(n4507), .Z(n4501) );
  XNOR U4473 ( .A(p_input[1039]), .B(p_input[207]), .Z(n4507) );
  XOR U4474 ( .A(n4498), .B(n4506), .Z(n4532) );
  XOR U4475 ( .A(n4533), .B(n4503), .Z(n4506) );
  XOR U4476 ( .A(p_input[1037]), .B(p_input[205]), .Z(n4503) );
  XNOR U4477 ( .A(p_input[1038]), .B(p_input[206]), .Z(n4533) );
  XOR U4478 ( .A(p_input[1033]), .B(p_input[201]), .Z(n4498) );
  XNOR U4479 ( .A(n4514), .B(n4513), .Z(n4496) );
  XNOR U4480 ( .A(n4534), .B(n4519), .Z(n4513) );
  XOR U4481 ( .A(p_input[1032]), .B(p_input[200]), .Z(n4519) );
  XOR U4482 ( .A(n4510), .B(n4518), .Z(n4534) );
  XOR U4483 ( .A(n4535), .B(n4515), .Z(n4518) );
  XOR U4484 ( .A(p_input[1030]), .B(p_input[198]), .Z(n4515) );
  XNOR U4485 ( .A(p_input[1031]), .B(p_input[199]), .Z(n4535) );
  XOR U4486 ( .A(p_input[1026]), .B(p_input[194]), .Z(n4510) );
  XNOR U4487 ( .A(n4524), .B(n4523), .Z(n4514) );
  XOR U4488 ( .A(n4536), .B(n4520), .Z(n4523) );
  XOR U4489 ( .A(p_input[1027]), .B(p_input[195]), .Z(n4520) );
  XNOR U4490 ( .A(p_input[1028]), .B(p_input[196]), .Z(n4536) );
  XOR U4491 ( .A(p_input[1029]), .B(p_input[197]), .Z(n4524) );
  XOR U4492 ( .A(n4537), .B(n4538), .Z(n4425) );
  AND U4493 ( .A(n55), .B(n4539), .Z(n4538) );
  XNOR U4494 ( .A(n4540), .B(n4537), .Z(n4539) );
  XNOR U4495 ( .A(n4541), .B(n4542), .Z(n55) );
  AND U4496 ( .A(n4543), .B(n4544), .Z(n4542) );
  XOR U4497 ( .A(n4438), .B(n4541), .Z(n4544) );
  AND U4498 ( .A(n4545), .B(n4546), .Z(n4438) );
  XNOR U4499 ( .A(n4435), .B(n4541), .Z(n4543) );
  XOR U4500 ( .A(n4547), .B(n4548), .Z(n4435) );
  AND U4501 ( .A(n59), .B(n4549), .Z(n4548) );
  XOR U4502 ( .A(n4550), .B(n4547), .Z(n4549) );
  XOR U4503 ( .A(n4551), .B(n4552), .Z(n4541) );
  AND U4504 ( .A(n4553), .B(n4554), .Z(n4552) );
  XNOR U4505 ( .A(n4551), .B(n4545), .Z(n4554) );
  IV U4506 ( .A(n4453), .Z(n4545) );
  XOR U4507 ( .A(n4555), .B(n4556), .Z(n4453) );
  XOR U4508 ( .A(n4557), .B(n4546), .Z(n4556) );
  AND U4509 ( .A(n4480), .B(n4558), .Z(n4546) );
  AND U4510 ( .A(n4559), .B(n4560), .Z(n4557) );
  XOR U4511 ( .A(n4561), .B(n4555), .Z(n4559) );
  XNOR U4512 ( .A(n4450), .B(n4551), .Z(n4553) );
  XOR U4513 ( .A(n4562), .B(n4563), .Z(n4450) );
  AND U4514 ( .A(n59), .B(n4564), .Z(n4563) );
  XOR U4515 ( .A(n4565), .B(n4562), .Z(n4564) );
  XOR U4516 ( .A(n4566), .B(n4567), .Z(n4551) );
  AND U4517 ( .A(n4568), .B(n4569), .Z(n4567) );
  XNOR U4518 ( .A(n4566), .B(n4480), .Z(n4569) );
  XOR U4519 ( .A(n4570), .B(n4560), .Z(n4480) );
  XNOR U4520 ( .A(n4571), .B(n4555), .Z(n4560) );
  XOR U4521 ( .A(n4572), .B(n4573), .Z(n4555) );
  AND U4522 ( .A(n4574), .B(n4575), .Z(n4573) );
  XOR U4523 ( .A(n4576), .B(n4572), .Z(n4574) );
  XNOR U4524 ( .A(n4577), .B(n4578), .Z(n4571) );
  AND U4525 ( .A(n4579), .B(n4580), .Z(n4578) );
  XOR U4526 ( .A(n4577), .B(n4581), .Z(n4579) );
  XNOR U4527 ( .A(n4561), .B(n4558), .Z(n4570) );
  AND U4528 ( .A(n4582), .B(n4583), .Z(n4558) );
  XOR U4529 ( .A(n4584), .B(n4585), .Z(n4561) );
  AND U4530 ( .A(n4586), .B(n4587), .Z(n4585) );
  XOR U4531 ( .A(n4584), .B(n4588), .Z(n4586) );
  XNOR U4532 ( .A(n4477), .B(n4566), .Z(n4568) );
  XOR U4533 ( .A(n4589), .B(n4590), .Z(n4477) );
  AND U4534 ( .A(n59), .B(n4591), .Z(n4590) );
  XNOR U4535 ( .A(n4592), .B(n4589), .Z(n4591) );
  XOR U4536 ( .A(n4593), .B(n4594), .Z(n4566) );
  AND U4537 ( .A(n4595), .B(n4596), .Z(n4594) );
  XNOR U4538 ( .A(n4593), .B(n4582), .Z(n4596) );
  IV U4539 ( .A(n4528), .Z(n4582) );
  XNOR U4540 ( .A(n4597), .B(n4575), .Z(n4528) );
  XNOR U4541 ( .A(n4598), .B(n4581), .Z(n4575) );
  XOR U4542 ( .A(n4599), .B(n4600), .Z(n4581) );
  NOR U4543 ( .A(n4601), .B(n4602), .Z(n4600) );
  XNOR U4544 ( .A(n4599), .B(n4603), .Z(n4601) );
  XNOR U4545 ( .A(n4580), .B(n4572), .Z(n4598) );
  XOR U4546 ( .A(n4604), .B(n4605), .Z(n4572) );
  AND U4547 ( .A(n4606), .B(n4607), .Z(n4605) );
  XNOR U4548 ( .A(n4604), .B(n4608), .Z(n4606) );
  XNOR U4549 ( .A(n4609), .B(n4577), .Z(n4580) );
  XOR U4550 ( .A(n4610), .B(n4611), .Z(n4577) );
  AND U4551 ( .A(n4612), .B(n4613), .Z(n4611) );
  XOR U4552 ( .A(n4610), .B(n4614), .Z(n4612) );
  XNOR U4553 ( .A(n4615), .B(n4616), .Z(n4609) );
  NOR U4554 ( .A(n4617), .B(n4618), .Z(n4616) );
  XOR U4555 ( .A(n4615), .B(n4619), .Z(n4617) );
  XNOR U4556 ( .A(n4576), .B(n4583), .Z(n4597) );
  NOR U4557 ( .A(n4540), .B(n4620), .Z(n4583) );
  XOR U4558 ( .A(n4588), .B(n4587), .Z(n4576) );
  XNOR U4559 ( .A(n4621), .B(n4584), .Z(n4587) );
  XOR U4560 ( .A(n4622), .B(n4623), .Z(n4584) );
  AND U4561 ( .A(n4624), .B(n4625), .Z(n4623) );
  XOR U4562 ( .A(n4622), .B(n4626), .Z(n4624) );
  XNOR U4563 ( .A(n4627), .B(n4628), .Z(n4621) );
  NOR U4564 ( .A(n4629), .B(n4630), .Z(n4628) );
  XNOR U4565 ( .A(n4627), .B(n4631), .Z(n4629) );
  XOR U4566 ( .A(n4632), .B(n4633), .Z(n4588) );
  NOR U4567 ( .A(n4634), .B(n4635), .Z(n4633) );
  XNOR U4568 ( .A(n4632), .B(n4636), .Z(n4634) );
  XNOR U4569 ( .A(n4525), .B(n4593), .Z(n4595) );
  XOR U4570 ( .A(n4637), .B(n4638), .Z(n4525) );
  AND U4571 ( .A(n59), .B(n4639), .Z(n4638) );
  XOR U4572 ( .A(n4640), .B(n4637), .Z(n4639) );
  AND U4573 ( .A(n4537), .B(n4540), .Z(n4593) );
  XOR U4574 ( .A(n4641), .B(n4620), .Z(n4540) );
  XNOR U4575 ( .A(p_input[1024]), .B(p_input[208]), .Z(n4620) );
  XOR U4576 ( .A(n4608), .B(n4607), .Z(n4641) );
  XNOR U4577 ( .A(n4642), .B(n4614), .Z(n4607) );
  XNOR U4578 ( .A(n4603), .B(n4602), .Z(n4614) );
  XOR U4579 ( .A(n4643), .B(n4599), .Z(n4602) );
  XOR U4580 ( .A(p_input[1034]), .B(p_input[218]), .Z(n4599) );
  XNOR U4581 ( .A(p_input[1035]), .B(p_input[219]), .Z(n4643) );
  XOR U4582 ( .A(p_input[1036]), .B(p_input[220]), .Z(n4603) );
  XNOR U4583 ( .A(n4613), .B(n4604), .Z(n4642) );
  XNOR U4584 ( .A(n3298), .B(p_input[209]), .Z(n4604) );
  XOR U4585 ( .A(n4644), .B(n4619), .Z(n4613) );
  XNOR U4586 ( .A(p_input[1039]), .B(p_input[223]), .Z(n4619) );
  XOR U4587 ( .A(n4610), .B(n4618), .Z(n4644) );
  XOR U4588 ( .A(n4645), .B(n4615), .Z(n4618) );
  XOR U4589 ( .A(p_input[1037]), .B(p_input[221]), .Z(n4615) );
  XNOR U4590 ( .A(p_input[1038]), .B(p_input[222]), .Z(n4645) );
  XOR U4591 ( .A(p_input[1033]), .B(p_input[217]), .Z(n4610) );
  XNOR U4592 ( .A(n4626), .B(n4625), .Z(n4608) );
  XNOR U4593 ( .A(n4646), .B(n4631), .Z(n4625) );
  XOR U4594 ( .A(p_input[1032]), .B(p_input[216]), .Z(n4631) );
  XOR U4595 ( .A(n4622), .B(n4630), .Z(n4646) );
  XOR U4596 ( .A(n4647), .B(n4627), .Z(n4630) );
  XOR U4597 ( .A(p_input[1030]), .B(p_input[214]), .Z(n4627) );
  XNOR U4598 ( .A(p_input[1031]), .B(p_input[215]), .Z(n4647) );
  XOR U4599 ( .A(p_input[1026]), .B(p_input[210]), .Z(n4622) );
  XNOR U4600 ( .A(n4636), .B(n4635), .Z(n4626) );
  XOR U4601 ( .A(n4648), .B(n4632), .Z(n4635) );
  XOR U4602 ( .A(p_input[1027]), .B(p_input[211]), .Z(n4632) );
  XNOR U4603 ( .A(p_input[1028]), .B(p_input[212]), .Z(n4648) );
  XOR U4604 ( .A(p_input[1029]), .B(p_input[213]), .Z(n4636) );
  XOR U4605 ( .A(n4649), .B(n4650), .Z(n4537) );
  AND U4606 ( .A(n59), .B(n4651), .Z(n4650) );
  XNOR U4607 ( .A(n4652), .B(n4649), .Z(n4651) );
  XNOR U4608 ( .A(n4653), .B(n4654), .Z(n59) );
  AND U4609 ( .A(n4655), .B(n4656), .Z(n4654) );
  XOR U4610 ( .A(n4550), .B(n4653), .Z(n4656) );
  AND U4611 ( .A(n4657), .B(n4658), .Z(n4550) );
  XNOR U4612 ( .A(n4547), .B(n4653), .Z(n4655) );
  XOR U4613 ( .A(n4659), .B(n4660), .Z(n4547) );
  AND U4614 ( .A(n63), .B(n4661), .Z(n4660) );
  XOR U4615 ( .A(n4662), .B(n4659), .Z(n4661) );
  XOR U4616 ( .A(n4663), .B(n4664), .Z(n4653) );
  AND U4617 ( .A(n4665), .B(n4666), .Z(n4664) );
  XNOR U4618 ( .A(n4663), .B(n4657), .Z(n4666) );
  IV U4619 ( .A(n4565), .Z(n4657) );
  XOR U4620 ( .A(n4667), .B(n4668), .Z(n4565) );
  XOR U4621 ( .A(n4669), .B(n4658), .Z(n4668) );
  AND U4622 ( .A(n4592), .B(n4670), .Z(n4658) );
  AND U4623 ( .A(n4671), .B(n4672), .Z(n4669) );
  XOR U4624 ( .A(n4673), .B(n4667), .Z(n4671) );
  XNOR U4625 ( .A(n4562), .B(n4663), .Z(n4665) );
  XOR U4626 ( .A(n4674), .B(n4675), .Z(n4562) );
  AND U4627 ( .A(n63), .B(n4676), .Z(n4675) );
  XOR U4628 ( .A(n4677), .B(n4674), .Z(n4676) );
  XOR U4629 ( .A(n4678), .B(n4679), .Z(n4663) );
  AND U4630 ( .A(n4680), .B(n4681), .Z(n4679) );
  XNOR U4631 ( .A(n4678), .B(n4592), .Z(n4681) );
  XOR U4632 ( .A(n4682), .B(n4672), .Z(n4592) );
  XNOR U4633 ( .A(n4683), .B(n4667), .Z(n4672) );
  XOR U4634 ( .A(n4684), .B(n4685), .Z(n4667) );
  AND U4635 ( .A(n4686), .B(n4687), .Z(n4685) );
  XOR U4636 ( .A(n4688), .B(n4684), .Z(n4686) );
  XNOR U4637 ( .A(n4689), .B(n4690), .Z(n4683) );
  AND U4638 ( .A(n4691), .B(n4692), .Z(n4690) );
  XOR U4639 ( .A(n4689), .B(n4693), .Z(n4691) );
  XNOR U4640 ( .A(n4673), .B(n4670), .Z(n4682) );
  AND U4641 ( .A(n4694), .B(n4695), .Z(n4670) );
  XOR U4642 ( .A(n4696), .B(n4697), .Z(n4673) );
  AND U4643 ( .A(n4698), .B(n4699), .Z(n4697) );
  XOR U4644 ( .A(n4696), .B(n4700), .Z(n4698) );
  XNOR U4645 ( .A(n4589), .B(n4678), .Z(n4680) );
  XOR U4646 ( .A(n4701), .B(n4702), .Z(n4589) );
  AND U4647 ( .A(n63), .B(n4703), .Z(n4702) );
  XNOR U4648 ( .A(n4704), .B(n4701), .Z(n4703) );
  XOR U4649 ( .A(n4705), .B(n4706), .Z(n4678) );
  AND U4650 ( .A(n4707), .B(n4708), .Z(n4706) );
  XNOR U4651 ( .A(n4705), .B(n4694), .Z(n4708) );
  IV U4652 ( .A(n4640), .Z(n4694) );
  XNOR U4653 ( .A(n4709), .B(n4687), .Z(n4640) );
  XNOR U4654 ( .A(n4710), .B(n4693), .Z(n4687) );
  XOR U4655 ( .A(n4711), .B(n4712), .Z(n4693) );
  NOR U4656 ( .A(n4713), .B(n4714), .Z(n4712) );
  XNOR U4657 ( .A(n4711), .B(n4715), .Z(n4713) );
  XNOR U4658 ( .A(n4692), .B(n4684), .Z(n4710) );
  XOR U4659 ( .A(n4716), .B(n4717), .Z(n4684) );
  AND U4660 ( .A(n4718), .B(n4719), .Z(n4717) );
  XNOR U4661 ( .A(n4716), .B(n4720), .Z(n4718) );
  XNOR U4662 ( .A(n4721), .B(n4689), .Z(n4692) );
  XOR U4663 ( .A(n4722), .B(n4723), .Z(n4689) );
  AND U4664 ( .A(n4724), .B(n4725), .Z(n4723) );
  XOR U4665 ( .A(n4722), .B(n4726), .Z(n4724) );
  XNOR U4666 ( .A(n4727), .B(n4728), .Z(n4721) );
  NOR U4667 ( .A(n4729), .B(n4730), .Z(n4728) );
  XOR U4668 ( .A(n4727), .B(n4731), .Z(n4729) );
  XNOR U4669 ( .A(n4688), .B(n4695), .Z(n4709) );
  NOR U4670 ( .A(n4652), .B(n4732), .Z(n4695) );
  XOR U4671 ( .A(n4700), .B(n4699), .Z(n4688) );
  XNOR U4672 ( .A(n4733), .B(n4696), .Z(n4699) );
  XOR U4673 ( .A(n4734), .B(n4735), .Z(n4696) );
  AND U4674 ( .A(n4736), .B(n4737), .Z(n4735) );
  XOR U4675 ( .A(n4734), .B(n4738), .Z(n4736) );
  XNOR U4676 ( .A(n4739), .B(n4740), .Z(n4733) );
  NOR U4677 ( .A(n4741), .B(n4742), .Z(n4740) );
  XNOR U4678 ( .A(n4739), .B(n4743), .Z(n4741) );
  XOR U4679 ( .A(n4744), .B(n4745), .Z(n4700) );
  NOR U4680 ( .A(n4746), .B(n4747), .Z(n4745) );
  XNOR U4681 ( .A(n4744), .B(n4748), .Z(n4746) );
  XNOR U4682 ( .A(n4637), .B(n4705), .Z(n4707) );
  XOR U4683 ( .A(n4749), .B(n4750), .Z(n4637) );
  AND U4684 ( .A(n63), .B(n4751), .Z(n4750) );
  XOR U4685 ( .A(n4752), .B(n4749), .Z(n4751) );
  AND U4686 ( .A(n4649), .B(n4652), .Z(n4705) );
  XOR U4687 ( .A(n4753), .B(n4732), .Z(n4652) );
  XNOR U4688 ( .A(p_input[1024]), .B(p_input[224]), .Z(n4732) );
  XOR U4689 ( .A(n4720), .B(n4719), .Z(n4753) );
  XNOR U4690 ( .A(n4754), .B(n4726), .Z(n4719) );
  XNOR U4691 ( .A(n4715), .B(n4714), .Z(n4726) );
  XOR U4692 ( .A(n4755), .B(n4711), .Z(n4714) );
  XOR U4693 ( .A(p_input[1034]), .B(p_input[234]), .Z(n4711) );
  XNOR U4694 ( .A(p_input[1035]), .B(p_input[235]), .Z(n4755) );
  XOR U4695 ( .A(p_input[1036]), .B(p_input[236]), .Z(n4715) );
  XNOR U4696 ( .A(n4725), .B(n4716), .Z(n4754) );
  XNOR U4697 ( .A(n3298), .B(p_input[225]), .Z(n4716) );
  XOR U4698 ( .A(n4756), .B(n4731), .Z(n4725) );
  XNOR U4699 ( .A(p_input[1039]), .B(p_input[239]), .Z(n4731) );
  XOR U4700 ( .A(n4722), .B(n4730), .Z(n4756) );
  XOR U4701 ( .A(n4757), .B(n4727), .Z(n4730) );
  XOR U4702 ( .A(p_input[1037]), .B(p_input[237]), .Z(n4727) );
  XNOR U4703 ( .A(p_input[1038]), .B(p_input[238]), .Z(n4757) );
  XOR U4704 ( .A(p_input[1033]), .B(p_input[233]), .Z(n4722) );
  XNOR U4705 ( .A(n4738), .B(n4737), .Z(n4720) );
  XNOR U4706 ( .A(n4758), .B(n4743), .Z(n4737) );
  XOR U4707 ( .A(p_input[1032]), .B(p_input[232]), .Z(n4743) );
  XOR U4708 ( .A(n4734), .B(n4742), .Z(n4758) );
  XOR U4709 ( .A(n4759), .B(n4739), .Z(n4742) );
  XOR U4710 ( .A(p_input[1030]), .B(p_input[230]), .Z(n4739) );
  XNOR U4711 ( .A(p_input[1031]), .B(p_input[231]), .Z(n4759) );
  XOR U4712 ( .A(p_input[1026]), .B(p_input[226]), .Z(n4734) );
  XNOR U4713 ( .A(n4748), .B(n4747), .Z(n4738) );
  XOR U4714 ( .A(n4760), .B(n4744), .Z(n4747) );
  XOR U4715 ( .A(p_input[1027]), .B(p_input[227]), .Z(n4744) );
  XNOR U4716 ( .A(p_input[1028]), .B(p_input[228]), .Z(n4760) );
  XOR U4717 ( .A(p_input[1029]), .B(p_input[229]), .Z(n4748) );
  XOR U4718 ( .A(n4761), .B(n4762), .Z(n4649) );
  AND U4719 ( .A(n63), .B(n4763), .Z(n4762) );
  XNOR U4720 ( .A(n4764), .B(n4761), .Z(n4763) );
  XNOR U4721 ( .A(n4765), .B(n4766), .Z(n63) );
  AND U4722 ( .A(n4767), .B(n4768), .Z(n4766) );
  XOR U4723 ( .A(n4662), .B(n4765), .Z(n4768) );
  AND U4724 ( .A(n4769), .B(n4770), .Z(n4662) );
  XNOR U4725 ( .A(n4659), .B(n4765), .Z(n4767) );
  XOR U4726 ( .A(n4771), .B(n4772), .Z(n4659) );
  AND U4727 ( .A(n67), .B(n4773), .Z(n4772) );
  XOR U4728 ( .A(n4774), .B(n4771), .Z(n4773) );
  XOR U4729 ( .A(n4775), .B(n4776), .Z(n4765) );
  AND U4730 ( .A(n4777), .B(n4778), .Z(n4776) );
  XNOR U4731 ( .A(n4775), .B(n4769), .Z(n4778) );
  IV U4732 ( .A(n4677), .Z(n4769) );
  XOR U4733 ( .A(n4779), .B(n4780), .Z(n4677) );
  XOR U4734 ( .A(n4781), .B(n4770), .Z(n4780) );
  AND U4735 ( .A(n4704), .B(n4782), .Z(n4770) );
  AND U4736 ( .A(n4783), .B(n4784), .Z(n4781) );
  XOR U4737 ( .A(n4785), .B(n4779), .Z(n4783) );
  XNOR U4738 ( .A(n4674), .B(n4775), .Z(n4777) );
  XOR U4739 ( .A(n4786), .B(n4787), .Z(n4674) );
  AND U4740 ( .A(n67), .B(n4788), .Z(n4787) );
  XOR U4741 ( .A(n4789), .B(n4786), .Z(n4788) );
  XOR U4742 ( .A(n4790), .B(n4791), .Z(n4775) );
  AND U4743 ( .A(n4792), .B(n4793), .Z(n4791) );
  XNOR U4744 ( .A(n4790), .B(n4704), .Z(n4793) );
  XOR U4745 ( .A(n4794), .B(n4784), .Z(n4704) );
  XNOR U4746 ( .A(n4795), .B(n4779), .Z(n4784) );
  XOR U4747 ( .A(n4796), .B(n4797), .Z(n4779) );
  AND U4748 ( .A(n4798), .B(n4799), .Z(n4797) );
  XOR U4749 ( .A(n4800), .B(n4796), .Z(n4798) );
  XNOR U4750 ( .A(n4801), .B(n4802), .Z(n4795) );
  AND U4751 ( .A(n4803), .B(n4804), .Z(n4802) );
  XOR U4752 ( .A(n4801), .B(n4805), .Z(n4803) );
  XNOR U4753 ( .A(n4785), .B(n4782), .Z(n4794) );
  AND U4754 ( .A(n4806), .B(n4807), .Z(n4782) );
  XOR U4755 ( .A(n4808), .B(n4809), .Z(n4785) );
  AND U4756 ( .A(n4810), .B(n4811), .Z(n4809) );
  XOR U4757 ( .A(n4808), .B(n4812), .Z(n4810) );
  XNOR U4758 ( .A(n4701), .B(n4790), .Z(n4792) );
  XOR U4759 ( .A(n4813), .B(n4814), .Z(n4701) );
  AND U4760 ( .A(n67), .B(n4815), .Z(n4814) );
  XNOR U4761 ( .A(n4816), .B(n4813), .Z(n4815) );
  XOR U4762 ( .A(n4817), .B(n4818), .Z(n4790) );
  AND U4763 ( .A(n4819), .B(n4820), .Z(n4818) );
  XNOR U4764 ( .A(n4817), .B(n4806), .Z(n4820) );
  IV U4765 ( .A(n4752), .Z(n4806) );
  XNOR U4766 ( .A(n4821), .B(n4799), .Z(n4752) );
  XNOR U4767 ( .A(n4822), .B(n4805), .Z(n4799) );
  XOR U4768 ( .A(n4823), .B(n4824), .Z(n4805) );
  NOR U4769 ( .A(n4825), .B(n4826), .Z(n4824) );
  XNOR U4770 ( .A(n4823), .B(n4827), .Z(n4825) );
  XNOR U4771 ( .A(n4804), .B(n4796), .Z(n4822) );
  XOR U4772 ( .A(n4828), .B(n4829), .Z(n4796) );
  AND U4773 ( .A(n4830), .B(n4831), .Z(n4829) );
  XNOR U4774 ( .A(n4828), .B(n4832), .Z(n4830) );
  XNOR U4775 ( .A(n4833), .B(n4801), .Z(n4804) );
  XOR U4776 ( .A(n4834), .B(n4835), .Z(n4801) );
  AND U4777 ( .A(n4836), .B(n4837), .Z(n4835) );
  XOR U4778 ( .A(n4834), .B(n4838), .Z(n4836) );
  XNOR U4779 ( .A(n4839), .B(n4840), .Z(n4833) );
  NOR U4780 ( .A(n4841), .B(n4842), .Z(n4840) );
  XOR U4781 ( .A(n4839), .B(n4843), .Z(n4841) );
  XNOR U4782 ( .A(n4800), .B(n4807), .Z(n4821) );
  NOR U4783 ( .A(n4764), .B(n4844), .Z(n4807) );
  XOR U4784 ( .A(n4812), .B(n4811), .Z(n4800) );
  XNOR U4785 ( .A(n4845), .B(n4808), .Z(n4811) );
  XOR U4786 ( .A(n4846), .B(n4847), .Z(n4808) );
  AND U4787 ( .A(n4848), .B(n4849), .Z(n4847) );
  XOR U4788 ( .A(n4846), .B(n4850), .Z(n4848) );
  XNOR U4789 ( .A(n4851), .B(n4852), .Z(n4845) );
  NOR U4790 ( .A(n4853), .B(n4854), .Z(n4852) );
  XNOR U4791 ( .A(n4851), .B(n4855), .Z(n4853) );
  XOR U4792 ( .A(n4856), .B(n4857), .Z(n4812) );
  NOR U4793 ( .A(n4858), .B(n4859), .Z(n4857) );
  XNOR U4794 ( .A(n4856), .B(n4860), .Z(n4858) );
  XNOR U4795 ( .A(n4749), .B(n4817), .Z(n4819) );
  XOR U4796 ( .A(n4861), .B(n4862), .Z(n4749) );
  AND U4797 ( .A(n67), .B(n4863), .Z(n4862) );
  XOR U4798 ( .A(n4864), .B(n4861), .Z(n4863) );
  AND U4799 ( .A(n4761), .B(n4764), .Z(n4817) );
  XOR U4800 ( .A(n4865), .B(n4844), .Z(n4764) );
  XNOR U4801 ( .A(p_input[1024]), .B(p_input[240]), .Z(n4844) );
  XOR U4802 ( .A(n4832), .B(n4831), .Z(n4865) );
  XNOR U4803 ( .A(n4866), .B(n4838), .Z(n4831) );
  XNOR U4804 ( .A(n4827), .B(n4826), .Z(n4838) );
  XOR U4805 ( .A(n4867), .B(n4823), .Z(n4826) );
  XOR U4806 ( .A(p_input[1034]), .B(p_input[250]), .Z(n4823) );
  XNOR U4807 ( .A(p_input[1035]), .B(p_input[251]), .Z(n4867) );
  XOR U4808 ( .A(p_input[1036]), .B(p_input[252]), .Z(n4827) );
  XNOR U4809 ( .A(n4837), .B(n4828), .Z(n4866) );
  XNOR U4810 ( .A(n3298), .B(p_input[241]), .Z(n4828) );
  XOR U4811 ( .A(n4868), .B(n4843), .Z(n4837) );
  XNOR U4812 ( .A(p_input[1039]), .B(p_input[255]), .Z(n4843) );
  XOR U4813 ( .A(n4834), .B(n4842), .Z(n4868) );
  XOR U4814 ( .A(n4869), .B(n4839), .Z(n4842) );
  XOR U4815 ( .A(p_input[1037]), .B(p_input[253]), .Z(n4839) );
  XNOR U4816 ( .A(p_input[1038]), .B(p_input[254]), .Z(n4869) );
  XOR U4817 ( .A(p_input[1033]), .B(p_input[249]), .Z(n4834) );
  XNOR U4818 ( .A(n4850), .B(n4849), .Z(n4832) );
  XNOR U4819 ( .A(n4870), .B(n4855), .Z(n4849) );
  XOR U4820 ( .A(p_input[1032]), .B(p_input[248]), .Z(n4855) );
  XOR U4821 ( .A(n4846), .B(n4854), .Z(n4870) );
  XOR U4822 ( .A(n4871), .B(n4851), .Z(n4854) );
  XOR U4823 ( .A(p_input[1030]), .B(p_input[246]), .Z(n4851) );
  XNOR U4824 ( .A(p_input[1031]), .B(p_input[247]), .Z(n4871) );
  XOR U4825 ( .A(p_input[1026]), .B(p_input[242]), .Z(n4846) );
  XNOR U4826 ( .A(n4860), .B(n4859), .Z(n4850) );
  XOR U4827 ( .A(n4872), .B(n4856), .Z(n4859) );
  XOR U4828 ( .A(p_input[1027]), .B(p_input[243]), .Z(n4856) );
  XNOR U4829 ( .A(p_input[1028]), .B(p_input[244]), .Z(n4872) );
  XOR U4830 ( .A(p_input[1029]), .B(p_input[245]), .Z(n4860) );
  XOR U4831 ( .A(n4873), .B(n4874), .Z(n4761) );
  AND U4832 ( .A(n67), .B(n4875), .Z(n4874) );
  XNOR U4833 ( .A(n4876), .B(n4873), .Z(n4875) );
  XNOR U4834 ( .A(n4877), .B(n4878), .Z(n67) );
  AND U4835 ( .A(n4879), .B(n4880), .Z(n4878) );
  XOR U4836 ( .A(n4774), .B(n4877), .Z(n4880) );
  AND U4837 ( .A(n4881), .B(n4882), .Z(n4774) );
  XNOR U4838 ( .A(n4771), .B(n4877), .Z(n4879) );
  XOR U4839 ( .A(n4883), .B(n4884), .Z(n4771) );
  AND U4840 ( .A(n71), .B(n4885), .Z(n4884) );
  XOR U4841 ( .A(n4886), .B(n4883), .Z(n4885) );
  XOR U4842 ( .A(n4887), .B(n4888), .Z(n4877) );
  AND U4843 ( .A(n4889), .B(n4890), .Z(n4888) );
  XNOR U4844 ( .A(n4887), .B(n4881), .Z(n4890) );
  IV U4845 ( .A(n4789), .Z(n4881) );
  XOR U4846 ( .A(n4891), .B(n4892), .Z(n4789) );
  XOR U4847 ( .A(n4893), .B(n4882), .Z(n4892) );
  AND U4848 ( .A(n4816), .B(n4894), .Z(n4882) );
  AND U4849 ( .A(n4895), .B(n4896), .Z(n4893) );
  XOR U4850 ( .A(n4897), .B(n4891), .Z(n4895) );
  XNOR U4851 ( .A(n4786), .B(n4887), .Z(n4889) );
  XOR U4852 ( .A(n4898), .B(n4899), .Z(n4786) );
  AND U4853 ( .A(n71), .B(n4900), .Z(n4899) );
  XOR U4854 ( .A(n4901), .B(n4898), .Z(n4900) );
  XOR U4855 ( .A(n4902), .B(n4903), .Z(n4887) );
  AND U4856 ( .A(n4904), .B(n4905), .Z(n4903) );
  XNOR U4857 ( .A(n4902), .B(n4816), .Z(n4905) );
  XOR U4858 ( .A(n4906), .B(n4896), .Z(n4816) );
  XNOR U4859 ( .A(n4907), .B(n4891), .Z(n4896) );
  XOR U4860 ( .A(n4908), .B(n4909), .Z(n4891) );
  AND U4861 ( .A(n4910), .B(n4911), .Z(n4909) );
  XOR U4862 ( .A(n4912), .B(n4908), .Z(n4910) );
  XNOR U4863 ( .A(n4913), .B(n4914), .Z(n4907) );
  AND U4864 ( .A(n4915), .B(n4916), .Z(n4914) );
  XOR U4865 ( .A(n4913), .B(n4917), .Z(n4915) );
  XNOR U4866 ( .A(n4897), .B(n4894), .Z(n4906) );
  AND U4867 ( .A(n4918), .B(n4919), .Z(n4894) );
  XOR U4868 ( .A(n4920), .B(n4921), .Z(n4897) );
  AND U4869 ( .A(n4922), .B(n4923), .Z(n4921) );
  XOR U4870 ( .A(n4920), .B(n4924), .Z(n4922) );
  XNOR U4871 ( .A(n4813), .B(n4902), .Z(n4904) );
  XOR U4872 ( .A(n4925), .B(n4926), .Z(n4813) );
  AND U4873 ( .A(n71), .B(n4927), .Z(n4926) );
  XNOR U4874 ( .A(n4928), .B(n4925), .Z(n4927) );
  XOR U4875 ( .A(n4929), .B(n4930), .Z(n4902) );
  AND U4876 ( .A(n4931), .B(n4932), .Z(n4930) );
  XNOR U4877 ( .A(n4929), .B(n4918), .Z(n4932) );
  IV U4878 ( .A(n4864), .Z(n4918) );
  XNOR U4879 ( .A(n4933), .B(n4911), .Z(n4864) );
  XNOR U4880 ( .A(n4934), .B(n4917), .Z(n4911) );
  XOR U4881 ( .A(n4935), .B(n4936), .Z(n4917) );
  NOR U4882 ( .A(n4937), .B(n4938), .Z(n4936) );
  XNOR U4883 ( .A(n4935), .B(n4939), .Z(n4937) );
  XNOR U4884 ( .A(n4916), .B(n4908), .Z(n4934) );
  XOR U4885 ( .A(n4940), .B(n4941), .Z(n4908) );
  AND U4886 ( .A(n4942), .B(n4943), .Z(n4941) );
  XNOR U4887 ( .A(n4940), .B(n4944), .Z(n4942) );
  XNOR U4888 ( .A(n4945), .B(n4913), .Z(n4916) );
  XOR U4889 ( .A(n4946), .B(n4947), .Z(n4913) );
  AND U4890 ( .A(n4948), .B(n4949), .Z(n4947) );
  XOR U4891 ( .A(n4946), .B(n4950), .Z(n4948) );
  XNOR U4892 ( .A(n4951), .B(n4952), .Z(n4945) );
  NOR U4893 ( .A(n4953), .B(n4954), .Z(n4952) );
  XOR U4894 ( .A(n4951), .B(n4955), .Z(n4953) );
  XNOR U4895 ( .A(n4912), .B(n4919), .Z(n4933) );
  NOR U4896 ( .A(n4876), .B(n4956), .Z(n4919) );
  XOR U4897 ( .A(n4924), .B(n4923), .Z(n4912) );
  XNOR U4898 ( .A(n4957), .B(n4920), .Z(n4923) );
  XOR U4899 ( .A(n4958), .B(n4959), .Z(n4920) );
  AND U4900 ( .A(n4960), .B(n4961), .Z(n4959) );
  XOR U4901 ( .A(n4958), .B(n4962), .Z(n4960) );
  XNOR U4902 ( .A(n4963), .B(n4964), .Z(n4957) );
  NOR U4903 ( .A(n4965), .B(n4966), .Z(n4964) );
  XNOR U4904 ( .A(n4963), .B(n4967), .Z(n4965) );
  XOR U4905 ( .A(n4968), .B(n4969), .Z(n4924) );
  NOR U4906 ( .A(n4970), .B(n4971), .Z(n4969) );
  XNOR U4907 ( .A(n4968), .B(n4972), .Z(n4970) );
  XNOR U4908 ( .A(n4861), .B(n4929), .Z(n4931) );
  XOR U4909 ( .A(n4973), .B(n4974), .Z(n4861) );
  AND U4910 ( .A(n71), .B(n4975), .Z(n4974) );
  XOR U4911 ( .A(n4976), .B(n4973), .Z(n4975) );
  AND U4912 ( .A(n4873), .B(n4876), .Z(n4929) );
  XOR U4913 ( .A(n4977), .B(n4956), .Z(n4876) );
  XNOR U4914 ( .A(p_input[1024]), .B(p_input[256]), .Z(n4956) );
  XOR U4915 ( .A(n4944), .B(n4943), .Z(n4977) );
  XNOR U4916 ( .A(n4978), .B(n4950), .Z(n4943) );
  XNOR U4917 ( .A(n4939), .B(n4938), .Z(n4950) );
  XOR U4918 ( .A(n4979), .B(n4935), .Z(n4938) );
  XOR U4919 ( .A(p_input[1034]), .B(p_input[266]), .Z(n4935) );
  XNOR U4920 ( .A(p_input[1035]), .B(p_input[267]), .Z(n4979) );
  XOR U4921 ( .A(p_input[1036]), .B(p_input[268]), .Z(n4939) );
  XNOR U4922 ( .A(n4949), .B(n4940), .Z(n4978) );
  XNOR U4923 ( .A(n3298), .B(p_input[257]), .Z(n4940) );
  XOR U4924 ( .A(n4980), .B(n4955), .Z(n4949) );
  XNOR U4925 ( .A(p_input[1039]), .B(p_input[271]), .Z(n4955) );
  XOR U4926 ( .A(n4946), .B(n4954), .Z(n4980) );
  XOR U4927 ( .A(n4981), .B(n4951), .Z(n4954) );
  XOR U4928 ( .A(p_input[1037]), .B(p_input[269]), .Z(n4951) );
  XNOR U4929 ( .A(p_input[1038]), .B(p_input[270]), .Z(n4981) );
  XOR U4930 ( .A(p_input[1033]), .B(p_input[265]), .Z(n4946) );
  XNOR U4931 ( .A(n4962), .B(n4961), .Z(n4944) );
  XNOR U4932 ( .A(n4982), .B(n4967), .Z(n4961) );
  XOR U4933 ( .A(p_input[1032]), .B(p_input[264]), .Z(n4967) );
  XOR U4934 ( .A(n4958), .B(n4966), .Z(n4982) );
  XOR U4935 ( .A(n4983), .B(n4963), .Z(n4966) );
  XOR U4936 ( .A(p_input[1030]), .B(p_input[262]), .Z(n4963) );
  XNOR U4937 ( .A(p_input[1031]), .B(p_input[263]), .Z(n4983) );
  XOR U4938 ( .A(p_input[1026]), .B(p_input[258]), .Z(n4958) );
  XNOR U4939 ( .A(n4972), .B(n4971), .Z(n4962) );
  XOR U4940 ( .A(n4984), .B(n4968), .Z(n4971) );
  XOR U4941 ( .A(p_input[1027]), .B(p_input[259]), .Z(n4968) );
  XNOR U4942 ( .A(p_input[1028]), .B(p_input[260]), .Z(n4984) );
  XOR U4943 ( .A(p_input[1029]), .B(p_input[261]), .Z(n4972) );
  XOR U4944 ( .A(n4985), .B(n4986), .Z(n4873) );
  AND U4945 ( .A(n71), .B(n4987), .Z(n4986) );
  XNOR U4946 ( .A(n4988), .B(n4985), .Z(n4987) );
  XNOR U4947 ( .A(n4989), .B(n4990), .Z(n71) );
  AND U4948 ( .A(n4991), .B(n4992), .Z(n4990) );
  XOR U4949 ( .A(n4886), .B(n4989), .Z(n4992) );
  AND U4950 ( .A(n4993), .B(n4994), .Z(n4886) );
  XNOR U4951 ( .A(n4883), .B(n4989), .Z(n4991) );
  XOR U4952 ( .A(n4995), .B(n4996), .Z(n4883) );
  AND U4953 ( .A(n75), .B(n4997), .Z(n4996) );
  XOR U4954 ( .A(n4998), .B(n4995), .Z(n4997) );
  XOR U4955 ( .A(n4999), .B(n5000), .Z(n4989) );
  AND U4956 ( .A(n5001), .B(n5002), .Z(n5000) );
  XNOR U4957 ( .A(n4999), .B(n4993), .Z(n5002) );
  IV U4958 ( .A(n4901), .Z(n4993) );
  XOR U4959 ( .A(n5003), .B(n5004), .Z(n4901) );
  XOR U4960 ( .A(n5005), .B(n4994), .Z(n5004) );
  AND U4961 ( .A(n4928), .B(n5006), .Z(n4994) );
  AND U4962 ( .A(n5007), .B(n5008), .Z(n5005) );
  XOR U4963 ( .A(n5009), .B(n5003), .Z(n5007) );
  XNOR U4964 ( .A(n4898), .B(n4999), .Z(n5001) );
  XOR U4965 ( .A(n5010), .B(n5011), .Z(n4898) );
  AND U4966 ( .A(n75), .B(n5012), .Z(n5011) );
  XOR U4967 ( .A(n5013), .B(n5010), .Z(n5012) );
  XOR U4968 ( .A(n5014), .B(n5015), .Z(n4999) );
  AND U4969 ( .A(n5016), .B(n5017), .Z(n5015) );
  XNOR U4970 ( .A(n5014), .B(n4928), .Z(n5017) );
  XOR U4971 ( .A(n5018), .B(n5008), .Z(n4928) );
  XNOR U4972 ( .A(n5019), .B(n5003), .Z(n5008) );
  XOR U4973 ( .A(n5020), .B(n5021), .Z(n5003) );
  AND U4974 ( .A(n5022), .B(n5023), .Z(n5021) );
  XOR U4975 ( .A(n5024), .B(n5020), .Z(n5022) );
  XNOR U4976 ( .A(n5025), .B(n5026), .Z(n5019) );
  AND U4977 ( .A(n5027), .B(n5028), .Z(n5026) );
  XOR U4978 ( .A(n5025), .B(n5029), .Z(n5027) );
  XNOR U4979 ( .A(n5009), .B(n5006), .Z(n5018) );
  AND U4980 ( .A(n5030), .B(n5031), .Z(n5006) );
  XOR U4981 ( .A(n5032), .B(n5033), .Z(n5009) );
  AND U4982 ( .A(n5034), .B(n5035), .Z(n5033) );
  XOR U4983 ( .A(n5032), .B(n5036), .Z(n5034) );
  XNOR U4984 ( .A(n4925), .B(n5014), .Z(n5016) );
  XOR U4985 ( .A(n5037), .B(n5038), .Z(n4925) );
  AND U4986 ( .A(n75), .B(n5039), .Z(n5038) );
  XNOR U4987 ( .A(n5040), .B(n5037), .Z(n5039) );
  XOR U4988 ( .A(n5041), .B(n5042), .Z(n5014) );
  AND U4989 ( .A(n5043), .B(n5044), .Z(n5042) );
  XNOR U4990 ( .A(n5041), .B(n5030), .Z(n5044) );
  IV U4991 ( .A(n4976), .Z(n5030) );
  XNOR U4992 ( .A(n5045), .B(n5023), .Z(n4976) );
  XNOR U4993 ( .A(n5046), .B(n5029), .Z(n5023) );
  XOR U4994 ( .A(n5047), .B(n5048), .Z(n5029) );
  NOR U4995 ( .A(n5049), .B(n5050), .Z(n5048) );
  XNOR U4996 ( .A(n5047), .B(n5051), .Z(n5049) );
  XNOR U4997 ( .A(n5028), .B(n5020), .Z(n5046) );
  XOR U4998 ( .A(n5052), .B(n5053), .Z(n5020) );
  AND U4999 ( .A(n5054), .B(n5055), .Z(n5053) );
  XNOR U5000 ( .A(n5052), .B(n5056), .Z(n5054) );
  XNOR U5001 ( .A(n5057), .B(n5025), .Z(n5028) );
  XOR U5002 ( .A(n5058), .B(n5059), .Z(n5025) );
  AND U5003 ( .A(n5060), .B(n5061), .Z(n5059) );
  XOR U5004 ( .A(n5058), .B(n5062), .Z(n5060) );
  XNOR U5005 ( .A(n5063), .B(n5064), .Z(n5057) );
  NOR U5006 ( .A(n5065), .B(n5066), .Z(n5064) );
  XOR U5007 ( .A(n5063), .B(n5067), .Z(n5065) );
  XNOR U5008 ( .A(n5024), .B(n5031), .Z(n5045) );
  NOR U5009 ( .A(n4988), .B(n5068), .Z(n5031) );
  XOR U5010 ( .A(n5036), .B(n5035), .Z(n5024) );
  XNOR U5011 ( .A(n5069), .B(n5032), .Z(n5035) );
  XOR U5012 ( .A(n5070), .B(n5071), .Z(n5032) );
  AND U5013 ( .A(n5072), .B(n5073), .Z(n5071) );
  XOR U5014 ( .A(n5070), .B(n5074), .Z(n5072) );
  XNOR U5015 ( .A(n5075), .B(n5076), .Z(n5069) );
  NOR U5016 ( .A(n5077), .B(n5078), .Z(n5076) );
  XNOR U5017 ( .A(n5075), .B(n5079), .Z(n5077) );
  XOR U5018 ( .A(n5080), .B(n5081), .Z(n5036) );
  NOR U5019 ( .A(n5082), .B(n5083), .Z(n5081) );
  XNOR U5020 ( .A(n5080), .B(n5084), .Z(n5082) );
  XNOR U5021 ( .A(n4973), .B(n5041), .Z(n5043) );
  XOR U5022 ( .A(n5085), .B(n5086), .Z(n4973) );
  AND U5023 ( .A(n75), .B(n5087), .Z(n5086) );
  XOR U5024 ( .A(n5088), .B(n5085), .Z(n5087) );
  AND U5025 ( .A(n4985), .B(n4988), .Z(n5041) );
  XOR U5026 ( .A(n5089), .B(n5068), .Z(n4988) );
  XNOR U5027 ( .A(p_input[1024]), .B(p_input[272]), .Z(n5068) );
  XOR U5028 ( .A(n5056), .B(n5055), .Z(n5089) );
  XNOR U5029 ( .A(n5090), .B(n5062), .Z(n5055) );
  XNOR U5030 ( .A(n5051), .B(n5050), .Z(n5062) );
  XOR U5031 ( .A(n5091), .B(n5047), .Z(n5050) );
  XOR U5032 ( .A(p_input[1034]), .B(p_input[282]), .Z(n5047) );
  XNOR U5033 ( .A(p_input[1035]), .B(p_input[283]), .Z(n5091) );
  XOR U5034 ( .A(p_input[1036]), .B(p_input[284]), .Z(n5051) );
  XNOR U5035 ( .A(n5061), .B(n5052), .Z(n5090) );
  XNOR U5036 ( .A(n3298), .B(p_input[273]), .Z(n5052) );
  XOR U5037 ( .A(n5092), .B(n5067), .Z(n5061) );
  XNOR U5038 ( .A(p_input[1039]), .B(p_input[287]), .Z(n5067) );
  XOR U5039 ( .A(n5058), .B(n5066), .Z(n5092) );
  XOR U5040 ( .A(n5093), .B(n5063), .Z(n5066) );
  XOR U5041 ( .A(p_input[1037]), .B(p_input[285]), .Z(n5063) );
  XNOR U5042 ( .A(p_input[1038]), .B(p_input[286]), .Z(n5093) );
  XOR U5043 ( .A(p_input[1033]), .B(p_input[281]), .Z(n5058) );
  XNOR U5044 ( .A(n5074), .B(n5073), .Z(n5056) );
  XNOR U5045 ( .A(n5094), .B(n5079), .Z(n5073) );
  XOR U5046 ( .A(p_input[1032]), .B(p_input[280]), .Z(n5079) );
  XOR U5047 ( .A(n5070), .B(n5078), .Z(n5094) );
  XOR U5048 ( .A(n5095), .B(n5075), .Z(n5078) );
  XOR U5049 ( .A(p_input[1030]), .B(p_input[278]), .Z(n5075) );
  XNOR U5050 ( .A(p_input[1031]), .B(p_input[279]), .Z(n5095) );
  XOR U5051 ( .A(p_input[1026]), .B(p_input[274]), .Z(n5070) );
  XNOR U5052 ( .A(n5084), .B(n5083), .Z(n5074) );
  XOR U5053 ( .A(n5096), .B(n5080), .Z(n5083) );
  XOR U5054 ( .A(p_input[1027]), .B(p_input[275]), .Z(n5080) );
  XNOR U5055 ( .A(p_input[1028]), .B(p_input[276]), .Z(n5096) );
  XOR U5056 ( .A(p_input[1029]), .B(p_input[277]), .Z(n5084) );
  XOR U5057 ( .A(n5097), .B(n5098), .Z(n4985) );
  AND U5058 ( .A(n75), .B(n5099), .Z(n5098) );
  XNOR U5059 ( .A(n5100), .B(n5097), .Z(n5099) );
  XNOR U5060 ( .A(n5101), .B(n5102), .Z(n75) );
  AND U5061 ( .A(n5103), .B(n5104), .Z(n5102) );
  XOR U5062 ( .A(n4998), .B(n5101), .Z(n5104) );
  AND U5063 ( .A(n5105), .B(n5106), .Z(n4998) );
  XNOR U5064 ( .A(n4995), .B(n5101), .Z(n5103) );
  XOR U5065 ( .A(n5107), .B(n5108), .Z(n4995) );
  AND U5066 ( .A(n79), .B(n5109), .Z(n5108) );
  XOR U5067 ( .A(n5110), .B(n5107), .Z(n5109) );
  XOR U5068 ( .A(n5111), .B(n5112), .Z(n5101) );
  AND U5069 ( .A(n5113), .B(n5114), .Z(n5112) );
  XNOR U5070 ( .A(n5111), .B(n5105), .Z(n5114) );
  IV U5071 ( .A(n5013), .Z(n5105) );
  XOR U5072 ( .A(n5115), .B(n5116), .Z(n5013) );
  XOR U5073 ( .A(n5117), .B(n5106), .Z(n5116) );
  AND U5074 ( .A(n5040), .B(n5118), .Z(n5106) );
  AND U5075 ( .A(n5119), .B(n5120), .Z(n5117) );
  XOR U5076 ( .A(n5121), .B(n5115), .Z(n5119) );
  XNOR U5077 ( .A(n5010), .B(n5111), .Z(n5113) );
  XOR U5078 ( .A(n5122), .B(n5123), .Z(n5010) );
  AND U5079 ( .A(n79), .B(n5124), .Z(n5123) );
  XOR U5080 ( .A(n5125), .B(n5122), .Z(n5124) );
  XOR U5081 ( .A(n5126), .B(n5127), .Z(n5111) );
  AND U5082 ( .A(n5128), .B(n5129), .Z(n5127) );
  XNOR U5083 ( .A(n5126), .B(n5040), .Z(n5129) );
  XOR U5084 ( .A(n5130), .B(n5120), .Z(n5040) );
  XNOR U5085 ( .A(n5131), .B(n5115), .Z(n5120) );
  XOR U5086 ( .A(n5132), .B(n5133), .Z(n5115) );
  AND U5087 ( .A(n5134), .B(n5135), .Z(n5133) );
  XOR U5088 ( .A(n5136), .B(n5132), .Z(n5134) );
  XNOR U5089 ( .A(n5137), .B(n5138), .Z(n5131) );
  AND U5090 ( .A(n5139), .B(n5140), .Z(n5138) );
  XOR U5091 ( .A(n5137), .B(n5141), .Z(n5139) );
  XNOR U5092 ( .A(n5121), .B(n5118), .Z(n5130) );
  AND U5093 ( .A(n5142), .B(n5143), .Z(n5118) );
  XOR U5094 ( .A(n5144), .B(n5145), .Z(n5121) );
  AND U5095 ( .A(n5146), .B(n5147), .Z(n5145) );
  XOR U5096 ( .A(n5144), .B(n5148), .Z(n5146) );
  XNOR U5097 ( .A(n5037), .B(n5126), .Z(n5128) );
  XOR U5098 ( .A(n5149), .B(n5150), .Z(n5037) );
  AND U5099 ( .A(n79), .B(n5151), .Z(n5150) );
  XNOR U5100 ( .A(n5152), .B(n5149), .Z(n5151) );
  XOR U5101 ( .A(n5153), .B(n5154), .Z(n5126) );
  AND U5102 ( .A(n5155), .B(n5156), .Z(n5154) );
  XNOR U5103 ( .A(n5153), .B(n5142), .Z(n5156) );
  IV U5104 ( .A(n5088), .Z(n5142) );
  XNOR U5105 ( .A(n5157), .B(n5135), .Z(n5088) );
  XNOR U5106 ( .A(n5158), .B(n5141), .Z(n5135) );
  XOR U5107 ( .A(n5159), .B(n5160), .Z(n5141) );
  NOR U5108 ( .A(n5161), .B(n5162), .Z(n5160) );
  XNOR U5109 ( .A(n5159), .B(n5163), .Z(n5161) );
  XNOR U5110 ( .A(n5140), .B(n5132), .Z(n5158) );
  XOR U5111 ( .A(n5164), .B(n5165), .Z(n5132) );
  AND U5112 ( .A(n5166), .B(n5167), .Z(n5165) );
  XNOR U5113 ( .A(n5164), .B(n5168), .Z(n5166) );
  XNOR U5114 ( .A(n5169), .B(n5137), .Z(n5140) );
  XOR U5115 ( .A(n5170), .B(n5171), .Z(n5137) );
  AND U5116 ( .A(n5172), .B(n5173), .Z(n5171) );
  XOR U5117 ( .A(n5170), .B(n5174), .Z(n5172) );
  XNOR U5118 ( .A(n5175), .B(n5176), .Z(n5169) );
  NOR U5119 ( .A(n5177), .B(n5178), .Z(n5176) );
  XOR U5120 ( .A(n5175), .B(n5179), .Z(n5177) );
  XNOR U5121 ( .A(n5136), .B(n5143), .Z(n5157) );
  NOR U5122 ( .A(n5100), .B(n5180), .Z(n5143) );
  XOR U5123 ( .A(n5148), .B(n5147), .Z(n5136) );
  XNOR U5124 ( .A(n5181), .B(n5144), .Z(n5147) );
  XOR U5125 ( .A(n5182), .B(n5183), .Z(n5144) );
  AND U5126 ( .A(n5184), .B(n5185), .Z(n5183) );
  XOR U5127 ( .A(n5182), .B(n5186), .Z(n5184) );
  XNOR U5128 ( .A(n5187), .B(n5188), .Z(n5181) );
  NOR U5129 ( .A(n5189), .B(n5190), .Z(n5188) );
  XNOR U5130 ( .A(n5187), .B(n5191), .Z(n5189) );
  XOR U5131 ( .A(n5192), .B(n5193), .Z(n5148) );
  NOR U5132 ( .A(n5194), .B(n5195), .Z(n5193) );
  XNOR U5133 ( .A(n5192), .B(n5196), .Z(n5194) );
  XNOR U5134 ( .A(n5085), .B(n5153), .Z(n5155) );
  XOR U5135 ( .A(n5197), .B(n5198), .Z(n5085) );
  AND U5136 ( .A(n79), .B(n5199), .Z(n5198) );
  XOR U5137 ( .A(n5200), .B(n5197), .Z(n5199) );
  AND U5138 ( .A(n5097), .B(n5100), .Z(n5153) );
  XOR U5139 ( .A(n5201), .B(n5180), .Z(n5100) );
  XNOR U5140 ( .A(p_input[1024]), .B(p_input[288]), .Z(n5180) );
  XOR U5141 ( .A(n5168), .B(n5167), .Z(n5201) );
  XNOR U5142 ( .A(n5202), .B(n5174), .Z(n5167) );
  XNOR U5143 ( .A(n5163), .B(n5162), .Z(n5174) );
  XOR U5144 ( .A(n5203), .B(n5159), .Z(n5162) );
  XOR U5145 ( .A(p_input[1034]), .B(p_input[298]), .Z(n5159) );
  XNOR U5146 ( .A(p_input[1035]), .B(p_input[299]), .Z(n5203) );
  XOR U5147 ( .A(p_input[1036]), .B(p_input[300]), .Z(n5163) );
  XNOR U5148 ( .A(n5173), .B(n5164), .Z(n5202) );
  XNOR U5149 ( .A(n3298), .B(p_input[289]), .Z(n5164) );
  XOR U5150 ( .A(n5204), .B(n5179), .Z(n5173) );
  XNOR U5151 ( .A(p_input[1039]), .B(p_input[303]), .Z(n5179) );
  XOR U5152 ( .A(n5170), .B(n5178), .Z(n5204) );
  XOR U5153 ( .A(n5205), .B(n5175), .Z(n5178) );
  XOR U5154 ( .A(p_input[1037]), .B(p_input[301]), .Z(n5175) );
  XNOR U5155 ( .A(p_input[1038]), .B(p_input[302]), .Z(n5205) );
  XOR U5156 ( .A(p_input[1033]), .B(p_input[297]), .Z(n5170) );
  XNOR U5157 ( .A(n5186), .B(n5185), .Z(n5168) );
  XNOR U5158 ( .A(n5206), .B(n5191), .Z(n5185) );
  XOR U5159 ( .A(p_input[1032]), .B(p_input[296]), .Z(n5191) );
  XOR U5160 ( .A(n5182), .B(n5190), .Z(n5206) );
  XOR U5161 ( .A(n5207), .B(n5187), .Z(n5190) );
  XOR U5162 ( .A(p_input[1030]), .B(p_input[294]), .Z(n5187) );
  XNOR U5163 ( .A(p_input[1031]), .B(p_input[295]), .Z(n5207) );
  XOR U5164 ( .A(p_input[1026]), .B(p_input[290]), .Z(n5182) );
  XNOR U5165 ( .A(n5196), .B(n5195), .Z(n5186) );
  XOR U5166 ( .A(n5208), .B(n5192), .Z(n5195) );
  XOR U5167 ( .A(p_input[1027]), .B(p_input[291]), .Z(n5192) );
  XNOR U5168 ( .A(p_input[1028]), .B(p_input[292]), .Z(n5208) );
  XOR U5169 ( .A(p_input[1029]), .B(p_input[293]), .Z(n5196) );
  XOR U5170 ( .A(n5209), .B(n5210), .Z(n5097) );
  AND U5171 ( .A(n79), .B(n5211), .Z(n5210) );
  XNOR U5172 ( .A(n5212), .B(n5209), .Z(n5211) );
  XNOR U5173 ( .A(n5213), .B(n5214), .Z(n79) );
  AND U5174 ( .A(n5215), .B(n5216), .Z(n5214) );
  XOR U5175 ( .A(n5110), .B(n5213), .Z(n5216) );
  AND U5176 ( .A(n5217), .B(n5218), .Z(n5110) );
  XNOR U5177 ( .A(n5107), .B(n5213), .Z(n5215) );
  XOR U5178 ( .A(n5219), .B(n5220), .Z(n5107) );
  AND U5179 ( .A(n83), .B(n5221), .Z(n5220) );
  XOR U5180 ( .A(n5222), .B(n5219), .Z(n5221) );
  XOR U5181 ( .A(n5223), .B(n5224), .Z(n5213) );
  AND U5182 ( .A(n5225), .B(n5226), .Z(n5224) );
  XNOR U5183 ( .A(n5223), .B(n5217), .Z(n5226) );
  IV U5184 ( .A(n5125), .Z(n5217) );
  XOR U5185 ( .A(n5227), .B(n5228), .Z(n5125) );
  XOR U5186 ( .A(n5229), .B(n5218), .Z(n5228) );
  AND U5187 ( .A(n5152), .B(n5230), .Z(n5218) );
  AND U5188 ( .A(n5231), .B(n5232), .Z(n5229) );
  XOR U5189 ( .A(n5233), .B(n5227), .Z(n5231) );
  XNOR U5190 ( .A(n5122), .B(n5223), .Z(n5225) );
  XOR U5191 ( .A(n5234), .B(n5235), .Z(n5122) );
  AND U5192 ( .A(n83), .B(n5236), .Z(n5235) );
  XOR U5193 ( .A(n5237), .B(n5234), .Z(n5236) );
  XOR U5194 ( .A(n5238), .B(n5239), .Z(n5223) );
  AND U5195 ( .A(n5240), .B(n5241), .Z(n5239) );
  XNOR U5196 ( .A(n5238), .B(n5152), .Z(n5241) );
  XOR U5197 ( .A(n5242), .B(n5232), .Z(n5152) );
  XNOR U5198 ( .A(n5243), .B(n5227), .Z(n5232) );
  XOR U5199 ( .A(n5244), .B(n5245), .Z(n5227) );
  AND U5200 ( .A(n5246), .B(n5247), .Z(n5245) );
  XOR U5201 ( .A(n5248), .B(n5244), .Z(n5246) );
  XNOR U5202 ( .A(n5249), .B(n5250), .Z(n5243) );
  AND U5203 ( .A(n5251), .B(n5252), .Z(n5250) );
  XOR U5204 ( .A(n5249), .B(n5253), .Z(n5251) );
  XNOR U5205 ( .A(n5233), .B(n5230), .Z(n5242) );
  AND U5206 ( .A(n5254), .B(n5255), .Z(n5230) );
  XOR U5207 ( .A(n5256), .B(n5257), .Z(n5233) );
  AND U5208 ( .A(n5258), .B(n5259), .Z(n5257) );
  XOR U5209 ( .A(n5256), .B(n5260), .Z(n5258) );
  XNOR U5210 ( .A(n5149), .B(n5238), .Z(n5240) );
  XOR U5211 ( .A(n5261), .B(n5262), .Z(n5149) );
  AND U5212 ( .A(n83), .B(n5263), .Z(n5262) );
  XNOR U5213 ( .A(n5264), .B(n5261), .Z(n5263) );
  XOR U5214 ( .A(n5265), .B(n5266), .Z(n5238) );
  AND U5215 ( .A(n5267), .B(n5268), .Z(n5266) );
  XNOR U5216 ( .A(n5265), .B(n5254), .Z(n5268) );
  IV U5217 ( .A(n5200), .Z(n5254) );
  XNOR U5218 ( .A(n5269), .B(n5247), .Z(n5200) );
  XNOR U5219 ( .A(n5270), .B(n5253), .Z(n5247) );
  XOR U5220 ( .A(n5271), .B(n5272), .Z(n5253) );
  NOR U5221 ( .A(n5273), .B(n5274), .Z(n5272) );
  XNOR U5222 ( .A(n5271), .B(n5275), .Z(n5273) );
  XNOR U5223 ( .A(n5252), .B(n5244), .Z(n5270) );
  XOR U5224 ( .A(n5276), .B(n5277), .Z(n5244) );
  AND U5225 ( .A(n5278), .B(n5279), .Z(n5277) );
  XNOR U5226 ( .A(n5276), .B(n5280), .Z(n5278) );
  XNOR U5227 ( .A(n5281), .B(n5249), .Z(n5252) );
  XOR U5228 ( .A(n5282), .B(n5283), .Z(n5249) );
  AND U5229 ( .A(n5284), .B(n5285), .Z(n5283) );
  XOR U5230 ( .A(n5282), .B(n5286), .Z(n5284) );
  XNOR U5231 ( .A(n5287), .B(n5288), .Z(n5281) );
  NOR U5232 ( .A(n5289), .B(n5290), .Z(n5288) );
  XOR U5233 ( .A(n5287), .B(n5291), .Z(n5289) );
  XNOR U5234 ( .A(n5248), .B(n5255), .Z(n5269) );
  NOR U5235 ( .A(n5212), .B(n5292), .Z(n5255) );
  XOR U5236 ( .A(n5260), .B(n5259), .Z(n5248) );
  XNOR U5237 ( .A(n5293), .B(n5256), .Z(n5259) );
  XOR U5238 ( .A(n5294), .B(n5295), .Z(n5256) );
  AND U5239 ( .A(n5296), .B(n5297), .Z(n5295) );
  XOR U5240 ( .A(n5294), .B(n5298), .Z(n5296) );
  XNOR U5241 ( .A(n5299), .B(n5300), .Z(n5293) );
  NOR U5242 ( .A(n5301), .B(n5302), .Z(n5300) );
  XNOR U5243 ( .A(n5299), .B(n5303), .Z(n5301) );
  XOR U5244 ( .A(n5304), .B(n5305), .Z(n5260) );
  NOR U5245 ( .A(n5306), .B(n5307), .Z(n5305) );
  XNOR U5246 ( .A(n5304), .B(n5308), .Z(n5306) );
  XNOR U5247 ( .A(n5197), .B(n5265), .Z(n5267) );
  XOR U5248 ( .A(n5309), .B(n5310), .Z(n5197) );
  AND U5249 ( .A(n83), .B(n5311), .Z(n5310) );
  XOR U5250 ( .A(n5312), .B(n5309), .Z(n5311) );
  AND U5251 ( .A(n5209), .B(n5212), .Z(n5265) );
  XOR U5252 ( .A(n5313), .B(n5292), .Z(n5212) );
  XNOR U5253 ( .A(p_input[1024]), .B(p_input[304]), .Z(n5292) );
  XOR U5254 ( .A(n5280), .B(n5279), .Z(n5313) );
  XNOR U5255 ( .A(n5314), .B(n5286), .Z(n5279) );
  XNOR U5256 ( .A(n5275), .B(n5274), .Z(n5286) );
  XOR U5257 ( .A(n5315), .B(n5271), .Z(n5274) );
  XOR U5258 ( .A(p_input[1034]), .B(p_input[314]), .Z(n5271) );
  XNOR U5259 ( .A(p_input[1035]), .B(p_input[315]), .Z(n5315) );
  XOR U5260 ( .A(p_input[1036]), .B(p_input[316]), .Z(n5275) );
  XNOR U5261 ( .A(n5285), .B(n5276), .Z(n5314) );
  XNOR U5262 ( .A(n3298), .B(p_input[305]), .Z(n5276) );
  XOR U5263 ( .A(n5316), .B(n5291), .Z(n5285) );
  XNOR U5264 ( .A(p_input[1039]), .B(p_input[319]), .Z(n5291) );
  XOR U5265 ( .A(n5282), .B(n5290), .Z(n5316) );
  XOR U5266 ( .A(n5317), .B(n5287), .Z(n5290) );
  XOR U5267 ( .A(p_input[1037]), .B(p_input[317]), .Z(n5287) );
  XNOR U5268 ( .A(p_input[1038]), .B(p_input[318]), .Z(n5317) );
  XOR U5269 ( .A(p_input[1033]), .B(p_input[313]), .Z(n5282) );
  XNOR U5270 ( .A(n5298), .B(n5297), .Z(n5280) );
  XNOR U5271 ( .A(n5318), .B(n5303), .Z(n5297) );
  XOR U5272 ( .A(p_input[1032]), .B(p_input[312]), .Z(n5303) );
  XOR U5273 ( .A(n5294), .B(n5302), .Z(n5318) );
  XOR U5274 ( .A(n5319), .B(n5299), .Z(n5302) );
  XOR U5275 ( .A(p_input[1030]), .B(p_input[310]), .Z(n5299) );
  XNOR U5276 ( .A(p_input[1031]), .B(p_input[311]), .Z(n5319) );
  XOR U5277 ( .A(p_input[1026]), .B(p_input[306]), .Z(n5294) );
  XNOR U5278 ( .A(n5308), .B(n5307), .Z(n5298) );
  XOR U5279 ( .A(n5320), .B(n5304), .Z(n5307) );
  XOR U5280 ( .A(p_input[1027]), .B(p_input[307]), .Z(n5304) );
  XNOR U5281 ( .A(p_input[1028]), .B(p_input[308]), .Z(n5320) );
  XOR U5282 ( .A(p_input[1029]), .B(p_input[309]), .Z(n5308) );
  XOR U5283 ( .A(n5321), .B(n5322), .Z(n5209) );
  AND U5284 ( .A(n83), .B(n5323), .Z(n5322) );
  XNOR U5285 ( .A(n5324), .B(n5321), .Z(n5323) );
  XNOR U5286 ( .A(n5325), .B(n5326), .Z(n83) );
  AND U5287 ( .A(n5327), .B(n5328), .Z(n5326) );
  XOR U5288 ( .A(n5222), .B(n5325), .Z(n5328) );
  AND U5289 ( .A(n5329), .B(n5330), .Z(n5222) );
  XNOR U5290 ( .A(n5219), .B(n5325), .Z(n5327) );
  XOR U5291 ( .A(n5331), .B(n5332), .Z(n5219) );
  AND U5292 ( .A(n87), .B(n5333), .Z(n5332) );
  XOR U5293 ( .A(n5334), .B(n5331), .Z(n5333) );
  XOR U5294 ( .A(n5335), .B(n5336), .Z(n5325) );
  AND U5295 ( .A(n5337), .B(n5338), .Z(n5336) );
  XNOR U5296 ( .A(n5335), .B(n5329), .Z(n5338) );
  IV U5297 ( .A(n5237), .Z(n5329) );
  XOR U5298 ( .A(n5339), .B(n5340), .Z(n5237) );
  XOR U5299 ( .A(n5341), .B(n5330), .Z(n5340) );
  AND U5300 ( .A(n5264), .B(n5342), .Z(n5330) );
  AND U5301 ( .A(n5343), .B(n5344), .Z(n5341) );
  XOR U5302 ( .A(n5345), .B(n5339), .Z(n5343) );
  XNOR U5303 ( .A(n5234), .B(n5335), .Z(n5337) );
  XOR U5304 ( .A(n5346), .B(n5347), .Z(n5234) );
  AND U5305 ( .A(n87), .B(n5348), .Z(n5347) );
  XOR U5306 ( .A(n5349), .B(n5346), .Z(n5348) );
  XOR U5307 ( .A(n5350), .B(n5351), .Z(n5335) );
  AND U5308 ( .A(n5352), .B(n5353), .Z(n5351) );
  XNOR U5309 ( .A(n5350), .B(n5264), .Z(n5353) );
  XOR U5310 ( .A(n5354), .B(n5344), .Z(n5264) );
  XNOR U5311 ( .A(n5355), .B(n5339), .Z(n5344) );
  XOR U5312 ( .A(n5356), .B(n5357), .Z(n5339) );
  AND U5313 ( .A(n5358), .B(n5359), .Z(n5357) );
  XOR U5314 ( .A(n5360), .B(n5356), .Z(n5358) );
  XNOR U5315 ( .A(n5361), .B(n5362), .Z(n5355) );
  AND U5316 ( .A(n5363), .B(n5364), .Z(n5362) );
  XOR U5317 ( .A(n5361), .B(n5365), .Z(n5363) );
  XNOR U5318 ( .A(n5345), .B(n5342), .Z(n5354) );
  AND U5319 ( .A(n5366), .B(n5367), .Z(n5342) );
  XOR U5320 ( .A(n5368), .B(n5369), .Z(n5345) );
  AND U5321 ( .A(n5370), .B(n5371), .Z(n5369) );
  XOR U5322 ( .A(n5368), .B(n5372), .Z(n5370) );
  XNOR U5323 ( .A(n5261), .B(n5350), .Z(n5352) );
  XOR U5324 ( .A(n5373), .B(n5374), .Z(n5261) );
  AND U5325 ( .A(n87), .B(n5375), .Z(n5374) );
  XNOR U5326 ( .A(n5376), .B(n5373), .Z(n5375) );
  XOR U5327 ( .A(n5377), .B(n5378), .Z(n5350) );
  AND U5328 ( .A(n5379), .B(n5380), .Z(n5378) );
  XNOR U5329 ( .A(n5377), .B(n5366), .Z(n5380) );
  IV U5330 ( .A(n5312), .Z(n5366) );
  XNOR U5331 ( .A(n5381), .B(n5359), .Z(n5312) );
  XNOR U5332 ( .A(n5382), .B(n5365), .Z(n5359) );
  XOR U5333 ( .A(n5383), .B(n5384), .Z(n5365) );
  NOR U5334 ( .A(n5385), .B(n5386), .Z(n5384) );
  XNOR U5335 ( .A(n5383), .B(n5387), .Z(n5385) );
  XNOR U5336 ( .A(n5364), .B(n5356), .Z(n5382) );
  XOR U5337 ( .A(n5388), .B(n5389), .Z(n5356) );
  AND U5338 ( .A(n5390), .B(n5391), .Z(n5389) );
  XNOR U5339 ( .A(n5388), .B(n5392), .Z(n5390) );
  XNOR U5340 ( .A(n5393), .B(n5361), .Z(n5364) );
  XOR U5341 ( .A(n5394), .B(n5395), .Z(n5361) );
  AND U5342 ( .A(n5396), .B(n5397), .Z(n5395) );
  XOR U5343 ( .A(n5394), .B(n5398), .Z(n5396) );
  XNOR U5344 ( .A(n5399), .B(n5400), .Z(n5393) );
  NOR U5345 ( .A(n5401), .B(n5402), .Z(n5400) );
  XOR U5346 ( .A(n5399), .B(n5403), .Z(n5401) );
  XNOR U5347 ( .A(n5360), .B(n5367), .Z(n5381) );
  NOR U5348 ( .A(n5324), .B(n5404), .Z(n5367) );
  XOR U5349 ( .A(n5372), .B(n5371), .Z(n5360) );
  XNOR U5350 ( .A(n5405), .B(n5368), .Z(n5371) );
  XOR U5351 ( .A(n5406), .B(n5407), .Z(n5368) );
  AND U5352 ( .A(n5408), .B(n5409), .Z(n5407) );
  XOR U5353 ( .A(n5406), .B(n5410), .Z(n5408) );
  XNOR U5354 ( .A(n5411), .B(n5412), .Z(n5405) );
  NOR U5355 ( .A(n5413), .B(n5414), .Z(n5412) );
  XNOR U5356 ( .A(n5411), .B(n5415), .Z(n5413) );
  XOR U5357 ( .A(n5416), .B(n5417), .Z(n5372) );
  NOR U5358 ( .A(n5418), .B(n5419), .Z(n5417) );
  XNOR U5359 ( .A(n5416), .B(n5420), .Z(n5418) );
  XNOR U5360 ( .A(n5309), .B(n5377), .Z(n5379) );
  XOR U5361 ( .A(n5421), .B(n5422), .Z(n5309) );
  AND U5362 ( .A(n87), .B(n5423), .Z(n5422) );
  XOR U5363 ( .A(n5424), .B(n5421), .Z(n5423) );
  AND U5364 ( .A(n5321), .B(n5324), .Z(n5377) );
  XOR U5365 ( .A(n5425), .B(n5404), .Z(n5324) );
  XNOR U5366 ( .A(p_input[1024]), .B(p_input[320]), .Z(n5404) );
  XOR U5367 ( .A(n5392), .B(n5391), .Z(n5425) );
  XNOR U5368 ( .A(n5426), .B(n5398), .Z(n5391) );
  XNOR U5369 ( .A(n5387), .B(n5386), .Z(n5398) );
  XOR U5370 ( .A(n5427), .B(n5383), .Z(n5386) );
  XOR U5371 ( .A(p_input[1034]), .B(p_input[330]), .Z(n5383) );
  XNOR U5372 ( .A(p_input[1035]), .B(p_input[331]), .Z(n5427) );
  XOR U5373 ( .A(p_input[1036]), .B(p_input[332]), .Z(n5387) );
  XNOR U5374 ( .A(n5397), .B(n5388), .Z(n5426) );
  XNOR U5375 ( .A(n3298), .B(p_input[321]), .Z(n5388) );
  XOR U5376 ( .A(n5428), .B(n5403), .Z(n5397) );
  XNOR U5377 ( .A(p_input[1039]), .B(p_input[335]), .Z(n5403) );
  XOR U5378 ( .A(n5394), .B(n5402), .Z(n5428) );
  XOR U5379 ( .A(n5429), .B(n5399), .Z(n5402) );
  XOR U5380 ( .A(p_input[1037]), .B(p_input[333]), .Z(n5399) );
  XNOR U5381 ( .A(p_input[1038]), .B(p_input[334]), .Z(n5429) );
  XOR U5382 ( .A(p_input[1033]), .B(p_input[329]), .Z(n5394) );
  XNOR U5383 ( .A(n5410), .B(n5409), .Z(n5392) );
  XNOR U5384 ( .A(n5430), .B(n5415), .Z(n5409) );
  XOR U5385 ( .A(p_input[1032]), .B(p_input[328]), .Z(n5415) );
  XOR U5386 ( .A(n5406), .B(n5414), .Z(n5430) );
  XOR U5387 ( .A(n5431), .B(n5411), .Z(n5414) );
  XOR U5388 ( .A(p_input[1030]), .B(p_input[326]), .Z(n5411) );
  XNOR U5389 ( .A(p_input[1031]), .B(p_input[327]), .Z(n5431) );
  XOR U5390 ( .A(p_input[1026]), .B(p_input[322]), .Z(n5406) );
  XNOR U5391 ( .A(n5420), .B(n5419), .Z(n5410) );
  XOR U5392 ( .A(n5432), .B(n5416), .Z(n5419) );
  XOR U5393 ( .A(p_input[1027]), .B(p_input[323]), .Z(n5416) );
  XNOR U5394 ( .A(p_input[1028]), .B(p_input[324]), .Z(n5432) );
  XOR U5395 ( .A(p_input[1029]), .B(p_input[325]), .Z(n5420) );
  XOR U5396 ( .A(n5433), .B(n5434), .Z(n5321) );
  AND U5397 ( .A(n87), .B(n5435), .Z(n5434) );
  XNOR U5398 ( .A(n5436), .B(n5433), .Z(n5435) );
  XNOR U5399 ( .A(n5437), .B(n5438), .Z(n87) );
  AND U5400 ( .A(n5439), .B(n5440), .Z(n5438) );
  XOR U5401 ( .A(n5334), .B(n5437), .Z(n5440) );
  AND U5402 ( .A(n5441), .B(n5442), .Z(n5334) );
  XNOR U5403 ( .A(n5331), .B(n5437), .Z(n5439) );
  XOR U5404 ( .A(n5443), .B(n5444), .Z(n5331) );
  AND U5405 ( .A(n91), .B(n5445), .Z(n5444) );
  XOR U5406 ( .A(n5446), .B(n5443), .Z(n5445) );
  XOR U5407 ( .A(n5447), .B(n5448), .Z(n5437) );
  AND U5408 ( .A(n5449), .B(n5450), .Z(n5448) );
  XNOR U5409 ( .A(n5447), .B(n5441), .Z(n5450) );
  IV U5410 ( .A(n5349), .Z(n5441) );
  XOR U5411 ( .A(n5451), .B(n5452), .Z(n5349) );
  XOR U5412 ( .A(n5453), .B(n5442), .Z(n5452) );
  AND U5413 ( .A(n5376), .B(n5454), .Z(n5442) );
  AND U5414 ( .A(n5455), .B(n5456), .Z(n5453) );
  XOR U5415 ( .A(n5457), .B(n5451), .Z(n5455) );
  XNOR U5416 ( .A(n5346), .B(n5447), .Z(n5449) );
  XOR U5417 ( .A(n5458), .B(n5459), .Z(n5346) );
  AND U5418 ( .A(n91), .B(n5460), .Z(n5459) );
  XOR U5419 ( .A(n5461), .B(n5458), .Z(n5460) );
  XOR U5420 ( .A(n5462), .B(n5463), .Z(n5447) );
  AND U5421 ( .A(n5464), .B(n5465), .Z(n5463) );
  XNOR U5422 ( .A(n5462), .B(n5376), .Z(n5465) );
  XOR U5423 ( .A(n5466), .B(n5456), .Z(n5376) );
  XNOR U5424 ( .A(n5467), .B(n5451), .Z(n5456) );
  XOR U5425 ( .A(n5468), .B(n5469), .Z(n5451) );
  AND U5426 ( .A(n5470), .B(n5471), .Z(n5469) );
  XOR U5427 ( .A(n5472), .B(n5468), .Z(n5470) );
  XNOR U5428 ( .A(n5473), .B(n5474), .Z(n5467) );
  AND U5429 ( .A(n5475), .B(n5476), .Z(n5474) );
  XOR U5430 ( .A(n5473), .B(n5477), .Z(n5475) );
  XNOR U5431 ( .A(n5457), .B(n5454), .Z(n5466) );
  AND U5432 ( .A(n5478), .B(n5479), .Z(n5454) );
  XOR U5433 ( .A(n5480), .B(n5481), .Z(n5457) );
  AND U5434 ( .A(n5482), .B(n5483), .Z(n5481) );
  XOR U5435 ( .A(n5480), .B(n5484), .Z(n5482) );
  XNOR U5436 ( .A(n5373), .B(n5462), .Z(n5464) );
  XOR U5437 ( .A(n5485), .B(n5486), .Z(n5373) );
  AND U5438 ( .A(n91), .B(n5487), .Z(n5486) );
  XNOR U5439 ( .A(n5488), .B(n5485), .Z(n5487) );
  XOR U5440 ( .A(n5489), .B(n5490), .Z(n5462) );
  AND U5441 ( .A(n5491), .B(n5492), .Z(n5490) );
  XNOR U5442 ( .A(n5489), .B(n5478), .Z(n5492) );
  IV U5443 ( .A(n5424), .Z(n5478) );
  XNOR U5444 ( .A(n5493), .B(n5471), .Z(n5424) );
  XNOR U5445 ( .A(n5494), .B(n5477), .Z(n5471) );
  XOR U5446 ( .A(n5495), .B(n5496), .Z(n5477) );
  NOR U5447 ( .A(n5497), .B(n5498), .Z(n5496) );
  XNOR U5448 ( .A(n5495), .B(n5499), .Z(n5497) );
  XNOR U5449 ( .A(n5476), .B(n5468), .Z(n5494) );
  XOR U5450 ( .A(n5500), .B(n5501), .Z(n5468) );
  AND U5451 ( .A(n5502), .B(n5503), .Z(n5501) );
  XNOR U5452 ( .A(n5500), .B(n5504), .Z(n5502) );
  XNOR U5453 ( .A(n5505), .B(n5473), .Z(n5476) );
  XOR U5454 ( .A(n5506), .B(n5507), .Z(n5473) );
  AND U5455 ( .A(n5508), .B(n5509), .Z(n5507) );
  XOR U5456 ( .A(n5506), .B(n5510), .Z(n5508) );
  XNOR U5457 ( .A(n5511), .B(n5512), .Z(n5505) );
  NOR U5458 ( .A(n5513), .B(n5514), .Z(n5512) );
  XOR U5459 ( .A(n5511), .B(n5515), .Z(n5513) );
  XNOR U5460 ( .A(n5472), .B(n5479), .Z(n5493) );
  NOR U5461 ( .A(n5436), .B(n5516), .Z(n5479) );
  XOR U5462 ( .A(n5484), .B(n5483), .Z(n5472) );
  XNOR U5463 ( .A(n5517), .B(n5480), .Z(n5483) );
  XOR U5464 ( .A(n5518), .B(n5519), .Z(n5480) );
  AND U5465 ( .A(n5520), .B(n5521), .Z(n5519) );
  XOR U5466 ( .A(n5518), .B(n5522), .Z(n5520) );
  XNOR U5467 ( .A(n5523), .B(n5524), .Z(n5517) );
  NOR U5468 ( .A(n5525), .B(n5526), .Z(n5524) );
  XNOR U5469 ( .A(n5523), .B(n5527), .Z(n5525) );
  XOR U5470 ( .A(n5528), .B(n5529), .Z(n5484) );
  NOR U5471 ( .A(n5530), .B(n5531), .Z(n5529) );
  XNOR U5472 ( .A(n5528), .B(n5532), .Z(n5530) );
  XNOR U5473 ( .A(n5421), .B(n5489), .Z(n5491) );
  XOR U5474 ( .A(n5533), .B(n5534), .Z(n5421) );
  AND U5475 ( .A(n91), .B(n5535), .Z(n5534) );
  XOR U5476 ( .A(n5536), .B(n5533), .Z(n5535) );
  AND U5477 ( .A(n5433), .B(n5436), .Z(n5489) );
  XOR U5478 ( .A(n5537), .B(n5516), .Z(n5436) );
  XNOR U5479 ( .A(p_input[1024]), .B(p_input[336]), .Z(n5516) );
  XOR U5480 ( .A(n5504), .B(n5503), .Z(n5537) );
  XNOR U5481 ( .A(n5538), .B(n5510), .Z(n5503) );
  XNOR U5482 ( .A(n5499), .B(n5498), .Z(n5510) );
  XOR U5483 ( .A(n5539), .B(n5495), .Z(n5498) );
  XOR U5484 ( .A(p_input[1034]), .B(p_input[346]), .Z(n5495) );
  XNOR U5485 ( .A(p_input[1035]), .B(p_input[347]), .Z(n5539) );
  XOR U5486 ( .A(p_input[1036]), .B(p_input[348]), .Z(n5499) );
  XNOR U5487 ( .A(n5509), .B(n5500), .Z(n5538) );
  XNOR U5488 ( .A(n3298), .B(p_input[337]), .Z(n5500) );
  XOR U5489 ( .A(n5540), .B(n5515), .Z(n5509) );
  XNOR U5490 ( .A(p_input[1039]), .B(p_input[351]), .Z(n5515) );
  XOR U5491 ( .A(n5506), .B(n5514), .Z(n5540) );
  XOR U5492 ( .A(n5541), .B(n5511), .Z(n5514) );
  XOR U5493 ( .A(p_input[1037]), .B(p_input[349]), .Z(n5511) );
  XNOR U5494 ( .A(p_input[1038]), .B(p_input[350]), .Z(n5541) );
  XOR U5495 ( .A(p_input[1033]), .B(p_input[345]), .Z(n5506) );
  XNOR U5496 ( .A(n5522), .B(n5521), .Z(n5504) );
  XNOR U5497 ( .A(n5542), .B(n5527), .Z(n5521) );
  XOR U5498 ( .A(p_input[1032]), .B(p_input[344]), .Z(n5527) );
  XOR U5499 ( .A(n5518), .B(n5526), .Z(n5542) );
  XOR U5500 ( .A(n5543), .B(n5523), .Z(n5526) );
  XOR U5501 ( .A(p_input[1030]), .B(p_input[342]), .Z(n5523) );
  XNOR U5502 ( .A(p_input[1031]), .B(p_input[343]), .Z(n5543) );
  XOR U5503 ( .A(p_input[1026]), .B(p_input[338]), .Z(n5518) );
  XNOR U5504 ( .A(n5532), .B(n5531), .Z(n5522) );
  XOR U5505 ( .A(n5544), .B(n5528), .Z(n5531) );
  XOR U5506 ( .A(p_input[1027]), .B(p_input[339]), .Z(n5528) );
  XNOR U5507 ( .A(p_input[1028]), .B(p_input[340]), .Z(n5544) );
  XOR U5508 ( .A(p_input[1029]), .B(p_input[341]), .Z(n5532) );
  XOR U5509 ( .A(n5545), .B(n5546), .Z(n5433) );
  AND U5510 ( .A(n91), .B(n5547), .Z(n5546) );
  XNOR U5511 ( .A(n5548), .B(n5545), .Z(n5547) );
  XNOR U5512 ( .A(n5549), .B(n5550), .Z(n91) );
  AND U5513 ( .A(n5551), .B(n5552), .Z(n5550) );
  XOR U5514 ( .A(n5446), .B(n5549), .Z(n5552) );
  AND U5515 ( .A(n5553), .B(n5554), .Z(n5446) );
  XNOR U5516 ( .A(n5443), .B(n5549), .Z(n5551) );
  XOR U5517 ( .A(n5555), .B(n5556), .Z(n5443) );
  AND U5518 ( .A(n95), .B(n5557), .Z(n5556) );
  XOR U5519 ( .A(n5558), .B(n5555), .Z(n5557) );
  XOR U5520 ( .A(n5559), .B(n5560), .Z(n5549) );
  AND U5521 ( .A(n5561), .B(n5562), .Z(n5560) );
  XNOR U5522 ( .A(n5559), .B(n5553), .Z(n5562) );
  IV U5523 ( .A(n5461), .Z(n5553) );
  XOR U5524 ( .A(n5563), .B(n5564), .Z(n5461) );
  XOR U5525 ( .A(n5565), .B(n5554), .Z(n5564) );
  AND U5526 ( .A(n5488), .B(n5566), .Z(n5554) );
  AND U5527 ( .A(n5567), .B(n5568), .Z(n5565) );
  XOR U5528 ( .A(n5569), .B(n5563), .Z(n5567) );
  XNOR U5529 ( .A(n5458), .B(n5559), .Z(n5561) );
  XOR U5530 ( .A(n5570), .B(n5571), .Z(n5458) );
  AND U5531 ( .A(n95), .B(n5572), .Z(n5571) );
  XOR U5532 ( .A(n5573), .B(n5570), .Z(n5572) );
  XOR U5533 ( .A(n5574), .B(n5575), .Z(n5559) );
  AND U5534 ( .A(n5576), .B(n5577), .Z(n5575) );
  XNOR U5535 ( .A(n5574), .B(n5488), .Z(n5577) );
  XOR U5536 ( .A(n5578), .B(n5568), .Z(n5488) );
  XNOR U5537 ( .A(n5579), .B(n5563), .Z(n5568) );
  XOR U5538 ( .A(n5580), .B(n5581), .Z(n5563) );
  AND U5539 ( .A(n5582), .B(n5583), .Z(n5581) );
  XOR U5540 ( .A(n5584), .B(n5580), .Z(n5582) );
  XNOR U5541 ( .A(n5585), .B(n5586), .Z(n5579) );
  AND U5542 ( .A(n5587), .B(n5588), .Z(n5586) );
  XOR U5543 ( .A(n5585), .B(n5589), .Z(n5587) );
  XNOR U5544 ( .A(n5569), .B(n5566), .Z(n5578) );
  AND U5545 ( .A(n5590), .B(n5591), .Z(n5566) );
  XOR U5546 ( .A(n5592), .B(n5593), .Z(n5569) );
  AND U5547 ( .A(n5594), .B(n5595), .Z(n5593) );
  XOR U5548 ( .A(n5592), .B(n5596), .Z(n5594) );
  XNOR U5549 ( .A(n5485), .B(n5574), .Z(n5576) );
  XOR U5550 ( .A(n5597), .B(n5598), .Z(n5485) );
  AND U5551 ( .A(n95), .B(n5599), .Z(n5598) );
  XNOR U5552 ( .A(n5600), .B(n5597), .Z(n5599) );
  XOR U5553 ( .A(n5601), .B(n5602), .Z(n5574) );
  AND U5554 ( .A(n5603), .B(n5604), .Z(n5602) );
  XNOR U5555 ( .A(n5601), .B(n5590), .Z(n5604) );
  IV U5556 ( .A(n5536), .Z(n5590) );
  XNOR U5557 ( .A(n5605), .B(n5583), .Z(n5536) );
  XNOR U5558 ( .A(n5606), .B(n5589), .Z(n5583) );
  XOR U5559 ( .A(n5607), .B(n5608), .Z(n5589) );
  NOR U5560 ( .A(n5609), .B(n5610), .Z(n5608) );
  XNOR U5561 ( .A(n5607), .B(n5611), .Z(n5609) );
  XNOR U5562 ( .A(n5588), .B(n5580), .Z(n5606) );
  XOR U5563 ( .A(n5612), .B(n5613), .Z(n5580) );
  AND U5564 ( .A(n5614), .B(n5615), .Z(n5613) );
  XNOR U5565 ( .A(n5612), .B(n5616), .Z(n5614) );
  XNOR U5566 ( .A(n5617), .B(n5585), .Z(n5588) );
  XOR U5567 ( .A(n5618), .B(n5619), .Z(n5585) );
  AND U5568 ( .A(n5620), .B(n5621), .Z(n5619) );
  XOR U5569 ( .A(n5618), .B(n5622), .Z(n5620) );
  XNOR U5570 ( .A(n5623), .B(n5624), .Z(n5617) );
  NOR U5571 ( .A(n5625), .B(n5626), .Z(n5624) );
  XOR U5572 ( .A(n5623), .B(n5627), .Z(n5625) );
  XNOR U5573 ( .A(n5584), .B(n5591), .Z(n5605) );
  NOR U5574 ( .A(n5548), .B(n5628), .Z(n5591) );
  XOR U5575 ( .A(n5596), .B(n5595), .Z(n5584) );
  XNOR U5576 ( .A(n5629), .B(n5592), .Z(n5595) );
  XOR U5577 ( .A(n5630), .B(n5631), .Z(n5592) );
  AND U5578 ( .A(n5632), .B(n5633), .Z(n5631) );
  XOR U5579 ( .A(n5630), .B(n5634), .Z(n5632) );
  XNOR U5580 ( .A(n5635), .B(n5636), .Z(n5629) );
  NOR U5581 ( .A(n5637), .B(n5638), .Z(n5636) );
  XNOR U5582 ( .A(n5635), .B(n5639), .Z(n5637) );
  XOR U5583 ( .A(n5640), .B(n5641), .Z(n5596) );
  NOR U5584 ( .A(n5642), .B(n5643), .Z(n5641) );
  XNOR U5585 ( .A(n5640), .B(n5644), .Z(n5642) );
  XNOR U5586 ( .A(n5533), .B(n5601), .Z(n5603) );
  XOR U5587 ( .A(n5645), .B(n5646), .Z(n5533) );
  AND U5588 ( .A(n95), .B(n5647), .Z(n5646) );
  XOR U5589 ( .A(n5648), .B(n5645), .Z(n5647) );
  AND U5590 ( .A(n5545), .B(n5548), .Z(n5601) );
  XOR U5591 ( .A(n5649), .B(n5628), .Z(n5548) );
  XNOR U5592 ( .A(p_input[1024]), .B(p_input[352]), .Z(n5628) );
  XOR U5593 ( .A(n5616), .B(n5615), .Z(n5649) );
  XNOR U5594 ( .A(n5650), .B(n5622), .Z(n5615) );
  XNOR U5595 ( .A(n5611), .B(n5610), .Z(n5622) );
  XOR U5596 ( .A(n5651), .B(n5607), .Z(n5610) );
  XOR U5597 ( .A(p_input[1034]), .B(p_input[362]), .Z(n5607) );
  XNOR U5598 ( .A(p_input[1035]), .B(p_input[363]), .Z(n5651) );
  XOR U5599 ( .A(p_input[1036]), .B(p_input[364]), .Z(n5611) );
  XNOR U5600 ( .A(n5621), .B(n5612), .Z(n5650) );
  XNOR U5601 ( .A(n3298), .B(p_input[353]), .Z(n5612) );
  XOR U5602 ( .A(n5652), .B(n5627), .Z(n5621) );
  XNOR U5603 ( .A(p_input[1039]), .B(p_input[367]), .Z(n5627) );
  XOR U5604 ( .A(n5618), .B(n5626), .Z(n5652) );
  XOR U5605 ( .A(n5653), .B(n5623), .Z(n5626) );
  XOR U5606 ( .A(p_input[1037]), .B(p_input[365]), .Z(n5623) );
  XNOR U5607 ( .A(p_input[1038]), .B(p_input[366]), .Z(n5653) );
  XOR U5608 ( .A(p_input[1033]), .B(p_input[361]), .Z(n5618) );
  XNOR U5609 ( .A(n5634), .B(n5633), .Z(n5616) );
  XNOR U5610 ( .A(n5654), .B(n5639), .Z(n5633) );
  XOR U5611 ( .A(p_input[1032]), .B(p_input[360]), .Z(n5639) );
  XOR U5612 ( .A(n5630), .B(n5638), .Z(n5654) );
  XOR U5613 ( .A(n5655), .B(n5635), .Z(n5638) );
  XOR U5614 ( .A(p_input[1030]), .B(p_input[358]), .Z(n5635) );
  XNOR U5615 ( .A(p_input[1031]), .B(p_input[359]), .Z(n5655) );
  XOR U5616 ( .A(p_input[1026]), .B(p_input[354]), .Z(n5630) );
  XNOR U5617 ( .A(n5644), .B(n5643), .Z(n5634) );
  XOR U5618 ( .A(n5656), .B(n5640), .Z(n5643) );
  XOR U5619 ( .A(p_input[1027]), .B(p_input[355]), .Z(n5640) );
  XNOR U5620 ( .A(p_input[1028]), .B(p_input[356]), .Z(n5656) );
  XOR U5621 ( .A(p_input[1029]), .B(p_input[357]), .Z(n5644) );
  XOR U5622 ( .A(n5657), .B(n5658), .Z(n5545) );
  AND U5623 ( .A(n95), .B(n5659), .Z(n5658) );
  XNOR U5624 ( .A(n5660), .B(n5657), .Z(n5659) );
  XNOR U5625 ( .A(n5661), .B(n5662), .Z(n95) );
  AND U5626 ( .A(n5663), .B(n5664), .Z(n5662) );
  XOR U5627 ( .A(n5558), .B(n5661), .Z(n5664) );
  AND U5628 ( .A(n5665), .B(n5666), .Z(n5558) );
  XNOR U5629 ( .A(n5555), .B(n5661), .Z(n5663) );
  XOR U5630 ( .A(n5667), .B(n5668), .Z(n5555) );
  AND U5631 ( .A(n99), .B(n5669), .Z(n5668) );
  XOR U5632 ( .A(n5670), .B(n5667), .Z(n5669) );
  XOR U5633 ( .A(n5671), .B(n5672), .Z(n5661) );
  AND U5634 ( .A(n5673), .B(n5674), .Z(n5672) );
  XNOR U5635 ( .A(n5671), .B(n5665), .Z(n5674) );
  IV U5636 ( .A(n5573), .Z(n5665) );
  XOR U5637 ( .A(n5675), .B(n5676), .Z(n5573) );
  XOR U5638 ( .A(n5677), .B(n5666), .Z(n5676) );
  AND U5639 ( .A(n5600), .B(n5678), .Z(n5666) );
  AND U5640 ( .A(n5679), .B(n5680), .Z(n5677) );
  XOR U5641 ( .A(n5681), .B(n5675), .Z(n5679) );
  XNOR U5642 ( .A(n5570), .B(n5671), .Z(n5673) );
  XOR U5643 ( .A(n5682), .B(n5683), .Z(n5570) );
  AND U5644 ( .A(n99), .B(n5684), .Z(n5683) );
  XOR U5645 ( .A(n5685), .B(n5682), .Z(n5684) );
  XOR U5646 ( .A(n5686), .B(n5687), .Z(n5671) );
  AND U5647 ( .A(n5688), .B(n5689), .Z(n5687) );
  XNOR U5648 ( .A(n5686), .B(n5600), .Z(n5689) );
  XOR U5649 ( .A(n5690), .B(n5680), .Z(n5600) );
  XNOR U5650 ( .A(n5691), .B(n5675), .Z(n5680) );
  XOR U5651 ( .A(n5692), .B(n5693), .Z(n5675) );
  AND U5652 ( .A(n5694), .B(n5695), .Z(n5693) );
  XOR U5653 ( .A(n5696), .B(n5692), .Z(n5694) );
  XNOR U5654 ( .A(n5697), .B(n5698), .Z(n5691) );
  AND U5655 ( .A(n5699), .B(n5700), .Z(n5698) );
  XOR U5656 ( .A(n5697), .B(n5701), .Z(n5699) );
  XNOR U5657 ( .A(n5681), .B(n5678), .Z(n5690) );
  AND U5658 ( .A(n5702), .B(n5703), .Z(n5678) );
  XOR U5659 ( .A(n5704), .B(n5705), .Z(n5681) );
  AND U5660 ( .A(n5706), .B(n5707), .Z(n5705) );
  XOR U5661 ( .A(n5704), .B(n5708), .Z(n5706) );
  XNOR U5662 ( .A(n5597), .B(n5686), .Z(n5688) );
  XOR U5663 ( .A(n5709), .B(n5710), .Z(n5597) );
  AND U5664 ( .A(n99), .B(n5711), .Z(n5710) );
  XNOR U5665 ( .A(n5712), .B(n5709), .Z(n5711) );
  XOR U5666 ( .A(n5713), .B(n5714), .Z(n5686) );
  AND U5667 ( .A(n5715), .B(n5716), .Z(n5714) );
  XNOR U5668 ( .A(n5713), .B(n5702), .Z(n5716) );
  IV U5669 ( .A(n5648), .Z(n5702) );
  XNOR U5670 ( .A(n5717), .B(n5695), .Z(n5648) );
  XNOR U5671 ( .A(n5718), .B(n5701), .Z(n5695) );
  XOR U5672 ( .A(n5719), .B(n5720), .Z(n5701) );
  NOR U5673 ( .A(n5721), .B(n5722), .Z(n5720) );
  XNOR U5674 ( .A(n5719), .B(n5723), .Z(n5721) );
  XNOR U5675 ( .A(n5700), .B(n5692), .Z(n5718) );
  XOR U5676 ( .A(n5724), .B(n5725), .Z(n5692) );
  AND U5677 ( .A(n5726), .B(n5727), .Z(n5725) );
  XNOR U5678 ( .A(n5724), .B(n5728), .Z(n5726) );
  XNOR U5679 ( .A(n5729), .B(n5697), .Z(n5700) );
  XOR U5680 ( .A(n5730), .B(n5731), .Z(n5697) );
  AND U5681 ( .A(n5732), .B(n5733), .Z(n5731) );
  XOR U5682 ( .A(n5730), .B(n5734), .Z(n5732) );
  XNOR U5683 ( .A(n5735), .B(n5736), .Z(n5729) );
  NOR U5684 ( .A(n5737), .B(n5738), .Z(n5736) );
  XOR U5685 ( .A(n5735), .B(n5739), .Z(n5737) );
  XNOR U5686 ( .A(n5696), .B(n5703), .Z(n5717) );
  NOR U5687 ( .A(n5660), .B(n5740), .Z(n5703) );
  XOR U5688 ( .A(n5708), .B(n5707), .Z(n5696) );
  XNOR U5689 ( .A(n5741), .B(n5704), .Z(n5707) );
  XOR U5690 ( .A(n5742), .B(n5743), .Z(n5704) );
  AND U5691 ( .A(n5744), .B(n5745), .Z(n5743) );
  XOR U5692 ( .A(n5742), .B(n5746), .Z(n5744) );
  XNOR U5693 ( .A(n5747), .B(n5748), .Z(n5741) );
  NOR U5694 ( .A(n5749), .B(n5750), .Z(n5748) );
  XNOR U5695 ( .A(n5747), .B(n5751), .Z(n5749) );
  XOR U5696 ( .A(n5752), .B(n5753), .Z(n5708) );
  NOR U5697 ( .A(n5754), .B(n5755), .Z(n5753) );
  XNOR U5698 ( .A(n5752), .B(n5756), .Z(n5754) );
  XNOR U5699 ( .A(n5645), .B(n5713), .Z(n5715) );
  XOR U5700 ( .A(n5757), .B(n5758), .Z(n5645) );
  AND U5701 ( .A(n99), .B(n5759), .Z(n5758) );
  XOR U5702 ( .A(n5760), .B(n5757), .Z(n5759) );
  AND U5703 ( .A(n5657), .B(n5660), .Z(n5713) );
  XOR U5704 ( .A(n5761), .B(n5740), .Z(n5660) );
  XNOR U5705 ( .A(p_input[1024]), .B(p_input[368]), .Z(n5740) );
  XOR U5706 ( .A(n5728), .B(n5727), .Z(n5761) );
  XNOR U5707 ( .A(n5762), .B(n5734), .Z(n5727) );
  XNOR U5708 ( .A(n5723), .B(n5722), .Z(n5734) );
  XOR U5709 ( .A(n5763), .B(n5719), .Z(n5722) );
  XOR U5710 ( .A(p_input[1034]), .B(p_input[378]), .Z(n5719) );
  XNOR U5711 ( .A(p_input[1035]), .B(p_input[379]), .Z(n5763) );
  XOR U5712 ( .A(p_input[1036]), .B(p_input[380]), .Z(n5723) );
  XNOR U5713 ( .A(n5733), .B(n5724), .Z(n5762) );
  XNOR U5714 ( .A(n3298), .B(p_input[369]), .Z(n5724) );
  XOR U5715 ( .A(n5764), .B(n5739), .Z(n5733) );
  XNOR U5716 ( .A(p_input[1039]), .B(p_input[383]), .Z(n5739) );
  XOR U5717 ( .A(n5730), .B(n5738), .Z(n5764) );
  XOR U5718 ( .A(n5765), .B(n5735), .Z(n5738) );
  XOR U5719 ( .A(p_input[1037]), .B(p_input[381]), .Z(n5735) );
  XNOR U5720 ( .A(p_input[1038]), .B(p_input[382]), .Z(n5765) );
  XOR U5721 ( .A(p_input[1033]), .B(p_input[377]), .Z(n5730) );
  XNOR U5722 ( .A(n5746), .B(n5745), .Z(n5728) );
  XNOR U5723 ( .A(n5766), .B(n5751), .Z(n5745) );
  XOR U5724 ( .A(p_input[1032]), .B(p_input[376]), .Z(n5751) );
  XOR U5725 ( .A(n5742), .B(n5750), .Z(n5766) );
  XOR U5726 ( .A(n5767), .B(n5747), .Z(n5750) );
  XOR U5727 ( .A(p_input[1030]), .B(p_input[374]), .Z(n5747) );
  XNOR U5728 ( .A(p_input[1031]), .B(p_input[375]), .Z(n5767) );
  XOR U5729 ( .A(p_input[1026]), .B(p_input[370]), .Z(n5742) );
  XNOR U5730 ( .A(n5756), .B(n5755), .Z(n5746) );
  XOR U5731 ( .A(n5768), .B(n5752), .Z(n5755) );
  XOR U5732 ( .A(p_input[1027]), .B(p_input[371]), .Z(n5752) );
  XNOR U5733 ( .A(p_input[1028]), .B(p_input[372]), .Z(n5768) );
  XOR U5734 ( .A(p_input[1029]), .B(p_input[373]), .Z(n5756) );
  XOR U5735 ( .A(n5769), .B(n5770), .Z(n5657) );
  AND U5736 ( .A(n99), .B(n5771), .Z(n5770) );
  XNOR U5737 ( .A(n5772), .B(n5769), .Z(n5771) );
  XNOR U5738 ( .A(n5773), .B(n5774), .Z(n99) );
  AND U5739 ( .A(n5775), .B(n5776), .Z(n5774) );
  XOR U5740 ( .A(n5670), .B(n5773), .Z(n5776) );
  AND U5741 ( .A(n5777), .B(n5778), .Z(n5670) );
  XNOR U5742 ( .A(n5667), .B(n5773), .Z(n5775) );
  XOR U5743 ( .A(n5779), .B(n5780), .Z(n5667) );
  AND U5744 ( .A(n103), .B(n5781), .Z(n5780) );
  XOR U5745 ( .A(n5782), .B(n5779), .Z(n5781) );
  XOR U5746 ( .A(n5783), .B(n5784), .Z(n5773) );
  AND U5747 ( .A(n5785), .B(n5786), .Z(n5784) );
  XNOR U5748 ( .A(n5783), .B(n5777), .Z(n5786) );
  IV U5749 ( .A(n5685), .Z(n5777) );
  XOR U5750 ( .A(n5787), .B(n5788), .Z(n5685) );
  XOR U5751 ( .A(n5789), .B(n5778), .Z(n5788) );
  AND U5752 ( .A(n5712), .B(n5790), .Z(n5778) );
  AND U5753 ( .A(n5791), .B(n5792), .Z(n5789) );
  XOR U5754 ( .A(n5793), .B(n5787), .Z(n5791) );
  XNOR U5755 ( .A(n5682), .B(n5783), .Z(n5785) );
  XOR U5756 ( .A(n5794), .B(n5795), .Z(n5682) );
  AND U5757 ( .A(n103), .B(n5796), .Z(n5795) );
  XOR U5758 ( .A(n5797), .B(n5794), .Z(n5796) );
  XOR U5759 ( .A(n5798), .B(n5799), .Z(n5783) );
  AND U5760 ( .A(n5800), .B(n5801), .Z(n5799) );
  XNOR U5761 ( .A(n5798), .B(n5712), .Z(n5801) );
  XOR U5762 ( .A(n5802), .B(n5792), .Z(n5712) );
  XNOR U5763 ( .A(n5803), .B(n5787), .Z(n5792) );
  XOR U5764 ( .A(n5804), .B(n5805), .Z(n5787) );
  AND U5765 ( .A(n5806), .B(n5807), .Z(n5805) );
  XOR U5766 ( .A(n5808), .B(n5804), .Z(n5806) );
  XNOR U5767 ( .A(n5809), .B(n5810), .Z(n5803) );
  AND U5768 ( .A(n5811), .B(n5812), .Z(n5810) );
  XOR U5769 ( .A(n5809), .B(n5813), .Z(n5811) );
  XNOR U5770 ( .A(n5793), .B(n5790), .Z(n5802) );
  AND U5771 ( .A(n5814), .B(n5815), .Z(n5790) );
  XOR U5772 ( .A(n5816), .B(n5817), .Z(n5793) );
  AND U5773 ( .A(n5818), .B(n5819), .Z(n5817) );
  XOR U5774 ( .A(n5816), .B(n5820), .Z(n5818) );
  XNOR U5775 ( .A(n5709), .B(n5798), .Z(n5800) );
  XOR U5776 ( .A(n5821), .B(n5822), .Z(n5709) );
  AND U5777 ( .A(n103), .B(n5823), .Z(n5822) );
  XNOR U5778 ( .A(n5824), .B(n5821), .Z(n5823) );
  XOR U5779 ( .A(n5825), .B(n5826), .Z(n5798) );
  AND U5780 ( .A(n5827), .B(n5828), .Z(n5826) );
  XNOR U5781 ( .A(n5825), .B(n5814), .Z(n5828) );
  IV U5782 ( .A(n5760), .Z(n5814) );
  XNOR U5783 ( .A(n5829), .B(n5807), .Z(n5760) );
  XNOR U5784 ( .A(n5830), .B(n5813), .Z(n5807) );
  XOR U5785 ( .A(n5831), .B(n5832), .Z(n5813) );
  NOR U5786 ( .A(n5833), .B(n5834), .Z(n5832) );
  XNOR U5787 ( .A(n5831), .B(n5835), .Z(n5833) );
  XNOR U5788 ( .A(n5812), .B(n5804), .Z(n5830) );
  XOR U5789 ( .A(n5836), .B(n5837), .Z(n5804) );
  AND U5790 ( .A(n5838), .B(n5839), .Z(n5837) );
  XNOR U5791 ( .A(n5836), .B(n5840), .Z(n5838) );
  XNOR U5792 ( .A(n5841), .B(n5809), .Z(n5812) );
  XOR U5793 ( .A(n5842), .B(n5843), .Z(n5809) );
  AND U5794 ( .A(n5844), .B(n5845), .Z(n5843) );
  XOR U5795 ( .A(n5842), .B(n5846), .Z(n5844) );
  XNOR U5796 ( .A(n5847), .B(n5848), .Z(n5841) );
  NOR U5797 ( .A(n5849), .B(n5850), .Z(n5848) );
  XOR U5798 ( .A(n5847), .B(n5851), .Z(n5849) );
  XNOR U5799 ( .A(n5808), .B(n5815), .Z(n5829) );
  NOR U5800 ( .A(n5772), .B(n5852), .Z(n5815) );
  XOR U5801 ( .A(n5820), .B(n5819), .Z(n5808) );
  XNOR U5802 ( .A(n5853), .B(n5816), .Z(n5819) );
  XOR U5803 ( .A(n5854), .B(n5855), .Z(n5816) );
  AND U5804 ( .A(n5856), .B(n5857), .Z(n5855) );
  XOR U5805 ( .A(n5854), .B(n5858), .Z(n5856) );
  XNOR U5806 ( .A(n5859), .B(n5860), .Z(n5853) );
  NOR U5807 ( .A(n5861), .B(n5862), .Z(n5860) );
  XNOR U5808 ( .A(n5859), .B(n5863), .Z(n5861) );
  XOR U5809 ( .A(n5864), .B(n5865), .Z(n5820) );
  NOR U5810 ( .A(n5866), .B(n5867), .Z(n5865) );
  XNOR U5811 ( .A(n5864), .B(n5868), .Z(n5866) );
  XNOR U5812 ( .A(n5757), .B(n5825), .Z(n5827) );
  XOR U5813 ( .A(n5869), .B(n5870), .Z(n5757) );
  AND U5814 ( .A(n103), .B(n5871), .Z(n5870) );
  XOR U5815 ( .A(n5872), .B(n5869), .Z(n5871) );
  AND U5816 ( .A(n5769), .B(n5772), .Z(n5825) );
  XOR U5817 ( .A(n5873), .B(n5852), .Z(n5772) );
  XNOR U5818 ( .A(p_input[1024]), .B(p_input[384]), .Z(n5852) );
  XOR U5819 ( .A(n5840), .B(n5839), .Z(n5873) );
  XNOR U5820 ( .A(n5874), .B(n5846), .Z(n5839) );
  XNOR U5821 ( .A(n5835), .B(n5834), .Z(n5846) );
  XOR U5822 ( .A(n5875), .B(n5831), .Z(n5834) );
  XOR U5823 ( .A(p_input[1034]), .B(p_input[394]), .Z(n5831) );
  XNOR U5824 ( .A(p_input[1035]), .B(p_input[395]), .Z(n5875) );
  XOR U5825 ( .A(p_input[1036]), .B(p_input[396]), .Z(n5835) );
  XNOR U5826 ( .A(n5845), .B(n5836), .Z(n5874) );
  XNOR U5827 ( .A(n3298), .B(p_input[385]), .Z(n5836) );
  XOR U5828 ( .A(n5876), .B(n5851), .Z(n5845) );
  XNOR U5829 ( .A(p_input[1039]), .B(p_input[399]), .Z(n5851) );
  XOR U5830 ( .A(n5842), .B(n5850), .Z(n5876) );
  XOR U5831 ( .A(n5877), .B(n5847), .Z(n5850) );
  XOR U5832 ( .A(p_input[1037]), .B(p_input[397]), .Z(n5847) );
  XNOR U5833 ( .A(p_input[1038]), .B(p_input[398]), .Z(n5877) );
  XOR U5834 ( .A(p_input[1033]), .B(p_input[393]), .Z(n5842) );
  XNOR U5835 ( .A(n5858), .B(n5857), .Z(n5840) );
  XNOR U5836 ( .A(n5878), .B(n5863), .Z(n5857) );
  XOR U5837 ( .A(p_input[1032]), .B(p_input[392]), .Z(n5863) );
  XOR U5838 ( .A(n5854), .B(n5862), .Z(n5878) );
  XOR U5839 ( .A(n5879), .B(n5859), .Z(n5862) );
  XOR U5840 ( .A(p_input[1030]), .B(p_input[390]), .Z(n5859) );
  XNOR U5841 ( .A(p_input[1031]), .B(p_input[391]), .Z(n5879) );
  XOR U5842 ( .A(p_input[1026]), .B(p_input[386]), .Z(n5854) );
  XNOR U5843 ( .A(n5868), .B(n5867), .Z(n5858) );
  XOR U5844 ( .A(n5880), .B(n5864), .Z(n5867) );
  XOR U5845 ( .A(p_input[1027]), .B(p_input[387]), .Z(n5864) );
  XNOR U5846 ( .A(p_input[1028]), .B(p_input[388]), .Z(n5880) );
  XOR U5847 ( .A(p_input[1029]), .B(p_input[389]), .Z(n5868) );
  XOR U5848 ( .A(n5881), .B(n5882), .Z(n5769) );
  AND U5849 ( .A(n103), .B(n5883), .Z(n5882) );
  XNOR U5850 ( .A(n5884), .B(n5881), .Z(n5883) );
  XNOR U5851 ( .A(n5885), .B(n5886), .Z(n103) );
  AND U5852 ( .A(n5887), .B(n5888), .Z(n5886) );
  XOR U5853 ( .A(n5782), .B(n5885), .Z(n5888) );
  AND U5854 ( .A(n5889), .B(n5890), .Z(n5782) );
  XNOR U5855 ( .A(n5779), .B(n5885), .Z(n5887) );
  XOR U5856 ( .A(n5891), .B(n5892), .Z(n5779) );
  AND U5857 ( .A(n107), .B(n5893), .Z(n5892) );
  XOR U5858 ( .A(n5894), .B(n5891), .Z(n5893) );
  XOR U5859 ( .A(n5895), .B(n5896), .Z(n5885) );
  AND U5860 ( .A(n5897), .B(n5898), .Z(n5896) );
  XNOR U5861 ( .A(n5895), .B(n5889), .Z(n5898) );
  IV U5862 ( .A(n5797), .Z(n5889) );
  XOR U5863 ( .A(n5899), .B(n5900), .Z(n5797) );
  XOR U5864 ( .A(n5901), .B(n5890), .Z(n5900) );
  AND U5865 ( .A(n5824), .B(n5902), .Z(n5890) );
  AND U5866 ( .A(n5903), .B(n5904), .Z(n5901) );
  XOR U5867 ( .A(n5905), .B(n5899), .Z(n5903) );
  XNOR U5868 ( .A(n5794), .B(n5895), .Z(n5897) );
  XOR U5869 ( .A(n5906), .B(n5907), .Z(n5794) );
  AND U5870 ( .A(n107), .B(n5908), .Z(n5907) );
  XOR U5871 ( .A(n5909), .B(n5906), .Z(n5908) );
  XOR U5872 ( .A(n5910), .B(n5911), .Z(n5895) );
  AND U5873 ( .A(n5912), .B(n5913), .Z(n5911) );
  XNOR U5874 ( .A(n5910), .B(n5824), .Z(n5913) );
  XOR U5875 ( .A(n5914), .B(n5904), .Z(n5824) );
  XNOR U5876 ( .A(n5915), .B(n5899), .Z(n5904) );
  XOR U5877 ( .A(n5916), .B(n5917), .Z(n5899) );
  AND U5878 ( .A(n5918), .B(n5919), .Z(n5917) );
  XOR U5879 ( .A(n5920), .B(n5916), .Z(n5918) );
  XNOR U5880 ( .A(n5921), .B(n5922), .Z(n5915) );
  AND U5881 ( .A(n5923), .B(n5924), .Z(n5922) );
  XOR U5882 ( .A(n5921), .B(n5925), .Z(n5923) );
  XNOR U5883 ( .A(n5905), .B(n5902), .Z(n5914) );
  AND U5884 ( .A(n5926), .B(n5927), .Z(n5902) );
  XOR U5885 ( .A(n5928), .B(n5929), .Z(n5905) );
  AND U5886 ( .A(n5930), .B(n5931), .Z(n5929) );
  XOR U5887 ( .A(n5928), .B(n5932), .Z(n5930) );
  XNOR U5888 ( .A(n5821), .B(n5910), .Z(n5912) );
  XOR U5889 ( .A(n5933), .B(n5934), .Z(n5821) );
  AND U5890 ( .A(n107), .B(n5935), .Z(n5934) );
  XNOR U5891 ( .A(n5936), .B(n5933), .Z(n5935) );
  XOR U5892 ( .A(n5937), .B(n5938), .Z(n5910) );
  AND U5893 ( .A(n5939), .B(n5940), .Z(n5938) );
  XNOR U5894 ( .A(n5937), .B(n5926), .Z(n5940) );
  IV U5895 ( .A(n5872), .Z(n5926) );
  XNOR U5896 ( .A(n5941), .B(n5919), .Z(n5872) );
  XNOR U5897 ( .A(n5942), .B(n5925), .Z(n5919) );
  XOR U5898 ( .A(n5943), .B(n5944), .Z(n5925) );
  NOR U5899 ( .A(n5945), .B(n5946), .Z(n5944) );
  XNOR U5900 ( .A(n5943), .B(n5947), .Z(n5945) );
  XNOR U5901 ( .A(n5924), .B(n5916), .Z(n5942) );
  XOR U5902 ( .A(n5948), .B(n5949), .Z(n5916) );
  AND U5903 ( .A(n5950), .B(n5951), .Z(n5949) );
  XNOR U5904 ( .A(n5948), .B(n5952), .Z(n5950) );
  XNOR U5905 ( .A(n5953), .B(n5921), .Z(n5924) );
  XOR U5906 ( .A(n5954), .B(n5955), .Z(n5921) );
  AND U5907 ( .A(n5956), .B(n5957), .Z(n5955) );
  XOR U5908 ( .A(n5954), .B(n5958), .Z(n5956) );
  XNOR U5909 ( .A(n5959), .B(n5960), .Z(n5953) );
  NOR U5910 ( .A(n5961), .B(n5962), .Z(n5960) );
  XOR U5911 ( .A(n5959), .B(n5963), .Z(n5961) );
  XNOR U5912 ( .A(n5920), .B(n5927), .Z(n5941) );
  NOR U5913 ( .A(n5884), .B(n5964), .Z(n5927) );
  XOR U5914 ( .A(n5932), .B(n5931), .Z(n5920) );
  XNOR U5915 ( .A(n5965), .B(n5928), .Z(n5931) );
  XOR U5916 ( .A(n5966), .B(n5967), .Z(n5928) );
  AND U5917 ( .A(n5968), .B(n5969), .Z(n5967) );
  XOR U5918 ( .A(n5966), .B(n5970), .Z(n5968) );
  XNOR U5919 ( .A(n5971), .B(n5972), .Z(n5965) );
  NOR U5920 ( .A(n5973), .B(n5974), .Z(n5972) );
  XNOR U5921 ( .A(n5971), .B(n5975), .Z(n5973) );
  XOR U5922 ( .A(n5976), .B(n5977), .Z(n5932) );
  NOR U5923 ( .A(n5978), .B(n5979), .Z(n5977) );
  XNOR U5924 ( .A(n5976), .B(n5980), .Z(n5978) );
  XNOR U5925 ( .A(n5869), .B(n5937), .Z(n5939) );
  XOR U5926 ( .A(n5981), .B(n5982), .Z(n5869) );
  AND U5927 ( .A(n107), .B(n5983), .Z(n5982) );
  XOR U5928 ( .A(n5984), .B(n5981), .Z(n5983) );
  AND U5929 ( .A(n5881), .B(n5884), .Z(n5937) );
  XOR U5930 ( .A(n5985), .B(n5964), .Z(n5884) );
  XNOR U5931 ( .A(p_input[1024]), .B(p_input[400]), .Z(n5964) );
  XOR U5932 ( .A(n5952), .B(n5951), .Z(n5985) );
  XNOR U5933 ( .A(n5986), .B(n5958), .Z(n5951) );
  XNOR U5934 ( .A(n5947), .B(n5946), .Z(n5958) );
  XOR U5935 ( .A(n5987), .B(n5943), .Z(n5946) );
  XOR U5936 ( .A(p_input[1034]), .B(p_input[410]), .Z(n5943) );
  XNOR U5937 ( .A(p_input[1035]), .B(p_input[411]), .Z(n5987) );
  XOR U5938 ( .A(p_input[1036]), .B(p_input[412]), .Z(n5947) );
  XNOR U5939 ( .A(n5957), .B(n5948), .Z(n5986) );
  XNOR U5940 ( .A(n3298), .B(p_input[401]), .Z(n5948) );
  XOR U5941 ( .A(n5988), .B(n5963), .Z(n5957) );
  XNOR U5942 ( .A(p_input[1039]), .B(p_input[415]), .Z(n5963) );
  XOR U5943 ( .A(n5954), .B(n5962), .Z(n5988) );
  XOR U5944 ( .A(n5989), .B(n5959), .Z(n5962) );
  XOR U5945 ( .A(p_input[1037]), .B(p_input[413]), .Z(n5959) );
  XNOR U5946 ( .A(p_input[1038]), .B(p_input[414]), .Z(n5989) );
  XOR U5947 ( .A(p_input[1033]), .B(p_input[409]), .Z(n5954) );
  XNOR U5948 ( .A(n5970), .B(n5969), .Z(n5952) );
  XNOR U5949 ( .A(n5990), .B(n5975), .Z(n5969) );
  XOR U5950 ( .A(p_input[1032]), .B(p_input[408]), .Z(n5975) );
  XOR U5951 ( .A(n5966), .B(n5974), .Z(n5990) );
  XOR U5952 ( .A(n5991), .B(n5971), .Z(n5974) );
  XOR U5953 ( .A(p_input[1030]), .B(p_input[406]), .Z(n5971) );
  XNOR U5954 ( .A(p_input[1031]), .B(p_input[407]), .Z(n5991) );
  XOR U5955 ( .A(p_input[1026]), .B(p_input[402]), .Z(n5966) );
  XNOR U5956 ( .A(n5980), .B(n5979), .Z(n5970) );
  XOR U5957 ( .A(n5992), .B(n5976), .Z(n5979) );
  XOR U5958 ( .A(p_input[1027]), .B(p_input[403]), .Z(n5976) );
  XNOR U5959 ( .A(p_input[1028]), .B(p_input[404]), .Z(n5992) );
  XOR U5960 ( .A(p_input[1029]), .B(p_input[405]), .Z(n5980) );
  XOR U5961 ( .A(n5993), .B(n5994), .Z(n5881) );
  AND U5962 ( .A(n107), .B(n5995), .Z(n5994) );
  XNOR U5963 ( .A(n5996), .B(n5993), .Z(n5995) );
  XNOR U5964 ( .A(n5997), .B(n5998), .Z(n107) );
  AND U5965 ( .A(n5999), .B(n6000), .Z(n5998) );
  XOR U5966 ( .A(n5894), .B(n5997), .Z(n6000) );
  AND U5967 ( .A(n6001), .B(n6002), .Z(n5894) );
  XNOR U5968 ( .A(n5891), .B(n5997), .Z(n5999) );
  XOR U5969 ( .A(n6003), .B(n6004), .Z(n5891) );
  AND U5970 ( .A(n111), .B(n6005), .Z(n6004) );
  XOR U5971 ( .A(n6006), .B(n6003), .Z(n6005) );
  XOR U5972 ( .A(n6007), .B(n6008), .Z(n5997) );
  AND U5973 ( .A(n6009), .B(n6010), .Z(n6008) );
  XNOR U5974 ( .A(n6007), .B(n6001), .Z(n6010) );
  IV U5975 ( .A(n5909), .Z(n6001) );
  XOR U5976 ( .A(n6011), .B(n6012), .Z(n5909) );
  XOR U5977 ( .A(n6013), .B(n6002), .Z(n6012) );
  AND U5978 ( .A(n5936), .B(n6014), .Z(n6002) );
  AND U5979 ( .A(n6015), .B(n6016), .Z(n6013) );
  XOR U5980 ( .A(n6017), .B(n6011), .Z(n6015) );
  XNOR U5981 ( .A(n5906), .B(n6007), .Z(n6009) );
  XOR U5982 ( .A(n6018), .B(n6019), .Z(n5906) );
  AND U5983 ( .A(n111), .B(n6020), .Z(n6019) );
  XOR U5984 ( .A(n6021), .B(n6018), .Z(n6020) );
  XOR U5985 ( .A(n6022), .B(n6023), .Z(n6007) );
  AND U5986 ( .A(n6024), .B(n6025), .Z(n6023) );
  XNOR U5987 ( .A(n6022), .B(n5936), .Z(n6025) );
  XOR U5988 ( .A(n6026), .B(n6016), .Z(n5936) );
  XNOR U5989 ( .A(n6027), .B(n6011), .Z(n6016) );
  XOR U5990 ( .A(n6028), .B(n6029), .Z(n6011) );
  AND U5991 ( .A(n6030), .B(n6031), .Z(n6029) );
  XOR U5992 ( .A(n6032), .B(n6028), .Z(n6030) );
  XNOR U5993 ( .A(n6033), .B(n6034), .Z(n6027) );
  AND U5994 ( .A(n6035), .B(n6036), .Z(n6034) );
  XOR U5995 ( .A(n6033), .B(n6037), .Z(n6035) );
  XNOR U5996 ( .A(n6017), .B(n6014), .Z(n6026) );
  AND U5997 ( .A(n6038), .B(n6039), .Z(n6014) );
  XOR U5998 ( .A(n6040), .B(n6041), .Z(n6017) );
  AND U5999 ( .A(n6042), .B(n6043), .Z(n6041) );
  XOR U6000 ( .A(n6040), .B(n6044), .Z(n6042) );
  XNOR U6001 ( .A(n5933), .B(n6022), .Z(n6024) );
  XOR U6002 ( .A(n6045), .B(n6046), .Z(n5933) );
  AND U6003 ( .A(n111), .B(n6047), .Z(n6046) );
  XNOR U6004 ( .A(n6048), .B(n6045), .Z(n6047) );
  XOR U6005 ( .A(n6049), .B(n6050), .Z(n6022) );
  AND U6006 ( .A(n6051), .B(n6052), .Z(n6050) );
  XNOR U6007 ( .A(n6049), .B(n6038), .Z(n6052) );
  IV U6008 ( .A(n5984), .Z(n6038) );
  XNOR U6009 ( .A(n6053), .B(n6031), .Z(n5984) );
  XNOR U6010 ( .A(n6054), .B(n6037), .Z(n6031) );
  XOR U6011 ( .A(n6055), .B(n6056), .Z(n6037) );
  NOR U6012 ( .A(n6057), .B(n6058), .Z(n6056) );
  XNOR U6013 ( .A(n6055), .B(n6059), .Z(n6057) );
  XNOR U6014 ( .A(n6036), .B(n6028), .Z(n6054) );
  XOR U6015 ( .A(n6060), .B(n6061), .Z(n6028) );
  AND U6016 ( .A(n6062), .B(n6063), .Z(n6061) );
  XNOR U6017 ( .A(n6060), .B(n6064), .Z(n6062) );
  XNOR U6018 ( .A(n6065), .B(n6033), .Z(n6036) );
  XOR U6019 ( .A(n6066), .B(n6067), .Z(n6033) );
  AND U6020 ( .A(n6068), .B(n6069), .Z(n6067) );
  XOR U6021 ( .A(n6066), .B(n6070), .Z(n6068) );
  XNOR U6022 ( .A(n6071), .B(n6072), .Z(n6065) );
  NOR U6023 ( .A(n6073), .B(n6074), .Z(n6072) );
  XOR U6024 ( .A(n6071), .B(n6075), .Z(n6073) );
  XNOR U6025 ( .A(n6032), .B(n6039), .Z(n6053) );
  NOR U6026 ( .A(n5996), .B(n6076), .Z(n6039) );
  XOR U6027 ( .A(n6044), .B(n6043), .Z(n6032) );
  XNOR U6028 ( .A(n6077), .B(n6040), .Z(n6043) );
  XOR U6029 ( .A(n6078), .B(n6079), .Z(n6040) );
  AND U6030 ( .A(n6080), .B(n6081), .Z(n6079) );
  XOR U6031 ( .A(n6078), .B(n6082), .Z(n6080) );
  XNOR U6032 ( .A(n6083), .B(n6084), .Z(n6077) );
  NOR U6033 ( .A(n6085), .B(n6086), .Z(n6084) );
  XNOR U6034 ( .A(n6083), .B(n6087), .Z(n6085) );
  XOR U6035 ( .A(n6088), .B(n6089), .Z(n6044) );
  NOR U6036 ( .A(n6090), .B(n6091), .Z(n6089) );
  XNOR U6037 ( .A(n6088), .B(n6092), .Z(n6090) );
  XNOR U6038 ( .A(n5981), .B(n6049), .Z(n6051) );
  XOR U6039 ( .A(n6093), .B(n6094), .Z(n5981) );
  AND U6040 ( .A(n111), .B(n6095), .Z(n6094) );
  XOR U6041 ( .A(n6096), .B(n6093), .Z(n6095) );
  AND U6042 ( .A(n5993), .B(n5996), .Z(n6049) );
  XOR U6043 ( .A(n6097), .B(n6076), .Z(n5996) );
  XNOR U6044 ( .A(p_input[1024]), .B(p_input[416]), .Z(n6076) );
  XOR U6045 ( .A(n6064), .B(n6063), .Z(n6097) );
  XNOR U6046 ( .A(n6098), .B(n6070), .Z(n6063) );
  XNOR U6047 ( .A(n6059), .B(n6058), .Z(n6070) );
  XOR U6048 ( .A(n6099), .B(n6055), .Z(n6058) );
  XOR U6049 ( .A(p_input[1034]), .B(p_input[426]), .Z(n6055) );
  XNOR U6050 ( .A(p_input[1035]), .B(p_input[427]), .Z(n6099) );
  XOR U6051 ( .A(p_input[1036]), .B(p_input[428]), .Z(n6059) );
  XNOR U6052 ( .A(n6069), .B(n6060), .Z(n6098) );
  XNOR U6053 ( .A(n3298), .B(p_input[417]), .Z(n6060) );
  XOR U6054 ( .A(n6100), .B(n6075), .Z(n6069) );
  XNOR U6055 ( .A(p_input[1039]), .B(p_input[431]), .Z(n6075) );
  XOR U6056 ( .A(n6066), .B(n6074), .Z(n6100) );
  XOR U6057 ( .A(n6101), .B(n6071), .Z(n6074) );
  XOR U6058 ( .A(p_input[1037]), .B(p_input[429]), .Z(n6071) );
  XNOR U6059 ( .A(p_input[1038]), .B(p_input[430]), .Z(n6101) );
  XOR U6060 ( .A(p_input[1033]), .B(p_input[425]), .Z(n6066) );
  XNOR U6061 ( .A(n6082), .B(n6081), .Z(n6064) );
  XNOR U6062 ( .A(n6102), .B(n6087), .Z(n6081) );
  XOR U6063 ( .A(p_input[1032]), .B(p_input[424]), .Z(n6087) );
  XOR U6064 ( .A(n6078), .B(n6086), .Z(n6102) );
  XOR U6065 ( .A(n6103), .B(n6083), .Z(n6086) );
  XOR U6066 ( .A(p_input[1030]), .B(p_input[422]), .Z(n6083) );
  XNOR U6067 ( .A(p_input[1031]), .B(p_input[423]), .Z(n6103) );
  XOR U6068 ( .A(p_input[1026]), .B(p_input[418]), .Z(n6078) );
  XNOR U6069 ( .A(n6092), .B(n6091), .Z(n6082) );
  XOR U6070 ( .A(n6104), .B(n6088), .Z(n6091) );
  XOR U6071 ( .A(p_input[1027]), .B(p_input[419]), .Z(n6088) );
  XNOR U6072 ( .A(p_input[1028]), .B(p_input[420]), .Z(n6104) );
  XOR U6073 ( .A(p_input[1029]), .B(p_input[421]), .Z(n6092) );
  XOR U6074 ( .A(n6105), .B(n6106), .Z(n5993) );
  AND U6075 ( .A(n111), .B(n6107), .Z(n6106) );
  XNOR U6076 ( .A(n6108), .B(n6105), .Z(n6107) );
  XNOR U6077 ( .A(n6109), .B(n6110), .Z(n111) );
  AND U6078 ( .A(n6111), .B(n6112), .Z(n6110) );
  XOR U6079 ( .A(n6006), .B(n6109), .Z(n6112) );
  AND U6080 ( .A(n6113), .B(n6114), .Z(n6006) );
  XNOR U6081 ( .A(n6003), .B(n6109), .Z(n6111) );
  XOR U6082 ( .A(n6115), .B(n6116), .Z(n6003) );
  AND U6083 ( .A(n115), .B(n6117), .Z(n6116) );
  XOR U6084 ( .A(n6118), .B(n6115), .Z(n6117) );
  XOR U6085 ( .A(n6119), .B(n6120), .Z(n6109) );
  AND U6086 ( .A(n6121), .B(n6122), .Z(n6120) );
  XNOR U6087 ( .A(n6119), .B(n6113), .Z(n6122) );
  IV U6088 ( .A(n6021), .Z(n6113) );
  XOR U6089 ( .A(n6123), .B(n6124), .Z(n6021) );
  XOR U6090 ( .A(n6125), .B(n6114), .Z(n6124) );
  AND U6091 ( .A(n6048), .B(n6126), .Z(n6114) );
  AND U6092 ( .A(n6127), .B(n6128), .Z(n6125) );
  XOR U6093 ( .A(n6129), .B(n6123), .Z(n6127) );
  XNOR U6094 ( .A(n6018), .B(n6119), .Z(n6121) );
  XOR U6095 ( .A(n6130), .B(n6131), .Z(n6018) );
  AND U6096 ( .A(n115), .B(n6132), .Z(n6131) );
  XOR U6097 ( .A(n6133), .B(n6130), .Z(n6132) );
  XOR U6098 ( .A(n6134), .B(n6135), .Z(n6119) );
  AND U6099 ( .A(n6136), .B(n6137), .Z(n6135) );
  XNOR U6100 ( .A(n6134), .B(n6048), .Z(n6137) );
  XOR U6101 ( .A(n6138), .B(n6128), .Z(n6048) );
  XNOR U6102 ( .A(n6139), .B(n6123), .Z(n6128) );
  XOR U6103 ( .A(n6140), .B(n6141), .Z(n6123) );
  AND U6104 ( .A(n6142), .B(n6143), .Z(n6141) );
  XOR U6105 ( .A(n6144), .B(n6140), .Z(n6142) );
  XNOR U6106 ( .A(n6145), .B(n6146), .Z(n6139) );
  AND U6107 ( .A(n6147), .B(n6148), .Z(n6146) );
  XOR U6108 ( .A(n6145), .B(n6149), .Z(n6147) );
  XNOR U6109 ( .A(n6129), .B(n6126), .Z(n6138) );
  AND U6110 ( .A(n6150), .B(n6151), .Z(n6126) );
  XOR U6111 ( .A(n6152), .B(n6153), .Z(n6129) );
  AND U6112 ( .A(n6154), .B(n6155), .Z(n6153) );
  XOR U6113 ( .A(n6152), .B(n6156), .Z(n6154) );
  XNOR U6114 ( .A(n6045), .B(n6134), .Z(n6136) );
  XOR U6115 ( .A(n6157), .B(n6158), .Z(n6045) );
  AND U6116 ( .A(n115), .B(n6159), .Z(n6158) );
  XNOR U6117 ( .A(n6160), .B(n6157), .Z(n6159) );
  XOR U6118 ( .A(n6161), .B(n6162), .Z(n6134) );
  AND U6119 ( .A(n6163), .B(n6164), .Z(n6162) );
  XNOR U6120 ( .A(n6161), .B(n6150), .Z(n6164) );
  IV U6121 ( .A(n6096), .Z(n6150) );
  XNOR U6122 ( .A(n6165), .B(n6143), .Z(n6096) );
  XNOR U6123 ( .A(n6166), .B(n6149), .Z(n6143) );
  XOR U6124 ( .A(n6167), .B(n6168), .Z(n6149) );
  NOR U6125 ( .A(n6169), .B(n6170), .Z(n6168) );
  XNOR U6126 ( .A(n6167), .B(n6171), .Z(n6169) );
  XNOR U6127 ( .A(n6148), .B(n6140), .Z(n6166) );
  XOR U6128 ( .A(n6172), .B(n6173), .Z(n6140) );
  AND U6129 ( .A(n6174), .B(n6175), .Z(n6173) );
  XNOR U6130 ( .A(n6172), .B(n6176), .Z(n6174) );
  XNOR U6131 ( .A(n6177), .B(n6145), .Z(n6148) );
  XOR U6132 ( .A(n6178), .B(n6179), .Z(n6145) );
  AND U6133 ( .A(n6180), .B(n6181), .Z(n6179) );
  XOR U6134 ( .A(n6178), .B(n6182), .Z(n6180) );
  XNOR U6135 ( .A(n6183), .B(n6184), .Z(n6177) );
  NOR U6136 ( .A(n6185), .B(n6186), .Z(n6184) );
  XOR U6137 ( .A(n6183), .B(n6187), .Z(n6185) );
  XNOR U6138 ( .A(n6144), .B(n6151), .Z(n6165) );
  NOR U6139 ( .A(n6108), .B(n6188), .Z(n6151) );
  XOR U6140 ( .A(n6156), .B(n6155), .Z(n6144) );
  XNOR U6141 ( .A(n6189), .B(n6152), .Z(n6155) );
  XOR U6142 ( .A(n6190), .B(n6191), .Z(n6152) );
  AND U6143 ( .A(n6192), .B(n6193), .Z(n6191) );
  XOR U6144 ( .A(n6190), .B(n6194), .Z(n6192) );
  XNOR U6145 ( .A(n6195), .B(n6196), .Z(n6189) );
  NOR U6146 ( .A(n6197), .B(n6198), .Z(n6196) );
  XNOR U6147 ( .A(n6195), .B(n6199), .Z(n6197) );
  XOR U6148 ( .A(n6200), .B(n6201), .Z(n6156) );
  NOR U6149 ( .A(n6202), .B(n6203), .Z(n6201) );
  XNOR U6150 ( .A(n6200), .B(n6204), .Z(n6202) );
  XNOR U6151 ( .A(n6093), .B(n6161), .Z(n6163) );
  XOR U6152 ( .A(n6205), .B(n6206), .Z(n6093) );
  AND U6153 ( .A(n115), .B(n6207), .Z(n6206) );
  XOR U6154 ( .A(n6208), .B(n6205), .Z(n6207) );
  AND U6155 ( .A(n6105), .B(n6108), .Z(n6161) );
  XOR U6156 ( .A(n6209), .B(n6188), .Z(n6108) );
  XNOR U6157 ( .A(p_input[1024]), .B(p_input[432]), .Z(n6188) );
  XOR U6158 ( .A(n6176), .B(n6175), .Z(n6209) );
  XNOR U6159 ( .A(n6210), .B(n6182), .Z(n6175) );
  XNOR U6160 ( .A(n6171), .B(n6170), .Z(n6182) );
  XOR U6161 ( .A(n6211), .B(n6167), .Z(n6170) );
  XOR U6162 ( .A(p_input[1034]), .B(p_input[442]), .Z(n6167) );
  XNOR U6163 ( .A(p_input[1035]), .B(p_input[443]), .Z(n6211) );
  XOR U6164 ( .A(p_input[1036]), .B(p_input[444]), .Z(n6171) );
  XNOR U6165 ( .A(n6181), .B(n6172), .Z(n6210) );
  XNOR U6166 ( .A(n3298), .B(p_input[433]), .Z(n6172) );
  XOR U6167 ( .A(n6212), .B(n6187), .Z(n6181) );
  XNOR U6168 ( .A(p_input[1039]), .B(p_input[447]), .Z(n6187) );
  XOR U6169 ( .A(n6178), .B(n6186), .Z(n6212) );
  XOR U6170 ( .A(n6213), .B(n6183), .Z(n6186) );
  XOR U6171 ( .A(p_input[1037]), .B(p_input[445]), .Z(n6183) );
  XNOR U6172 ( .A(p_input[1038]), .B(p_input[446]), .Z(n6213) );
  XOR U6173 ( .A(p_input[1033]), .B(p_input[441]), .Z(n6178) );
  XNOR U6174 ( .A(n6194), .B(n6193), .Z(n6176) );
  XNOR U6175 ( .A(n6214), .B(n6199), .Z(n6193) );
  XOR U6176 ( .A(p_input[1032]), .B(p_input[440]), .Z(n6199) );
  XOR U6177 ( .A(n6190), .B(n6198), .Z(n6214) );
  XOR U6178 ( .A(n6215), .B(n6195), .Z(n6198) );
  XOR U6179 ( .A(p_input[1030]), .B(p_input[438]), .Z(n6195) );
  XNOR U6180 ( .A(p_input[1031]), .B(p_input[439]), .Z(n6215) );
  XOR U6181 ( .A(p_input[1026]), .B(p_input[434]), .Z(n6190) );
  XNOR U6182 ( .A(n6204), .B(n6203), .Z(n6194) );
  XOR U6183 ( .A(n6216), .B(n6200), .Z(n6203) );
  XOR U6184 ( .A(p_input[1027]), .B(p_input[435]), .Z(n6200) );
  XNOR U6185 ( .A(p_input[1028]), .B(p_input[436]), .Z(n6216) );
  XOR U6186 ( .A(p_input[1029]), .B(p_input[437]), .Z(n6204) );
  XOR U6187 ( .A(n6217), .B(n6218), .Z(n6105) );
  AND U6188 ( .A(n115), .B(n6219), .Z(n6218) );
  XNOR U6189 ( .A(n6220), .B(n6217), .Z(n6219) );
  XNOR U6190 ( .A(n6221), .B(n6222), .Z(n115) );
  AND U6191 ( .A(n6223), .B(n6224), .Z(n6222) );
  XOR U6192 ( .A(n6118), .B(n6221), .Z(n6224) );
  AND U6193 ( .A(n6225), .B(n6226), .Z(n6118) );
  XNOR U6194 ( .A(n6115), .B(n6221), .Z(n6223) );
  XOR U6195 ( .A(n6227), .B(n6228), .Z(n6115) );
  AND U6196 ( .A(n119), .B(n6229), .Z(n6228) );
  XOR U6197 ( .A(n6230), .B(n6227), .Z(n6229) );
  XOR U6198 ( .A(n6231), .B(n6232), .Z(n6221) );
  AND U6199 ( .A(n6233), .B(n6234), .Z(n6232) );
  XNOR U6200 ( .A(n6231), .B(n6225), .Z(n6234) );
  IV U6201 ( .A(n6133), .Z(n6225) );
  XOR U6202 ( .A(n6235), .B(n6236), .Z(n6133) );
  XOR U6203 ( .A(n6237), .B(n6226), .Z(n6236) );
  AND U6204 ( .A(n6160), .B(n6238), .Z(n6226) );
  AND U6205 ( .A(n6239), .B(n6240), .Z(n6237) );
  XOR U6206 ( .A(n6241), .B(n6235), .Z(n6239) );
  XNOR U6207 ( .A(n6130), .B(n6231), .Z(n6233) );
  XOR U6208 ( .A(n6242), .B(n6243), .Z(n6130) );
  AND U6209 ( .A(n119), .B(n6244), .Z(n6243) );
  XOR U6210 ( .A(n6245), .B(n6242), .Z(n6244) );
  XOR U6211 ( .A(n6246), .B(n6247), .Z(n6231) );
  AND U6212 ( .A(n6248), .B(n6249), .Z(n6247) );
  XNOR U6213 ( .A(n6246), .B(n6160), .Z(n6249) );
  XOR U6214 ( .A(n6250), .B(n6240), .Z(n6160) );
  XNOR U6215 ( .A(n6251), .B(n6235), .Z(n6240) );
  XOR U6216 ( .A(n6252), .B(n6253), .Z(n6235) );
  AND U6217 ( .A(n6254), .B(n6255), .Z(n6253) );
  XOR U6218 ( .A(n6256), .B(n6252), .Z(n6254) );
  XNOR U6219 ( .A(n6257), .B(n6258), .Z(n6251) );
  AND U6220 ( .A(n6259), .B(n6260), .Z(n6258) );
  XOR U6221 ( .A(n6257), .B(n6261), .Z(n6259) );
  XNOR U6222 ( .A(n6241), .B(n6238), .Z(n6250) );
  AND U6223 ( .A(n6262), .B(n6263), .Z(n6238) );
  XOR U6224 ( .A(n6264), .B(n6265), .Z(n6241) );
  AND U6225 ( .A(n6266), .B(n6267), .Z(n6265) );
  XOR U6226 ( .A(n6264), .B(n6268), .Z(n6266) );
  XNOR U6227 ( .A(n6157), .B(n6246), .Z(n6248) );
  XOR U6228 ( .A(n6269), .B(n6270), .Z(n6157) );
  AND U6229 ( .A(n119), .B(n6271), .Z(n6270) );
  XNOR U6230 ( .A(n6272), .B(n6269), .Z(n6271) );
  XOR U6231 ( .A(n6273), .B(n6274), .Z(n6246) );
  AND U6232 ( .A(n6275), .B(n6276), .Z(n6274) );
  XNOR U6233 ( .A(n6273), .B(n6262), .Z(n6276) );
  IV U6234 ( .A(n6208), .Z(n6262) );
  XNOR U6235 ( .A(n6277), .B(n6255), .Z(n6208) );
  XNOR U6236 ( .A(n6278), .B(n6261), .Z(n6255) );
  XOR U6237 ( .A(n6279), .B(n6280), .Z(n6261) );
  NOR U6238 ( .A(n6281), .B(n6282), .Z(n6280) );
  XNOR U6239 ( .A(n6279), .B(n6283), .Z(n6281) );
  XNOR U6240 ( .A(n6260), .B(n6252), .Z(n6278) );
  XOR U6241 ( .A(n6284), .B(n6285), .Z(n6252) );
  AND U6242 ( .A(n6286), .B(n6287), .Z(n6285) );
  XNOR U6243 ( .A(n6284), .B(n6288), .Z(n6286) );
  XNOR U6244 ( .A(n6289), .B(n6257), .Z(n6260) );
  XOR U6245 ( .A(n6290), .B(n6291), .Z(n6257) );
  AND U6246 ( .A(n6292), .B(n6293), .Z(n6291) );
  XOR U6247 ( .A(n6290), .B(n6294), .Z(n6292) );
  XNOR U6248 ( .A(n6295), .B(n6296), .Z(n6289) );
  NOR U6249 ( .A(n6297), .B(n6298), .Z(n6296) );
  XOR U6250 ( .A(n6295), .B(n6299), .Z(n6297) );
  XNOR U6251 ( .A(n6256), .B(n6263), .Z(n6277) );
  NOR U6252 ( .A(n6220), .B(n6300), .Z(n6263) );
  XOR U6253 ( .A(n6268), .B(n6267), .Z(n6256) );
  XNOR U6254 ( .A(n6301), .B(n6264), .Z(n6267) );
  XOR U6255 ( .A(n6302), .B(n6303), .Z(n6264) );
  AND U6256 ( .A(n6304), .B(n6305), .Z(n6303) );
  XOR U6257 ( .A(n6302), .B(n6306), .Z(n6304) );
  XNOR U6258 ( .A(n6307), .B(n6308), .Z(n6301) );
  NOR U6259 ( .A(n6309), .B(n6310), .Z(n6308) );
  XNOR U6260 ( .A(n6307), .B(n6311), .Z(n6309) );
  XOR U6261 ( .A(n6312), .B(n6313), .Z(n6268) );
  NOR U6262 ( .A(n6314), .B(n6315), .Z(n6313) );
  XNOR U6263 ( .A(n6312), .B(n6316), .Z(n6314) );
  XNOR U6264 ( .A(n6205), .B(n6273), .Z(n6275) );
  XOR U6265 ( .A(n6317), .B(n6318), .Z(n6205) );
  AND U6266 ( .A(n119), .B(n6319), .Z(n6318) );
  XOR U6267 ( .A(n6320), .B(n6317), .Z(n6319) );
  AND U6268 ( .A(n6217), .B(n6220), .Z(n6273) );
  XOR U6269 ( .A(n6321), .B(n6300), .Z(n6220) );
  XNOR U6270 ( .A(p_input[1024]), .B(p_input[448]), .Z(n6300) );
  XOR U6271 ( .A(n6288), .B(n6287), .Z(n6321) );
  XNOR U6272 ( .A(n6322), .B(n6294), .Z(n6287) );
  XNOR U6273 ( .A(n6283), .B(n6282), .Z(n6294) );
  XOR U6274 ( .A(n6323), .B(n6279), .Z(n6282) );
  XOR U6275 ( .A(p_input[1034]), .B(p_input[458]), .Z(n6279) );
  XNOR U6276 ( .A(p_input[1035]), .B(p_input[459]), .Z(n6323) );
  XOR U6277 ( .A(p_input[1036]), .B(p_input[460]), .Z(n6283) );
  XNOR U6278 ( .A(n6293), .B(n6284), .Z(n6322) );
  XNOR U6279 ( .A(n3298), .B(p_input[449]), .Z(n6284) );
  XOR U6280 ( .A(n6324), .B(n6299), .Z(n6293) );
  XNOR U6281 ( .A(p_input[1039]), .B(p_input[463]), .Z(n6299) );
  XOR U6282 ( .A(n6290), .B(n6298), .Z(n6324) );
  XOR U6283 ( .A(n6325), .B(n6295), .Z(n6298) );
  XOR U6284 ( .A(p_input[1037]), .B(p_input[461]), .Z(n6295) );
  XNOR U6285 ( .A(p_input[1038]), .B(p_input[462]), .Z(n6325) );
  XOR U6286 ( .A(p_input[1033]), .B(p_input[457]), .Z(n6290) );
  XNOR U6287 ( .A(n6306), .B(n6305), .Z(n6288) );
  XNOR U6288 ( .A(n6326), .B(n6311), .Z(n6305) );
  XOR U6289 ( .A(p_input[1032]), .B(p_input[456]), .Z(n6311) );
  XOR U6290 ( .A(n6302), .B(n6310), .Z(n6326) );
  XOR U6291 ( .A(n6327), .B(n6307), .Z(n6310) );
  XOR U6292 ( .A(p_input[1030]), .B(p_input[454]), .Z(n6307) );
  XNOR U6293 ( .A(p_input[1031]), .B(p_input[455]), .Z(n6327) );
  XOR U6294 ( .A(p_input[1026]), .B(p_input[450]), .Z(n6302) );
  XNOR U6295 ( .A(n6316), .B(n6315), .Z(n6306) );
  XOR U6296 ( .A(n6328), .B(n6312), .Z(n6315) );
  XOR U6297 ( .A(p_input[1027]), .B(p_input[451]), .Z(n6312) );
  XNOR U6298 ( .A(p_input[1028]), .B(p_input[452]), .Z(n6328) );
  XOR U6299 ( .A(p_input[1029]), .B(p_input[453]), .Z(n6316) );
  XOR U6300 ( .A(n6329), .B(n6330), .Z(n6217) );
  AND U6301 ( .A(n119), .B(n6331), .Z(n6330) );
  XNOR U6302 ( .A(n6332), .B(n6329), .Z(n6331) );
  XNOR U6303 ( .A(n6333), .B(n6334), .Z(n119) );
  AND U6304 ( .A(n6335), .B(n6336), .Z(n6334) );
  XOR U6305 ( .A(n6230), .B(n6333), .Z(n6336) );
  AND U6306 ( .A(n6337), .B(n6338), .Z(n6230) );
  XNOR U6307 ( .A(n6227), .B(n6333), .Z(n6335) );
  XOR U6308 ( .A(n6339), .B(n6340), .Z(n6227) );
  AND U6309 ( .A(n123), .B(n6341), .Z(n6340) );
  XOR U6310 ( .A(n6342), .B(n6339), .Z(n6341) );
  XOR U6311 ( .A(n6343), .B(n6344), .Z(n6333) );
  AND U6312 ( .A(n6345), .B(n6346), .Z(n6344) );
  XNOR U6313 ( .A(n6343), .B(n6337), .Z(n6346) );
  IV U6314 ( .A(n6245), .Z(n6337) );
  XOR U6315 ( .A(n6347), .B(n6348), .Z(n6245) );
  XOR U6316 ( .A(n6349), .B(n6338), .Z(n6348) );
  AND U6317 ( .A(n6272), .B(n6350), .Z(n6338) );
  AND U6318 ( .A(n6351), .B(n6352), .Z(n6349) );
  XOR U6319 ( .A(n6353), .B(n6347), .Z(n6351) );
  XNOR U6320 ( .A(n6242), .B(n6343), .Z(n6345) );
  XOR U6321 ( .A(n6354), .B(n6355), .Z(n6242) );
  AND U6322 ( .A(n123), .B(n6356), .Z(n6355) );
  XOR U6323 ( .A(n6357), .B(n6354), .Z(n6356) );
  XOR U6324 ( .A(n6358), .B(n6359), .Z(n6343) );
  AND U6325 ( .A(n6360), .B(n6361), .Z(n6359) );
  XNOR U6326 ( .A(n6358), .B(n6272), .Z(n6361) );
  XOR U6327 ( .A(n6362), .B(n6352), .Z(n6272) );
  XNOR U6328 ( .A(n6363), .B(n6347), .Z(n6352) );
  XOR U6329 ( .A(n6364), .B(n6365), .Z(n6347) );
  AND U6330 ( .A(n6366), .B(n6367), .Z(n6365) );
  XOR U6331 ( .A(n6368), .B(n6364), .Z(n6366) );
  XNOR U6332 ( .A(n6369), .B(n6370), .Z(n6363) );
  AND U6333 ( .A(n6371), .B(n6372), .Z(n6370) );
  XOR U6334 ( .A(n6369), .B(n6373), .Z(n6371) );
  XNOR U6335 ( .A(n6353), .B(n6350), .Z(n6362) );
  AND U6336 ( .A(n6374), .B(n6375), .Z(n6350) );
  XOR U6337 ( .A(n6376), .B(n6377), .Z(n6353) );
  AND U6338 ( .A(n6378), .B(n6379), .Z(n6377) );
  XOR U6339 ( .A(n6376), .B(n6380), .Z(n6378) );
  XNOR U6340 ( .A(n6269), .B(n6358), .Z(n6360) );
  XOR U6341 ( .A(n6381), .B(n6382), .Z(n6269) );
  AND U6342 ( .A(n123), .B(n6383), .Z(n6382) );
  XNOR U6343 ( .A(n6384), .B(n6381), .Z(n6383) );
  XOR U6344 ( .A(n6385), .B(n6386), .Z(n6358) );
  AND U6345 ( .A(n6387), .B(n6388), .Z(n6386) );
  XNOR U6346 ( .A(n6385), .B(n6374), .Z(n6388) );
  IV U6347 ( .A(n6320), .Z(n6374) );
  XNOR U6348 ( .A(n6389), .B(n6367), .Z(n6320) );
  XNOR U6349 ( .A(n6390), .B(n6373), .Z(n6367) );
  XOR U6350 ( .A(n6391), .B(n6392), .Z(n6373) );
  NOR U6351 ( .A(n6393), .B(n6394), .Z(n6392) );
  XNOR U6352 ( .A(n6391), .B(n6395), .Z(n6393) );
  XNOR U6353 ( .A(n6372), .B(n6364), .Z(n6390) );
  XOR U6354 ( .A(n6396), .B(n6397), .Z(n6364) );
  AND U6355 ( .A(n6398), .B(n6399), .Z(n6397) );
  XNOR U6356 ( .A(n6396), .B(n6400), .Z(n6398) );
  XNOR U6357 ( .A(n6401), .B(n6369), .Z(n6372) );
  XOR U6358 ( .A(n6402), .B(n6403), .Z(n6369) );
  AND U6359 ( .A(n6404), .B(n6405), .Z(n6403) );
  XOR U6360 ( .A(n6402), .B(n6406), .Z(n6404) );
  XNOR U6361 ( .A(n6407), .B(n6408), .Z(n6401) );
  NOR U6362 ( .A(n6409), .B(n6410), .Z(n6408) );
  XOR U6363 ( .A(n6407), .B(n6411), .Z(n6409) );
  XNOR U6364 ( .A(n6368), .B(n6375), .Z(n6389) );
  NOR U6365 ( .A(n6332), .B(n6412), .Z(n6375) );
  XOR U6366 ( .A(n6380), .B(n6379), .Z(n6368) );
  XNOR U6367 ( .A(n6413), .B(n6376), .Z(n6379) );
  XOR U6368 ( .A(n6414), .B(n6415), .Z(n6376) );
  AND U6369 ( .A(n6416), .B(n6417), .Z(n6415) );
  XOR U6370 ( .A(n6414), .B(n6418), .Z(n6416) );
  XNOR U6371 ( .A(n6419), .B(n6420), .Z(n6413) );
  NOR U6372 ( .A(n6421), .B(n6422), .Z(n6420) );
  XNOR U6373 ( .A(n6419), .B(n6423), .Z(n6421) );
  XOR U6374 ( .A(n6424), .B(n6425), .Z(n6380) );
  NOR U6375 ( .A(n6426), .B(n6427), .Z(n6425) );
  XNOR U6376 ( .A(n6424), .B(n6428), .Z(n6426) );
  XNOR U6377 ( .A(n6317), .B(n6385), .Z(n6387) );
  XOR U6378 ( .A(n6429), .B(n6430), .Z(n6317) );
  AND U6379 ( .A(n123), .B(n6431), .Z(n6430) );
  XOR U6380 ( .A(n6432), .B(n6429), .Z(n6431) );
  AND U6381 ( .A(n6329), .B(n6332), .Z(n6385) );
  XOR U6382 ( .A(n6433), .B(n6412), .Z(n6332) );
  XNOR U6383 ( .A(p_input[1024]), .B(p_input[464]), .Z(n6412) );
  XOR U6384 ( .A(n6400), .B(n6399), .Z(n6433) );
  XNOR U6385 ( .A(n6434), .B(n6406), .Z(n6399) );
  XNOR U6386 ( .A(n6395), .B(n6394), .Z(n6406) );
  XOR U6387 ( .A(n6435), .B(n6391), .Z(n6394) );
  XOR U6388 ( .A(p_input[1034]), .B(p_input[474]), .Z(n6391) );
  XNOR U6389 ( .A(p_input[1035]), .B(p_input[475]), .Z(n6435) );
  XOR U6390 ( .A(p_input[1036]), .B(p_input[476]), .Z(n6395) );
  XNOR U6391 ( .A(n6405), .B(n6396), .Z(n6434) );
  XNOR U6392 ( .A(n3298), .B(p_input[465]), .Z(n6396) );
  XOR U6393 ( .A(n6436), .B(n6411), .Z(n6405) );
  XNOR U6394 ( .A(p_input[1039]), .B(p_input[479]), .Z(n6411) );
  XOR U6395 ( .A(n6402), .B(n6410), .Z(n6436) );
  XOR U6396 ( .A(n6437), .B(n6407), .Z(n6410) );
  XOR U6397 ( .A(p_input[1037]), .B(p_input[477]), .Z(n6407) );
  XNOR U6398 ( .A(p_input[1038]), .B(p_input[478]), .Z(n6437) );
  XOR U6399 ( .A(p_input[1033]), .B(p_input[473]), .Z(n6402) );
  XNOR U6400 ( .A(n6418), .B(n6417), .Z(n6400) );
  XNOR U6401 ( .A(n6438), .B(n6423), .Z(n6417) );
  XOR U6402 ( .A(p_input[1032]), .B(p_input[472]), .Z(n6423) );
  XOR U6403 ( .A(n6414), .B(n6422), .Z(n6438) );
  XOR U6404 ( .A(n6439), .B(n6419), .Z(n6422) );
  XOR U6405 ( .A(p_input[1030]), .B(p_input[470]), .Z(n6419) );
  XNOR U6406 ( .A(p_input[1031]), .B(p_input[471]), .Z(n6439) );
  XOR U6407 ( .A(p_input[1026]), .B(p_input[466]), .Z(n6414) );
  XNOR U6408 ( .A(n6428), .B(n6427), .Z(n6418) );
  XOR U6409 ( .A(n6440), .B(n6424), .Z(n6427) );
  XOR U6410 ( .A(p_input[1027]), .B(p_input[467]), .Z(n6424) );
  XNOR U6411 ( .A(p_input[1028]), .B(p_input[468]), .Z(n6440) );
  XOR U6412 ( .A(p_input[1029]), .B(p_input[469]), .Z(n6428) );
  XOR U6413 ( .A(n6441), .B(n6442), .Z(n6329) );
  AND U6414 ( .A(n123), .B(n6443), .Z(n6442) );
  XNOR U6415 ( .A(n6444), .B(n6441), .Z(n6443) );
  XNOR U6416 ( .A(n6445), .B(n6446), .Z(n123) );
  AND U6417 ( .A(n6447), .B(n6448), .Z(n6446) );
  XOR U6418 ( .A(n6342), .B(n6445), .Z(n6448) );
  AND U6419 ( .A(n6449), .B(n6450), .Z(n6342) );
  XNOR U6420 ( .A(n6339), .B(n6445), .Z(n6447) );
  XOR U6421 ( .A(n6451), .B(n6452), .Z(n6339) );
  AND U6422 ( .A(n127), .B(n6453), .Z(n6452) );
  XOR U6423 ( .A(n6454), .B(n6451), .Z(n6453) );
  XOR U6424 ( .A(n6455), .B(n6456), .Z(n6445) );
  AND U6425 ( .A(n6457), .B(n6458), .Z(n6456) );
  XNOR U6426 ( .A(n6455), .B(n6449), .Z(n6458) );
  IV U6427 ( .A(n6357), .Z(n6449) );
  XOR U6428 ( .A(n6459), .B(n6460), .Z(n6357) );
  XOR U6429 ( .A(n6461), .B(n6450), .Z(n6460) );
  AND U6430 ( .A(n6384), .B(n6462), .Z(n6450) );
  AND U6431 ( .A(n6463), .B(n6464), .Z(n6461) );
  XOR U6432 ( .A(n6465), .B(n6459), .Z(n6463) );
  XNOR U6433 ( .A(n6354), .B(n6455), .Z(n6457) );
  XOR U6434 ( .A(n6466), .B(n6467), .Z(n6354) );
  AND U6435 ( .A(n127), .B(n6468), .Z(n6467) );
  XOR U6436 ( .A(n6469), .B(n6466), .Z(n6468) );
  XOR U6437 ( .A(n6470), .B(n6471), .Z(n6455) );
  AND U6438 ( .A(n6472), .B(n6473), .Z(n6471) );
  XNOR U6439 ( .A(n6470), .B(n6384), .Z(n6473) );
  XOR U6440 ( .A(n6474), .B(n6464), .Z(n6384) );
  XNOR U6441 ( .A(n6475), .B(n6459), .Z(n6464) );
  XOR U6442 ( .A(n6476), .B(n6477), .Z(n6459) );
  AND U6443 ( .A(n6478), .B(n6479), .Z(n6477) );
  XOR U6444 ( .A(n6480), .B(n6476), .Z(n6478) );
  XNOR U6445 ( .A(n6481), .B(n6482), .Z(n6475) );
  AND U6446 ( .A(n6483), .B(n6484), .Z(n6482) );
  XOR U6447 ( .A(n6481), .B(n6485), .Z(n6483) );
  XNOR U6448 ( .A(n6465), .B(n6462), .Z(n6474) );
  AND U6449 ( .A(n6486), .B(n6487), .Z(n6462) );
  XOR U6450 ( .A(n6488), .B(n6489), .Z(n6465) );
  AND U6451 ( .A(n6490), .B(n6491), .Z(n6489) );
  XOR U6452 ( .A(n6488), .B(n6492), .Z(n6490) );
  XNOR U6453 ( .A(n6381), .B(n6470), .Z(n6472) );
  XOR U6454 ( .A(n6493), .B(n6494), .Z(n6381) );
  AND U6455 ( .A(n127), .B(n6495), .Z(n6494) );
  XNOR U6456 ( .A(n6496), .B(n6493), .Z(n6495) );
  XOR U6457 ( .A(n6497), .B(n6498), .Z(n6470) );
  AND U6458 ( .A(n6499), .B(n6500), .Z(n6498) );
  XNOR U6459 ( .A(n6497), .B(n6486), .Z(n6500) );
  IV U6460 ( .A(n6432), .Z(n6486) );
  XNOR U6461 ( .A(n6501), .B(n6479), .Z(n6432) );
  XNOR U6462 ( .A(n6502), .B(n6485), .Z(n6479) );
  XOR U6463 ( .A(n6503), .B(n6504), .Z(n6485) );
  NOR U6464 ( .A(n6505), .B(n6506), .Z(n6504) );
  XNOR U6465 ( .A(n6503), .B(n6507), .Z(n6505) );
  XNOR U6466 ( .A(n6484), .B(n6476), .Z(n6502) );
  XOR U6467 ( .A(n6508), .B(n6509), .Z(n6476) );
  AND U6468 ( .A(n6510), .B(n6511), .Z(n6509) );
  XNOR U6469 ( .A(n6508), .B(n6512), .Z(n6510) );
  XNOR U6470 ( .A(n6513), .B(n6481), .Z(n6484) );
  XOR U6471 ( .A(n6514), .B(n6515), .Z(n6481) );
  AND U6472 ( .A(n6516), .B(n6517), .Z(n6515) );
  XOR U6473 ( .A(n6514), .B(n6518), .Z(n6516) );
  XNOR U6474 ( .A(n6519), .B(n6520), .Z(n6513) );
  NOR U6475 ( .A(n6521), .B(n6522), .Z(n6520) );
  XOR U6476 ( .A(n6519), .B(n6523), .Z(n6521) );
  XNOR U6477 ( .A(n6480), .B(n6487), .Z(n6501) );
  NOR U6478 ( .A(n6444), .B(n6524), .Z(n6487) );
  XOR U6479 ( .A(n6492), .B(n6491), .Z(n6480) );
  XNOR U6480 ( .A(n6525), .B(n6488), .Z(n6491) );
  XOR U6481 ( .A(n6526), .B(n6527), .Z(n6488) );
  AND U6482 ( .A(n6528), .B(n6529), .Z(n6527) );
  XOR U6483 ( .A(n6526), .B(n6530), .Z(n6528) );
  XNOR U6484 ( .A(n6531), .B(n6532), .Z(n6525) );
  NOR U6485 ( .A(n6533), .B(n6534), .Z(n6532) );
  XNOR U6486 ( .A(n6531), .B(n6535), .Z(n6533) );
  XOR U6487 ( .A(n6536), .B(n6537), .Z(n6492) );
  NOR U6488 ( .A(n6538), .B(n6539), .Z(n6537) );
  XNOR U6489 ( .A(n6536), .B(n6540), .Z(n6538) );
  XNOR U6490 ( .A(n6429), .B(n6497), .Z(n6499) );
  XOR U6491 ( .A(n6541), .B(n6542), .Z(n6429) );
  AND U6492 ( .A(n127), .B(n6543), .Z(n6542) );
  XOR U6493 ( .A(n6544), .B(n6541), .Z(n6543) );
  AND U6494 ( .A(n6441), .B(n6444), .Z(n6497) );
  XOR U6495 ( .A(n6545), .B(n6524), .Z(n6444) );
  XNOR U6496 ( .A(p_input[1024]), .B(p_input[480]), .Z(n6524) );
  XOR U6497 ( .A(n6512), .B(n6511), .Z(n6545) );
  XNOR U6498 ( .A(n6546), .B(n6518), .Z(n6511) );
  XNOR U6499 ( .A(n6507), .B(n6506), .Z(n6518) );
  XOR U6500 ( .A(n6547), .B(n6503), .Z(n6506) );
  XOR U6501 ( .A(p_input[1034]), .B(p_input[490]), .Z(n6503) );
  XNOR U6502 ( .A(p_input[1035]), .B(p_input[491]), .Z(n6547) );
  XOR U6503 ( .A(p_input[1036]), .B(p_input[492]), .Z(n6507) );
  XNOR U6504 ( .A(n6517), .B(n6508), .Z(n6546) );
  XNOR U6505 ( .A(n3298), .B(p_input[481]), .Z(n6508) );
  XOR U6506 ( .A(n6548), .B(n6523), .Z(n6517) );
  XNOR U6507 ( .A(p_input[1039]), .B(p_input[495]), .Z(n6523) );
  XOR U6508 ( .A(n6514), .B(n6522), .Z(n6548) );
  XOR U6509 ( .A(n6549), .B(n6519), .Z(n6522) );
  XOR U6510 ( .A(p_input[1037]), .B(p_input[493]), .Z(n6519) );
  XNOR U6511 ( .A(p_input[1038]), .B(p_input[494]), .Z(n6549) );
  XOR U6512 ( .A(p_input[1033]), .B(p_input[489]), .Z(n6514) );
  XNOR U6513 ( .A(n6530), .B(n6529), .Z(n6512) );
  XNOR U6514 ( .A(n6550), .B(n6535), .Z(n6529) );
  XOR U6515 ( .A(p_input[1032]), .B(p_input[488]), .Z(n6535) );
  XOR U6516 ( .A(n6526), .B(n6534), .Z(n6550) );
  XOR U6517 ( .A(n6551), .B(n6531), .Z(n6534) );
  XOR U6518 ( .A(p_input[1030]), .B(p_input[486]), .Z(n6531) );
  XNOR U6519 ( .A(p_input[1031]), .B(p_input[487]), .Z(n6551) );
  XOR U6520 ( .A(p_input[1026]), .B(p_input[482]), .Z(n6526) );
  XNOR U6521 ( .A(n6540), .B(n6539), .Z(n6530) );
  XOR U6522 ( .A(n6552), .B(n6536), .Z(n6539) );
  XOR U6523 ( .A(p_input[1027]), .B(p_input[483]), .Z(n6536) );
  XNOR U6524 ( .A(p_input[1028]), .B(p_input[484]), .Z(n6552) );
  XOR U6525 ( .A(p_input[1029]), .B(p_input[485]), .Z(n6540) );
  XOR U6526 ( .A(n6553), .B(n6554), .Z(n6441) );
  AND U6527 ( .A(n127), .B(n6555), .Z(n6554) );
  XNOR U6528 ( .A(n6556), .B(n6553), .Z(n6555) );
  XNOR U6529 ( .A(n6557), .B(n6558), .Z(n127) );
  AND U6530 ( .A(n6559), .B(n6560), .Z(n6558) );
  XOR U6531 ( .A(n6454), .B(n6557), .Z(n6560) );
  AND U6532 ( .A(n6561), .B(n6562), .Z(n6454) );
  XNOR U6533 ( .A(n6451), .B(n6557), .Z(n6559) );
  XOR U6534 ( .A(n6563), .B(n6564), .Z(n6451) );
  AND U6535 ( .A(n131), .B(n6565), .Z(n6564) );
  XOR U6536 ( .A(n6566), .B(n6563), .Z(n6565) );
  XOR U6537 ( .A(n6567), .B(n6568), .Z(n6557) );
  AND U6538 ( .A(n6569), .B(n6570), .Z(n6568) );
  XNOR U6539 ( .A(n6567), .B(n6561), .Z(n6570) );
  IV U6540 ( .A(n6469), .Z(n6561) );
  XOR U6541 ( .A(n6571), .B(n6572), .Z(n6469) );
  XOR U6542 ( .A(n6573), .B(n6562), .Z(n6572) );
  AND U6543 ( .A(n6496), .B(n6574), .Z(n6562) );
  AND U6544 ( .A(n6575), .B(n6576), .Z(n6573) );
  XOR U6545 ( .A(n6577), .B(n6571), .Z(n6575) );
  XNOR U6546 ( .A(n6466), .B(n6567), .Z(n6569) );
  XOR U6547 ( .A(n6578), .B(n6579), .Z(n6466) );
  AND U6548 ( .A(n131), .B(n6580), .Z(n6579) );
  XOR U6549 ( .A(n6581), .B(n6578), .Z(n6580) );
  XOR U6550 ( .A(n6582), .B(n6583), .Z(n6567) );
  AND U6551 ( .A(n6584), .B(n6585), .Z(n6583) );
  XNOR U6552 ( .A(n6582), .B(n6496), .Z(n6585) );
  XOR U6553 ( .A(n6586), .B(n6576), .Z(n6496) );
  XNOR U6554 ( .A(n6587), .B(n6571), .Z(n6576) );
  XOR U6555 ( .A(n6588), .B(n6589), .Z(n6571) );
  AND U6556 ( .A(n6590), .B(n6591), .Z(n6589) );
  XOR U6557 ( .A(n6592), .B(n6588), .Z(n6590) );
  XNOR U6558 ( .A(n6593), .B(n6594), .Z(n6587) );
  AND U6559 ( .A(n6595), .B(n6596), .Z(n6594) );
  XOR U6560 ( .A(n6593), .B(n6597), .Z(n6595) );
  XNOR U6561 ( .A(n6577), .B(n6574), .Z(n6586) );
  AND U6562 ( .A(n6598), .B(n6599), .Z(n6574) );
  XOR U6563 ( .A(n6600), .B(n6601), .Z(n6577) );
  AND U6564 ( .A(n6602), .B(n6603), .Z(n6601) );
  XOR U6565 ( .A(n6600), .B(n6604), .Z(n6602) );
  XNOR U6566 ( .A(n6493), .B(n6582), .Z(n6584) );
  XOR U6567 ( .A(n6605), .B(n6606), .Z(n6493) );
  AND U6568 ( .A(n131), .B(n6607), .Z(n6606) );
  XNOR U6569 ( .A(n6608), .B(n6605), .Z(n6607) );
  XOR U6570 ( .A(n6609), .B(n6610), .Z(n6582) );
  AND U6571 ( .A(n6611), .B(n6612), .Z(n6610) );
  XNOR U6572 ( .A(n6609), .B(n6598), .Z(n6612) );
  IV U6573 ( .A(n6544), .Z(n6598) );
  XNOR U6574 ( .A(n6613), .B(n6591), .Z(n6544) );
  XNOR U6575 ( .A(n6614), .B(n6597), .Z(n6591) );
  XOR U6576 ( .A(n6615), .B(n6616), .Z(n6597) );
  NOR U6577 ( .A(n6617), .B(n6618), .Z(n6616) );
  XNOR U6578 ( .A(n6615), .B(n6619), .Z(n6617) );
  XNOR U6579 ( .A(n6596), .B(n6588), .Z(n6614) );
  XOR U6580 ( .A(n6620), .B(n6621), .Z(n6588) );
  AND U6581 ( .A(n6622), .B(n6623), .Z(n6621) );
  XNOR U6582 ( .A(n6620), .B(n6624), .Z(n6622) );
  XNOR U6583 ( .A(n6625), .B(n6593), .Z(n6596) );
  XOR U6584 ( .A(n6626), .B(n6627), .Z(n6593) );
  AND U6585 ( .A(n6628), .B(n6629), .Z(n6627) );
  XOR U6586 ( .A(n6626), .B(n6630), .Z(n6628) );
  XNOR U6587 ( .A(n6631), .B(n6632), .Z(n6625) );
  NOR U6588 ( .A(n6633), .B(n6634), .Z(n6632) );
  XOR U6589 ( .A(n6631), .B(n6635), .Z(n6633) );
  XNOR U6590 ( .A(n6592), .B(n6599), .Z(n6613) );
  NOR U6591 ( .A(n6556), .B(n6636), .Z(n6599) );
  XOR U6592 ( .A(n6604), .B(n6603), .Z(n6592) );
  XNOR U6593 ( .A(n6637), .B(n6600), .Z(n6603) );
  XOR U6594 ( .A(n6638), .B(n6639), .Z(n6600) );
  AND U6595 ( .A(n6640), .B(n6641), .Z(n6639) );
  XOR U6596 ( .A(n6638), .B(n6642), .Z(n6640) );
  XNOR U6597 ( .A(n6643), .B(n6644), .Z(n6637) );
  NOR U6598 ( .A(n6645), .B(n6646), .Z(n6644) );
  XNOR U6599 ( .A(n6643), .B(n6647), .Z(n6645) );
  XOR U6600 ( .A(n6648), .B(n6649), .Z(n6604) );
  NOR U6601 ( .A(n6650), .B(n6651), .Z(n6649) );
  XNOR U6602 ( .A(n6648), .B(n6652), .Z(n6650) );
  XNOR U6603 ( .A(n6541), .B(n6609), .Z(n6611) );
  XOR U6604 ( .A(n6653), .B(n6654), .Z(n6541) );
  AND U6605 ( .A(n131), .B(n6655), .Z(n6654) );
  XOR U6606 ( .A(n6656), .B(n6653), .Z(n6655) );
  AND U6607 ( .A(n6553), .B(n6556), .Z(n6609) );
  XOR U6608 ( .A(n6657), .B(n6636), .Z(n6556) );
  XNOR U6609 ( .A(p_input[1024]), .B(p_input[496]), .Z(n6636) );
  XOR U6610 ( .A(n6624), .B(n6623), .Z(n6657) );
  XNOR U6611 ( .A(n6658), .B(n6630), .Z(n6623) );
  XNOR U6612 ( .A(n6619), .B(n6618), .Z(n6630) );
  XOR U6613 ( .A(n6659), .B(n6615), .Z(n6618) );
  XOR U6614 ( .A(p_input[1034]), .B(p_input[506]), .Z(n6615) );
  XNOR U6615 ( .A(p_input[1035]), .B(p_input[507]), .Z(n6659) );
  XOR U6616 ( .A(p_input[1036]), .B(p_input[508]), .Z(n6619) );
  XNOR U6617 ( .A(n6629), .B(n6620), .Z(n6658) );
  XNOR U6618 ( .A(n3298), .B(p_input[497]), .Z(n6620) );
  XOR U6619 ( .A(n6660), .B(n6635), .Z(n6629) );
  XNOR U6620 ( .A(p_input[1039]), .B(p_input[511]), .Z(n6635) );
  XOR U6621 ( .A(n6626), .B(n6634), .Z(n6660) );
  XOR U6622 ( .A(n6661), .B(n6631), .Z(n6634) );
  XOR U6623 ( .A(p_input[1037]), .B(p_input[509]), .Z(n6631) );
  XNOR U6624 ( .A(p_input[1038]), .B(p_input[510]), .Z(n6661) );
  XOR U6625 ( .A(p_input[1033]), .B(p_input[505]), .Z(n6626) );
  XNOR U6626 ( .A(n6642), .B(n6641), .Z(n6624) );
  XNOR U6627 ( .A(n6662), .B(n6647), .Z(n6641) );
  XOR U6628 ( .A(p_input[1032]), .B(p_input[504]), .Z(n6647) );
  XOR U6629 ( .A(n6638), .B(n6646), .Z(n6662) );
  XOR U6630 ( .A(n6663), .B(n6643), .Z(n6646) );
  XOR U6631 ( .A(p_input[1030]), .B(p_input[502]), .Z(n6643) );
  XNOR U6632 ( .A(p_input[1031]), .B(p_input[503]), .Z(n6663) );
  XOR U6633 ( .A(p_input[1026]), .B(p_input[498]), .Z(n6638) );
  XNOR U6634 ( .A(n6652), .B(n6651), .Z(n6642) );
  XOR U6635 ( .A(n6664), .B(n6648), .Z(n6651) );
  XOR U6636 ( .A(p_input[1027]), .B(p_input[499]), .Z(n6648) );
  XNOR U6637 ( .A(p_input[1028]), .B(p_input[500]), .Z(n6664) );
  XOR U6638 ( .A(p_input[1029]), .B(p_input[501]), .Z(n6652) );
  XOR U6639 ( .A(n6665), .B(n6666), .Z(n6553) );
  AND U6640 ( .A(n131), .B(n6667), .Z(n6666) );
  XNOR U6641 ( .A(n6668), .B(n6665), .Z(n6667) );
  XNOR U6642 ( .A(n6669), .B(n6670), .Z(n131) );
  AND U6643 ( .A(n6671), .B(n6672), .Z(n6670) );
  XOR U6644 ( .A(n6566), .B(n6669), .Z(n6672) );
  AND U6645 ( .A(n6673), .B(n6674), .Z(n6566) );
  XNOR U6646 ( .A(n6563), .B(n6669), .Z(n6671) );
  XOR U6647 ( .A(n6675), .B(n6676), .Z(n6563) );
  AND U6648 ( .A(n135), .B(n6677), .Z(n6676) );
  XOR U6649 ( .A(n6678), .B(n6675), .Z(n6677) );
  XOR U6650 ( .A(n6679), .B(n6680), .Z(n6669) );
  AND U6651 ( .A(n6681), .B(n6682), .Z(n6680) );
  XNOR U6652 ( .A(n6679), .B(n6673), .Z(n6682) );
  IV U6653 ( .A(n6581), .Z(n6673) );
  XOR U6654 ( .A(n6683), .B(n6684), .Z(n6581) );
  XOR U6655 ( .A(n6685), .B(n6674), .Z(n6684) );
  AND U6656 ( .A(n6608), .B(n6686), .Z(n6674) );
  AND U6657 ( .A(n6687), .B(n6688), .Z(n6685) );
  XOR U6658 ( .A(n6689), .B(n6683), .Z(n6687) );
  XNOR U6659 ( .A(n6578), .B(n6679), .Z(n6681) );
  XOR U6660 ( .A(n6690), .B(n6691), .Z(n6578) );
  AND U6661 ( .A(n135), .B(n6692), .Z(n6691) );
  XOR U6662 ( .A(n6693), .B(n6690), .Z(n6692) );
  XOR U6663 ( .A(n6694), .B(n6695), .Z(n6679) );
  AND U6664 ( .A(n6696), .B(n6697), .Z(n6695) );
  XNOR U6665 ( .A(n6694), .B(n6608), .Z(n6697) );
  XOR U6666 ( .A(n6698), .B(n6688), .Z(n6608) );
  XNOR U6667 ( .A(n6699), .B(n6683), .Z(n6688) );
  XOR U6668 ( .A(n6700), .B(n6701), .Z(n6683) );
  AND U6669 ( .A(n6702), .B(n6703), .Z(n6701) );
  XOR U6670 ( .A(n6704), .B(n6700), .Z(n6702) );
  XNOR U6671 ( .A(n6705), .B(n6706), .Z(n6699) );
  AND U6672 ( .A(n6707), .B(n6708), .Z(n6706) );
  XOR U6673 ( .A(n6705), .B(n6709), .Z(n6707) );
  XNOR U6674 ( .A(n6689), .B(n6686), .Z(n6698) );
  AND U6675 ( .A(n6710), .B(n6711), .Z(n6686) );
  XOR U6676 ( .A(n6712), .B(n6713), .Z(n6689) );
  AND U6677 ( .A(n6714), .B(n6715), .Z(n6713) );
  XOR U6678 ( .A(n6712), .B(n6716), .Z(n6714) );
  XNOR U6679 ( .A(n6605), .B(n6694), .Z(n6696) );
  XOR U6680 ( .A(n6717), .B(n6718), .Z(n6605) );
  AND U6681 ( .A(n135), .B(n6719), .Z(n6718) );
  XNOR U6682 ( .A(n6720), .B(n6717), .Z(n6719) );
  XOR U6683 ( .A(n6721), .B(n6722), .Z(n6694) );
  AND U6684 ( .A(n6723), .B(n6724), .Z(n6722) );
  XNOR U6685 ( .A(n6721), .B(n6710), .Z(n6724) );
  IV U6686 ( .A(n6656), .Z(n6710) );
  XNOR U6687 ( .A(n6725), .B(n6703), .Z(n6656) );
  XNOR U6688 ( .A(n6726), .B(n6709), .Z(n6703) );
  XOR U6689 ( .A(n6727), .B(n6728), .Z(n6709) );
  NOR U6690 ( .A(n6729), .B(n6730), .Z(n6728) );
  XNOR U6691 ( .A(n6727), .B(n6731), .Z(n6729) );
  XNOR U6692 ( .A(n6708), .B(n6700), .Z(n6726) );
  XOR U6693 ( .A(n6732), .B(n6733), .Z(n6700) );
  AND U6694 ( .A(n6734), .B(n6735), .Z(n6733) );
  XNOR U6695 ( .A(n6732), .B(n6736), .Z(n6734) );
  XNOR U6696 ( .A(n6737), .B(n6705), .Z(n6708) );
  XOR U6697 ( .A(n6738), .B(n6739), .Z(n6705) );
  AND U6698 ( .A(n6740), .B(n6741), .Z(n6739) );
  XOR U6699 ( .A(n6738), .B(n6742), .Z(n6740) );
  XNOR U6700 ( .A(n6743), .B(n6744), .Z(n6737) );
  NOR U6701 ( .A(n6745), .B(n6746), .Z(n6744) );
  XOR U6702 ( .A(n6743), .B(n6747), .Z(n6745) );
  XNOR U6703 ( .A(n6704), .B(n6711), .Z(n6725) );
  NOR U6704 ( .A(n6668), .B(n6748), .Z(n6711) );
  XOR U6705 ( .A(n6716), .B(n6715), .Z(n6704) );
  XNOR U6706 ( .A(n6749), .B(n6712), .Z(n6715) );
  XOR U6707 ( .A(n6750), .B(n6751), .Z(n6712) );
  AND U6708 ( .A(n6752), .B(n6753), .Z(n6751) );
  XOR U6709 ( .A(n6750), .B(n6754), .Z(n6752) );
  XNOR U6710 ( .A(n6755), .B(n6756), .Z(n6749) );
  NOR U6711 ( .A(n6757), .B(n6758), .Z(n6756) );
  XNOR U6712 ( .A(n6755), .B(n6759), .Z(n6757) );
  XOR U6713 ( .A(n6760), .B(n6761), .Z(n6716) );
  NOR U6714 ( .A(n6762), .B(n6763), .Z(n6761) );
  XNOR U6715 ( .A(n6760), .B(n6764), .Z(n6762) );
  XNOR U6716 ( .A(n6653), .B(n6721), .Z(n6723) );
  XOR U6717 ( .A(n6765), .B(n6766), .Z(n6653) );
  AND U6718 ( .A(n135), .B(n6767), .Z(n6766) );
  XOR U6719 ( .A(n6768), .B(n6765), .Z(n6767) );
  AND U6720 ( .A(n6665), .B(n6668), .Z(n6721) );
  XOR U6721 ( .A(n6769), .B(n6748), .Z(n6668) );
  XNOR U6722 ( .A(p_input[1024]), .B(p_input[512]), .Z(n6748) );
  XOR U6723 ( .A(n6736), .B(n6735), .Z(n6769) );
  XNOR U6724 ( .A(n6770), .B(n6742), .Z(n6735) );
  XNOR U6725 ( .A(n6731), .B(n6730), .Z(n6742) );
  XOR U6726 ( .A(n6771), .B(n6727), .Z(n6730) );
  XOR U6727 ( .A(p_input[1034]), .B(p_input[522]), .Z(n6727) );
  XNOR U6728 ( .A(p_input[1035]), .B(p_input[523]), .Z(n6771) );
  XOR U6729 ( .A(p_input[1036]), .B(p_input[524]), .Z(n6731) );
  XNOR U6730 ( .A(n6741), .B(n6732), .Z(n6770) );
  XNOR U6731 ( .A(n3298), .B(p_input[513]), .Z(n6732) );
  XOR U6732 ( .A(n6772), .B(n6747), .Z(n6741) );
  XNOR U6733 ( .A(p_input[1039]), .B(p_input[527]), .Z(n6747) );
  XOR U6734 ( .A(n6738), .B(n6746), .Z(n6772) );
  XOR U6735 ( .A(n6773), .B(n6743), .Z(n6746) );
  XOR U6736 ( .A(p_input[1037]), .B(p_input[525]), .Z(n6743) );
  XNOR U6737 ( .A(p_input[1038]), .B(p_input[526]), .Z(n6773) );
  XOR U6738 ( .A(p_input[1033]), .B(p_input[521]), .Z(n6738) );
  XNOR U6739 ( .A(n6754), .B(n6753), .Z(n6736) );
  XNOR U6740 ( .A(n6774), .B(n6759), .Z(n6753) );
  XOR U6741 ( .A(p_input[1032]), .B(p_input[520]), .Z(n6759) );
  XOR U6742 ( .A(n6750), .B(n6758), .Z(n6774) );
  XOR U6743 ( .A(n6775), .B(n6755), .Z(n6758) );
  XOR U6744 ( .A(p_input[1030]), .B(p_input[518]), .Z(n6755) );
  XNOR U6745 ( .A(p_input[1031]), .B(p_input[519]), .Z(n6775) );
  XOR U6746 ( .A(p_input[1026]), .B(p_input[514]), .Z(n6750) );
  XNOR U6747 ( .A(n6764), .B(n6763), .Z(n6754) );
  XOR U6748 ( .A(n6776), .B(n6760), .Z(n6763) );
  XOR U6749 ( .A(p_input[1027]), .B(p_input[515]), .Z(n6760) );
  XNOR U6750 ( .A(p_input[1028]), .B(p_input[516]), .Z(n6776) );
  XOR U6751 ( .A(p_input[1029]), .B(p_input[517]), .Z(n6764) );
  XOR U6752 ( .A(n6777), .B(n6778), .Z(n6665) );
  AND U6753 ( .A(n135), .B(n6779), .Z(n6778) );
  XNOR U6754 ( .A(n6780), .B(n6777), .Z(n6779) );
  XNOR U6755 ( .A(n6781), .B(n6782), .Z(n135) );
  AND U6756 ( .A(n6783), .B(n6784), .Z(n6782) );
  XOR U6757 ( .A(n6678), .B(n6781), .Z(n6784) );
  AND U6758 ( .A(n6785), .B(n6786), .Z(n6678) );
  XNOR U6759 ( .A(n6675), .B(n6781), .Z(n6783) );
  XOR U6760 ( .A(n6787), .B(n6788), .Z(n6675) );
  AND U6761 ( .A(n139), .B(n6789), .Z(n6788) );
  XOR U6762 ( .A(n6790), .B(n6787), .Z(n6789) );
  XOR U6763 ( .A(n6791), .B(n6792), .Z(n6781) );
  AND U6764 ( .A(n6793), .B(n6794), .Z(n6792) );
  XNOR U6765 ( .A(n6791), .B(n6785), .Z(n6794) );
  IV U6766 ( .A(n6693), .Z(n6785) );
  XOR U6767 ( .A(n6795), .B(n6796), .Z(n6693) );
  XOR U6768 ( .A(n6797), .B(n6786), .Z(n6796) );
  AND U6769 ( .A(n6720), .B(n6798), .Z(n6786) );
  AND U6770 ( .A(n6799), .B(n6800), .Z(n6797) );
  XOR U6771 ( .A(n6801), .B(n6795), .Z(n6799) );
  XNOR U6772 ( .A(n6690), .B(n6791), .Z(n6793) );
  XOR U6773 ( .A(n6802), .B(n6803), .Z(n6690) );
  AND U6774 ( .A(n139), .B(n6804), .Z(n6803) );
  XOR U6775 ( .A(n6805), .B(n6802), .Z(n6804) );
  XOR U6776 ( .A(n6806), .B(n6807), .Z(n6791) );
  AND U6777 ( .A(n6808), .B(n6809), .Z(n6807) );
  XNOR U6778 ( .A(n6806), .B(n6720), .Z(n6809) );
  XOR U6779 ( .A(n6810), .B(n6800), .Z(n6720) );
  XNOR U6780 ( .A(n6811), .B(n6795), .Z(n6800) );
  XOR U6781 ( .A(n6812), .B(n6813), .Z(n6795) );
  AND U6782 ( .A(n6814), .B(n6815), .Z(n6813) );
  XOR U6783 ( .A(n6816), .B(n6812), .Z(n6814) );
  XNOR U6784 ( .A(n6817), .B(n6818), .Z(n6811) );
  AND U6785 ( .A(n6819), .B(n6820), .Z(n6818) );
  XOR U6786 ( .A(n6817), .B(n6821), .Z(n6819) );
  XNOR U6787 ( .A(n6801), .B(n6798), .Z(n6810) );
  AND U6788 ( .A(n6822), .B(n6823), .Z(n6798) );
  XOR U6789 ( .A(n6824), .B(n6825), .Z(n6801) );
  AND U6790 ( .A(n6826), .B(n6827), .Z(n6825) );
  XOR U6791 ( .A(n6824), .B(n6828), .Z(n6826) );
  XNOR U6792 ( .A(n6717), .B(n6806), .Z(n6808) );
  XOR U6793 ( .A(n6829), .B(n6830), .Z(n6717) );
  AND U6794 ( .A(n139), .B(n6831), .Z(n6830) );
  XNOR U6795 ( .A(n6832), .B(n6829), .Z(n6831) );
  XOR U6796 ( .A(n6833), .B(n6834), .Z(n6806) );
  AND U6797 ( .A(n6835), .B(n6836), .Z(n6834) );
  XNOR U6798 ( .A(n6833), .B(n6822), .Z(n6836) );
  IV U6799 ( .A(n6768), .Z(n6822) );
  XNOR U6800 ( .A(n6837), .B(n6815), .Z(n6768) );
  XNOR U6801 ( .A(n6838), .B(n6821), .Z(n6815) );
  XOR U6802 ( .A(n6839), .B(n6840), .Z(n6821) );
  NOR U6803 ( .A(n6841), .B(n6842), .Z(n6840) );
  XNOR U6804 ( .A(n6839), .B(n6843), .Z(n6841) );
  XNOR U6805 ( .A(n6820), .B(n6812), .Z(n6838) );
  XOR U6806 ( .A(n6844), .B(n6845), .Z(n6812) );
  AND U6807 ( .A(n6846), .B(n6847), .Z(n6845) );
  XNOR U6808 ( .A(n6844), .B(n6848), .Z(n6846) );
  XNOR U6809 ( .A(n6849), .B(n6817), .Z(n6820) );
  XOR U6810 ( .A(n6850), .B(n6851), .Z(n6817) );
  AND U6811 ( .A(n6852), .B(n6853), .Z(n6851) );
  XOR U6812 ( .A(n6850), .B(n6854), .Z(n6852) );
  XNOR U6813 ( .A(n6855), .B(n6856), .Z(n6849) );
  NOR U6814 ( .A(n6857), .B(n6858), .Z(n6856) );
  XOR U6815 ( .A(n6855), .B(n6859), .Z(n6857) );
  XNOR U6816 ( .A(n6816), .B(n6823), .Z(n6837) );
  NOR U6817 ( .A(n6780), .B(n6860), .Z(n6823) );
  XOR U6818 ( .A(n6828), .B(n6827), .Z(n6816) );
  XNOR U6819 ( .A(n6861), .B(n6824), .Z(n6827) );
  XOR U6820 ( .A(n6862), .B(n6863), .Z(n6824) );
  AND U6821 ( .A(n6864), .B(n6865), .Z(n6863) );
  XOR U6822 ( .A(n6862), .B(n6866), .Z(n6864) );
  XNOR U6823 ( .A(n6867), .B(n6868), .Z(n6861) );
  NOR U6824 ( .A(n6869), .B(n6870), .Z(n6868) );
  XNOR U6825 ( .A(n6867), .B(n6871), .Z(n6869) );
  XOR U6826 ( .A(n6872), .B(n6873), .Z(n6828) );
  NOR U6827 ( .A(n6874), .B(n6875), .Z(n6873) );
  XNOR U6828 ( .A(n6872), .B(n6876), .Z(n6874) );
  XNOR U6829 ( .A(n6765), .B(n6833), .Z(n6835) );
  XOR U6830 ( .A(n6877), .B(n6878), .Z(n6765) );
  AND U6831 ( .A(n139), .B(n6879), .Z(n6878) );
  XOR U6832 ( .A(n6880), .B(n6877), .Z(n6879) );
  AND U6833 ( .A(n6777), .B(n6780), .Z(n6833) );
  XOR U6834 ( .A(n6881), .B(n6860), .Z(n6780) );
  XNOR U6835 ( .A(p_input[1024]), .B(p_input[528]), .Z(n6860) );
  XOR U6836 ( .A(n6848), .B(n6847), .Z(n6881) );
  XNOR U6837 ( .A(n6882), .B(n6854), .Z(n6847) );
  XNOR U6838 ( .A(n6843), .B(n6842), .Z(n6854) );
  XOR U6839 ( .A(n6883), .B(n6839), .Z(n6842) );
  XOR U6840 ( .A(p_input[1034]), .B(p_input[538]), .Z(n6839) );
  XNOR U6841 ( .A(p_input[1035]), .B(p_input[539]), .Z(n6883) );
  XOR U6842 ( .A(p_input[1036]), .B(p_input[540]), .Z(n6843) );
  XNOR U6843 ( .A(n6853), .B(n6844), .Z(n6882) );
  XNOR U6844 ( .A(n3298), .B(p_input[529]), .Z(n6844) );
  XOR U6845 ( .A(n6884), .B(n6859), .Z(n6853) );
  XNOR U6846 ( .A(p_input[1039]), .B(p_input[543]), .Z(n6859) );
  XOR U6847 ( .A(n6850), .B(n6858), .Z(n6884) );
  XOR U6848 ( .A(n6885), .B(n6855), .Z(n6858) );
  XOR U6849 ( .A(p_input[1037]), .B(p_input[541]), .Z(n6855) );
  XNOR U6850 ( .A(p_input[1038]), .B(p_input[542]), .Z(n6885) );
  XOR U6851 ( .A(p_input[1033]), .B(p_input[537]), .Z(n6850) );
  XNOR U6852 ( .A(n6866), .B(n6865), .Z(n6848) );
  XNOR U6853 ( .A(n6886), .B(n6871), .Z(n6865) );
  XOR U6854 ( .A(p_input[1032]), .B(p_input[536]), .Z(n6871) );
  XOR U6855 ( .A(n6862), .B(n6870), .Z(n6886) );
  XOR U6856 ( .A(n6887), .B(n6867), .Z(n6870) );
  XOR U6857 ( .A(p_input[1030]), .B(p_input[534]), .Z(n6867) );
  XNOR U6858 ( .A(p_input[1031]), .B(p_input[535]), .Z(n6887) );
  XOR U6859 ( .A(p_input[1026]), .B(p_input[530]), .Z(n6862) );
  XNOR U6860 ( .A(n6876), .B(n6875), .Z(n6866) );
  XOR U6861 ( .A(n6888), .B(n6872), .Z(n6875) );
  XOR U6862 ( .A(p_input[1027]), .B(p_input[531]), .Z(n6872) );
  XNOR U6863 ( .A(p_input[1028]), .B(p_input[532]), .Z(n6888) );
  XOR U6864 ( .A(p_input[1029]), .B(p_input[533]), .Z(n6876) );
  XOR U6865 ( .A(n6889), .B(n6890), .Z(n6777) );
  AND U6866 ( .A(n139), .B(n6891), .Z(n6890) );
  XNOR U6867 ( .A(n6892), .B(n6889), .Z(n6891) );
  XNOR U6868 ( .A(n6893), .B(n6894), .Z(n139) );
  AND U6869 ( .A(n6895), .B(n6896), .Z(n6894) );
  XOR U6870 ( .A(n6790), .B(n6893), .Z(n6896) );
  AND U6871 ( .A(n6897), .B(n6898), .Z(n6790) );
  XNOR U6872 ( .A(n6787), .B(n6893), .Z(n6895) );
  XOR U6873 ( .A(n6899), .B(n6900), .Z(n6787) );
  AND U6874 ( .A(n143), .B(n6901), .Z(n6900) );
  XOR U6875 ( .A(n6902), .B(n6899), .Z(n6901) );
  XOR U6876 ( .A(n6903), .B(n6904), .Z(n6893) );
  AND U6877 ( .A(n6905), .B(n6906), .Z(n6904) );
  XNOR U6878 ( .A(n6903), .B(n6897), .Z(n6906) );
  IV U6879 ( .A(n6805), .Z(n6897) );
  XOR U6880 ( .A(n6907), .B(n6908), .Z(n6805) );
  XOR U6881 ( .A(n6909), .B(n6898), .Z(n6908) );
  AND U6882 ( .A(n6832), .B(n6910), .Z(n6898) );
  AND U6883 ( .A(n6911), .B(n6912), .Z(n6909) );
  XOR U6884 ( .A(n6913), .B(n6907), .Z(n6911) );
  XNOR U6885 ( .A(n6802), .B(n6903), .Z(n6905) );
  XOR U6886 ( .A(n6914), .B(n6915), .Z(n6802) );
  AND U6887 ( .A(n143), .B(n6916), .Z(n6915) );
  XOR U6888 ( .A(n6917), .B(n6914), .Z(n6916) );
  XOR U6889 ( .A(n6918), .B(n6919), .Z(n6903) );
  AND U6890 ( .A(n6920), .B(n6921), .Z(n6919) );
  XNOR U6891 ( .A(n6918), .B(n6832), .Z(n6921) );
  XOR U6892 ( .A(n6922), .B(n6912), .Z(n6832) );
  XNOR U6893 ( .A(n6923), .B(n6907), .Z(n6912) );
  XOR U6894 ( .A(n6924), .B(n6925), .Z(n6907) );
  AND U6895 ( .A(n6926), .B(n6927), .Z(n6925) );
  XOR U6896 ( .A(n6928), .B(n6924), .Z(n6926) );
  XNOR U6897 ( .A(n6929), .B(n6930), .Z(n6923) );
  AND U6898 ( .A(n6931), .B(n6932), .Z(n6930) );
  XOR U6899 ( .A(n6929), .B(n6933), .Z(n6931) );
  XNOR U6900 ( .A(n6913), .B(n6910), .Z(n6922) );
  AND U6901 ( .A(n6934), .B(n6935), .Z(n6910) );
  XOR U6902 ( .A(n6936), .B(n6937), .Z(n6913) );
  AND U6903 ( .A(n6938), .B(n6939), .Z(n6937) );
  XOR U6904 ( .A(n6936), .B(n6940), .Z(n6938) );
  XNOR U6905 ( .A(n6829), .B(n6918), .Z(n6920) );
  XOR U6906 ( .A(n6941), .B(n6942), .Z(n6829) );
  AND U6907 ( .A(n143), .B(n6943), .Z(n6942) );
  XNOR U6908 ( .A(n6944), .B(n6941), .Z(n6943) );
  XOR U6909 ( .A(n6945), .B(n6946), .Z(n6918) );
  AND U6910 ( .A(n6947), .B(n6948), .Z(n6946) );
  XNOR U6911 ( .A(n6945), .B(n6934), .Z(n6948) );
  IV U6912 ( .A(n6880), .Z(n6934) );
  XNOR U6913 ( .A(n6949), .B(n6927), .Z(n6880) );
  XNOR U6914 ( .A(n6950), .B(n6933), .Z(n6927) );
  XOR U6915 ( .A(n6951), .B(n6952), .Z(n6933) );
  NOR U6916 ( .A(n6953), .B(n6954), .Z(n6952) );
  XNOR U6917 ( .A(n6951), .B(n6955), .Z(n6953) );
  XNOR U6918 ( .A(n6932), .B(n6924), .Z(n6950) );
  XOR U6919 ( .A(n6956), .B(n6957), .Z(n6924) );
  AND U6920 ( .A(n6958), .B(n6959), .Z(n6957) );
  XNOR U6921 ( .A(n6956), .B(n6960), .Z(n6958) );
  XNOR U6922 ( .A(n6961), .B(n6929), .Z(n6932) );
  XOR U6923 ( .A(n6962), .B(n6963), .Z(n6929) );
  AND U6924 ( .A(n6964), .B(n6965), .Z(n6963) );
  XOR U6925 ( .A(n6962), .B(n6966), .Z(n6964) );
  XNOR U6926 ( .A(n6967), .B(n6968), .Z(n6961) );
  NOR U6927 ( .A(n6969), .B(n6970), .Z(n6968) );
  XOR U6928 ( .A(n6967), .B(n6971), .Z(n6969) );
  XNOR U6929 ( .A(n6928), .B(n6935), .Z(n6949) );
  NOR U6930 ( .A(n6892), .B(n6972), .Z(n6935) );
  XOR U6931 ( .A(n6940), .B(n6939), .Z(n6928) );
  XNOR U6932 ( .A(n6973), .B(n6936), .Z(n6939) );
  XOR U6933 ( .A(n6974), .B(n6975), .Z(n6936) );
  AND U6934 ( .A(n6976), .B(n6977), .Z(n6975) );
  XOR U6935 ( .A(n6974), .B(n6978), .Z(n6976) );
  XNOR U6936 ( .A(n6979), .B(n6980), .Z(n6973) );
  NOR U6937 ( .A(n6981), .B(n6982), .Z(n6980) );
  XNOR U6938 ( .A(n6979), .B(n6983), .Z(n6981) );
  XOR U6939 ( .A(n6984), .B(n6985), .Z(n6940) );
  NOR U6940 ( .A(n6986), .B(n6987), .Z(n6985) );
  XNOR U6941 ( .A(n6984), .B(n6988), .Z(n6986) );
  XNOR U6942 ( .A(n6877), .B(n6945), .Z(n6947) );
  XOR U6943 ( .A(n6989), .B(n6990), .Z(n6877) );
  AND U6944 ( .A(n143), .B(n6991), .Z(n6990) );
  XOR U6945 ( .A(n6992), .B(n6989), .Z(n6991) );
  AND U6946 ( .A(n6889), .B(n6892), .Z(n6945) );
  XOR U6947 ( .A(n6993), .B(n6972), .Z(n6892) );
  XNOR U6948 ( .A(p_input[1024]), .B(p_input[544]), .Z(n6972) );
  XOR U6949 ( .A(n6960), .B(n6959), .Z(n6993) );
  XNOR U6950 ( .A(n6994), .B(n6966), .Z(n6959) );
  XNOR U6951 ( .A(n6955), .B(n6954), .Z(n6966) );
  XOR U6952 ( .A(n6995), .B(n6951), .Z(n6954) );
  XOR U6953 ( .A(p_input[1034]), .B(p_input[554]), .Z(n6951) );
  XNOR U6954 ( .A(p_input[1035]), .B(p_input[555]), .Z(n6995) );
  XOR U6955 ( .A(p_input[1036]), .B(p_input[556]), .Z(n6955) );
  XNOR U6956 ( .A(n6965), .B(n6956), .Z(n6994) );
  XNOR U6957 ( .A(n3298), .B(p_input[545]), .Z(n6956) );
  XOR U6958 ( .A(n6996), .B(n6971), .Z(n6965) );
  XNOR U6959 ( .A(p_input[1039]), .B(p_input[559]), .Z(n6971) );
  XOR U6960 ( .A(n6962), .B(n6970), .Z(n6996) );
  XOR U6961 ( .A(n6997), .B(n6967), .Z(n6970) );
  XOR U6962 ( .A(p_input[1037]), .B(p_input[557]), .Z(n6967) );
  XNOR U6963 ( .A(p_input[1038]), .B(p_input[558]), .Z(n6997) );
  XOR U6964 ( .A(p_input[1033]), .B(p_input[553]), .Z(n6962) );
  XNOR U6965 ( .A(n6978), .B(n6977), .Z(n6960) );
  XNOR U6966 ( .A(n6998), .B(n6983), .Z(n6977) );
  XOR U6967 ( .A(p_input[1032]), .B(p_input[552]), .Z(n6983) );
  XOR U6968 ( .A(n6974), .B(n6982), .Z(n6998) );
  XOR U6969 ( .A(n6999), .B(n6979), .Z(n6982) );
  XOR U6970 ( .A(p_input[1030]), .B(p_input[550]), .Z(n6979) );
  XNOR U6971 ( .A(p_input[1031]), .B(p_input[551]), .Z(n6999) );
  XOR U6972 ( .A(p_input[1026]), .B(p_input[546]), .Z(n6974) );
  XNOR U6973 ( .A(n6988), .B(n6987), .Z(n6978) );
  XOR U6974 ( .A(n7000), .B(n6984), .Z(n6987) );
  XOR U6975 ( .A(p_input[1027]), .B(p_input[547]), .Z(n6984) );
  XNOR U6976 ( .A(p_input[1028]), .B(p_input[548]), .Z(n7000) );
  XOR U6977 ( .A(p_input[1029]), .B(p_input[549]), .Z(n6988) );
  XOR U6978 ( .A(n7001), .B(n7002), .Z(n6889) );
  AND U6979 ( .A(n143), .B(n7003), .Z(n7002) );
  XNOR U6980 ( .A(n7004), .B(n7001), .Z(n7003) );
  XNOR U6981 ( .A(n7005), .B(n7006), .Z(n143) );
  AND U6982 ( .A(n7007), .B(n7008), .Z(n7006) );
  XOR U6983 ( .A(n6902), .B(n7005), .Z(n7008) );
  AND U6984 ( .A(n7009), .B(n7010), .Z(n6902) );
  XNOR U6985 ( .A(n6899), .B(n7005), .Z(n7007) );
  XOR U6986 ( .A(n7011), .B(n7012), .Z(n6899) );
  AND U6987 ( .A(n147), .B(n7013), .Z(n7012) );
  XOR U6988 ( .A(n7014), .B(n7011), .Z(n7013) );
  XOR U6989 ( .A(n7015), .B(n7016), .Z(n7005) );
  AND U6990 ( .A(n7017), .B(n7018), .Z(n7016) );
  XNOR U6991 ( .A(n7015), .B(n7009), .Z(n7018) );
  IV U6992 ( .A(n6917), .Z(n7009) );
  XOR U6993 ( .A(n7019), .B(n7020), .Z(n6917) );
  XOR U6994 ( .A(n7021), .B(n7010), .Z(n7020) );
  AND U6995 ( .A(n6944), .B(n7022), .Z(n7010) );
  AND U6996 ( .A(n7023), .B(n7024), .Z(n7021) );
  XOR U6997 ( .A(n7025), .B(n7019), .Z(n7023) );
  XNOR U6998 ( .A(n6914), .B(n7015), .Z(n7017) );
  XOR U6999 ( .A(n7026), .B(n7027), .Z(n6914) );
  AND U7000 ( .A(n147), .B(n7028), .Z(n7027) );
  XOR U7001 ( .A(n7029), .B(n7026), .Z(n7028) );
  XOR U7002 ( .A(n7030), .B(n7031), .Z(n7015) );
  AND U7003 ( .A(n7032), .B(n7033), .Z(n7031) );
  XNOR U7004 ( .A(n7030), .B(n6944), .Z(n7033) );
  XOR U7005 ( .A(n7034), .B(n7024), .Z(n6944) );
  XNOR U7006 ( .A(n7035), .B(n7019), .Z(n7024) );
  XOR U7007 ( .A(n7036), .B(n7037), .Z(n7019) );
  AND U7008 ( .A(n7038), .B(n7039), .Z(n7037) );
  XOR U7009 ( .A(n7040), .B(n7036), .Z(n7038) );
  XNOR U7010 ( .A(n7041), .B(n7042), .Z(n7035) );
  AND U7011 ( .A(n7043), .B(n7044), .Z(n7042) );
  XOR U7012 ( .A(n7041), .B(n7045), .Z(n7043) );
  XNOR U7013 ( .A(n7025), .B(n7022), .Z(n7034) );
  AND U7014 ( .A(n7046), .B(n7047), .Z(n7022) );
  XOR U7015 ( .A(n7048), .B(n7049), .Z(n7025) );
  AND U7016 ( .A(n7050), .B(n7051), .Z(n7049) );
  XOR U7017 ( .A(n7048), .B(n7052), .Z(n7050) );
  XNOR U7018 ( .A(n6941), .B(n7030), .Z(n7032) );
  XOR U7019 ( .A(n7053), .B(n7054), .Z(n6941) );
  AND U7020 ( .A(n147), .B(n7055), .Z(n7054) );
  XNOR U7021 ( .A(n7056), .B(n7053), .Z(n7055) );
  XOR U7022 ( .A(n7057), .B(n7058), .Z(n7030) );
  AND U7023 ( .A(n7059), .B(n7060), .Z(n7058) );
  XNOR U7024 ( .A(n7057), .B(n7046), .Z(n7060) );
  IV U7025 ( .A(n6992), .Z(n7046) );
  XNOR U7026 ( .A(n7061), .B(n7039), .Z(n6992) );
  XNOR U7027 ( .A(n7062), .B(n7045), .Z(n7039) );
  XOR U7028 ( .A(n7063), .B(n7064), .Z(n7045) );
  NOR U7029 ( .A(n7065), .B(n7066), .Z(n7064) );
  XNOR U7030 ( .A(n7063), .B(n7067), .Z(n7065) );
  XNOR U7031 ( .A(n7044), .B(n7036), .Z(n7062) );
  XOR U7032 ( .A(n7068), .B(n7069), .Z(n7036) );
  AND U7033 ( .A(n7070), .B(n7071), .Z(n7069) );
  XNOR U7034 ( .A(n7068), .B(n7072), .Z(n7070) );
  XNOR U7035 ( .A(n7073), .B(n7041), .Z(n7044) );
  XOR U7036 ( .A(n7074), .B(n7075), .Z(n7041) );
  AND U7037 ( .A(n7076), .B(n7077), .Z(n7075) );
  XOR U7038 ( .A(n7074), .B(n7078), .Z(n7076) );
  XNOR U7039 ( .A(n7079), .B(n7080), .Z(n7073) );
  NOR U7040 ( .A(n7081), .B(n7082), .Z(n7080) );
  XOR U7041 ( .A(n7079), .B(n7083), .Z(n7081) );
  XNOR U7042 ( .A(n7040), .B(n7047), .Z(n7061) );
  NOR U7043 ( .A(n7004), .B(n7084), .Z(n7047) );
  XOR U7044 ( .A(n7052), .B(n7051), .Z(n7040) );
  XNOR U7045 ( .A(n7085), .B(n7048), .Z(n7051) );
  XOR U7046 ( .A(n7086), .B(n7087), .Z(n7048) );
  AND U7047 ( .A(n7088), .B(n7089), .Z(n7087) );
  XOR U7048 ( .A(n7086), .B(n7090), .Z(n7088) );
  XNOR U7049 ( .A(n7091), .B(n7092), .Z(n7085) );
  NOR U7050 ( .A(n7093), .B(n7094), .Z(n7092) );
  XNOR U7051 ( .A(n7091), .B(n7095), .Z(n7093) );
  XOR U7052 ( .A(n7096), .B(n7097), .Z(n7052) );
  NOR U7053 ( .A(n7098), .B(n7099), .Z(n7097) );
  XNOR U7054 ( .A(n7096), .B(n7100), .Z(n7098) );
  XNOR U7055 ( .A(n6989), .B(n7057), .Z(n7059) );
  XOR U7056 ( .A(n7101), .B(n7102), .Z(n6989) );
  AND U7057 ( .A(n147), .B(n7103), .Z(n7102) );
  XOR U7058 ( .A(n7104), .B(n7101), .Z(n7103) );
  AND U7059 ( .A(n7001), .B(n7004), .Z(n7057) );
  XOR U7060 ( .A(n7105), .B(n7084), .Z(n7004) );
  XNOR U7061 ( .A(p_input[1024]), .B(p_input[560]), .Z(n7084) );
  XOR U7062 ( .A(n7072), .B(n7071), .Z(n7105) );
  XNOR U7063 ( .A(n7106), .B(n7078), .Z(n7071) );
  XNOR U7064 ( .A(n7067), .B(n7066), .Z(n7078) );
  XOR U7065 ( .A(n7107), .B(n7063), .Z(n7066) );
  XOR U7066 ( .A(p_input[1034]), .B(p_input[570]), .Z(n7063) );
  XNOR U7067 ( .A(p_input[1035]), .B(p_input[571]), .Z(n7107) );
  XOR U7068 ( .A(p_input[1036]), .B(p_input[572]), .Z(n7067) );
  XNOR U7069 ( .A(n7077), .B(n7068), .Z(n7106) );
  XNOR U7070 ( .A(n3298), .B(p_input[561]), .Z(n7068) );
  XOR U7071 ( .A(n7108), .B(n7083), .Z(n7077) );
  XNOR U7072 ( .A(p_input[1039]), .B(p_input[575]), .Z(n7083) );
  XOR U7073 ( .A(n7074), .B(n7082), .Z(n7108) );
  XOR U7074 ( .A(n7109), .B(n7079), .Z(n7082) );
  XOR U7075 ( .A(p_input[1037]), .B(p_input[573]), .Z(n7079) );
  XNOR U7076 ( .A(p_input[1038]), .B(p_input[574]), .Z(n7109) );
  XOR U7077 ( .A(p_input[1033]), .B(p_input[569]), .Z(n7074) );
  XNOR U7078 ( .A(n7090), .B(n7089), .Z(n7072) );
  XNOR U7079 ( .A(n7110), .B(n7095), .Z(n7089) );
  XOR U7080 ( .A(p_input[1032]), .B(p_input[568]), .Z(n7095) );
  XOR U7081 ( .A(n7086), .B(n7094), .Z(n7110) );
  XOR U7082 ( .A(n7111), .B(n7091), .Z(n7094) );
  XOR U7083 ( .A(p_input[1030]), .B(p_input[566]), .Z(n7091) );
  XNOR U7084 ( .A(p_input[1031]), .B(p_input[567]), .Z(n7111) );
  XOR U7085 ( .A(p_input[1026]), .B(p_input[562]), .Z(n7086) );
  XNOR U7086 ( .A(n7100), .B(n7099), .Z(n7090) );
  XOR U7087 ( .A(n7112), .B(n7096), .Z(n7099) );
  XOR U7088 ( .A(p_input[1027]), .B(p_input[563]), .Z(n7096) );
  XNOR U7089 ( .A(p_input[1028]), .B(p_input[564]), .Z(n7112) );
  XOR U7090 ( .A(p_input[1029]), .B(p_input[565]), .Z(n7100) );
  XOR U7091 ( .A(n7113), .B(n7114), .Z(n7001) );
  AND U7092 ( .A(n147), .B(n7115), .Z(n7114) );
  XNOR U7093 ( .A(n7116), .B(n7113), .Z(n7115) );
  XNOR U7094 ( .A(n7117), .B(n7118), .Z(n147) );
  AND U7095 ( .A(n7119), .B(n7120), .Z(n7118) );
  XOR U7096 ( .A(n7014), .B(n7117), .Z(n7120) );
  AND U7097 ( .A(n7121), .B(n7122), .Z(n7014) );
  XNOR U7098 ( .A(n7011), .B(n7117), .Z(n7119) );
  XOR U7099 ( .A(n7123), .B(n7124), .Z(n7011) );
  AND U7100 ( .A(n151), .B(n7125), .Z(n7124) );
  XOR U7101 ( .A(n7126), .B(n7123), .Z(n7125) );
  XOR U7102 ( .A(n7127), .B(n7128), .Z(n7117) );
  AND U7103 ( .A(n7129), .B(n7130), .Z(n7128) );
  XNOR U7104 ( .A(n7127), .B(n7121), .Z(n7130) );
  IV U7105 ( .A(n7029), .Z(n7121) );
  XOR U7106 ( .A(n7131), .B(n7132), .Z(n7029) );
  XOR U7107 ( .A(n7133), .B(n7122), .Z(n7132) );
  AND U7108 ( .A(n7056), .B(n7134), .Z(n7122) );
  AND U7109 ( .A(n7135), .B(n7136), .Z(n7133) );
  XOR U7110 ( .A(n7137), .B(n7131), .Z(n7135) );
  XNOR U7111 ( .A(n7026), .B(n7127), .Z(n7129) );
  XOR U7112 ( .A(n7138), .B(n7139), .Z(n7026) );
  AND U7113 ( .A(n151), .B(n7140), .Z(n7139) );
  XOR U7114 ( .A(n7141), .B(n7138), .Z(n7140) );
  XOR U7115 ( .A(n7142), .B(n7143), .Z(n7127) );
  AND U7116 ( .A(n7144), .B(n7145), .Z(n7143) );
  XNOR U7117 ( .A(n7142), .B(n7056), .Z(n7145) );
  XOR U7118 ( .A(n7146), .B(n7136), .Z(n7056) );
  XNOR U7119 ( .A(n7147), .B(n7131), .Z(n7136) );
  XOR U7120 ( .A(n7148), .B(n7149), .Z(n7131) );
  AND U7121 ( .A(n7150), .B(n7151), .Z(n7149) );
  XOR U7122 ( .A(n7152), .B(n7148), .Z(n7150) );
  XNOR U7123 ( .A(n7153), .B(n7154), .Z(n7147) );
  AND U7124 ( .A(n7155), .B(n7156), .Z(n7154) );
  XOR U7125 ( .A(n7153), .B(n7157), .Z(n7155) );
  XNOR U7126 ( .A(n7137), .B(n7134), .Z(n7146) );
  AND U7127 ( .A(n7158), .B(n7159), .Z(n7134) );
  XOR U7128 ( .A(n7160), .B(n7161), .Z(n7137) );
  AND U7129 ( .A(n7162), .B(n7163), .Z(n7161) );
  XOR U7130 ( .A(n7160), .B(n7164), .Z(n7162) );
  XNOR U7131 ( .A(n7053), .B(n7142), .Z(n7144) );
  XOR U7132 ( .A(n7165), .B(n7166), .Z(n7053) );
  AND U7133 ( .A(n151), .B(n7167), .Z(n7166) );
  XNOR U7134 ( .A(n7168), .B(n7165), .Z(n7167) );
  XOR U7135 ( .A(n7169), .B(n7170), .Z(n7142) );
  AND U7136 ( .A(n7171), .B(n7172), .Z(n7170) );
  XNOR U7137 ( .A(n7169), .B(n7158), .Z(n7172) );
  IV U7138 ( .A(n7104), .Z(n7158) );
  XNOR U7139 ( .A(n7173), .B(n7151), .Z(n7104) );
  XNOR U7140 ( .A(n7174), .B(n7157), .Z(n7151) );
  XOR U7141 ( .A(n7175), .B(n7176), .Z(n7157) );
  NOR U7142 ( .A(n7177), .B(n7178), .Z(n7176) );
  XNOR U7143 ( .A(n7175), .B(n7179), .Z(n7177) );
  XNOR U7144 ( .A(n7156), .B(n7148), .Z(n7174) );
  XOR U7145 ( .A(n7180), .B(n7181), .Z(n7148) );
  AND U7146 ( .A(n7182), .B(n7183), .Z(n7181) );
  XNOR U7147 ( .A(n7180), .B(n7184), .Z(n7182) );
  XNOR U7148 ( .A(n7185), .B(n7153), .Z(n7156) );
  XOR U7149 ( .A(n7186), .B(n7187), .Z(n7153) );
  AND U7150 ( .A(n7188), .B(n7189), .Z(n7187) );
  XOR U7151 ( .A(n7186), .B(n7190), .Z(n7188) );
  XNOR U7152 ( .A(n7191), .B(n7192), .Z(n7185) );
  NOR U7153 ( .A(n7193), .B(n7194), .Z(n7192) );
  XOR U7154 ( .A(n7191), .B(n7195), .Z(n7193) );
  XNOR U7155 ( .A(n7152), .B(n7159), .Z(n7173) );
  NOR U7156 ( .A(n7116), .B(n7196), .Z(n7159) );
  XOR U7157 ( .A(n7164), .B(n7163), .Z(n7152) );
  XNOR U7158 ( .A(n7197), .B(n7160), .Z(n7163) );
  XOR U7159 ( .A(n7198), .B(n7199), .Z(n7160) );
  AND U7160 ( .A(n7200), .B(n7201), .Z(n7199) );
  XOR U7161 ( .A(n7198), .B(n7202), .Z(n7200) );
  XNOR U7162 ( .A(n7203), .B(n7204), .Z(n7197) );
  NOR U7163 ( .A(n7205), .B(n7206), .Z(n7204) );
  XNOR U7164 ( .A(n7203), .B(n7207), .Z(n7205) );
  XOR U7165 ( .A(n7208), .B(n7209), .Z(n7164) );
  NOR U7166 ( .A(n7210), .B(n7211), .Z(n7209) );
  XNOR U7167 ( .A(n7208), .B(n7212), .Z(n7210) );
  XNOR U7168 ( .A(n7101), .B(n7169), .Z(n7171) );
  XOR U7169 ( .A(n7213), .B(n7214), .Z(n7101) );
  AND U7170 ( .A(n151), .B(n7215), .Z(n7214) );
  XOR U7171 ( .A(n7216), .B(n7213), .Z(n7215) );
  AND U7172 ( .A(n7113), .B(n7116), .Z(n7169) );
  XOR U7173 ( .A(n7217), .B(n7196), .Z(n7116) );
  XNOR U7174 ( .A(p_input[1024]), .B(p_input[576]), .Z(n7196) );
  XOR U7175 ( .A(n7184), .B(n7183), .Z(n7217) );
  XNOR U7176 ( .A(n7218), .B(n7190), .Z(n7183) );
  XNOR U7177 ( .A(n7179), .B(n7178), .Z(n7190) );
  XOR U7178 ( .A(n7219), .B(n7175), .Z(n7178) );
  XOR U7179 ( .A(p_input[1034]), .B(p_input[586]), .Z(n7175) );
  XNOR U7180 ( .A(p_input[1035]), .B(p_input[587]), .Z(n7219) );
  XOR U7181 ( .A(p_input[1036]), .B(p_input[588]), .Z(n7179) );
  XNOR U7182 ( .A(n7189), .B(n7180), .Z(n7218) );
  XNOR U7183 ( .A(n3298), .B(p_input[577]), .Z(n7180) );
  XOR U7184 ( .A(n7220), .B(n7195), .Z(n7189) );
  XNOR U7185 ( .A(p_input[1039]), .B(p_input[591]), .Z(n7195) );
  XOR U7186 ( .A(n7186), .B(n7194), .Z(n7220) );
  XOR U7187 ( .A(n7221), .B(n7191), .Z(n7194) );
  XOR U7188 ( .A(p_input[1037]), .B(p_input[589]), .Z(n7191) );
  XNOR U7189 ( .A(p_input[1038]), .B(p_input[590]), .Z(n7221) );
  XOR U7190 ( .A(p_input[1033]), .B(p_input[585]), .Z(n7186) );
  XNOR U7191 ( .A(n7202), .B(n7201), .Z(n7184) );
  XNOR U7192 ( .A(n7222), .B(n7207), .Z(n7201) );
  XOR U7193 ( .A(p_input[1032]), .B(p_input[584]), .Z(n7207) );
  XOR U7194 ( .A(n7198), .B(n7206), .Z(n7222) );
  XOR U7195 ( .A(n7223), .B(n7203), .Z(n7206) );
  XOR U7196 ( .A(p_input[1030]), .B(p_input[582]), .Z(n7203) );
  XNOR U7197 ( .A(p_input[1031]), .B(p_input[583]), .Z(n7223) );
  XOR U7198 ( .A(p_input[1026]), .B(p_input[578]), .Z(n7198) );
  XNOR U7199 ( .A(n7212), .B(n7211), .Z(n7202) );
  XOR U7200 ( .A(n7224), .B(n7208), .Z(n7211) );
  XOR U7201 ( .A(p_input[1027]), .B(p_input[579]), .Z(n7208) );
  XNOR U7202 ( .A(p_input[1028]), .B(p_input[580]), .Z(n7224) );
  XOR U7203 ( .A(p_input[1029]), .B(p_input[581]), .Z(n7212) );
  XOR U7204 ( .A(n7225), .B(n7226), .Z(n7113) );
  AND U7205 ( .A(n151), .B(n7227), .Z(n7226) );
  XNOR U7206 ( .A(n7228), .B(n7225), .Z(n7227) );
  XNOR U7207 ( .A(n7229), .B(n7230), .Z(n151) );
  AND U7208 ( .A(n7231), .B(n7232), .Z(n7230) );
  XOR U7209 ( .A(n7126), .B(n7229), .Z(n7232) );
  AND U7210 ( .A(n7233), .B(n7234), .Z(n7126) );
  XNOR U7211 ( .A(n7123), .B(n7229), .Z(n7231) );
  XOR U7212 ( .A(n7235), .B(n7236), .Z(n7123) );
  AND U7213 ( .A(n155), .B(n7237), .Z(n7236) );
  XOR U7214 ( .A(n7238), .B(n7235), .Z(n7237) );
  XOR U7215 ( .A(n7239), .B(n7240), .Z(n7229) );
  AND U7216 ( .A(n7241), .B(n7242), .Z(n7240) );
  XNOR U7217 ( .A(n7239), .B(n7233), .Z(n7242) );
  IV U7218 ( .A(n7141), .Z(n7233) );
  XOR U7219 ( .A(n7243), .B(n7244), .Z(n7141) );
  XOR U7220 ( .A(n7245), .B(n7234), .Z(n7244) );
  AND U7221 ( .A(n7168), .B(n7246), .Z(n7234) );
  AND U7222 ( .A(n7247), .B(n7248), .Z(n7245) );
  XOR U7223 ( .A(n7249), .B(n7243), .Z(n7247) );
  XNOR U7224 ( .A(n7138), .B(n7239), .Z(n7241) );
  XOR U7225 ( .A(n7250), .B(n7251), .Z(n7138) );
  AND U7226 ( .A(n155), .B(n7252), .Z(n7251) );
  XOR U7227 ( .A(n7253), .B(n7250), .Z(n7252) );
  XOR U7228 ( .A(n7254), .B(n7255), .Z(n7239) );
  AND U7229 ( .A(n7256), .B(n7257), .Z(n7255) );
  XNOR U7230 ( .A(n7254), .B(n7168), .Z(n7257) );
  XOR U7231 ( .A(n7258), .B(n7248), .Z(n7168) );
  XNOR U7232 ( .A(n7259), .B(n7243), .Z(n7248) );
  XOR U7233 ( .A(n7260), .B(n7261), .Z(n7243) );
  AND U7234 ( .A(n7262), .B(n7263), .Z(n7261) );
  XOR U7235 ( .A(n7264), .B(n7260), .Z(n7262) );
  XNOR U7236 ( .A(n7265), .B(n7266), .Z(n7259) );
  AND U7237 ( .A(n7267), .B(n7268), .Z(n7266) );
  XOR U7238 ( .A(n7265), .B(n7269), .Z(n7267) );
  XNOR U7239 ( .A(n7249), .B(n7246), .Z(n7258) );
  AND U7240 ( .A(n7270), .B(n7271), .Z(n7246) );
  XOR U7241 ( .A(n7272), .B(n7273), .Z(n7249) );
  AND U7242 ( .A(n7274), .B(n7275), .Z(n7273) );
  XOR U7243 ( .A(n7272), .B(n7276), .Z(n7274) );
  XNOR U7244 ( .A(n7165), .B(n7254), .Z(n7256) );
  XOR U7245 ( .A(n7277), .B(n7278), .Z(n7165) );
  AND U7246 ( .A(n155), .B(n7279), .Z(n7278) );
  XNOR U7247 ( .A(n7280), .B(n7277), .Z(n7279) );
  XOR U7248 ( .A(n7281), .B(n7282), .Z(n7254) );
  AND U7249 ( .A(n7283), .B(n7284), .Z(n7282) );
  XNOR U7250 ( .A(n7281), .B(n7270), .Z(n7284) );
  IV U7251 ( .A(n7216), .Z(n7270) );
  XNOR U7252 ( .A(n7285), .B(n7263), .Z(n7216) );
  XNOR U7253 ( .A(n7286), .B(n7269), .Z(n7263) );
  XOR U7254 ( .A(n7287), .B(n7288), .Z(n7269) );
  NOR U7255 ( .A(n7289), .B(n7290), .Z(n7288) );
  XNOR U7256 ( .A(n7287), .B(n7291), .Z(n7289) );
  XNOR U7257 ( .A(n7268), .B(n7260), .Z(n7286) );
  XOR U7258 ( .A(n7292), .B(n7293), .Z(n7260) );
  AND U7259 ( .A(n7294), .B(n7295), .Z(n7293) );
  XNOR U7260 ( .A(n7292), .B(n7296), .Z(n7294) );
  XNOR U7261 ( .A(n7297), .B(n7265), .Z(n7268) );
  XOR U7262 ( .A(n7298), .B(n7299), .Z(n7265) );
  AND U7263 ( .A(n7300), .B(n7301), .Z(n7299) );
  XOR U7264 ( .A(n7298), .B(n7302), .Z(n7300) );
  XNOR U7265 ( .A(n7303), .B(n7304), .Z(n7297) );
  NOR U7266 ( .A(n7305), .B(n7306), .Z(n7304) );
  XOR U7267 ( .A(n7303), .B(n7307), .Z(n7305) );
  XNOR U7268 ( .A(n7264), .B(n7271), .Z(n7285) );
  NOR U7269 ( .A(n7228), .B(n7308), .Z(n7271) );
  XOR U7270 ( .A(n7276), .B(n7275), .Z(n7264) );
  XNOR U7271 ( .A(n7309), .B(n7272), .Z(n7275) );
  XOR U7272 ( .A(n7310), .B(n7311), .Z(n7272) );
  AND U7273 ( .A(n7312), .B(n7313), .Z(n7311) );
  XOR U7274 ( .A(n7310), .B(n7314), .Z(n7312) );
  XNOR U7275 ( .A(n7315), .B(n7316), .Z(n7309) );
  NOR U7276 ( .A(n7317), .B(n7318), .Z(n7316) );
  XNOR U7277 ( .A(n7315), .B(n7319), .Z(n7317) );
  XOR U7278 ( .A(n7320), .B(n7321), .Z(n7276) );
  NOR U7279 ( .A(n7322), .B(n7323), .Z(n7321) );
  XNOR U7280 ( .A(n7320), .B(n7324), .Z(n7322) );
  XNOR U7281 ( .A(n7213), .B(n7281), .Z(n7283) );
  XOR U7282 ( .A(n7325), .B(n7326), .Z(n7213) );
  AND U7283 ( .A(n155), .B(n7327), .Z(n7326) );
  XOR U7284 ( .A(n7328), .B(n7325), .Z(n7327) );
  AND U7285 ( .A(n7225), .B(n7228), .Z(n7281) );
  XOR U7286 ( .A(n7329), .B(n7308), .Z(n7228) );
  XNOR U7287 ( .A(p_input[1024]), .B(p_input[592]), .Z(n7308) );
  XOR U7288 ( .A(n7296), .B(n7295), .Z(n7329) );
  XNOR U7289 ( .A(n7330), .B(n7302), .Z(n7295) );
  XNOR U7290 ( .A(n7291), .B(n7290), .Z(n7302) );
  XOR U7291 ( .A(n7331), .B(n7287), .Z(n7290) );
  XOR U7292 ( .A(p_input[1034]), .B(p_input[602]), .Z(n7287) );
  XNOR U7293 ( .A(p_input[1035]), .B(p_input[603]), .Z(n7331) );
  XOR U7294 ( .A(p_input[1036]), .B(p_input[604]), .Z(n7291) );
  XNOR U7295 ( .A(n7301), .B(n7292), .Z(n7330) );
  XNOR U7296 ( .A(n3298), .B(p_input[593]), .Z(n7292) );
  XOR U7297 ( .A(n7332), .B(n7307), .Z(n7301) );
  XNOR U7298 ( .A(p_input[1039]), .B(p_input[607]), .Z(n7307) );
  XOR U7299 ( .A(n7298), .B(n7306), .Z(n7332) );
  XOR U7300 ( .A(n7333), .B(n7303), .Z(n7306) );
  XOR U7301 ( .A(p_input[1037]), .B(p_input[605]), .Z(n7303) );
  XNOR U7302 ( .A(p_input[1038]), .B(p_input[606]), .Z(n7333) );
  XOR U7303 ( .A(p_input[1033]), .B(p_input[601]), .Z(n7298) );
  XNOR U7304 ( .A(n7314), .B(n7313), .Z(n7296) );
  XNOR U7305 ( .A(n7334), .B(n7319), .Z(n7313) );
  XOR U7306 ( .A(p_input[1032]), .B(p_input[600]), .Z(n7319) );
  XOR U7307 ( .A(n7310), .B(n7318), .Z(n7334) );
  XOR U7308 ( .A(n7335), .B(n7315), .Z(n7318) );
  XOR U7309 ( .A(p_input[1030]), .B(p_input[598]), .Z(n7315) );
  XNOR U7310 ( .A(p_input[1031]), .B(p_input[599]), .Z(n7335) );
  XOR U7311 ( .A(p_input[1026]), .B(p_input[594]), .Z(n7310) );
  XNOR U7312 ( .A(n7324), .B(n7323), .Z(n7314) );
  XOR U7313 ( .A(n7336), .B(n7320), .Z(n7323) );
  XOR U7314 ( .A(p_input[1027]), .B(p_input[595]), .Z(n7320) );
  XNOR U7315 ( .A(p_input[1028]), .B(p_input[596]), .Z(n7336) );
  XOR U7316 ( .A(p_input[1029]), .B(p_input[597]), .Z(n7324) );
  XOR U7317 ( .A(n7337), .B(n7338), .Z(n7225) );
  AND U7318 ( .A(n155), .B(n7339), .Z(n7338) );
  XNOR U7319 ( .A(n7340), .B(n7337), .Z(n7339) );
  XNOR U7320 ( .A(n7341), .B(n7342), .Z(n155) );
  AND U7321 ( .A(n7343), .B(n7344), .Z(n7342) );
  XOR U7322 ( .A(n7238), .B(n7341), .Z(n7344) );
  AND U7323 ( .A(n7345), .B(n7346), .Z(n7238) );
  XNOR U7324 ( .A(n7235), .B(n7341), .Z(n7343) );
  XOR U7325 ( .A(n7347), .B(n7348), .Z(n7235) );
  AND U7326 ( .A(n159), .B(n7349), .Z(n7348) );
  XOR U7327 ( .A(n7350), .B(n7347), .Z(n7349) );
  XOR U7328 ( .A(n7351), .B(n7352), .Z(n7341) );
  AND U7329 ( .A(n7353), .B(n7354), .Z(n7352) );
  XNOR U7330 ( .A(n7351), .B(n7345), .Z(n7354) );
  IV U7331 ( .A(n7253), .Z(n7345) );
  XOR U7332 ( .A(n7355), .B(n7356), .Z(n7253) );
  XOR U7333 ( .A(n7357), .B(n7346), .Z(n7356) );
  AND U7334 ( .A(n7280), .B(n7358), .Z(n7346) );
  AND U7335 ( .A(n7359), .B(n7360), .Z(n7357) );
  XOR U7336 ( .A(n7361), .B(n7355), .Z(n7359) );
  XNOR U7337 ( .A(n7250), .B(n7351), .Z(n7353) );
  XOR U7338 ( .A(n7362), .B(n7363), .Z(n7250) );
  AND U7339 ( .A(n159), .B(n7364), .Z(n7363) );
  XOR U7340 ( .A(n7365), .B(n7362), .Z(n7364) );
  XOR U7341 ( .A(n7366), .B(n7367), .Z(n7351) );
  AND U7342 ( .A(n7368), .B(n7369), .Z(n7367) );
  XNOR U7343 ( .A(n7366), .B(n7280), .Z(n7369) );
  XOR U7344 ( .A(n7370), .B(n7360), .Z(n7280) );
  XNOR U7345 ( .A(n7371), .B(n7355), .Z(n7360) );
  XOR U7346 ( .A(n7372), .B(n7373), .Z(n7355) );
  AND U7347 ( .A(n7374), .B(n7375), .Z(n7373) );
  XOR U7348 ( .A(n7376), .B(n7372), .Z(n7374) );
  XNOR U7349 ( .A(n7377), .B(n7378), .Z(n7371) );
  AND U7350 ( .A(n7379), .B(n7380), .Z(n7378) );
  XOR U7351 ( .A(n7377), .B(n7381), .Z(n7379) );
  XNOR U7352 ( .A(n7361), .B(n7358), .Z(n7370) );
  AND U7353 ( .A(n7382), .B(n7383), .Z(n7358) );
  XOR U7354 ( .A(n7384), .B(n7385), .Z(n7361) );
  AND U7355 ( .A(n7386), .B(n7387), .Z(n7385) );
  XOR U7356 ( .A(n7384), .B(n7388), .Z(n7386) );
  XNOR U7357 ( .A(n7277), .B(n7366), .Z(n7368) );
  XOR U7358 ( .A(n7389), .B(n7390), .Z(n7277) );
  AND U7359 ( .A(n159), .B(n7391), .Z(n7390) );
  XNOR U7360 ( .A(n7392), .B(n7389), .Z(n7391) );
  XOR U7361 ( .A(n7393), .B(n7394), .Z(n7366) );
  AND U7362 ( .A(n7395), .B(n7396), .Z(n7394) );
  XNOR U7363 ( .A(n7393), .B(n7382), .Z(n7396) );
  IV U7364 ( .A(n7328), .Z(n7382) );
  XNOR U7365 ( .A(n7397), .B(n7375), .Z(n7328) );
  XNOR U7366 ( .A(n7398), .B(n7381), .Z(n7375) );
  XOR U7367 ( .A(n7399), .B(n7400), .Z(n7381) );
  NOR U7368 ( .A(n7401), .B(n7402), .Z(n7400) );
  XNOR U7369 ( .A(n7399), .B(n7403), .Z(n7401) );
  XNOR U7370 ( .A(n7380), .B(n7372), .Z(n7398) );
  XOR U7371 ( .A(n7404), .B(n7405), .Z(n7372) );
  AND U7372 ( .A(n7406), .B(n7407), .Z(n7405) );
  XNOR U7373 ( .A(n7404), .B(n7408), .Z(n7406) );
  XNOR U7374 ( .A(n7409), .B(n7377), .Z(n7380) );
  XOR U7375 ( .A(n7410), .B(n7411), .Z(n7377) );
  AND U7376 ( .A(n7412), .B(n7413), .Z(n7411) );
  XOR U7377 ( .A(n7410), .B(n7414), .Z(n7412) );
  XNOR U7378 ( .A(n7415), .B(n7416), .Z(n7409) );
  NOR U7379 ( .A(n7417), .B(n7418), .Z(n7416) );
  XOR U7380 ( .A(n7415), .B(n7419), .Z(n7417) );
  XNOR U7381 ( .A(n7376), .B(n7383), .Z(n7397) );
  NOR U7382 ( .A(n7340), .B(n7420), .Z(n7383) );
  XOR U7383 ( .A(n7388), .B(n7387), .Z(n7376) );
  XNOR U7384 ( .A(n7421), .B(n7384), .Z(n7387) );
  XOR U7385 ( .A(n7422), .B(n7423), .Z(n7384) );
  AND U7386 ( .A(n7424), .B(n7425), .Z(n7423) );
  XOR U7387 ( .A(n7422), .B(n7426), .Z(n7424) );
  XNOR U7388 ( .A(n7427), .B(n7428), .Z(n7421) );
  NOR U7389 ( .A(n7429), .B(n7430), .Z(n7428) );
  XNOR U7390 ( .A(n7427), .B(n7431), .Z(n7429) );
  XOR U7391 ( .A(n7432), .B(n7433), .Z(n7388) );
  NOR U7392 ( .A(n7434), .B(n7435), .Z(n7433) );
  XNOR U7393 ( .A(n7432), .B(n7436), .Z(n7434) );
  XNOR U7394 ( .A(n7325), .B(n7393), .Z(n7395) );
  XOR U7395 ( .A(n7437), .B(n7438), .Z(n7325) );
  AND U7396 ( .A(n159), .B(n7439), .Z(n7438) );
  XOR U7397 ( .A(n7440), .B(n7437), .Z(n7439) );
  AND U7398 ( .A(n7337), .B(n7340), .Z(n7393) );
  XOR U7399 ( .A(n7441), .B(n7420), .Z(n7340) );
  XNOR U7400 ( .A(p_input[1024]), .B(p_input[608]), .Z(n7420) );
  XOR U7401 ( .A(n7408), .B(n7407), .Z(n7441) );
  XNOR U7402 ( .A(n7442), .B(n7414), .Z(n7407) );
  XNOR U7403 ( .A(n7403), .B(n7402), .Z(n7414) );
  XOR U7404 ( .A(n7443), .B(n7399), .Z(n7402) );
  XOR U7405 ( .A(p_input[1034]), .B(p_input[618]), .Z(n7399) );
  XNOR U7406 ( .A(p_input[1035]), .B(p_input[619]), .Z(n7443) );
  XOR U7407 ( .A(p_input[1036]), .B(p_input[620]), .Z(n7403) );
  XNOR U7408 ( .A(n7413), .B(n7404), .Z(n7442) );
  XNOR U7409 ( .A(n3298), .B(p_input[609]), .Z(n7404) );
  XOR U7410 ( .A(n7444), .B(n7419), .Z(n7413) );
  XNOR U7411 ( .A(p_input[1039]), .B(p_input[623]), .Z(n7419) );
  XOR U7412 ( .A(n7410), .B(n7418), .Z(n7444) );
  XOR U7413 ( .A(n7445), .B(n7415), .Z(n7418) );
  XOR U7414 ( .A(p_input[1037]), .B(p_input[621]), .Z(n7415) );
  XNOR U7415 ( .A(p_input[1038]), .B(p_input[622]), .Z(n7445) );
  XOR U7416 ( .A(p_input[1033]), .B(p_input[617]), .Z(n7410) );
  XNOR U7417 ( .A(n7426), .B(n7425), .Z(n7408) );
  XNOR U7418 ( .A(n7446), .B(n7431), .Z(n7425) );
  XOR U7419 ( .A(p_input[1032]), .B(p_input[616]), .Z(n7431) );
  XOR U7420 ( .A(n7422), .B(n7430), .Z(n7446) );
  XOR U7421 ( .A(n7447), .B(n7427), .Z(n7430) );
  XOR U7422 ( .A(p_input[1030]), .B(p_input[614]), .Z(n7427) );
  XNOR U7423 ( .A(p_input[1031]), .B(p_input[615]), .Z(n7447) );
  XOR U7424 ( .A(p_input[1026]), .B(p_input[610]), .Z(n7422) );
  XNOR U7425 ( .A(n7436), .B(n7435), .Z(n7426) );
  XOR U7426 ( .A(n7448), .B(n7432), .Z(n7435) );
  XOR U7427 ( .A(p_input[1027]), .B(p_input[611]), .Z(n7432) );
  XNOR U7428 ( .A(p_input[1028]), .B(p_input[612]), .Z(n7448) );
  XOR U7429 ( .A(p_input[1029]), .B(p_input[613]), .Z(n7436) );
  XOR U7430 ( .A(n7449), .B(n7450), .Z(n7337) );
  AND U7431 ( .A(n159), .B(n7451), .Z(n7450) );
  XNOR U7432 ( .A(n7452), .B(n7449), .Z(n7451) );
  XNOR U7433 ( .A(n7453), .B(n7454), .Z(n159) );
  AND U7434 ( .A(n7455), .B(n7456), .Z(n7454) );
  XOR U7435 ( .A(n7350), .B(n7453), .Z(n7456) );
  AND U7436 ( .A(n7457), .B(n7458), .Z(n7350) );
  XNOR U7437 ( .A(n7347), .B(n7453), .Z(n7455) );
  XOR U7438 ( .A(n7459), .B(n7460), .Z(n7347) );
  AND U7439 ( .A(n163), .B(n7461), .Z(n7460) );
  XOR U7440 ( .A(n7462), .B(n7459), .Z(n7461) );
  XOR U7441 ( .A(n7463), .B(n7464), .Z(n7453) );
  AND U7442 ( .A(n7465), .B(n7466), .Z(n7464) );
  XNOR U7443 ( .A(n7463), .B(n7457), .Z(n7466) );
  IV U7444 ( .A(n7365), .Z(n7457) );
  XOR U7445 ( .A(n7467), .B(n7468), .Z(n7365) );
  XOR U7446 ( .A(n7469), .B(n7458), .Z(n7468) );
  AND U7447 ( .A(n7392), .B(n7470), .Z(n7458) );
  AND U7448 ( .A(n7471), .B(n7472), .Z(n7469) );
  XOR U7449 ( .A(n7473), .B(n7467), .Z(n7471) );
  XNOR U7450 ( .A(n7362), .B(n7463), .Z(n7465) );
  XOR U7451 ( .A(n7474), .B(n7475), .Z(n7362) );
  AND U7452 ( .A(n163), .B(n7476), .Z(n7475) );
  XOR U7453 ( .A(n7477), .B(n7474), .Z(n7476) );
  XOR U7454 ( .A(n7478), .B(n7479), .Z(n7463) );
  AND U7455 ( .A(n7480), .B(n7481), .Z(n7479) );
  XNOR U7456 ( .A(n7478), .B(n7392), .Z(n7481) );
  XOR U7457 ( .A(n7482), .B(n7472), .Z(n7392) );
  XNOR U7458 ( .A(n7483), .B(n7467), .Z(n7472) );
  XOR U7459 ( .A(n7484), .B(n7485), .Z(n7467) );
  AND U7460 ( .A(n7486), .B(n7487), .Z(n7485) );
  XOR U7461 ( .A(n7488), .B(n7484), .Z(n7486) );
  XNOR U7462 ( .A(n7489), .B(n7490), .Z(n7483) );
  AND U7463 ( .A(n7491), .B(n7492), .Z(n7490) );
  XOR U7464 ( .A(n7489), .B(n7493), .Z(n7491) );
  XNOR U7465 ( .A(n7473), .B(n7470), .Z(n7482) );
  AND U7466 ( .A(n7494), .B(n7495), .Z(n7470) );
  XOR U7467 ( .A(n7496), .B(n7497), .Z(n7473) );
  AND U7468 ( .A(n7498), .B(n7499), .Z(n7497) );
  XOR U7469 ( .A(n7496), .B(n7500), .Z(n7498) );
  XNOR U7470 ( .A(n7389), .B(n7478), .Z(n7480) );
  XOR U7471 ( .A(n7501), .B(n7502), .Z(n7389) );
  AND U7472 ( .A(n163), .B(n7503), .Z(n7502) );
  XNOR U7473 ( .A(n7504), .B(n7501), .Z(n7503) );
  XOR U7474 ( .A(n7505), .B(n7506), .Z(n7478) );
  AND U7475 ( .A(n7507), .B(n7508), .Z(n7506) );
  XNOR U7476 ( .A(n7505), .B(n7494), .Z(n7508) );
  IV U7477 ( .A(n7440), .Z(n7494) );
  XNOR U7478 ( .A(n7509), .B(n7487), .Z(n7440) );
  XNOR U7479 ( .A(n7510), .B(n7493), .Z(n7487) );
  XOR U7480 ( .A(n7511), .B(n7512), .Z(n7493) );
  NOR U7481 ( .A(n7513), .B(n7514), .Z(n7512) );
  XNOR U7482 ( .A(n7511), .B(n7515), .Z(n7513) );
  XNOR U7483 ( .A(n7492), .B(n7484), .Z(n7510) );
  XOR U7484 ( .A(n7516), .B(n7517), .Z(n7484) );
  AND U7485 ( .A(n7518), .B(n7519), .Z(n7517) );
  XNOR U7486 ( .A(n7516), .B(n7520), .Z(n7518) );
  XNOR U7487 ( .A(n7521), .B(n7489), .Z(n7492) );
  XOR U7488 ( .A(n7522), .B(n7523), .Z(n7489) );
  AND U7489 ( .A(n7524), .B(n7525), .Z(n7523) );
  XOR U7490 ( .A(n7522), .B(n7526), .Z(n7524) );
  XNOR U7491 ( .A(n7527), .B(n7528), .Z(n7521) );
  NOR U7492 ( .A(n7529), .B(n7530), .Z(n7528) );
  XOR U7493 ( .A(n7527), .B(n7531), .Z(n7529) );
  XNOR U7494 ( .A(n7488), .B(n7495), .Z(n7509) );
  NOR U7495 ( .A(n7452), .B(n7532), .Z(n7495) );
  XOR U7496 ( .A(n7500), .B(n7499), .Z(n7488) );
  XNOR U7497 ( .A(n7533), .B(n7496), .Z(n7499) );
  XOR U7498 ( .A(n7534), .B(n7535), .Z(n7496) );
  AND U7499 ( .A(n7536), .B(n7537), .Z(n7535) );
  XOR U7500 ( .A(n7534), .B(n7538), .Z(n7536) );
  XNOR U7501 ( .A(n7539), .B(n7540), .Z(n7533) );
  NOR U7502 ( .A(n7541), .B(n7542), .Z(n7540) );
  XNOR U7503 ( .A(n7539), .B(n7543), .Z(n7541) );
  XOR U7504 ( .A(n7544), .B(n7545), .Z(n7500) );
  NOR U7505 ( .A(n7546), .B(n7547), .Z(n7545) );
  XNOR U7506 ( .A(n7544), .B(n7548), .Z(n7546) );
  XNOR U7507 ( .A(n7437), .B(n7505), .Z(n7507) );
  XOR U7508 ( .A(n7549), .B(n7550), .Z(n7437) );
  AND U7509 ( .A(n163), .B(n7551), .Z(n7550) );
  XOR U7510 ( .A(n7552), .B(n7549), .Z(n7551) );
  AND U7511 ( .A(n7449), .B(n7452), .Z(n7505) );
  XOR U7512 ( .A(n7553), .B(n7532), .Z(n7452) );
  XNOR U7513 ( .A(p_input[1024]), .B(p_input[624]), .Z(n7532) );
  XOR U7514 ( .A(n7520), .B(n7519), .Z(n7553) );
  XNOR U7515 ( .A(n7554), .B(n7526), .Z(n7519) );
  XNOR U7516 ( .A(n7515), .B(n7514), .Z(n7526) );
  XOR U7517 ( .A(n7555), .B(n7511), .Z(n7514) );
  XOR U7518 ( .A(p_input[1034]), .B(p_input[634]), .Z(n7511) );
  XNOR U7519 ( .A(p_input[1035]), .B(p_input[635]), .Z(n7555) );
  XOR U7520 ( .A(p_input[1036]), .B(p_input[636]), .Z(n7515) );
  XNOR U7521 ( .A(n7525), .B(n7516), .Z(n7554) );
  XNOR U7522 ( .A(n3298), .B(p_input[625]), .Z(n7516) );
  XOR U7523 ( .A(n7556), .B(n7531), .Z(n7525) );
  XNOR U7524 ( .A(p_input[1039]), .B(p_input[639]), .Z(n7531) );
  XOR U7525 ( .A(n7522), .B(n7530), .Z(n7556) );
  XOR U7526 ( .A(n7557), .B(n7527), .Z(n7530) );
  XOR U7527 ( .A(p_input[1037]), .B(p_input[637]), .Z(n7527) );
  XNOR U7528 ( .A(p_input[1038]), .B(p_input[638]), .Z(n7557) );
  XOR U7529 ( .A(p_input[1033]), .B(p_input[633]), .Z(n7522) );
  XNOR U7530 ( .A(n7538), .B(n7537), .Z(n7520) );
  XNOR U7531 ( .A(n7558), .B(n7543), .Z(n7537) );
  XOR U7532 ( .A(p_input[1032]), .B(p_input[632]), .Z(n7543) );
  XOR U7533 ( .A(n7534), .B(n7542), .Z(n7558) );
  XOR U7534 ( .A(n7559), .B(n7539), .Z(n7542) );
  XOR U7535 ( .A(p_input[1030]), .B(p_input[630]), .Z(n7539) );
  XNOR U7536 ( .A(p_input[1031]), .B(p_input[631]), .Z(n7559) );
  XOR U7537 ( .A(p_input[1026]), .B(p_input[626]), .Z(n7534) );
  XNOR U7538 ( .A(n7548), .B(n7547), .Z(n7538) );
  XOR U7539 ( .A(n7560), .B(n7544), .Z(n7547) );
  XOR U7540 ( .A(p_input[1027]), .B(p_input[627]), .Z(n7544) );
  XNOR U7541 ( .A(p_input[1028]), .B(p_input[628]), .Z(n7560) );
  XOR U7542 ( .A(p_input[1029]), .B(p_input[629]), .Z(n7548) );
  XOR U7543 ( .A(n7561), .B(n7562), .Z(n7449) );
  AND U7544 ( .A(n163), .B(n7563), .Z(n7562) );
  XNOR U7545 ( .A(n7564), .B(n7561), .Z(n7563) );
  XNOR U7546 ( .A(n7565), .B(n7566), .Z(n163) );
  AND U7547 ( .A(n7567), .B(n7568), .Z(n7566) );
  XOR U7548 ( .A(n7462), .B(n7565), .Z(n7568) );
  AND U7549 ( .A(n7569), .B(n7570), .Z(n7462) );
  XNOR U7550 ( .A(n7459), .B(n7565), .Z(n7567) );
  XOR U7551 ( .A(n7571), .B(n7572), .Z(n7459) );
  AND U7552 ( .A(n167), .B(n7573), .Z(n7572) );
  XOR U7553 ( .A(n7574), .B(n7571), .Z(n7573) );
  XOR U7554 ( .A(n7575), .B(n7576), .Z(n7565) );
  AND U7555 ( .A(n7577), .B(n7578), .Z(n7576) );
  XNOR U7556 ( .A(n7575), .B(n7569), .Z(n7578) );
  IV U7557 ( .A(n7477), .Z(n7569) );
  XOR U7558 ( .A(n7579), .B(n7580), .Z(n7477) );
  XOR U7559 ( .A(n7581), .B(n7570), .Z(n7580) );
  AND U7560 ( .A(n7504), .B(n7582), .Z(n7570) );
  AND U7561 ( .A(n7583), .B(n7584), .Z(n7581) );
  XOR U7562 ( .A(n7585), .B(n7579), .Z(n7583) );
  XNOR U7563 ( .A(n7474), .B(n7575), .Z(n7577) );
  XOR U7564 ( .A(n7586), .B(n7587), .Z(n7474) );
  AND U7565 ( .A(n167), .B(n7588), .Z(n7587) );
  XOR U7566 ( .A(n7589), .B(n7586), .Z(n7588) );
  XOR U7567 ( .A(n7590), .B(n7591), .Z(n7575) );
  AND U7568 ( .A(n7592), .B(n7593), .Z(n7591) );
  XNOR U7569 ( .A(n7590), .B(n7504), .Z(n7593) );
  XOR U7570 ( .A(n7594), .B(n7584), .Z(n7504) );
  XNOR U7571 ( .A(n7595), .B(n7579), .Z(n7584) );
  XOR U7572 ( .A(n7596), .B(n7597), .Z(n7579) );
  AND U7573 ( .A(n7598), .B(n7599), .Z(n7597) );
  XOR U7574 ( .A(n7600), .B(n7596), .Z(n7598) );
  XNOR U7575 ( .A(n7601), .B(n7602), .Z(n7595) );
  AND U7576 ( .A(n7603), .B(n7604), .Z(n7602) );
  XOR U7577 ( .A(n7601), .B(n7605), .Z(n7603) );
  XNOR U7578 ( .A(n7585), .B(n7582), .Z(n7594) );
  AND U7579 ( .A(n7606), .B(n7607), .Z(n7582) );
  XOR U7580 ( .A(n7608), .B(n7609), .Z(n7585) );
  AND U7581 ( .A(n7610), .B(n7611), .Z(n7609) );
  XOR U7582 ( .A(n7608), .B(n7612), .Z(n7610) );
  XNOR U7583 ( .A(n7501), .B(n7590), .Z(n7592) );
  XOR U7584 ( .A(n7613), .B(n7614), .Z(n7501) );
  AND U7585 ( .A(n167), .B(n7615), .Z(n7614) );
  XNOR U7586 ( .A(n7616), .B(n7613), .Z(n7615) );
  XOR U7587 ( .A(n7617), .B(n7618), .Z(n7590) );
  AND U7588 ( .A(n7619), .B(n7620), .Z(n7618) );
  XNOR U7589 ( .A(n7617), .B(n7606), .Z(n7620) );
  IV U7590 ( .A(n7552), .Z(n7606) );
  XNOR U7591 ( .A(n7621), .B(n7599), .Z(n7552) );
  XNOR U7592 ( .A(n7622), .B(n7605), .Z(n7599) );
  XOR U7593 ( .A(n7623), .B(n7624), .Z(n7605) );
  NOR U7594 ( .A(n7625), .B(n7626), .Z(n7624) );
  XNOR U7595 ( .A(n7623), .B(n7627), .Z(n7625) );
  XNOR U7596 ( .A(n7604), .B(n7596), .Z(n7622) );
  XOR U7597 ( .A(n7628), .B(n7629), .Z(n7596) );
  AND U7598 ( .A(n7630), .B(n7631), .Z(n7629) );
  XNOR U7599 ( .A(n7628), .B(n7632), .Z(n7630) );
  XNOR U7600 ( .A(n7633), .B(n7601), .Z(n7604) );
  XOR U7601 ( .A(n7634), .B(n7635), .Z(n7601) );
  AND U7602 ( .A(n7636), .B(n7637), .Z(n7635) );
  XOR U7603 ( .A(n7634), .B(n7638), .Z(n7636) );
  XNOR U7604 ( .A(n7639), .B(n7640), .Z(n7633) );
  NOR U7605 ( .A(n7641), .B(n7642), .Z(n7640) );
  XOR U7606 ( .A(n7639), .B(n7643), .Z(n7641) );
  XNOR U7607 ( .A(n7600), .B(n7607), .Z(n7621) );
  NOR U7608 ( .A(n7564), .B(n7644), .Z(n7607) );
  XOR U7609 ( .A(n7612), .B(n7611), .Z(n7600) );
  XNOR U7610 ( .A(n7645), .B(n7608), .Z(n7611) );
  XOR U7611 ( .A(n7646), .B(n7647), .Z(n7608) );
  AND U7612 ( .A(n7648), .B(n7649), .Z(n7647) );
  XOR U7613 ( .A(n7646), .B(n7650), .Z(n7648) );
  XNOR U7614 ( .A(n7651), .B(n7652), .Z(n7645) );
  NOR U7615 ( .A(n7653), .B(n7654), .Z(n7652) );
  XNOR U7616 ( .A(n7651), .B(n7655), .Z(n7653) );
  XOR U7617 ( .A(n7656), .B(n7657), .Z(n7612) );
  NOR U7618 ( .A(n7658), .B(n7659), .Z(n7657) );
  XNOR U7619 ( .A(n7656), .B(n7660), .Z(n7658) );
  XNOR U7620 ( .A(n7549), .B(n7617), .Z(n7619) );
  XOR U7621 ( .A(n7661), .B(n7662), .Z(n7549) );
  AND U7622 ( .A(n167), .B(n7663), .Z(n7662) );
  XOR U7623 ( .A(n7664), .B(n7661), .Z(n7663) );
  AND U7624 ( .A(n7561), .B(n7564), .Z(n7617) );
  XOR U7625 ( .A(n7665), .B(n7644), .Z(n7564) );
  XNOR U7626 ( .A(p_input[1024]), .B(p_input[640]), .Z(n7644) );
  XOR U7627 ( .A(n7632), .B(n7631), .Z(n7665) );
  XNOR U7628 ( .A(n7666), .B(n7638), .Z(n7631) );
  XNOR U7629 ( .A(n7627), .B(n7626), .Z(n7638) );
  XOR U7630 ( .A(n7667), .B(n7623), .Z(n7626) );
  XOR U7631 ( .A(p_input[1034]), .B(p_input[650]), .Z(n7623) );
  XNOR U7632 ( .A(p_input[1035]), .B(p_input[651]), .Z(n7667) );
  XOR U7633 ( .A(p_input[1036]), .B(p_input[652]), .Z(n7627) );
  XNOR U7634 ( .A(n7637), .B(n7628), .Z(n7666) );
  XNOR U7635 ( .A(n3298), .B(p_input[641]), .Z(n7628) );
  XOR U7636 ( .A(n7668), .B(n7643), .Z(n7637) );
  XNOR U7637 ( .A(p_input[1039]), .B(p_input[655]), .Z(n7643) );
  XOR U7638 ( .A(n7634), .B(n7642), .Z(n7668) );
  XOR U7639 ( .A(n7669), .B(n7639), .Z(n7642) );
  XOR U7640 ( .A(p_input[1037]), .B(p_input[653]), .Z(n7639) );
  XNOR U7641 ( .A(p_input[1038]), .B(p_input[654]), .Z(n7669) );
  XOR U7642 ( .A(p_input[1033]), .B(p_input[649]), .Z(n7634) );
  XNOR U7643 ( .A(n7650), .B(n7649), .Z(n7632) );
  XNOR U7644 ( .A(n7670), .B(n7655), .Z(n7649) );
  XOR U7645 ( .A(p_input[1032]), .B(p_input[648]), .Z(n7655) );
  XOR U7646 ( .A(n7646), .B(n7654), .Z(n7670) );
  XOR U7647 ( .A(n7671), .B(n7651), .Z(n7654) );
  XOR U7648 ( .A(p_input[1030]), .B(p_input[646]), .Z(n7651) );
  XNOR U7649 ( .A(p_input[1031]), .B(p_input[647]), .Z(n7671) );
  XOR U7650 ( .A(p_input[1026]), .B(p_input[642]), .Z(n7646) );
  XNOR U7651 ( .A(n7660), .B(n7659), .Z(n7650) );
  XOR U7652 ( .A(n7672), .B(n7656), .Z(n7659) );
  XOR U7653 ( .A(p_input[1027]), .B(p_input[643]), .Z(n7656) );
  XNOR U7654 ( .A(p_input[1028]), .B(p_input[644]), .Z(n7672) );
  XOR U7655 ( .A(p_input[1029]), .B(p_input[645]), .Z(n7660) );
  XOR U7656 ( .A(n7673), .B(n7674), .Z(n7561) );
  AND U7657 ( .A(n167), .B(n7675), .Z(n7674) );
  XNOR U7658 ( .A(n7676), .B(n7673), .Z(n7675) );
  XNOR U7659 ( .A(n7677), .B(n7678), .Z(n167) );
  AND U7660 ( .A(n7679), .B(n7680), .Z(n7678) );
  XOR U7661 ( .A(n7574), .B(n7677), .Z(n7680) );
  AND U7662 ( .A(n7681), .B(n7682), .Z(n7574) );
  XNOR U7663 ( .A(n7571), .B(n7677), .Z(n7679) );
  XOR U7664 ( .A(n7683), .B(n7684), .Z(n7571) );
  AND U7665 ( .A(n171), .B(n7685), .Z(n7684) );
  XOR U7666 ( .A(n7686), .B(n7683), .Z(n7685) );
  XOR U7667 ( .A(n7687), .B(n7688), .Z(n7677) );
  AND U7668 ( .A(n7689), .B(n7690), .Z(n7688) );
  XNOR U7669 ( .A(n7687), .B(n7681), .Z(n7690) );
  IV U7670 ( .A(n7589), .Z(n7681) );
  XOR U7671 ( .A(n7691), .B(n7692), .Z(n7589) );
  XOR U7672 ( .A(n7693), .B(n7682), .Z(n7692) );
  AND U7673 ( .A(n7616), .B(n7694), .Z(n7682) );
  AND U7674 ( .A(n7695), .B(n7696), .Z(n7693) );
  XOR U7675 ( .A(n7697), .B(n7691), .Z(n7695) );
  XNOR U7676 ( .A(n7586), .B(n7687), .Z(n7689) );
  XOR U7677 ( .A(n7698), .B(n7699), .Z(n7586) );
  AND U7678 ( .A(n171), .B(n7700), .Z(n7699) );
  XOR U7679 ( .A(n7701), .B(n7698), .Z(n7700) );
  XOR U7680 ( .A(n7702), .B(n7703), .Z(n7687) );
  AND U7681 ( .A(n7704), .B(n7705), .Z(n7703) );
  XNOR U7682 ( .A(n7702), .B(n7616), .Z(n7705) );
  XOR U7683 ( .A(n7706), .B(n7696), .Z(n7616) );
  XNOR U7684 ( .A(n7707), .B(n7691), .Z(n7696) );
  XOR U7685 ( .A(n7708), .B(n7709), .Z(n7691) );
  AND U7686 ( .A(n7710), .B(n7711), .Z(n7709) );
  XOR U7687 ( .A(n7712), .B(n7708), .Z(n7710) );
  XNOR U7688 ( .A(n7713), .B(n7714), .Z(n7707) );
  AND U7689 ( .A(n7715), .B(n7716), .Z(n7714) );
  XOR U7690 ( .A(n7713), .B(n7717), .Z(n7715) );
  XNOR U7691 ( .A(n7697), .B(n7694), .Z(n7706) );
  AND U7692 ( .A(n7718), .B(n7719), .Z(n7694) );
  XOR U7693 ( .A(n7720), .B(n7721), .Z(n7697) );
  AND U7694 ( .A(n7722), .B(n7723), .Z(n7721) );
  XOR U7695 ( .A(n7720), .B(n7724), .Z(n7722) );
  XNOR U7696 ( .A(n7613), .B(n7702), .Z(n7704) );
  XOR U7697 ( .A(n7725), .B(n7726), .Z(n7613) );
  AND U7698 ( .A(n171), .B(n7727), .Z(n7726) );
  XNOR U7699 ( .A(n7728), .B(n7725), .Z(n7727) );
  XOR U7700 ( .A(n7729), .B(n7730), .Z(n7702) );
  AND U7701 ( .A(n7731), .B(n7732), .Z(n7730) );
  XNOR U7702 ( .A(n7729), .B(n7718), .Z(n7732) );
  IV U7703 ( .A(n7664), .Z(n7718) );
  XNOR U7704 ( .A(n7733), .B(n7711), .Z(n7664) );
  XNOR U7705 ( .A(n7734), .B(n7717), .Z(n7711) );
  XOR U7706 ( .A(n7735), .B(n7736), .Z(n7717) );
  NOR U7707 ( .A(n7737), .B(n7738), .Z(n7736) );
  XNOR U7708 ( .A(n7735), .B(n7739), .Z(n7737) );
  XNOR U7709 ( .A(n7716), .B(n7708), .Z(n7734) );
  XOR U7710 ( .A(n7740), .B(n7741), .Z(n7708) );
  AND U7711 ( .A(n7742), .B(n7743), .Z(n7741) );
  XNOR U7712 ( .A(n7740), .B(n7744), .Z(n7742) );
  XNOR U7713 ( .A(n7745), .B(n7713), .Z(n7716) );
  XOR U7714 ( .A(n7746), .B(n7747), .Z(n7713) );
  AND U7715 ( .A(n7748), .B(n7749), .Z(n7747) );
  XOR U7716 ( .A(n7746), .B(n7750), .Z(n7748) );
  XNOR U7717 ( .A(n7751), .B(n7752), .Z(n7745) );
  NOR U7718 ( .A(n7753), .B(n7754), .Z(n7752) );
  XOR U7719 ( .A(n7751), .B(n7755), .Z(n7753) );
  XNOR U7720 ( .A(n7712), .B(n7719), .Z(n7733) );
  NOR U7721 ( .A(n7676), .B(n7756), .Z(n7719) );
  XOR U7722 ( .A(n7724), .B(n7723), .Z(n7712) );
  XNOR U7723 ( .A(n7757), .B(n7720), .Z(n7723) );
  XOR U7724 ( .A(n7758), .B(n7759), .Z(n7720) );
  AND U7725 ( .A(n7760), .B(n7761), .Z(n7759) );
  XOR U7726 ( .A(n7758), .B(n7762), .Z(n7760) );
  XNOR U7727 ( .A(n7763), .B(n7764), .Z(n7757) );
  NOR U7728 ( .A(n7765), .B(n7766), .Z(n7764) );
  XNOR U7729 ( .A(n7763), .B(n7767), .Z(n7765) );
  XOR U7730 ( .A(n7768), .B(n7769), .Z(n7724) );
  NOR U7731 ( .A(n7770), .B(n7771), .Z(n7769) );
  XNOR U7732 ( .A(n7768), .B(n7772), .Z(n7770) );
  XNOR U7733 ( .A(n7661), .B(n7729), .Z(n7731) );
  XOR U7734 ( .A(n7773), .B(n7774), .Z(n7661) );
  AND U7735 ( .A(n171), .B(n7775), .Z(n7774) );
  XOR U7736 ( .A(n7776), .B(n7773), .Z(n7775) );
  AND U7737 ( .A(n7673), .B(n7676), .Z(n7729) );
  XOR U7738 ( .A(n7777), .B(n7756), .Z(n7676) );
  XNOR U7739 ( .A(p_input[1024]), .B(p_input[656]), .Z(n7756) );
  XOR U7740 ( .A(n7744), .B(n7743), .Z(n7777) );
  XNOR U7741 ( .A(n7778), .B(n7750), .Z(n7743) );
  XNOR U7742 ( .A(n7739), .B(n7738), .Z(n7750) );
  XOR U7743 ( .A(n7779), .B(n7735), .Z(n7738) );
  XOR U7744 ( .A(p_input[1034]), .B(p_input[666]), .Z(n7735) );
  XNOR U7745 ( .A(p_input[1035]), .B(p_input[667]), .Z(n7779) );
  XOR U7746 ( .A(p_input[1036]), .B(p_input[668]), .Z(n7739) );
  XNOR U7747 ( .A(n7749), .B(n7740), .Z(n7778) );
  XNOR U7748 ( .A(n3298), .B(p_input[657]), .Z(n7740) );
  XOR U7749 ( .A(n7780), .B(n7755), .Z(n7749) );
  XNOR U7750 ( .A(p_input[1039]), .B(p_input[671]), .Z(n7755) );
  XOR U7751 ( .A(n7746), .B(n7754), .Z(n7780) );
  XOR U7752 ( .A(n7781), .B(n7751), .Z(n7754) );
  XOR U7753 ( .A(p_input[1037]), .B(p_input[669]), .Z(n7751) );
  XNOR U7754 ( .A(p_input[1038]), .B(p_input[670]), .Z(n7781) );
  XOR U7755 ( .A(p_input[1033]), .B(p_input[665]), .Z(n7746) );
  XNOR U7756 ( .A(n7762), .B(n7761), .Z(n7744) );
  XNOR U7757 ( .A(n7782), .B(n7767), .Z(n7761) );
  XOR U7758 ( .A(p_input[1032]), .B(p_input[664]), .Z(n7767) );
  XOR U7759 ( .A(n7758), .B(n7766), .Z(n7782) );
  XOR U7760 ( .A(n7783), .B(n7763), .Z(n7766) );
  XOR U7761 ( .A(p_input[1030]), .B(p_input[662]), .Z(n7763) );
  XNOR U7762 ( .A(p_input[1031]), .B(p_input[663]), .Z(n7783) );
  XOR U7763 ( .A(p_input[1026]), .B(p_input[658]), .Z(n7758) );
  XNOR U7764 ( .A(n7772), .B(n7771), .Z(n7762) );
  XOR U7765 ( .A(n7784), .B(n7768), .Z(n7771) );
  XOR U7766 ( .A(p_input[1027]), .B(p_input[659]), .Z(n7768) );
  XNOR U7767 ( .A(p_input[1028]), .B(p_input[660]), .Z(n7784) );
  XOR U7768 ( .A(p_input[1029]), .B(p_input[661]), .Z(n7772) );
  XOR U7769 ( .A(n7785), .B(n7786), .Z(n7673) );
  AND U7770 ( .A(n171), .B(n7787), .Z(n7786) );
  XNOR U7771 ( .A(n7788), .B(n7785), .Z(n7787) );
  XNOR U7772 ( .A(n7789), .B(n7790), .Z(n171) );
  AND U7773 ( .A(n7791), .B(n7792), .Z(n7790) );
  XOR U7774 ( .A(n7686), .B(n7789), .Z(n7792) );
  AND U7775 ( .A(n7793), .B(n7794), .Z(n7686) );
  XNOR U7776 ( .A(n7683), .B(n7789), .Z(n7791) );
  XOR U7777 ( .A(n7795), .B(n7796), .Z(n7683) );
  AND U7778 ( .A(n175), .B(n7797), .Z(n7796) );
  XOR U7779 ( .A(n7798), .B(n7795), .Z(n7797) );
  XOR U7780 ( .A(n7799), .B(n7800), .Z(n7789) );
  AND U7781 ( .A(n7801), .B(n7802), .Z(n7800) );
  XNOR U7782 ( .A(n7799), .B(n7793), .Z(n7802) );
  IV U7783 ( .A(n7701), .Z(n7793) );
  XOR U7784 ( .A(n7803), .B(n7804), .Z(n7701) );
  XOR U7785 ( .A(n7805), .B(n7794), .Z(n7804) );
  AND U7786 ( .A(n7728), .B(n7806), .Z(n7794) );
  AND U7787 ( .A(n7807), .B(n7808), .Z(n7805) );
  XOR U7788 ( .A(n7809), .B(n7803), .Z(n7807) );
  XNOR U7789 ( .A(n7698), .B(n7799), .Z(n7801) );
  XOR U7790 ( .A(n7810), .B(n7811), .Z(n7698) );
  AND U7791 ( .A(n175), .B(n7812), .Z(n7811) );
  XOR U7792 ( .A(n7813), .B(n7810), .Z(n7812) );
  XOR U7793 ( .A(n7814), .B(n7815), .Z(n7799) );
  AND U7794 ( .A(n7816), .B(n7817), .Z(n7815) );
  XNOR U7795 ( .A(n7814), .B(n7728), .Z(n7817) );
  XOR U7796 ( .A(n7818), .B(n7808), .Z(n7728) );
  XNOR U7797 ( .A(n7819), .B(n7803), .Z(n7808) );
  XOR U7798 ( .A(n7820), .B(n7821), .Z(n7803) );
  AND U7799 ( .A(n7822), .B(n7823), .Z(n7821) );
  XOR U7800 ( .A(n7824), .B(n7820), .Z(n7822) );
  XNOR U7801 ( .A(n7825), .B(n7826), .Z(n7819) );
  AND U7802 ( .A(n7827), .B(n7828), .Z(n7826) );
  XOR U7803 ( .A(n7825), .B(n7829), .Z(n7827) );
  XNOR U7804 ( .A(n7809), .B(n7806), .Z(n7818) );
  AND U7805 ( .A(n7830), .B(n7831), .Z(n7806) );
  XOR U7806 ( .A(n7832), .B(n7833), .Z(n7809) );
  AND U7807 ( .A(n7834), .B(n7835), .Z(n7833) );
  XOR U7808 ( .A(n7832), .B(n7836), .Z(n7834) );
  XNOR U7809 ( .A(n7725), .B(n7814), .Z(n7816) );
  XOR U7810 ( .A(n7837), .B(n7838), .Z(n7725) );
  AND U7811 ( .A(n175), .B(n7839), .Z(n7838) );
  XNOR U7812 ( .A(n7840), .B(n7837), .Z(n7839) );
  XOR U7813 ( .A(n7841), .B(n7842), .Z(n7814) );
  AND U7814 ( .A(n7843), .B(n7844), .Z(n7842) );
  XNOR U7815 ( .A(n7841), .B(n7830), .Z(n7844) );
  IV U7816 ( .A(n7776), .Z(n7830) );
  XNOR U7817 ( .A(n7845), .B(n7823), .Z(n7776) );
  XNOR U7818 ( .A(n7846), .B(n7829), .Z(n7823) );
  XOR U7819 ( .A(n7847), .B(n7848), .Z(n7829) );
  NOR U7820 ( .A(n7849), .B(n7850), .Z(n7848) );
  XNOR U7821 ( .A(n7847), .B(n7851), .Z(n7849) );
  XNOR U7822 ( .A(n7828), .B(n7820), .Z(n7846) );
  XOR U7823 ( .A(n7852), .B(n7853), .Z(n7820) );
  AND U7824 ( .A(n7854), .B(n7855), .Z(n7853) );
  XNOR U7825 ( .A(n7852), .B(n7856), .Z(n7854) );
  XNOR U7826 ( .A(n7857), .B(n7825), .Z(n7828) );
  XOR U7827 ( .A(n7858), .B(n7859), .Z(n7825) );
  AND U7828 ( .A(n7860), .B(n7861), .Z(n7859) );
  XOR U7829 ( .A(n7858), .B(n7862), .Z(n7860) );
  XNOR U7830 ( .A(n7863), .B(n7864), .Z(n7857) );
  NOR U7831 ( .A(n7865), .B(n7866), .Z(n7864) );
  XOR U7832 ( .A(n7863), .B(n7867), .Z(n7865) );
  XNOR U7833 ( .A(n7824), .B(n7831), .Z(n7845) );
  NOR U7834 ( .A(n7788), .B(n7868), .Z(n7831) );
  XOR U7835 ( .A(n7836), .B(n7835), .Z(n7824) );
  XNOR U7836 ( .A(n7869), .B(n7832), .Z(n7835) );
  XOR U7837 ( .A(n7870), .B(n7871), .Z(n7832) );
  AND U7838 ( .A(n7872), .B(n7873), .Z(n7871) );
  XOR U7839 ( .A(n7870), .B(n7874), .Z(n7872) );
  XNOR U7840 ( .A(n7875), .B(n7876), .Z(n7869) );
  NOR U7841 ( .A(n7877), .B(n7878), .Z(n7876) );
  XNOR U7842 ( .A(n7875), .B(n7879), .Z(n7877) );
  XOR U7843 ( .A(n7880), .B(n7881), .Z(n7836) );
  NOR U7844 ( .A(n7882), .B(n7883), .Z(n7881) );
  XNOR U7845 ( .A(n7880), .B(n7884), .Z(n7882) );
  XNOR U7846 ( .A(n7773), .B(n7841), .Z(n7843) );
  XOR U7847 ( .A(n7885), .B(n7886), .Z(n7773) );
  AND U7848 ( .A(n175), .B(n7887), .Z(n7886) );
  XOR U7849 ( .A(n7888), .B(n7885), .Z(n7887) );
  AND U7850 ( .A(n7785), .B(n7788), .Z(n7841) );
  XOR U7851 ( .A(n7889), .B(n7868), .Z(n7788) );
  XNOR U7852 ( .A(p_input[1024]), .B(p_input[672]), .Z(n7868) );
  XOR U7853 ( .A(n7856), .B(n7855), .Z(n7889) );
  XNOR U7854 ( .A(n7890), .B(n7862), .Z(n7855) );
  XNOR U7855 ( .A(n7851), .B(n7850), .Z(n7862) );
  XOR U7856 ( .A(n7891), .B(n7847), .Z(n7850) );
  XOR U7857 ( .A(p_input[1034]), .B(p_input[682]), .Z(n7847) );
  XNOR U7858 ( .A(p_input[1035]), .B(p_input[683]), .Z(n7891) );
  XOR U7859 ( .A(p_input[1036]), .B(p_input[684]), .Z(n7851) );
  XNOR U7860 ( .A(n7861), .B(n7852), .Z(n7890) );
  XNOR U7861 ( .A(n3298), .B(p_input[673]), .Z(n7852) );
  XOR U7862 ( .A(n7892), .B(n7867), .Z(n7861) );
  XNOR U7863 ( .A(p_input[1039]), .B(p_input[687]), .Z(n7867) );
  XOR U7864 ( .A(n7858), .B(n7866), .Z(n7892) );
  XOR U7865 ( .A(n7893), .B(n7863), .Z(n7866) );
  XOR U7866 ( .A(p_input[1037]), .B(p_input[685]), .Z(n7863) );
  XNOR U7867 ( .A(p_input[1038]), .B(p_input[686]), .Z(n7893) );
  XOR U7868 ( .A(p_input[1033]), .B(p_input[681]), .Z(n7858) );
  XNOR U7869 ( .A(n7874), .B(n7873), .Z(n7856) );
  XNOR U7870 ( .A(n7894), .B(n7879), .Z(n7873) );
  XOR U7871 ( .A(p_input[1032]), .B(p_input[680]), .Z(n7879) );
  XOR U7872 ( .A(n7870), .B(n7878), .Z(n7894) );
  XOR U7873 ( .A(n7895), .B(n7875), .Z(n7878) );
  XOR U7874 ( .A(p_input[1030]), .B(p_input[678]), .Z(n7875) );
  XNOR U7875 ( .A(p_input[1031]), .B(p_input[679]), .Z(n7895) );
  XOR U7876 ( .A(p_input[1026]), .B(p_input[674]), .Z(n7870) );
  XNOR U7877 ( .A(n7884), .B(n7883), .Z(n7874) );
  XOR U7878 ( .A(n7896), .B(n7880), .Z(n7883) );
  XOR U7879 ( .A(p_input[1027]), .B(p_input[675]), .Z(n7880) );
  XNOR U7880 ( .A(p_input[1028]), .B(p_input[676]), .Z(n7896) );
  XOR U7881 ( .A(p_input[1029]), .B(p_input[677]), .Z(n7884) );
  XOR U7882 ( .A(n7897), .B(n7898), .Z(n7785) );
  AND U7883 ( .A(n175), .B(n7899), .Z(n7898) );
  XNOR U7884 ( .A(n7900), .B(n7897), .Z(n7899) );
  XNOR U7885 ( .A(n7901), .B(n7902), .Z(n175) );
  AND U7886 ( .A(n7903), .B(n7904), .Z(n7902) );
  XOR U7887 ( .A(n7798), .B(n7901), .Z(n7904) );
  AND U7888 ( .A(n7905), .B(n7906), .Z(n7798) );
  XNOR U7889 ( .A(n7795), .B(n7901), .Z(n7903) );
  XOR U7890 ( .A(n7907), .B(n7908), .Z(n7795) );
  AND U7891 ( .A(n179), .B(n7909), .Z(n7908) );
  XOR U7892 ( .A(n7910), .B(n7907), .Z(n7909) );
  XOR U7893 ( .A(n7911), .B(n7912), .Z(n7901) );
  AND U7894 ( .A(n7913), .B(n7914), .Z(n7912) );
  XNOR U7895 ( .A(n7911), .B(n7905), .Z(n7914) );
  IV U7896 ( .A(n7813), .Z(n7905) );
  XOR U7897 ( .A(n7915), .B(n7916), .Z(n7813) );
  XOR U7898 ( .A(n7917), .B(n7906), .Z(n7916) );
  AND U7899 ( .A(n7840), .B(n7918), .Z(n7906) );
  AND U7900 ( .A(n7919), .B(n7920), .Z(n7917) );
  XOR U7901 ( .A(n7921), .B(n7915), .Z(n7919) );
  XNOR U7902 ( .A(n7810), .B(n7911), .Z(n7913) );
  XOR U7903 ( .A(n7922), .B(n7923), .Z(n7810) );
  AND U7904 ( .A(n179), .B(n7924), .Z(n7923) );
  XOR U7905 ( .A(n7925), .B(n7922), .Z(n7924) );
  XOR U7906 ( .A(n7926), .B(n7927), .Z(n7911) );
  AND U7907 ( .A(n7928), .B(n7929), .Z(n7927) );
  XNOR U7908 ( .A(n7926), .B(n7840), .Z(n7929) );
  XOR U7909 ( .A(n7930), .B(n7920), .Z(n7840) );
  XNOR U7910 ( .A(n7931), .B(n7915), .Z(n7920) );
  XOR U7911 ( .A(n7932), .B(n7933), .Z(n7915) );
  AND U7912 ( .A(n7934), .B(n7935), .Z(n7933) );
  XOR U7913 ( .A(n7936), .B(n7932), .Z(n7934) );
  XNOR U7914 ( .A(n7937), .B(n7938), .Z(n7931) );
  AND U7915 ( .A(n7939), .B(n7940), .Z(n7938) );
  XOR U7916 ( .A(n7937), .B(n7941), .Z(n7939) );
  XNOR U7917 ( .A(n7921), .B(n7918), .Z(n7930) );
  AND U7918 ( .A(n7942), .B(n7943), .Z(n7918) );
  XOR U7919 ( .A(n7944), .B(n7945), .Z(n7921) );
  AND U7920 ( .A(n7946), .B(n7947), .Z(n7945) );
  XOR U7921 ( .A(n7944), .B(n7948), .Z(n7946) );
  XNOR U7922 ( .A(n7837), .B(n7926), .Z(n7928) );
  XOR U7923 ( .A(n7949), .B(n7950), .Z(n7837) );
  AND U7924 ( .A(n179), .B(n7951), .Z(n7950) );
  XNOR U7925 ( .A(n7952), .B(n7949), .Z(n7951) );
  XOR U7926 ( .A(n7953), .B(n7954), .Z(n7926) );
  AND U7927 ( .A(n7955), .B(n7956), .Z(n7954) );
  XNOR U7928 ( .A(n7953), .B(n7942), .Z(n7956) );
  IV U7929 ( .A(n7888), .Z(n7942) );
  XNOR U7930 ( .A(n7957), .B(n7935), .Z(n7888) );
  XNOR U7931 ( .A(n7958), .B(n7941), .Z(n7935) );
  XOR U7932 ( .A(n7959), .B(n7960), .Z(n7941) );
  NOR U7933 ( .A(n7961), .B(n7962), .Z(n7960) );
  XNOR U7934 ( .A(n7959), .B(n7963), .Z(n7961) );
  XNOR U7935 ( .A(n7940), .B(n7932), .Z(n7958) );
  XOR U7936 ( .A(n7964), .B(n7965), .Z(n7932) );
  AND U7937 ( .A(n7966), .B(n7967), .Z(n7965) );
  XNOR U7938 ( .A(n7964), .B(n7968), .Z(n7966) );
  XNOR U7939 ( .A(n7969), .B(n7937), .Z(n7940) );
  XOR U7940 ( .A(n7970), .B(n7971), .Z(n7937) );
  AND U7941 ( .A(n7972), .B(n7973), .Z(n7971) );
  XOR U7942 ( .A(n7970), .B(n7974), .Z(n7972) );
  XNOR U7943 ( .A(n7975), .B(n7976), .Z(n7969) );
  NOR U7944 ( .A(n7977), .B(n7978), .Z(n7976) );
  XOR U7945 ( .A(n7975), .B(n7979), .Z(n7977) );
  XNOR U7946 ( .A(n7936), .B(n7943), .Z(n7957) );
  NOR U7947 ( .A(n7900), .B(n7980), .Z(n7943) );
  XOR U7948 ( .A(n7948), .B(n7947), .Z(n7936) );
  XNOR U7949 ( .A(n7981), .B(n7944), .Z(n7947) );
  XOR U7950 ( .A(n7982), .B(n7983), .Z(n7944) );
  AND U7951 ( .A(n7984), .B(n7985), .Z(n7983) );
  XOR U7952 ( .A(n7982), .B(n7986), .Z(n7984) );
  XNOR U7953 ( .A(n7987), .B(n7988), .Z(n7981) );
  NOR U7954 ( .A(n7989), .B(n7990), .Z(n7988) );
  XNOR U7955 ( .A(n7987), .B(n7991), .Z(n7989) );
  XOR U7956 ( .A(n7992), .B(n7993), .Z(n7948) );
  NOR U7957 ( .A(n7994), .B(n7995), .Z(n7993) );
  XNOR U7958 ( .A(n7992), .B(n7996), .Z(n7994) );
  XNOR U7959 ( .A(n7885), .B(n7953), .Z(n7955) );
  XOR U7960 ( .A(n7997), .B(n7998), .Z(n7885) );
  AND U7961 ( .A(n179), .B(n7999), .Z(n7998) );
  XOR U7962 ( .A(n8000), .B(n7997), .Z(n7999) );
  AND U7963 ( .A(n7897), .B(n7900), .Z(n7953) );
  XOR U7964 ( .A(n8001), .B(n7980), .Z(n7900) );
  XNOR U7965 ( .A(p_input[1024]), .B(p_input[688]), .Z(n7980) );
  XOR U7966 ( .A(n7968), .B(n7967), .Z(n8001) );
  XNOR U7967 ( .A(n8002), .B(n7974), .Z(n7967) );
  XNOR U7968 ( .A(n7963), .B(n7962), .Z(n7974) );
  XOR U7969 ( .A(n8003), .B(n7959), .Z(n7962) );
  XOR U7970 ( .A(p_input[1034]), .B(p_input[698]), .Z(n7959) );
  XNOR U7971 ( .A(p_input[1035]), .B(p_input[699]), .Z(n8003) );
  XOR U7972 ( .A(p_input[1036]), .B(p_input[700]), .Z(n7963) );
  XNOR U7973 ( .A(n7973), .B(n7964), .Z(n8002) );
  XNOR U7974 ( .A(n3298), .B(p_input[689]), .Z(n7964) );
  XOR U7975 ( .A(n8004), .B(n7979), .Z(n7973) );
  XNOR U7976 ( .A(p_input[1039]), .B(p_input[703]), .Z(n7979) );
  XOR U7977 ( .A(n7970), .B(n7978), .Z(n8004) );
  XOR U7978 ( .A(n8005), .B(n7975), .Z(n7978) );
  XOR U7979 ( .A(p_input[1037]), .B(p_input[701]), .Z(n7975) );
  XNOR U7980 ( .A(p_input[1038]), .B(p_input[702]), .Z(n8005) );
  XOR U7981 ( .A(p_input[1033]), .B(p_input[697]), .Z(n7970) );
  XNOR U7982 ( .A(n7986), .B(n7985), .Z(n7968) );
  XNOR U7983 ( .A(n8006), .B(n7991), .Z(n7985) );
  XOR U7984 ( .A(p_input[1032]), .B(p_input[696]), .Z(n7991) );
  XOR U7985 ( .A(n7982), .B(n7990), .Z(n8006) );
  XOR U7986 ( .A(n8007), .B(n7987), .Z(n7990) );
  XOR U7987 ( .A(p_input[1030]), .B(p_input[694]), .Z(n7987) );
  XNOR U7988 ( .A(p_input[1031]), .B(p_input[695]), .Z(n8007) );
  XOR U7989 ( .A(p_input[1026]), .B(p_input[690]), .Z(n7982) );
  XNOR U7990 ( .A(n7996), .B(n7995), .Z(n7986) );
  XOR U7991 ( .A(n8008), .B(n7992), .Z(n7995) );
  XOR U7992 ( .A(p_input[1027]), .B(p_input[691]), .Z(n7992) );
  XNOR U7993 ( .A(p_input[1028]), .B(p_input[692]), .Z(n8008) );
  XOR U7994 ( .A(p_input[1029]), .B(p_input[693]), .Z(n7996) );
  XOR U7995 ( .A(n8009), .B(n8010), .Z(n7897) );
  AND U7996 ( .A(n179), .B(n8011), .Z(n8010) );
  XNOR U7997 ( .A(n8012), .B(n8009), .Z(n8011) );
  XNOR U7998 ( .A(n8013), .B(n8014), .Z(n179) );
  AND U7999 ( .A(n8015), .B(n8016), .Z(n8014) );
  XOR U8000 ( .A(n7910), .B(n8013), .Z(n8016) );
  AND U8001 ( .A(n8017), .B(n8018), .Z(n7910) );
  XNOR U8002 ( .A(n7907), .B(n8013), .Z(n8015) );
  XOR U8003 ( .A(n8019), .B(n8020), .Z(n7907) );
  AND U8004 ( .A(n183), .B(n8021), .Z(n8020) );
  XOR U8005 ( .A(n8022), .B(n8019), .Z(n8021) );
  XOR U8006 ( .A(n8023), .B(n8024), .Z(n8013) );
  AND U8007 ( .A(n8025), .B(n8026), .Z(n8024) );
  XNOR U8008 ( .A(n8023), .B(n8017), .Z(n8026) );
  IV U8009 ( .A(n7925), .Z(n8017) );
  XOR U8010 ( .A(n8027), .B(n8028), .Z(n7925) );
  XOR U8011 ( .A(n8029), .B(n8018), .Z(n8028) );
  AND U8012 ( .A(n7952), .B(n8030), .Z(n8018) );
  AND U8013 ( .A(n8031), .B(n8032), .Z(n8029) );
  XOR U8014 ( .A(n8033), .B(n8027), .Z(n8031) );
  XNOR U8015 ( .A(n7922), .B(n8023), .Z(n8025) );
  XOR U8016 ( .A(n8034), .B(n8035), .Z(n7922) );
  AND U8017 ( .A(n183), .B(n8036), .Z(n8035) );
  XOR U8018 ( .A(n8037), .B(n8034), .Z(n8036) );
  XOR U8019 ( .A(n8038), .B(n8039), .Z(n8023) );
  AND U8020 ( .A(n8040), .B(n8041), .Z(n8039) );
  XNOR U8021 ( .A(n8038), .B(n7952), .Z(n8041) );
  XOR U8022 ( .A(n8042), .B(n8032), .Z(n7952) );
  XNOR U8023 ( .A(n8043), .B(n8027), .Z(n8032) );
  XOR U8024 ( .A(n8044), .B(n8045), .Z(n8027) );
  AND U8025 ( .A(n8046), .B(n8047), .Z(n8045) );
  XOR U8026 ( .A(n8048), .B(n8044), .Z(n8046) );
  XNOR U8027 ( .A(n8049), .B(n8050), .Z(n8043) );
  AND U8028 ( .A(n8051), .B(n8052), .Z(n8050) );
  XOR U8029 ( .A(n8049), .B(n8053), .Z(n8051) );
  XNOR U8030 ( .A(n8033), .B(n8030), .Z(n8042) );
  AND U8031 ( .A(n8054), .B(n8055), .Z(n8030) );
  XOR U8032 ( .A(n8056), .B(n8057), .Z(n8033) );
  AND U8033 ( .A(n8058), .B(n8059), .Z(n8057) );
  XOR U8034 ( .A(n8056), .B(n8060), .Z(n8058) );
  XNOR U8035 ( .A(n7949), .B(n8038), .Z(n8040) );
  XOR U8036 ( .A(n8061), .B(n8062), .Z(n7949) );
  AND U8037 ( .A(n183), .B(n8063), .Z(n8062) );
  XNOR U8038 ( .A(n8064), .B(n8061), .Z(n8063) );
  XOR U8039 ( .A(n8065), .B(n8066), .Z(n8038) );
  AND U8040 ( .A(n8067), .B(n8068), .Z(n8066) );
  XNOR U8041 ( .A(n8065), .B(n8054), .Z(n8068) );
  IV U8042 ( .A(n8000), .Z(n8054) );
  XNOR U8043 ( .A(n8069), .B(n8047), .Z(n8000) );
  XNOR U8044 ( .A(n8070), .B(n8053), .Z(n8047) );
  XOR U8045 ( .A(n8071), .B(n8072), .Z(n8053) );
  NOR U8046 ( .A(n8073), .B(n8074), .Z(n8072) );
  XNOR U8047 ( .A(n8071), .B(n8075), .Z(n8073) );
  XNOR U8048 ( .A(n8052), .B(n8044), .Z(n8070) );
  XOR U8049 ( .A(n8076), .B(n8077), .Z(n8044) );
  AND U8050 ( .A(n8078), .B(n8079), .Z(n8077) );
  XNOR U8051 ( .A(n8076), .B(n8080), .Z(n8078) );
  XNOR U8052 ( .A(n8081), .B(n8049), .Z(n8052) );
  XOR U8053 ( .A(n8082), .B(n8083), .Z(n8049) );
  AND U8054 ( .A(n8084), .B(n8085), .Z(n8083) );
  XOR U8055 ( .A(n8082), .B(n8086), .Z(n8084) );
  XNOR U8056 ( .A(n8087), .B(n8088), .Z(n8081) );
  NOR U8057 ( .A(n8089), .B(n8090), .Z(n8088) );
  XOR U8058 ( .A(n8087), .B(n8091), .Z(n8089) );
  XNOR U8059 ( .A(n8048), .B(n8055), .Z(n8069) );
  NOR U8060 ( .A(n8012), .B(n8092), .Z(n8055) );
  XOR U8061 ( .A(n8060), .B(n8059), .Z(n8048) );
  XNOR U8062 ( .A(n8093), .B(n8056), .Z(n8059) );
  XOR U8063 ( .A(n8094), .B(n8095), .Z(n8056) );
  AND U8064 ( .A(n8096), .B(n8097), .Z(n8095) );
  XOR U8065 ( .A(n8094), .B(n8098), .Z(n8096) );
  XNOR U8066 ( .A(n8099), .B(n8100), .Z(n8093) );
  NOR U8067 ( .A(n8101), .B(n8102), .Z(n8100) );
  XNOR U8068 ( .A(n8099), .B(n8103), .Z(n8101) );
  XOR U8069 ( .A(n8104), .B(n8105), .Z(n8060) );
  NOR U8070 ( .A(n8106), .B(n8107), .Z(n8105) );
  XNOR U8071 ( .A(n8104), .B(n8108), .Z(n8106) );
  XNOR U8072 ( .A(n7997), .B(n8065), .Z(n8067) );
  XOR U8073 ( .A(n8109), .B(n8110), .Z(n7997) );
  AND U8074 ( .A(n183), .B(n8111), .Z(n8110) );
  XOR U8075 ( .A(n8112), .B(n8109), .Z(n8111) );
  AND U8076 ( .A(n8009), .B(n8012), .Z(n8065) );
  XOR U8077 ( .A(n8113), .B(n8092), .Z(n8012) );
  XNOR U8078 ( .A(p_input[1024]), .B(p_input[704]), .Z(n8092) );
  XOR U8079 ( .A(n8080), .B(n8079), .Z(n8113) );
  XNOR U8080 ( .A(n8114), .B(n8086), .Z(n8079) );
  XNOR U8081 ( .A(n8075), .B(n8074), .Z(n8086) );
  XOR U8082 ( .A(n8115), .B(n8071), .Z(n8074) );
  XOR U8083 ( .A(p_input[1034]), .B(p_input[714]), .Z(n8071) );
  XNOR U8084 ( .A(p_input[1035]), .B(p_input[715]), .Z(n8115) );
  XOR U8085 ( .A(p_input[1036]), .B(p_input[716]), .Z(n8075) );
  XNOR U8086 ( .A(n8085), .B(n8076), .Z(n8114) );
  XNOR U8087 ( .A(n3298), .B(p_input[705]), .Z(n8076) );
  XOR U8088 ( .A(n8116), .B(n8091), .Z(n8085) );
  XNOR U8089 ( .A(p_input[1039]), .B(p_input[719]), .Z(n8091) );
  XOR U8090 ( .A(n8082), .B(n8090), .Z(n8116) );
  XOR U8091 ( .A(n8117), .B(n8087), .Z(n8090) );
  XOR U8092 ( .A(p_input[1037]), .B(p_input[717]), .Z(n8087) );
  XNOR U8093 ( .A(p_input[1038]), .B(p_input[718]), .Z(n8117) );
  XOR U8094 ( .A(p_input[1033]), .B(p_input[713]), .Z(n8082) );
  XNOR U8095 ( .A(n8098), .B(n8097), .Z(n8080) );
  XNOR U8096 ( .A(n8118), .B(n8103), .Z(n8097) );
  XOR U8097 ( .A(p_input[1032]), .B(p_input[712]), .Z(n8103) );
  XOR U8098 ( .A(n8094), .B(n8102), .Z(n8118) );
  XOR U8099 ( .A(n8119), .B(n8099), .Z(n8102) );
  XOR U8100 ( .A(p_input[1030]), .B(p_input[710]), .Z(n8099) );
  XNOR U8101 ( .A(p_input[1031]), .B(p_input[711]), .Z(n8119) );
  XOR U8102 ( .A(p_input[1026]), .B(p_input[706]), .Z(n8094) );
  XNOR U8103 ( .A(n8108), .B(n8107), .Z(n8098) );
  XOR U8104 ( .A(n8120), .B(n8104), .Z(n8107) );
  XOR U8105 ( .A(p_input[1027]), .B(p_input[707]), .Z(n8104) );
  XNOR U8106 ( .A(p_input[1028]), .B(p_input[708]), .Z(n8120) );
  XOR U8107 ( .A(p_input[1029]), .B(p_input[709]), .Z(n8108) );
  XOR U8108 ( .A(n8121), .B(n8122), .Z(n8009) );
  AND U8109 ( .A(n183), .B(n8123), .Z(n8122) );
  XNOR U8110 ( .A(n8124), .B(n8121), .Z(n8123) );
  XNOR U8111 ( .A(n8125), .B(n8126), .Z(n183) );
  AND U8112 ( .A(n8127), .B(n8128), .Z(n8126) );
  XOR U8113 ( .A(n8022), .B(n8125), .Z(n8128) );
  AND U8114 ( .A(n8129), .B(n8130), .Z(n8022) );
  XNOR U8115 ( .A(n8019), .B(n8125), .Z(n8127) );
  XOR U8116 ( .A(n8131), .B(n8132), .Z(n8019) );
  AND U8117 ( .A(n187), .B(n8133), .Z(n8132) );
  XOR U8118 ( .A(n8134), .B(n8131), .Z(n8133) );
  XOR U8119 ( .A(n8135), .B(n8136), .Z(n8125) );
  AND U8120 ( .A(n8137), .B(n8138), .Z(n8136) );
  XNOR U8121 ( .A(n8135), .B(n8129), .Z(n8138) );
  IV U8122 ( .A(n8037), .Z(n8129) );
  XOR U8123 ( .A(n8139), .B(n8140), .Z(n8037) );
  XOR U8124 ( .A(n8141), .B(n8130), .Z(n8140) );
  AND U8125 ( .A(n8064), .B(n8142), .Z(n8130) );
  AND U8126 ( .A(n8143), .B(n8144), .Z(n8141) );
  XOR U8127 ( .A(n8145), .B(n8139), .Z(n8143) );
  XNOR U8128 ( .A(n8034), .B(n8135), .Z(n8137) );
  XOR U8129 ( .A(n8146), .B(n8147), .Z(n8034) );
  AND U8130 ( .A(n187), .B(n8148), .Z(n8147) );
  XOR U8131 ( .A(n8149), .B(n8146), .Z(n8148) );
  XOR U8132 ( .A(n8150), .B(n8151), .Z(n8135) );
  AND U8133 ( .A(n8152), .B(n8153), .Z(n8151) );
  XNOR U8134 ( .A(n8150), .B(n8064), .Z(n8153) );
  XOR U8135 ( .A(n8154), .B(n8144), .Z(n8064) );
  XNOR U8136 ( .A(n8155), .B(n8139), .Z(n8144) );
  XOR U8137 ( .A(n8156), .B(n8157), .Z(n8139) );
  AND U8138 ( .A(n8158), .B(n8159), .Z(n8157) );
  XOR U8139 ( .A(n8160), .B(n8156), .Z(n8158) );
  XNOR U8140 ( .A(n8161), .B(n8162), .Z(n8155) );
  AND U8141 ( .A(n8163), .B(n8164), .Z(n8162) );
  XOR U8142 ( .A(n8161), .B(n8165), .Z(n8163) );
  XNOR U8143 ( .A(n8145), .B(n8142), .Z(n8154) );
  AND U8144 ( .A(n8166), .B(n8167), .Z(n8142) );
  XOR U8145 ( .A(n8168), .B(n8169), .Z(n8145) );
  AND U8146 ( .A(n8170), .B(n8171), .Z(n8169) );
  XOR U8147 ( .A(n8168), .B(n8172), .Z(n8170) );
  XNOR U8148 ( .A(n8061), .B(n8150), .Z(n8152) );
  XOR U8149 ( .A(n8173), .B(n8174), .Z(n8061) );
  AND U8150 ( .A(n187), .B(n8175), .Z(n8174) );
  XNOR U8151 ( .A(n8176), .B(n8173), .Z(n8175) );
  XOR U8152 ( .A(n8177), .B(n8178), .Z(n8150) );
  AND U8153 ( .A(n8179), .B(n8180), .Z(n8178) );
  XNOR U8154 ( .A(n8177), .B(n8166), .Z(n8180) );
  IV U8155 ( .A(n8112), .Z(n8166) );
  XNOR U8156 ( .A(n8181), .B(n8159), .Z(n8112) );
  XNOR U8157 ( .A(n8182), .B(n8165), .Z(n8159) );
  XOR U8158 ( .A(n8183), .B(n8184), .Z(n8165) );
  NOR U8159 ( .A(n8185), .B(n8186), .Z(n8184) );
  XNOR U8160 ( .A(n8183), .B(n8187), .Z(n8185) );
  XNOR U8161 ( .A(n8164), .B(n8156), .Z(n8182) );
  XOR U8162 ( .A(n8188), .B(n8189), .Z(n8156) );
  AND U8163 ( .A(n8190), .B(n8191), .Z(n8189) );
  XNOR U8164 ( .A(n8188), .B(n8192), .Z(n8190) );
  XNOR U8165 ( .A(n8193), .B(n8161), .Z(n8164) );
  XOR U8166 ( .A(n8194), .B(n8195), .Z(n8161) );
  AND U8167 ( .A(n8196), .B(n8197), .Z(n8195) );
  XOR U8168 ( .A(n8194), .B(n8198), .Z(n8196) );
  XNOR U8169 ( .A(n8199), .B(n8200), .Z(n8193) );
  NOR U8170 ( .A(n8201), .B(n8202), .Z(n8200) );
  XOR U8171 ( .A(n8199), .B(n8203), .Z(n8201) );
  XNOR U8172 ( .A(n8160), .B(n8167), .Z(n8181) );
  NOR U8173 ( .A(n8124), .B(n8204), .Z(n8167) );
  XOR U8174 ( .A(n8172), .B(n8171), .Z(n8160) );
  XNOR U8175 ( .A(n8205), .B(n8168), .Z(n8171) );
  XOR U8176 ( .A(n8206), .B(n8207), .Z(n8168) );
  AND U8177 ( .A(n8208), .B(n8209), .Z(n8207) );
  XOR U8178 ( .A(n8206), .B(n8210), .Z(n8208) );
  XNOR U8179 ( .A(n8211), .B(n8212), .Z(n8205) );
  NOR U8180 ( .A(n8213), .B(n8214), .Z(n8212) );
  XNOR U8181 ( .A(n8211), .B(n8215), .Z(n8213) );
  XOR U8182 ( .A(n8216), .B(n8217), .Z(n8172) );
  NOR U8183 ( .A(n8218), .B(n8219), .Z(n8217) );
  XNOR U8184 ( .A(n8216), .B(n8220), .Z(n8218) );
  XNOR U8185 ( .A(n8109), .B(n8177), .Z(n8179) );
  XOR U8186 ( .A(n8221), .B(n8222), .Z(n8109) );
  AND U8187 ( .A(n187), .B(n8223), .Z(n8222) );
  XOR U8188 ( .A(n8224), .B(n8221), .Z(n8223) );
  AND U8189 ( .A(n8121), .B(n8124), .Z(n8177) );
  XOR U8190 ( .A(n8225), .B(n8204), .Z(n8124) );
  XNOR U8191 ( .A(p_input[1024]), .B(p_input[720]), .Z(n8204) );
  XOR U8192 ( .A(n8192), .B(n8191), .Z(n8225) );
  XNOR U8193 ( .A(n8226), .B(n8198), .Z(n8191) );
  XNOR U8194 ( .A(n8187), .B(n8186), .Z(n8198) );
  XOR U8195 ( .A(n8227), .B(n8183), .Z(n8186) );
  XOR U8196 ( .A(p_input[1034]), .B(p_input[730]), .Z(n8183) );
  XNOR U8197 ( .A(p_input[1035]), .B(p_input[731]), .Z(n8227) );
  XOR U8198 ( .A(p_input[1036]), .B(p_input[732]), .Z(n8187) );
  XNOR U8199 ( .A(n8197), .B(n8188), .Z(n8226) );
  XNOR U8200 ( .A(n3298), .B(p_input[721]), .Z(n8188) );
  XOR U8201 ( .A(n8228), .B(n8203), .Z(n8197) );
  XNOR U8202 ( .A(p_input[1039]), .B(p_input[735]), .Z(n8203) );
  XOR U8203 ( .A(n8194), .B(n8202), .Z(n8228) );
  XOR U8204 ( .A(n8229), .B(n8199), .Z(n8202) );
  XOR U8205 ( .A(p_input[1037]), .B(p_input[733]), .Z(n8199) );
  XNOR U8206 ( .A(p_input[1038]), .B(p_input[734]), .Z(n8229) );
  XOR U8207 ( .A(p_input[1033]), .B(p_input[729]), .Z(n8194) );
  XNOR U8208 ( .A(n8210), .B(n8209), .Z(n8192) );
  XNOR U8209 ( .A(n8230), .B(n8215), .Z(n8209) );
  XOR U8210 ( .A(p_input[1032]), .B(p_input[728]), .Z(n8215) );
  XOR U8211 ( .A(n8206), .B(n8214), .Z(n8230) );
  XOR U8212 ( .A(n8231), .B(n8211), .Z(n8214) );
  XOR U8213 ( .A(p_input[1030]), .B(p_input[726]), .Z(n8211) );
  XNOR U8214 ( .A(p_input[1031]), .B(p_input[727]), .Z(n8231) );
  XOR U8215 ( .A(p_input[1026]), .B(p_input[722]), .Z(n8206) );
  XNOR U8216 ( .A(n8220), .B(n8219), .Z(n8210) );
  XOR U8217 ( .A(n8232), .B(n8216), .Z(n8219) );
  XOR U8218 ( .A(p_input[1027]), .B(p_input[723]), .Z(n8216) );
  XNOR U8219 ( .A(p_input[1028]), .B(p_input[724]), .Z(n8232) );
  XOR U8220 ( .A(p_input[1029]), .B(p_input[725]), .Z(n8220) );
  XOR U8221 ( .A(n8233), .B(n8234), .Z(n8121) );
  AND U8222 ( .A(n187), .B(n8235), .Z(n8234) );
  XNOR U8223 ( .A(n8236), .B(n8233), .Z(n8235) );
  XNOR U8224 ( .A(n8237), .B(n8238), .Z(n187) );
  AND U8225 ( .A(n8239), .B(n8240), .Z(n8238) );
  XOR U8226 ( .A(n8134), .B(n8237), .Z(n8240) );
  AND U8227 ( .A(n8241), .B(n8242), .Z(n8134) );
  XNOR U8228 ( .A(n8131), .B(n8237), .Z(n8239) );
  XOR U8229 ( .A(n8243), .B(n8244), .Z(n8131) );
  AND U8230 ( .A(n191), .B(n8245), .Z(n8244) );
  XOR U8231 ( .A(n8246), .B(n8243), .Z(n8245) );
  XOR U8232 ( .A(n8247), .B(n8248), .Z(n8237) );
  AND U8233 ( .A(n8249), .B(n8250), .Z(n8248) );
  XNOR U8234 ( .A(n8247), .B(n8241), .Z(n8250) );
  IV U8235 ( .A(n8149), .Z(n8241) );
  XOR U8236 ( .A(n8251), .B(n8252), .Z(n8149) );
  XOR U8237 ( .A(n8253), .B(n8242), .Z(n8252) );
  AND U8238 ( .A(n8176), .B(n8254), .Z(n8242) );
  AND U8239 ( .A(n8255), .B(n8256), .Z(n8253) );
  XOR U8240 ( .A(n8257), .B(n8251), .Z(n8255) );
  XNOR U8241 ( .A(n8146), .B(n8247), .Z(n8249) );
  XOR U8242 ( .A(n8258), .B(n8259), .Z(n8146) );
  AND U8243 ( .A(n191), .B(n8260), .Z(n8259) );
  XOR U8244 ( .A(n8261), .B(n8258), .Z(n8260) );
  XOR U8245 ( .A(n8262), .B(n8263), .Z(n8247) );
  AND U8246 ( .A(n8264), .B(n8265), .Z(n8263) );
  XNOR U8247 ( .A(n8262), .B(n8176), .Z(n8265) );
  XOR U8248 ( .A(n8266), .B(n8256), .Z(n8176) );
  XNOR U8249 ( .A(n8267), .B(n8251), .Z(n8256) );
  XOR U8250 ( .A(n8268), .B(n8269), .Z(n8251) );
  AND U8251 ( .A(n8270), .B(n8271), .Z(n8269) );
  XOR U8252 ( .A(n8272), .B(n8268), .Z(n8270) );
  XNOR U8253 ( .A(n8273), .B(n8274), .Z(n8267) );
  AND U8254 ( .A(n8275), .B(n8276), .Z(n8274) );
  XOR U8255 ( .A(n8273), .B(n8277), .Z(n8275) );
  XNOR U8256 ( .A(n8257), .B(n8254), .Z(n8266) );
  AND U8257 ( .A(n8278), .B(n8279), .Z(n8254) );
  XOR U8258 ( .A(n8280), .B(n8281), .Z(n8257) );
  AND U8259 ( .A(n8282), .B(n8283), .Z(n8281) );
  XOR U8260 ( .A(n8280), .B(n8284), .Z(n8282) );
  XNOR U8261 ( .A(n8173), .B(n8262), .Z(n8264) );
  XOR U8262 ( .A(n8285), .B(n8286), .Z(n8173) );
  AND U8263 ( .A(n191), .B(n8287), .Z(n8286) );
  XNOR U8264 ( .A(n8288), .B(n8285), .Z(n8287) );
  XOR U8265 ( .A(n8289), .B(n8290), .Z(n8262) );
  AND U8266 ( .A(n8291), .B(n8292), .Z(n8290) );
  XNOR U8267 ( .A(n8289), .B(n8278), .Z(n8292) );
  IV U8268 ( .A(n8224), .Z(n8278) );
  XNOR U8269 ( .A(n8293), .B(n8271), .Z(n8224) );
  XNOR U8270 ( .A(n8294), .B(n8277), .Z(n8271) );
  XOR U8271 ( .A(n8295), .B(n8296), .Z(n8277) );
  NOR U8272 ( .A(n8297), .B(n8298), .Z(n8296) );
  XNOR U8273 ( .A(n8295), .B(n8299), .Z(n8297) );
  XNOR U8274 ( .A(n8276), .B(n8268), .Z(n8294) );
  XOR U8275 ( .A(n8300), .B(n8301), .Z(n8268) );
  AND U8276 ( .A(n8302), .B(n8303), .Z(n8301) );
  XNOR U8277 ( .A(n8300), .B(n8304), .Z(n8302) );
  XNOR U8278 ( .A(n8305), .B(n8273), .Z(n8276) );
  XOR U8279 ( .A(n8306), .B(n8307), .Z(n8273) );
  AND U8280 ( .A(n8308), .B(n8309), .Z(n8307) );
  XOR U8281 ( .A(n8306), .B(n8310), .Z(n8308) );
  XNOR U8282 ( .A(n8311), .B(n8312), .Z(n8305) );
  NOR U8283 ( .A(n8313), .B(n8314), .Z(n8312) );
  XOR U8284 ( .A(n8311), .B(n8315), .Z(n8313) );
  XNOR U8285 ( .A(n8272), .B(n8279), .Z(n8293) );
  NOR U8286 ( .A(n8236), .B(n8316), .Z(n8279) );
  XOR U8287 ( .A(n8284), .B(n8283), .Z(n8272) );
  XNOR U8288 ( .A(n8317), .B(n8280), .Z(n8283) );
  XOR U8289 ( .A(n8318), .B(n8319), .Z(n8280) );
  AND U8290 ( .A(n8320), .B(n8321), .Z(n8319) );
  XOR U8291 ( .A(n8318), .B(n8322), .Z(n8320) );
  XNOR U8292 ( .A(n8323), .B(n8324), .Z(n8317) );
  NOR U8293 ( .A(n8325), .B(n8326), .Z(n8324) );
  XNOR U8294 ( .A(n8323), .B(n8327), .Z(n8325) );
  XOR U8295 ( .A(n8328), .B(n8329), .Z(n8284) );
  NOR U8296 ( .A(n8330), .B(n8331), .Z(n8329) );
  XNOR U8297 ( .A(n8328), .B(n8332), .Z(n8330) );
  XNOR U8298 ( .A(n8221), .B(n8289), .Z(n8291) );
  XOR U8299 ( .A(n8333), .B(n8334), .Z(n8221) );
  AND U8300 ( .A(n191), .B(n8335), .Z(n8334) );
  XOR U8301 ( .A(n8336), .B(n8333), .Z(n8335) );
  AND U8302 ( .A(n8233), .B(n8236), .Z(n8289) );
  XOR U8303 ( .A(n8337), .B(n8316), .Z(n8236) );
  XNOR U8304 ( .A(p_input[1024]), .B(p_input[736]), .Z(n8316) );
  XOR U8305 ( .A(n8304), .B(n8303), .Z(n8337) );
  XNOR U8306 ( .A(n8338), .B(n8310), .Z(n8303) );
  XNOR U8307 ( .A(n8299), .B(n8298), .Z(n8310) );
  XOR U8308 ( .A(n8339), .B(n8295), .Z(n8298) );
  XOR U8309 ( .A(p_input[1034]), .B(p_input[746]), .Z(n8295) );
  XNOR U8310 ( .A(p_input[1035]), .B(p_input[747]), .Z(n8339) );
  XOR U8311 ( .A(p_input[1036]), .B(p_input[748]), .Z(n8299) );
  XNOR U8312 ( .A(n8309), .B(n8300), .Z(n8338) );
  XNOR U8313 ( .A(n3298), .B(p_input[737]), .Z(n8300) );
  XOR U8314 ( .A(n8340), .B(n8315), .Z(n8309) );
  XNOR U8315 ( .A(p_input[1039]), .B(p_input[751]), .Z(n8315) );
  XOR U8316 ( .A(n8306), .B(n8314), .Z(n8340) );
  XOR U8317 ( .A(n8341), .B(n8311), .Z(n8314) );
  XOR U8318 ( .A(p_input[1037]), .B(p_input[749]), .Z(n8311) );
  XNOR U8319 ( .A(p_input[1038]), .B(p_input[750]), .Z(n8341) );
  XOR U8320 ( .A(p_input[1033]), .B(p_input[745]), .Z(n8306) );
  XNOR U8321 ( .A(n8322), .B(n8321), .Z(n8304) );
  XNOR U8322 ( .A(n8342), .B(n8327), .Z(n8321) );
  XOR U8323 ( .A(p_input[1032]), .B(p_input[744]), .Z(n8327) );
  XOR U8324 ( .A(n8318), .B(n8326), .Z(n8342) );
  XOR U8325 ( .A(n8343), .B(n8323), .Z(n8326) );
  XOR U8326 ( .A(p_input[1030]), .B(p_input[742]), .Z(n8323) );
  XNOR U8327 ( .A(p_input[1031]), .B(p_input[743]), .Z(n8343) );
  XOR U8328 ( .A(p_input[1026]), .B(p_input[738]), .Z(n8318) );
  XNOR U8329 ( .A(n8332), .B(n8331), .Z(n8322) );
  XOR U8330 ( .A(n8344), .B(n8328), .Z(n8331) );
  XOR U8331 ( .A(p_input[1027]), .B(p_input[739]), .Z(n8328) );
  XNOR U8332 ( .A(p_input[1028]), .B(p_input[740]), .Z(n8344) );
  XOR U8333 ( .A(p_input[1029]), .B(p_input[741]), .Z(n8332) );
  XOR U8334 ( .A(n8345), .B(n8346), .Z(n8233) );
  AND U8335 ( .A(n191), .B(n8347), .Z(n8346) );
  XNOR U8336 ( .A(n8348), .B(n8345), .Z(n8347) );
  XNOR U8337 ( .A(n8349), .B(n8350), .Z(n191) );
  AND U8338 ( .A(n8351), .B(n8352), .Z(n8350) );
  XOR U8339 ( .A(n8246), .B(n8349), .Z(n8352) );
  AND U8340 ( .A(n8353), .B(n8354), .Z(n8246) );
  XNOR U8341 ( .A(n8243), .B(n8349), .Z(n8351) );
  XOR U8342 ( .A(n8355), .B(n8356), .Z(n8243) );
  AND U8343 ( .A(n195), .B(n8357), .Z(n8356) );
  XOR U8344 ( .A(n8358), .B(n8355), .Z(n8357) );
  XOR U8345 ( .A(n8359), .B(n8360), .Z(n8349) );
  AND U8346 ( .A(n8361), .B(n8362), .Z(n8360) );
  XNOR U8347 ( .A(n8359), .B(n8353), .Z(n8362) );
  IV U8348 ( .A(n8261), .Z(n8353) );
  XOR U8349 ( .A(n8363), .B(n8364), .Z(n8261) );
  XOR U8350 ( .A(n8365), .B(n8354), .Z(n8364) );
  AND U8351 ( .A(n8288), .B(n8366), .Z(n8354) );
  AND U8352 ( .A(n8367), .B(n8368), .Z(n8365) );
  XOR U8353 ( .A(n8369), .B(n8363), .Z(n8367) );
  XNOR U8354 ( .A(n8258), .B(n8359), .Z(n8361) );
  XOR U8355 ( .A(n8370), .B(n8371), .Z(n8258) );
  AND U8356 ( .A(n195), .B(n8372), .Z(n8371) );
  XOR U8357 ( .A(n8373), .B(n8370), .Z(n8372) );
  XOR U8358 ( .A(n8374), .B(n8375), .Z(n8359) );
  AND U8359 ( .A(n8376), .B(n8377), .Z(n8375) );
  XNOR U8360 ( .A(n8374), .B(n8288), .Z(n8377) );
  XOR U8361 ( .A(n8378), .B(n8368), .Z(n8288) );
  XNOR U8362 ( .A(n8379), .B(n8363), .Z(n8368) );
  XOR U8363 ( .A(n8380), .B(n8381), .Z(n8363) );
  AND U8364 ( .A(n8382), .B(n8383), .Z(n8381) );
  XOR U8365 ( .A(n8384), .B(n8380), .Z(n8382) );
  XNOR U8366 ( .A(n8385), .B(n8386), .Z(n8379) );
  AND U8367 ( .A(n8387), .B(n8388), .Z(n8386) );
  XOR U8368 ( .A(n8385), .B(n8389), .Z(n8387) );
  XNOR U8369 ( .A(n8369), .B(n8366), .Z(n8378) );
  AND U8370 ( .A(n8390), .B(n8391), .Z(n8366) );
  XOR U8371 ( .A(n8392), .B(n8393), .Z(n8369) );
  AND U8372 ( .A(n8394), .B(n8395), .Z(n8393) );
  XOR U8373 ( .A(n8392), .B(n8396), .Z(n8394) );
  XNOR U8374 ( .A(n8285), .B(n8374), .Z(n8376) );
  XOR U8375 ( .A(n8397), .B(n8398), .Z(n8285) );
  AND U8376 ( .A(n195), .B(n8399), .Z(n8398) );
  XNOR U8377 ( .A(n8400), .B(n8397), .Z(n8399) );
  XOR U8378 ( .A(n8401), .B(n8402), .Z(n8374) );
  AND U8379 ( .A(n8403), .B(n8404), .Z(n8402) );
  XNOR U8380 ( .A(n8401), .B(n8390), .Z(n8404) );
  IV U8381 ( .A(n8336), .Z(n8390) );
  XNOR U8382 ( .A(n8405), .B(n8383), .Z(n8336) );
  XNOR U8383 ( .A(n8406), .B(n8389), .Z(n8383) );
  XOR U8384 ( .A(n8407), .B(n8408), .Z(n8389) );
  NOR U8385 ( .A(n8409), .B(n8410), .Z(n8408) );
  XNOR U8386 ( .A(n8407), .B(n8411), .Z(n8409) );
  XNOR U8387 ( .A(n8388), .B(n8380), .Z(n8406) );
  XOR U8388 ( .A(n8412), .B(n8413), .Z(n8380) );
  AND U8389 ( .A(n8414), .B(n8415), .Z(n8413) );
  XNOR U8390 ( .A(n8412), .B(n8416), .Z(n8414) );
  XNOR U8391 ( .A(n8417), .B(n8385), .Z(n8388) );
  XOR U8392 ( .A(n8418), .B(n8419), .Z(n8385) );
  AND U8393 ( .A(n8420), .B(n8421), .Z(n8419) );
  XOR U8394 ( .A(n8418), .B(n8422), .Z(n8420) );
  XNOR U8395 ( .A(n8423), .B(n8424), .Z(n8417) );
  NOR U8396 ( .A(n8425), .B(n8426), .Z(n8424) );
  XOR U8397 ( .A(n8423), .B(n8427), .Z(n8425) );
  XNOR U8398 ( .A(n8384), .B(n8391), .Z(n8405) );
  NOR U8399 ( .A(n8348), .B(n8428), .Z(n8391) );
  XOR U8400 ( .A(n8396), .B(n8395), .Z(n8384) );
  XNOR U8401 ( .A(n8429), .B(n8392), .Z(n8395) );
  XOR U8402 ( .A(n8430), .B(n8431), .Z(n8392) );
  AND U8403 ( .A(n8432), .B(n8433), .Z(n8431) );
  XOR U8404 ( .A(n8430), .B(n8434), .Z(n8432) );
  XNOR U8405 ( .A(n8435), .B(n8436), .Z(n8429) );
  NOR U8406 ( .A(n8437), .B(n8438), .Z(n8436) );
  XNOR U8407 ( .A(n8435), .B(n8439), .Z(n8437) );
  XOR U8408 ( .A(n8440), .B(n8441), .Z(n8396) );
  NOR U8409 ( .A(n8442), .B(n8443), .Z(n8441) );
  XNOR U8410 ( .A(n8440), .B(n8444), .Z(n8442) );
  XNOR U8411 ( .A(n8333), .B(n8401), .Z(n8403) );
  XOR U8412 ( .A(n8445), .B(n8446), .Z(n8333) );
  AND U8413 ( .A(n195), .B(n8447), .Z(n8446) );
  XOR U8414 ( .A(n8448), .B(n8445), .Z(n8447) );
  AND U8415 ( .A(n8345), .B(n8348), .Z(n8401) );
  XOR U8416 ( .A(n8449), .B(n8428), .Z(n8348) );
  XNOR U8417 ( .A(p_input[1024]), .B(p_input[752]), .Z(n8428) );
  XOR U8418 ( .A(n8416), .B(n8415), .Z(n8449) );
  XNOR U8419 ( .A(n8450), .B(n8422), .Z(n8415) );
  XNOR U8420 ( .A(n8411), .B(n8410), .Z(n8422) );
  XOR U8421 ( .A(n8451), .B(n8407), .Z(n8410) );
  XOR U8422 ( .A(p_input[1034]), .B(p_input[762]), .Z(n8407) );
  XNOR U8423 ( .A(p_input[1035]), .B(p_input[763]), .Z(n8451) );
  XOR U8424 ( .A(p_input[1036]), .B(p_input[764]), .Z(n8411) );
  XNOR U8425 ( .A(n8421), .B(n8412), .Z(n8450) );
  XNOR U8426 ( .A(n3298), .B(p_input[753]), .Z(n8412) );
  XOR U8427 ( .A(n8452), .B(n8427), .Z(n8421) );
  XNOR U8428 ( .A(p_input[1039]), .B(p_input[767]), .Z(n8427) );
  XOR U8429 ( .A(n8418), .B(n8426), .Z(n8452) );
  XOR U8430 ( .A(n8453), .B(n8423), .Z(n8426) );
  XOR U8431 ( .A(p_input[1037]), .B(p_input[765]), .Z(n8423) );
  XNOR U8432 ( .A(p_input[1038]), .B(p_input[766]), .Z(n8453) );
  XOR U8433 ( .A(p_input[1033]), .B(p_input[761]), .Z(n8418) );
  XNOR U8434 ( .A(n8434), .B(n8433), .Z(n8416) );
  XNOR U8435 ( .A(n8454), .B(n8439), .Z(n8433) );
  XOR U8436 ( .A(p_input[1032]), .B(p_input[760]), .Z(n8439) );
  XOR U8437 ( .A(n8430), .B(n8438), .Z(n8454) );
  XOR U8438 ( .A(n8455), .B(n8435), .Z(n8438) );
  XOR U8439 ( .A(p_input[1030]), .B(p_input[758]), .Z(n8435) );
  XNOR U8440 ( .A(p_input[1031]), .B(p_input[759]), .Z(n8455) );
  XOR U8441 ( .A(p_input[1026]), .B(p_input[754]), .Z(n8430) );
  XNOR U8442 ( .A(n8444), .B(n8443), .Z(n8434) );
  XOR U8443 ( .A(n8456), .B(n8440), .Z(n8443) );
  XOR U8444 ( .A(p_input[1027]), .B(p_input[755]), .Z(n8440) );
  XNOR U8445 ( .A(p_input[1028]), .B(p_input[756]), .Z(n8456) );
  XOR U8446 ( .A(p_input[1029]), .B(p_input[757]), .Z(n8444) );
  XOR U8447 ( .A(n8457), .B(n8458), .Z(n8345) );
  AND U8448 ( .A(n195), .B(n8459), .Z(n8458) );
  XNOR U8449 ( .A(n8460), .B(n8457), .Z(n8459) );
  XNOR U8450 ( .A(n8461), .B(n8462), .Z(n195) );
  AND U8451 ( .A(n8463), .B(n8464), .Z(n8462) );
  XOR U8452 ( .A(n8358), .B(n8461), .Z(n8464) );
  AND U8453 ( .A(n8465), .B(n8466), .Z(n8358) );
  XNOR U8454 ( .A(n8355), .B(n8461), .Z(n8463) );
  XOR U8455 ( .A(n8467), .B(n8468), .Z(n8355) );
  AND U8456 ( .A(n199), .B(n8469), .Z(n8468) );
  XOR U8457 ( .A(n8470), .B(n8467), .Z(n8469) );
  XOR U8458 ( .A(n8471), .B(n8472), .Z(n8461) );
  AND U8459 ( .A(n8473), .B(n8474), .Z(n8472) );
  XNOR U8460 ( .A(n8471), .B(n8465), .Z(n8474) );
  IV U8461 ( .A(n8373), .Z(n8465) );
  XOR U8462 ( .A(n8475), .B(n8476), .Z(n8373) );
  XOR U8463 ( .A(n8477), .B(n8466), .Z(n8476) );
  AND U8464 ( .A(n8400), .B(n8478), .Z(n8466) );
  AND U8465 ( .A(n8479), .B(n8480), .Z(n8477) );
  XOR U8466 ( .A(n8481), .B(n8475), .Z(n8479) );
  XNOR U8467 ( .A(n8370), .B(n8471), .Z(n8473) );
  XOR U8468 ( .A(n8482), .B(n8483), .Z(n8370) );
  AND U8469 ( .A(n199), .B(n8484), .Z(n8483) );
  XOR U8470 ( .A(n8485), .B(n8482), .Z(n8484) );
  XOR U8471 ( .A(n8486), .B(n8487), .Z(n8471) );
  AND U8472 ( .A(n8488), .B(n8489), .Z(n8487) );
  XNOR U8473 ( .A(n8486), .B(n8400), .Z(n8489) );
  XOR U8474 ( .A(n8490), .B(n8480), .Z(n8400) );
  XNOR U8475 ( .A(n8491), .B(n8475), .Z(n8480) );
  XOR U8476 ( .A(n8492), .B(n8493), .Z(n8475) );
  AND U8477 ( .A(n8494), .B(n8495), .Z(n8493) );
  XOR U8478 ( .A(n8496), .B(n8492), .Z(n8494) );
  XNOR U8479 ( .A(n8497), .B(n8498), .Z(n8491) );
  AND U8480 ( .A(n8499), .B(n8500), .Z(n8498) );
  XOR U8481 ( .A(n8497), .B(n8501), .Z(n8499) );
  XNOR U8482 ( .A(n8481), .B(n8478), .Z(n8490) );
  AND U8483 ( .A(n8502), .B(n8503), .Z(n8478) );
  XOR U8484 ( .A(n8504), .B(n8505), .Z(n8481) );
  AND U8485 ( .A(n8506), .B(n8507), .Z(n8505) );
  XOR U8486 ( .A(n8504), .B(n8508), .Z(n8506) );
  XNOR U8487 ( .A(n8397), .B(n8486), .Z(n8488) );
  XOR U8488 ( .A(n8509), .B(n8510), .Z(n8397) );
  AND U8489 ( .A(n199), .B(n8511), .Z(n8510) );
  XNOR U8490 ( .A(n8512), .B(n8509), .Z(n8511) );
  XOR U8491 ( .A(n8513), .B(n8514), .Z(n8486) );
  AND U8492 ( .A(n8515), .B(n8516), .Z(n8514) );
  XNOR U8493 ( .A(n8513), .B(n8502), .Z(n8516) );
  IV U8494 ( .A(n8448), .Z(n8502) );
  XNOR U8495 ( .A(n8517), .B(n8495), .Z(n8448) );
  XNOR U8496 ( .A(n8518), .B(n8501), .Z(n8495) );
  XOR U8497 ( .A(n8519), .B(n8520), .Z(n8501) );
  NOR U8498 ( .A(n8521), .B(n8522), .Z(n8520) );
  XNOR U8499 ( .A(n8519), .B(n8523), .Z(n8521) );
  XNOR U8500 ( .A(n8500), .B(n8492), .Z(n8518) );
  XOR U8501 ( .A(n8524), .B(n8525), .Z(n8492) );
  AND U8502 ( .A(n8526), .B(n8527), .Z(n8525) );
  XNOR U8503 ( .A(n8524), .B(n8528), .Z(n8526) );
  XNOR U8504 ( .A(n8529), .B(n8497), .Z(n8500) );
  XOR U8505 ( .A(n8530), .B(n8531), .Z(n8497) );
  AND U8506 ( .A(n8532), .B(n8533), .Z(n8531) );
  XOR U8507 ( .A(n8530), .B(n8534), .Z(n8532) );
  XNOR U8508 ( .A(n8535), .B(n8536), .Z(n8529) );
  NOR U8509 ( .A(n8537), .B(n8538), .Z(n8536) );
  XOR U8510 ( .A(n8535), .B(n8539), .Z(n8537) );
  XNOR U8511 ( .A(n8496), .B(n8503), .Z(n8517) );
  NOR U8512 ( .A(n8460), .B(n8540), .Z(n8503) );
  XOR U8513 ( .A(n8508), .B(n8507), .Z(n8496) );
  XNOR U8514 ( .A(n8541), .B(n8504), .Z(n8507) );
  XOR U8515 ( .A(n8542), .B(n8543), .Z(n8504) );
  AND U8516 ( .A(n8544), .B(n8545), .Z(n8543) );
  XOR U8517 ( .A(n8542), .B(n8546), .Z(n8544) );
  XNOR U8518 ( .A(n8547), .B(n8548), .Z(n8541) );
  NOR U8519 ( .A(n8549), .B(n8550), .Z(n8548) );
  XNOR U8520 ( .A(n8547), .B(n8551), .Z(n8549) );
  XOR U8521 ( .A(n8552), .B(n8553), .Z(n8508) );
  NOR U8522 ( .A(n8554), .B(n8555), .Z(n8553) );
  XNOR U8523 ( .A(n8552), .B(n8556), .Z(n8554) );
  XNOR U8524 ( .A(n8445), .B(n8513), .Z(n8515) );
  XOR U8525 ( .A(n8557), .B(n8558), .Z(n8445) );
  AND U8526 ( .A(n199), .B(n8559), .Z(n8558) );
  XOR U8527 ( .A(n8560), .B(n8557), .Z(n8559) );
  AND U8528 ( .A(n8457), .B(n8460), .Z(n8513) );
  XOR U8529 ( .A(n8561), .B(n8540), .Z(n8460) );
  XNOR U8530 ( .A(p_input[1024]), .B(p_input[768]), .Z(n8540) );
  XOR U8531 ( .A(n8528), .B(n8527), .Z(n8561) );
  XNOR U8532 ( .A(n8562), .B(n8534), .Z(n8527) );
  XNOR U8533 ( .A(n8523), .B(n8522), .Z(n8534) );
  XOR U8534 ( .A(n8563), .B(n8519), .Z(n8522) );
  XOR U8535 ( .A(p_input[1034]), .B(p_input[778]), .Z(n8519) );
  XNOR U8536 ( .A(p_input[1035]), .B(p_input[779]), .Z(n8563) );
  XOR U8537 ( .A(p_input[1036]), .B(p_input[780]), .Z(n8523) );
  XNOR U8538 ( .A(n8533), .B(n8524), .Z(n8562) );
  XNOR U8539 ( .A(n3298), .B(p_input[769]), .Z(n8524) );
  XOR U8540 ( .A(n8564), .B(n8539), .Z(n8533) );
  XNOR U8541 ( .A(p_input[1039]), .B(p_input[783]), .Z(n8539) );
  XOR U8542 ( .A(n8530), .B(n8538), .Z(n8564) );
  XOR U8543 ( .A(n8565), .B(n8535), .Z(n8538) );
  XOR U8544 ( .A(p_input[1037]), .B(p_input[781]), .Z(n8535) );
  XNOR U8545 ( .A(p_input[1038]), .B(p_input[782]), .Z(n8565) );
  XOR U8546 ( .A(p_input[1033]), .B(p_input[777]), .Z(n8530) );
  XNOR U8547 ( .A(n8546), .B(n8545), .Z(n8528) );
  XNOR U8548 ( .A(n8566), .B(n8551), .Z(n8545) );
  XOR U8549 ( .A(p_input[1032]), .B(p_input[776]), .Z(n8551) );
  XOR U8550 ( .A(n8542), .B(n8550), .Z(n8566) );
  XOR U8551 ( .A(n8567), .B(n8547), .Z(n8550) );
  XOR U8552 ( .A(p_input[1030]), .B(p_input[774]), .Z(n8547) );
  XNOR U8553 ( .A(p_input[1031]), .B(p_input[775]), .Z(n8567) );
  XOR U8554 ( .A(p_input[1026]), .B(p_input[770]), .Z(n8542) );
  XNOR U8555 ( .A(n8556), .B(n8555), .Z(n8546) );
  XOR U8556 ( .A(n8568), .B(n8552), .Z(n8555) );
  XOR U8557 ( .A(p_input[1027]), .B(p_input[771]), .Z(n8552) );
  XNOR U8558 ( .A(p_input[1028]), .B(p_input[772]), .Z(n8568) );
  XOR U8559 ( .A(p_input[1029]), .B(p_input[773]), .Z(n8556) );
  XOR U8560 ( .A(n8569), .B(n8570), .Z(n8457) );
  AND U8561 ( .A(n199), .B(n8571), .Z(n8570) );
  XNOR U8562 ( .A(n8572), .B(n8569), .Z(n8571) );
  XNOR U8563 ( .A(n8573), .B(n8574), .Z(n199) );
  AND U8564 ( .A(n8575), .B(n8576), .Z(n8574) );
  XOR U8565 ( .A(n8470), .B(n8573), .Z(n8576) );
  AND U8566 ( .A(n8577), .B(n8578), .Z(n8470) );
  XNOR U8567 ( .A(n8467), .B(n8573), .Z(n8575) );
  XOR U8568 ( .A(n8579), .B(n8580), .Z(n8467) );
  AND U8569 ( .A(n203), .B(n8581), .Z(n8580) );
  XOR U8570 ( .A(n8582), .B(n8579), .Z(n8581) );
  XOR U8571 ( .A(n8583), .B(n8584), .Z(n8573) );
  AND U8572 ( .A(n8585), .B(n8586), .Z(n8584) );
  XNOR U8573 ( .A(n8583), .B(n8577), .Z(n8586) );
  IV U8574 ( .A(n8485), .Z(n8577) );
  XOR U8575 ( .A(n8587), .B(n8588), .Z(n8485) );
  XOR U8576 ( .A(n8589), .B(n8578), .Z(n8588) );
  AND U8577 ( .A(n8512), .B(n8590), .Z(n8578) );
  AND U8578 ( .A(n8591), .B(n8592), .Z(n8589) );
  XOR U8579 ( .A(n8593), .B(n8587), .Z(n8591) );
  XNOR U8580 ( .A(n8482), .B(n8583), .Z(n8585) );
  XOR U8581 ( .A(n8594), .B(n8595), .Z(n8482) );
  AND U8582 ( .A(n203), .B(n8596), .Z(n8595) );
  XOR U8583 ( .A(n8597), .B(n8594), .Z(n8596) );
  XOR U8584 ( .A(n8598), .B(n8599), .Z(n8583) );
  AND U8585 ( .A(n8600), .B(n8601), .Z(n8599) );
  XNOR U8586 ( .A(n8598), .B(n8512), .Z(n8601) );
  XOR U8587 ( .A(n8602), .B(n8592), .Z(n8512) );
  XNOR U8588 ( .A(n8603), .B(n8587), .Z(n8592) );
  XOR U8589 ( .A(n8604), .B(n8605), .Z(n8587) );
  AND U8590 ( .A(n8606), .B(n8607), .Z(n8605) );
  XOR U8591 ( .A(n8608), .B(n8604), .Z(n8606) );
  XNOR U8592 ( .A(n8609), .B(n8610), .Z(n8603) );
  AND U8593 ( .A(n8611), .B(n8612), .Z(n8610) );
  XOR U8594 ( .A(n8609), .B(n8613), .Z(n8611) );
  XNOR U8595 ( .A(n8593), .B(n8590), .Z(n8602) );
  AND U8596 ( .A(n8614), .B(n8615), .Z(n8590) );
  XOR U8597 ( .A(n8616), .B(n8617), .Z(n8593) );
  AND U8598 ( .A(n8618), .B(n8619), .Z(n8617) );
  XOR U8599 ( .A(n8616), .B(n8620), .Z(n8618) );
  XNOR U8600 ( .A(n8509), .B(n8598), .Z(n8600) );
  XOR U8601 ( .A(n8621), .B(n8622), .Z(n8509) );
  AND U8602 ( .A(n203), .B(n8623), .Z(n8622) );
  XNOR U8603 ( .A(n8624), .B(n8621), .Z(n8623) );
  XOR U8604 ( .A(n8625), .B(n8626), .Z(n8598) );
  AND U8605 ( .A(n8627), .B(n8628), .Z(n8626) );
  XNOR U8606 ( .A(n8625), .B(n8614), .Z(n8628) );
  IV U8607 ( .A(n8560), .Z(n8614) );
  XNOR U8608 ( .A(n8629), .B(n8607), .Z(n8560) );
  XNOR U8609 ( .A(n8630), .B(n8613), .Z(n8607) );
  XOR U8610 ( .A(n8631), .B(n8632), .Z(n8613) );
  NOR U8611 ( .A(n8633), .B(n8634), .Z(n8632) );
  XNOR U8612 ( .A(n8631), .B(n8635), .Z(n8633) );
  XNOR U8613 ( .A(n8612), .B(n8604), .Z(n8630) );
  XOR U8614 ( .A(n8636), .B(n8637), .Z(n8604) );
  AND U8615 ( .A(n8638), .B(n8639), .Z(n8637) );
  XNOR U8616 ( .A(n8636), .B(n8640), .Z(n8638) );
  XNOR U8617 ( .A(n8641), .B(n8609), .Z(n8612) );
  XOR U8618 ( .A(n8642), .B(n8643), .Z(n8609) );
  AND U8619 ( .A(n8644), .B(n8645), .Z(n8643) );
  XOR U8620 ( .A(n8642), .B(n8646), .Z(n8644) );
  XNOR U8621 ( .A(n8647), .B(n8648), .Z(n8641) );
  NOR U8622 ( .A(n8649), .B(n8650), .Z(n8648) );
  XOR U8623 ( .A(n8647), .B(n8651), .Z(n8649) );
  XNOR U8624 ( .A(n8608), .B(n8615), .Z(n8629) );
  NOR U8625 ( .A(n8572), .B(n8652), .Z(n8615) );
  XOR U8626 ( .A(n8620), .B(n8619), .Z(n8608) );
  XNOR U8627 ( .A(n8653), .B(n8616), .Z(n8619) );
  XOR U8628 ( .A(n8654), .B(n8655), .Z(n8616) );
  AND U8629 ( .A(n8656), .B(n8657), .Z(n8655) );
  XOR U8630 ( .A(n8654), .B(n8658), .Z(n8656) );
  XNOR U8631 ( .A(n8659), .B(n8660), .Z(n8653) );
  NOR U8632 ( .A(n8661), .B(n8662), .Z(n8660) );
  XNOR U8633 ( .A(n8659), .B(n8663), .Z(n8661) );
  XOR U8634 ( .A(n8664), .B(n8665), .Z(n8620) );
  NOR U8635 ( .A(n8666), .B(n8667), .Z(n8665) );
  XNOR U8636 ( .A(n8664), .B(n8668), .Z(n8666) );
  XNOR U8637 ( .A(n8557), .B(n8625), .Z(n8627) );
  XOR U8638 ( .A(n8669), .B(n8670), .Z(n8557) );
  AND U8639 ( .A(n203), .B(n8671), .Z(n8670) );
  XOR U8640 ( .A(n8672), .B(n8669), .Z(n8671) );
  AND U8641 ( .A(n8569), .B(n8572), .Z(n8625) );
  XOR U8642 ( .A(n8673), .B(n8652), .Z(n8572) );
  XNOR U8643 ( .A(p_input[1024]), .B(p_input[784]), .Z(n8652) );
  XOR U8644 ( .A(n8640), .B(n8639), .Z(n8673) );
  XNOR U8645 ( .A(n8674), .B(n8646), .Z(n8639) );
  XNOR U8646 ( .A(n8635), .B(n8634), .Z(n8646) );
  XOR U8647 ( .A(n8675), .B(n8631), .Z(n8634) );
  XOR U8648 ( .A(p_input[1034]), .B(p_input[794]), .Z(n8631) );
  XNOR U8649 ( .A(p_input[1035]), .B(p_input[795]), .Z(n8675) );
  XOR U8650 ( .A(p_input[1036]), .B(p_input[796]), .Z(n8635) );
  XNOR U8651 ( .A(n8645), .B(n8636), .Z(n8674) );
  XNOR U8652 ( .A(n3298), .B(p_input[785]), .Z(n8636) );
  XOR U8653 ( .A(n8676), .B(n8651), .Z(n8645) );
  XNOR U8654 ( .A(p_input[1039]), .B(p_input[799]), .Z(n8651) );
  XOR U8655 ( .A(n8642), .B(n8650), .Z(n8676) );
  XOR U8656 ( .A(n8677), .B(n8647), .Z(n8650) );
  XOR U8657 ( .A(p_input[1037]), .B(p_input[797]), .Z(n8647) );
  XNOR U8658 ( .A(p_input[1038]), .B(p_input[798]), .Z(n8677) );
  XOR U8659 ( .A(p_input[1033]), .B(p_input[793]), .Z(n8642) );
  XNOR U8660 ( .A(n8658), .B(n8657), .Z(n8640) );
  XNOR U8661 ( .A(n8678), .B(n8663), .Z(n8657) );
  XOR U8662 ( .A(p_input[1032]), .B(p_input[792]), .Z(n8663) );
  XOR U8663 ( .A(n8654), .B(n8662), .Z(n8678) );
  XOR U8664 ( .A(n8679), .B(n8659), .Z(n8662) );
  XOR U8665 ( .A(p_input[1030]), .B(p_input[790]), .Z(n8659) );
  XNOR U8666 ( .A(p_input[1031]), .B(p_input[791]), .Z(n8679) );
  XOR U8667 ( .A(p_input[1026]), .B(p_input[786]), .Z(n8654) );
  XNOR U8668 ( .A(n8668), .B(n8667), .Z(n8658) );
  XOR U8669 ( .A(n8680), .B(n8664), .Z(n8667) );
  XOR U8670 ( .A(p_input[1027]), .B(p_input[787]), .Z(n8664) );
  XNOR U8671 ( .A(p_input[1028]), .B(p_input[788]), .Z(n8680) );
  XOR U8672 ( .A(p_input[1029]), .B(p_input[789]), .Z(n8668) );
  XOR U8673 ( .A(n8681), .B(n8682), .Z(n8569) );
  AND U8674 ( .A(n203), .B(n8683), .Z(n8682) );
  XNOR U8675 ( .A(n8684), .B(n8681), .Z(n8683) );
  XNOR U8676 ( .A(n8685), .B(n8686), .Z(n203) );
  AND U8677 ( .A(n8687), .B(n8688), .Z(n8686) );
  XOR U8678 ( .A(n8582), .B(n8685), .Z(n8688) );
  AND U8679 ( .A(n8689), .B(n8690), .Z(n8582) );
  XNOR U8680 ( .A(n8579), .B(n8685), .Z(n8687) );
  XOR U8681 ( .A(n8691), .B(n8692), .Z(n8579) );
  AND U8682 ( .A(n207), .B(n8693), .Z(n8692) );
  XOR U8683 ( .A(n8694), .B(n8691), .Z(n8693) );
  XOR U8684 ( .A(n8695), .B(n8696), .Z(n8685) );
  AND U8685 ( .A(n8697), .B(n8698), .Z(n8696) );
  XNOR U8686 ( .A(n8695), .B(n8689), .Z(n8698) );
  IV U8687 ( .A(n8597), .Z(n8689) );
  XOR U8688 ( .A(n8699), .B(n8700), .Z(n8597) );
  XOR U8689 ( .A(n8701), .B(n8690), .Z(n8700) );
  AND U8690 ( .A(n8624), .B(n8702), .Z(n8690) );
  AND U8691 ( .A(n8703), .B(n8704), .Z(n8701) );
  XOR U8692 ( .A(n8705), .B(n8699), .Z(n8703) );
  XNOR U8693 ( .A(n8594), .B(n8695), .Z(n8697) );
  XOR U8694 ( .A(n8706), .B(n8707), .Z(n8594) );
  AND U8695 ( .A(n207), .B(n8708), .Z(n8707) );
  XOR U8696 ( .A(n8709), .B(n8706), .Z(n8708) );
  XOR U8697 ( .A(n8710), .B(n8711), .Z(n8695) );
  AND U8698 ( .A(n8712), .B(n8713), .Z(n8711) );
  XNOR U8699 ( .A(n8710), .B(n8624), .Z(n8713) );
  XOR U8700 ( .A(n8714), .B(n8704), .Z(n8624) );
  XNOR U8701 ( .A(n8715), .B(n8699), .Z(n8704) );
  XOR U8702 ( .A(n8716), .B(n8717), .Z(n8699) );
  AND U8703 ( .A(n8718), .B(n8719), .Z(n8717) );
  XOR U8704 ( .A(n8720), .B(n8716), .Z(n8718) );
  XNOR U8705 ( .A(n8721), .B(n8722), .Z(n8715) );
  AND U8706 ( .A(n8723), .B(n8724), .Z(n8722) );
  XOR U8707 ( .A(n8721), .B(n8725), .Z(n8723) );
  XNOR U8708 ( .A(n8705), .B(n8702), .Z(n8714) );
  AND U8709 ( .A(n8726), .B(n8727), .Z(n8702) );
  XOR U8710 ( .A(n8728), .B(n8729), .Z(n8705) );
  AND U8711 ( .A(n8730), .B(n8731), .Z(n8729) );
  XOR U8712 ( .A(n8728), .B(n8732), .Z(n8730) );
  XNOR U8713 ( .A(n8621), .B(n8710), .Z(n8712) );
  XOR U8714 ( .A(n8733), .B(n8734), .Z(n8621) );
  AND U8715 ( .A(n207), .B(n8735), .Z(n8734) );
  XNOR U8716 ( .A(n8736), .B(n8733), .Z(n8735) );
  XOR U8717 ( .A(n8737), .B(n8738), .Z(n8710) );
  AND U8718 ( .A(n8739), .B(n8740), .Z(n8738) );
  XNOR U8719 ( .A(n8737), .B(n8726), .Z(n8740) );
  IV U8720 ( .A(n8672), .Z(n8726) );
  XNOR U8721 ( .A(n8741), .B(n8719), .Z(n8672) );
  XNOR U8722 ( .A(n8742), .B(n8725), .Z(n8719) );
  XOR U8723 ( .A(n8743), .B(n8744), .Z(n8725) );
  NOR U8724 ( .A(n8745), .B(n8746), .Z(n8744) );
  XNOR U8725 ( .A(n8743), .B(n8747), .Z(n8745) );
  XNOR U8726 ( .A(n8724), .B(n8716), .Z(n8742) );
  XOR U8727 ( .A(n8748), .B(n8749), .Z(n8716) );
  AND U8728 ( .A(n8750), .B(n8751), .Z(n8749) );
  XNOR U8729 ( .A(n8748), .B(n8752), .Z(n8750) );
  XNOR U8730 ( .A(n8753), .B(n8721), .Z(n8724) );
  XOR U8731 ( .A(n8754), .B(n8755), .Z(n8721) );
  AND U8732 ( .A(n8756), .B(n8757), .Z(n8755) );
  XOR U8733 ( .A(n8754), .B(n8758), .Z(n8756) );
  XNOR U8734 ( .A(n8759), .B(n8760), .Z(n8753) );
  NOR U8735 ( .A(n8761), .B(n8762), .Z(n8760) );
  XOR U8736 ( .A(n8759), .B(n8763), .Z(n8761) );
  XNOR U8737 ( .A(n8720), .B(n8727), .Z(n8741) );
  NOR U8738 ( .A(n8684), .B(n8764), .Z(n8727) );
  XOR U8739 ( .A(n8732), .B(n8731), .Z(n8720) );
  XNOR U8740 ( .A(n8765), .B(n8728), .Z(n8731) );
  XOR U8741 ( .A(n8766), .B(n8767), .Z(n8728) );
  AND U8742 ( .A(n8768), .B(n8769), .Z(n8767) );
  XOR U8743 ( .A(n8766), .B(n8770), .Z(n8768) );
  XNOR U8744 ( .A(n8771), .B(n8772), .Z(n8765) );
  NOR U8745 ( .A(n8773), .B(n8774), .Z(n8772) );
  XNOR U8746 ( .A(n8771), .B(n8775), .Z(n8773) );
  XOR U8747 ( .A(n8776), .B(n8777), .Z(n8732) );
  NOR U8748 ( .A(n8778), .B(n8779), .Z(n8777) );
  XNOR U8749 ( .A(n8776), .B(n8780), .Z(n8778) );
  XNOR U8750 ( .A(n8669), .B(n8737), .Z(n8739) );
  XOR U8751 ( .A(n8781), .B(n8782), .Z(n8669) );
  AND U8752 ( .A(n207), .B(n8783), .Z(n8782) );
  XOR U8753 ( .A(n8784), .B(n8781), .Z(n8783) );
  AND U8754 ( .A(n8681), .B(n8684), .Z(n8737) );
  XOR U8755 ( .A(n8785), .B(n8764), .Z(n8684) );
  XNOR U8756 ( .A(p_input[1024]), .B(p_input[800]), .Z(n8764) );
  XOR U8757 ( .A(n8752), .B(n8751), .Z(n8785) );
  XNOR U8758 ( .A(n8786), .B(n8758), .Z(n8751) );
  XNOR U8759 ( .A(n8747), .B(n8746), .Z(n8758) );
  XOR U8760 ( .A(n8787), .B(n8743), .Z(n8746) );
  XOR U8761 ( .A(p_input[1034]), .B(p_input[810]), .Z(n8743) );
  XNOR U8762 ( .A(p_input[1035]), .B(p_input[811]), .Z(n8787) );
  XOR U8763 ( .A(p_input[1036]), .B(p_input[812]), .Z(n8747) );
  XNOR U8764 ( .A(n8757), .B(n8748), .Z(n8786) );
  XNOR U8765 ( .A(n3298), .B(p_input[801]), .Z(n8748) );
  XOR U8766 ( .A(n8788), .B(n8763), .Z(n8757) );
  XNOR U8767 ( .A(p_input[1039]), .B(p_input[815]), .Z(n8763) );
  XOR U8768 ( .A(n8754), .B(n8762), .Z(n8788) );
  XOR U8769 ( .A(n8789), .B(n8759), .Z(n8762) );
  XOR U8770 ( .A(p_input[1037]), .B(p_input[813]), .Z(n8759) );
  XNOR U8771 ( .A(p_input[1038]), .B(p_input[814]), .Z(n8789) );
  XOR U8772 ( .A(p_input[1033]), .B(p_input[809]), .Z(n8754) );
  XNOR U8773 ( .A(n8770), .B(n8769), .Z(n8752) );
  XNOR U8774 ( .A(n8790), .B(n8775), .Z(n8769) );
  XOR U8775 ( .A(p_input[1032]), .B(p_input[808]), .Z(n8775) );
  XOR U8776 ( .A(n8766), .B(n8774), .Z(n8790) );
  XOR U8777 ( .A(n8791), .B(n8771), .Z(n8774) );
  XOR U8778 ( .A(p_input[1030]), .B(p_input[806]), .Z(n8771) );
  XNOR U8779 ( .A(p_input[1031]), .B(p_input[807]), .Z(n8791) );
  XOR U8780 ( .A(p_input[1026]), .B(p_input[802]), .Z(n8766) );
  XNOR U8781 ( .A(n8780), .B(n8779), .Z(n8770) );
  XOR U8782 ( .A(n8792), .B(n8776), .Z(n8779) );
  XOR U8783 ( .A(p_input[1027]), .B(p_input[803]), .Z(n8776) );
  XNOR U8784 ( .A(p_input[1028]), .B(p_input[804]), .Z(n8792) );
  XOR U8785 ( .A(p_input[1029]), .B(p_input[805]), .Z(n8780) );
  XOR U8786 ( .A(n8793), .B(n8794), .Z(n8681) );
  AND U8787 ( .A(n207), .B(n8795), .Z(n8794) );
  XNOR U8788 ( .A(n8796), .B(n8793), .Z(n8795) );
  XNOR U8789 ( .A(n8797), .B(n8798), .Z(n207) );
  AND U8790 ( .A(n8799), .B(n8800), .Z(n8798) );
  XOR U8791 ( .A(n8694), .B(n8797), .Z(n8800) );
  AND U8792 ( .A(n8801), .B(n8802), .Z(n8694) );
  XNOR U8793 ( .A(n8691), .B(n8797), .Z(n8799) );
  XOR U8794 ( .A(n8803), .B(n8804), .Z(n8691) );
  AND U8795 ( .A(n211), .B(n8805), .Z(n8804) );
  XOR U8796 ( .A(n8806), .B(n8803), .Z(n8805) );
  XOR U8797 ( .A(n8807), .B(n8808), .Z(n8797) );
  AND U8798 ( .A(n8809), .B(n8810), .Z(n8808) );
  XNOR U8799 ( .A(n8807), .B(n8801), .Z(n8810) );
  IV U8800 ( .A(n8709), .Z(n8801) );
  XOR U8801 ( .A(n8811), .B(n8812), .Z(n8709) );
  XOR U8802 ( .A(n8813), .B(n8802), .Z(n8812) );
  AND U8803 ( .A(n8736), .B(n8814), .Z(n8802) );
  AND U8804 ( .A(n8815), .B(n8816), .Z(n8813) );
  XOR U8805 ( .A(n8817), .B(n8811), .Z(n8815) );
  XNOR U8806 ( .A(n8706), .B(n8807), .Z(n8809) );
  XOR U8807 ( .A(n8818), .B(n8819), .Z(n8706) );
  AND U8808 ( .A(n211), .B(n8820), .Z(n8819) );
  XOR U8809 ( .A(n8821), .B(n8818), .Z(n8820) );
  XOR U8810 ( .A(n8822), .B(n8823), .Z(n8807) );
  AND U8811 ( .A(n8824), .B(n8825), .Z(n8823) );
  XNOR U8812 ( .A(n8822), .B(n8736), .Z(n8825) );
  XOR U8813 ( .A(n8826), .B(n8816), .Z(n8736) );
  XNOR U8814 ( .A(n8827), .B(n8811), .Z(n8816) );
  XOR U8815 ( .A(n8828), .B(n8829), .Z(n8811) );
  AND U8816 ( .A(n8830), .B(n8831), .Z(n8829) );
  XOR U8817 ( .A(n8832), .B(n8828), .Z(n8830) );
  XNOR U8818 ( .A(n8833), .B(n8834), .Z(n8827) );
  AND U8819 ( .A(n8835), .B(n8836), .Z(n8834) );
  XOR U8820 ( .A(n8833), .B(n8837), .Z(n8835) );
  XNOR U8821 ( .A(n8817), .B(n8814), .Z(n8826) );
  AND U8822 ( .A(n8838), .B(n8839), .Z(n8814) );
  XOR U8823 ( .A(n8840), .B(n8841), .Z(n8817) );
  AND U8824 ( .A(n8842), .B(n8843), .Z(n8841) );
  XOR U8825 ( .A(n8840), .B(n8844), .Z(n8842) );
  XNOR U8826 ( .A(n8733), .B(n8822), .Z(n8824) );
  XOR U8827 ( .A(n8845), .B(n8846), .Z(n8733) );
  AND U8828 ( .A(n211), .B(n8847), .Z(n8846) );
  XNOR U8829 ( .A(n8848), .B(n8845), .Z(n8847) );
  XOR U8830 ( .A(n8849), .B(n8850), .Z(n8822) );
  AND U8831 ( .A(n8851), .B(n8852), .Z(n8850) );
  XNOR U8832 ( .A(n8849), .B(n8838), .Z(n8852) );
  IV U8833 ( .A(n8784), .Z(n8838) );
  XNOR U8834 ( .A(n8853), .B(n8831), .Z(n8784) );
  XNOR U8835 ( .A(n8854), .B(n8837), .Z(n8831) );
  XOR U8836 ( .A(n8855), .B(n8856), .Z(n8837) );
  NOR U8837 ( .A(n8857), .B(n8858), .Z(n8856) );
  XNOR U8838 ( .A(n8855), .B(n8859), .Z(n8857) );
  XNOR U8839 ( .A(n8836), .B(n8828), .Z(n8854) );
  XOR U8840 ( .A(n8860), .B(n8861), .Z(n8828) );
  AND U8841 ( .A(n8862), .B(n8863), .Z(n8861) );
  XNOR U8842 ( .A(n8860), .B(n8864), .Z(n8862) );
  XNOR U8843 ( .A(n8865), .B(n8833), .Z(n8836) );
  XOR U8844 ( .A(n8866), .B(n8867), .Z(n8833) );
  AND U8845 ( .A(n8868), .B(n8869), .Z(n8867) );
  XOR U8846 ( .A(n8866), .B(n8870), .Z(n8868) );
  XNOR U8847 ( .A(n8871), .B(n8872), .Z(n8865) );
  NOR U8848 ( .A(n8873), .B(n8874), .Z(n8872) );
  XOR U8849 ( .A(n8871), .B(n8875), .Z(n8873) );
  XNOR U8850 ( .A(n8832), .B(n8839), .Z(n8853) );
  NOR U8851 ( .A(n8796), .B(n8876), .Z(n8839) );
  XOR U8852 ( .A(n8844), .B(n8843), .Z(n8832) );
  XNOR U8853 ( .A(n8877), .B(n8840), .Z(n8843) );
  XOR U8854 ( .A(n8878), .B(n8879), .Z(n8840) );
  AND U8855 ( .A(n8880), .B(n8881), .Z(n8879) );
  XOR U8856 ( .A(n8878), .B(n8882), .Z(n8880) );
  XNOR U8857 ( .A(n8883), .B(n8884), .Z(n8877) );
  NOR U8858 ( .A(n8885), .B(n8886), .Z(n8884) );
  XNOR U8859 ( .A(n8883), .B(n8887), .Z(n8885) );
  XOR U8860 ( .A(n8888), .B(n8889), .Z(n8844) );
  NOR U8861 ( .A(n8890), .B(n8891), .Z(n8889) );
  XNOR U8862 ( .A(n8888), .B(n8892), .Z(n8890) );
  XNOR U8863 ( .A(n8781), .B(n8849), .Z(n8851) );
  XOR U8864 ( .A(n8893), .B(n8894), .Z(n8781) );
  AND U8865 ( .A(n211), .B(n8895), .Z(n8894) );
  XOR U8866 ( .A(n8896), .B(n8893), .Z(n8895) );
  AND U8867 ( .A(n8793), .B(n8796), .Z(n8849) );
  XOR U8868 ( .A(n8897), .B(n8876), .Z(n8796) );
  XNOR U8869 ( .A(p_input[1024]), .B(p_input[816]), .Z(n8876) );
  XOR U8870 ( .A(n8864), .B(n8863), .Z(n8897) );
  XNOR U8871 ( .A(n8898), .B(n8870), .Z(n8863) );
  XNOR U8872 ( .A(n8859), .B(n8858), .Z(n8870) );
  XOR U8873 ( .A(n8899), .B(n8855), .Z(n8858) );
  XOR U8874 ( .A(p_input[1034]), .B(p_input[826]), .Z(n8855) );
  XNOR U8875 ( .A(p_input[1035]), .B(p_input[827]), .Z(n8899) );
  XOR U8876 ( .A(p_input[1036]), .B(p_input[828]), .Z(n8859) );
  XNOR U8877 ( .A(n8869), .B(n8860), .Z(n8898) );
  XNOR U8878 ( .A(n3298), .B(p_input[817]), .Z(n8860) );
  XOR U8879 ( .A(n8900), .B(n8875), .Z(n8869) );
  XNOR U8880 ( .A(p_input[1039]), .B(p_input[831]), .Z(n8875) );
  XOR U8881 ( .A(n8866), .B(n8874), .Z(n8900) );
  XOR U8882 ( .A(n8901), .B(n8871), .Z(n8874) );
  XOR U8883 ( .A(p_input[1037]), .B(p_input[829]), .Z(n8871) );
  XNOR U8884 ( .A(p_input[1038]), .B(p_input[830]), .Z(n8901) );
  XOR U8885 ( .A(p_input[1033]), .B(p_input[825]), .Z(n8866) );
  XNOR U8886 ( .A(n8882), .B(n8881), .Z(n8864) );
  XNOR U8887 ( .A(n8902), .B(n8887), .Z(n8881) );
  XOR U8888 ( .A(p_input[1032]), .B(p_input[824]), .Z(n8887) );
  XOR U8889 ( .A(n8878), .B(n8886), .Z(n8902) );
  XOR U8890 ( .A(n8903), .B(n8883), .Z(n8886) );
  XOR U8891 ( .A(p_input[1030]), .B(p_input[822]), .Z(n8883) );
  XNOR U8892 ( .A(p_input[1031]), .B(p_input[823]), .Z(n8903) );
  XOR U8893 ( .A(p_input[1026]), .B(p_input[818]), .Z(n8878) );
  XNOR U8894 ( .A(n8892), .B(n8891), .Z(n8882) );
  XOR U8895 ( .A(n8904), .B(n8888), .Z(n8891) );
  XOR U8896 ( .A(p_input[1027]), .B(p_input[819]), .Z(n8888) );
  XNOR U8897 ( .A(p_input[1028]), .B(p_input[820]), .Z(n8904) );
  XOR U8898 ( .A(p_input[1029]), .B(p_input[821]), .Z(n8892) );
  XOR U8899 ( .A(n8905), .B(n8906), .Z(n8793) );
  AND U8900 ( .A(n211), .B(n8907), .Z(n8906) );
  XNOR U8901 ( .A(n8908), .B(n8905), .Z(n8907) );
  XNOR U8902 ( .A(n8909), .B(n8910), .Z(n211) );
  AND U8903 ( .A(n8911), .B(n8912), .Z(n8910) );
  XOR U8904 ( .A(n8806), .B(n8909), .Z(n8912) );
  AND U8905 ( .A(n8913), .B(n8914), .Z(n8806) );
  XNOR U8906 ( .A(n8803), .B(n8909), .Z(n8911) );
  XOR U8907 ( .A(n8915), .B(n8916), .Z(n8803) );
  AND U8908 ( .A(n8917), .B(n215), .Z(n8916) );
  AND U8909 ( .A(n8915), .B(n8918), .Z(n8917) );
  XOR U8910 ( .A(n8919), .B(n8920), .Z(n8909) );
  AND U8911 ( .A(n8921), .B(n8922), .Z(n8920) );
  XNOR U8912 ( .A(n8919), .B(n8913), .Z(n8922) );
  IV U8913 ( .A(n8821), .Z(n8913) );
  XOR U8914 ( .A(n8923), .B(n8924), .Z(n8821) );
  XOR U8915 ( .A(n8925), .B(n8914), .Z(n8924) );
  AND U8916 ( .A(n8848), .B(n8926), .Z(n8914) );
  AND U8917 ( .A(n8927), .B(n8928), .Z(n8925) );
  XOR U8918 ( .A(n8929), .B(n8923), .Z(n8927) );
  XNOR U8919 ( .A(n8818), .B(n8919), .Z(n8921) );
  XOR U8920 ( .A(n8930), .B(n8931), .Z(n8818) );
  AND U8921 ( .A(n215), .B(n8932), .Z(n8931) );
  XOR U8922 ( .A(n8933), .B(n8930), .Z(n8932) );
  XOR U8923 ( .A(n8934), .B(n8935), .Z(n8919) );
  AND U8924 ( .A(n8936), .B(n8937), .Z(n8935) );
  XNOR U8925 ( .A(n8934), .B(n8848), .Z(n8937) );
  XOR U8926 ( .A(n8938), .B(n8928), .Z(n8848) );
  XNOR U8927 ( .A(n8939), .B(n8923), .Z(n8928) );
  XOR U8928 ( .A(n8940), .B(n8941), .Z(n8923) );
  AND U8929 ( .A(n8942), .B(n8943), .Z(n8941) );
  XOR U8930 ( .A(n8944), .B(n8940), .Z(n8942) );
  XNOR U8931 ( .A(n8945), .B(n8946), .Z(n8939) );
  AND U8932 ( .A(n8947), .B(n8948), .Z(n8946) );
  XOR U8933 ( .A(n8945), .B(n8949), .Z(n8947) );
  XNOR U8934 ( .A(n8929), .B(n8926), .Z(n8938) );
  AND U8935 ( .A(n8950), .B(n8951), .Z(n8926) );
  XOR U8936 ( .A(n8952), .B(n8953), .Z(n8929) );
  AND U8937 ( .A(n8954), .B(n8955), .Z(n8953) );
  XOR U8938 ( .A(n8952), .B(n8956), .Z(n8954) );
  XNOR U8939 ( .A(n8845), .B(n8934), .Z(n8936) );
  XOR U8940 ( .A(n8957), .B(n8958), .Z(n8845) );
  AND U8941 ( .A(n215), .B(n8959), .Z(n8958) );
  XNOR U8942 ( .A(n8960), .B(n8957), .Z(n8959) );
  XOR U8943 ( .A(n8961), .B(n8962), .Z(n8934) );
  AND U8944 ( .A(n8963), .B(n8964), .Z(n8962) );
  XNOR U8945 ( .A(n8961), .B(n8950), .Z(n8964) );
  IV U8946 ( .A(n8896), .Z(n8950) );
  XNOR U8947 ( .A(n8965), .B(n8943), .Z(n8896) );
  XNOR U8948 ( .A(n8966), .B(n8949), .Z(n8943) );
  XOR U8949 ( .A(n8967), .B(n8968), .Z(n8949) );
  NOR U8950 ( .A(n8969), .B(n8970), .Z(n8968) );
  XNOR U8951 ( .A(n8967), .B(n8971), .Z(n8969) );
  XNOR U8952 ( .A(n8948), .B(n8940), .Z(n8966) );
  XOR U8953 ( .A(n8972), .B(n8973), .Z(n8940) );
  AND U8954 ( .A(n8974), .B(n8975), .Z(n8973) );
  XNOR U8955 ( .A(n8972), .B(n8976), .Z(n8974) );
  XNOR U8956 ( .A(n8977), .B(n8945), .Z(n8948) );
  XOR U8957 ( .A(n8978), .B(n8979), .Z(n8945) );
  AND U8958 ( .A(n8980), .B(n8981), .Z(n8979) );
  XOR U8959 ( .A(n8978), .B(n8982), .Z(n8980) );
  XNOR U8960 ( .A(n8983), .B(n8984), .Z(n8977) );
  NOR U8961 ( .A(n8985), .B(n8986), .Z(n8984) );
  XOR U8962 ( .A(n8983), .B(n8987), .Z(n8985) );
  XNOR U8963 ( .A(n8944), .B(n8951), .Z(n8965) );
  NOR U8964 ( .A(n8908), .B(n8988), .Z(n8951) );
  XOR U8965 ( .A(n8956), .B(n8955), .Z(n8944) );
  XNOR U8966 ( .A(n8989), .B(n8952), .Z(n8955) );
  XOR U8967 ( .A(n8990), .B(n8991), .Z(n8952) );
  AND U8968 ( .A(n8992), .B(n8993), .Z(n8991) );
  XOR U8969 ( .A(n8990), .B(n8994), .Z(n8992) );
  XNOR U8970 ( .A(n8995), .B(n8996), .Z(n8989) );
  NOR U8971 ( .A(n8997), .B(n8998), .Z(n8996) );
  XNOR U8972 ( .A(n8995), .B(n8999), .Z(n8997) );
  XOR U8973 ( .A(n9000), .B(n9001), .Z(n8956) );
  NOR U8974 ( .A(n9002), .B(n9003), .Z(n9001) );
  XNOR U8975 ( .A(n9000), .B(n9004), .Z(n9002) );
  XNOR U8976 ( .A(n8893), .B(n8961), .Z(n8963) );
  XOR U8977 ( .A(n9005), .B(n9006), .Z(n8893) );
  AND U8978 ( .A(n215), .B(n9007), .Z(n9006) );
  XOR U8979 ( .A(n9008), .B(n9005), .Z(n9007) );
  AND U8980 ( .A(n8905), .B(n8908), .Z(n8961) );
  XOR U8981 ( .A(n9009), .B(n8988), .Z(n8908) );
  XNOR U8982 ( .A(p_input[1024]), .B(p_input[832]), .Z(n8988) );
  XOR U8983 ( .A(n8976), .B(n8975), .Z(n9009) );
  XNOR U8984 ( .A(n9010), .B(n8982), .Z(n8975) );
  XNOR U8985 ( .A(n8971), .B(n8970), .Z(n8982) );
  XOR U8986 ( .A(n9011), .B(n8967), .Z(n8970) );
  XOR U8987 ( .A(p_input[1034]), .B(p_input[842]), .Z(n8967) );
  XNOR U8988 ( .A(p_input[1035]), .B(p_input[843]), .Z(n9011) );
  XOR U8989 ( .A(p_input[1036]), .B(p_input[844]), .Z(n8971) );
  XNOR U8990 ( .A(n8981), .B(n8972), .Z(n9010) );
  XNOR U8991 ( .A(n3298), .B(p_input[833]), .Z(n8972) );
  XOR U8992 ( .A(n9012), .B(n8987), .Z(n8981) );
  XNOR U8993 ( .A(p_input[1039]), .B(p_input[847]), .Z(n8987) );
  XOR U8994 ( .A(n8978), .B(n8986), .Z(n9012) );
  XOR U8995 ( .A(n9013), .B(n8983), .Z(n8986) );
  XOR U8996 ( .A(p_input[1037]), .B(p_input[845]), .Z(n8983) );
  XNOR U8997 ( .A(p_input[1038]), .B(p_input[846]), .Z(n9013) );
  XOR U8998 ( .A(p_input[1033]), .B(p_input[841]), .Z(n8978) );
  XNOR U8999 ( .A(n8994), .B(n8993), .Z(n8976) );
  XNOR U9000 ( .A(n9014), .B(n8999), .Z(n8993) );
  XOR U9001 ( .A(p_input[1032]), .B(p_input[840]), .Z(n8999) );
  XOR U9002 ( .A(n8990), .B(n8998), .Z(n9014) );
  XOR U9003 ( .A(n9015), .B(n8995), .Z(n8998) );
  XOR U9004 ( .A(p_input[1030]), .B(p_input[838]), .Z(n8995) );
  XNOR U9005 ( .A(p_input[1031]), .B(p_input[839]), .Z(n9015) );
  XOR U9006 ( .A(p_input[1026]), .B(p_input[834]), .Z(n8990) );
  XNOR U9007 ( .A(n9004), .B(n9003), .Z(n8994) );
  XOR U9008 ( .A(n9016), .B(n9000), .Z(n9003) );
  XOR U9009 ( .A(p_input[1027]), .B(p_input[835]), .Z(n9000) );
  XNOR U9010 ( .A(p_input[1028]), .B(p_input[836]), .Z(n9016) );
  XOR U9011 ( .A(p_input[1029]), .B(p_input[837]), .Z(n9004) );
  XOR U9012 ( .A(n9017), .B(n9018), .Z(n8905) );
  AND U9013 ( .A(n215), .B(n9019), .Z(n9018) );
  XNOR U9014 ( .A(n9020), .B(n9017), .Z(n9019) );
  XNOR U9015 ( .A(n9021), .B(n9022), .Z(n215) );
  AND U9016 ( .A(n9023), .B(n9024), .Z(n9022) );
  XNOR U9017 ( .A(n8918), .B(n9021), .Z(n9024) );
  IV U9018 ( .A(n9025), .Z(n8918) );
  AND U9019 ( .A(n9026), .B(n9027), .Z(n9025) );
  XNOR U9020 ( .A(n9021), .B(n8915), .Z(n9023) );
  AND U9021 ( .A(n9028), .B(n9029), .Z(n8915) );
  XOR U9022 ( .A(n9030), .B(n9031), .Z(n9021) );
  AND U9023 ( .A(n9032), .B(n9033), .Z(n9031) );
  XNOR U9024 ( .A(n9030), .B(n9026), .Z(n9033) );
  IV U9025 ( .A(n8933), .Z(n9026) );
  XOR U9026 ( .A(n9034), .B(n9035), .Z(n8933) );
  XOR U9027 ( .A(n9036), .B(n9027), .Z(n9035) );
  AND U9028 ( .A(n8960), .B(n9037), .Z(n9027) );
  AND U9029 ( .A(n9038), .B(n9039), .Z(n9036) );
  XOR U9030 ( .A(n9040), .B(n9034), .Z(n9038) );
  XNOR U9031 ( .A(n8930), .B(n9030), .Z(n9032) );
  XOR U9032 ( .A(n9041), .B(n9042), .Z(n8930) );
  AND U9033 ( .A(n219), .B(n9043), .Z(n9042) );
  XOR U9034 ( .A(n9044), .B(n9041), .Z(n9043) );
  XOR U9035 ( .A(n9045), .B(n9046), .Z(n9030) );
  AND U9036 ( .A(n9047), .B(n9048), .Z(n9046) );
  XNOR U9037 ( .A(n9045), .B(n8960), .Z(n9048) );
  XOR U9038 ( .A(n9049), .B(n9039), .Z(n8960) );
  XNOR U9039 ( .A(n9050), .B(n9034), .Z(n9039) );
  XOR U9040 ( .A(n9051), .B(n9052), .Z(n9034) );
  AND U9041 ( .A(n9053), .B(n9054), .Z(n9052) );
  XOR U9042 ( .A(n9055), .B(n9051), .Z(n9053) );
  XNOR U9043 ( .A(n9056), .B(n9057), .Z(n9050) );
  AND U9044 ( .A(n9058), .B(n9059), .Z(n9057) );
  XOR U9045 ( .A(n9056), .B(n9060), .Z(n9058) );
  XNOR U9046 ( .A(n9040), .B(n9037), .Z(n9049) );
  AND U9047 ( .A(n9061), .B(n9062), .Z(n9037) );
  XOR U9048 ( .A(n9063), .B(n9064), .Z(n9040) );
  AND U9049 ( .A(n9065), .B(n9066), .Z(n9064) );
  XOR U9050 ( .A(n9063), .B(n9067), .Z(n9065) );
  XNOR U9051 ( .A(n8957), .B(n9045), .Z(n9047) );
  XOR U9052 ( .A(n9068), .B(n9069), .Z(n8957) );
  AND U9053 ( .A(n219), .B(n9070), .Z(n9069) );
  XNOR U9054 ( .A(n9071), .B(n9068), .Z(n9070) );
  XOR U9055 ( .A(n9072), .B(n9073), .Z(n9045) );
  AND U9056 ( .A(n9074), .B(n9075), .Z(n9073) );
  XNOR U9057 ( .A(n9072), .B(n9061), .Z(n9075) );
  IV U9058 ( .A(n9008), .Z(n9061) );
  XNOR U9059 ( .A(n9076), .B(n9054), .Z(n9008) );
  XNOR U9060 ( .A(n9077), .B(n9060), .Z(n9054) );
  XOR U9061 ( .A(n9078), .B(n9079), .Z(n9060) );
  NOR U9062 ( .A(n9080), .B(n9081), .Z(n9079) );
  XNOR U9063 ( .A(n9078), .B(n9082), .Z(n9080) );
  XNOR U9064 ( .A(n9059), .B(n9051), .Z(n9077) );
  XOR U9065 ( .A(n9083), .B(n9084), .Z(n9051) );
  AND U9066 ( .A(n9085), .B(n9086), .Z(n9084) );
  XNOR U9067 ( .A(n9083), .B(n9087), .Z(n9085) );
  XNOR U9068 ( .A(n9088), .B(n9056), .Z(n9059) );
  XOR U9069 ( .A(n9089), .B(n9090), .Z(n9056) );
  AND U9070 ( .A(n9091), .B(n9092), .Z(n9090) );
  XOR U9071 ( .A(n9089), .B(n9093), .Z(n9091) );
  XNOR U9072 ( .A(n9094), .B(n9095), .Z(n9088) );
  NOR U9073 ( .A(n9096), .B(n9097), .Z(n9095) );
  XOR U9074 ( .A(n9094), .B(n9098), .Z(n9096) );
  XNOR U9075 ( .A(n9055), .B(n9062), .Z(n9076) );
  NOR U9076 ( .A(n9020), .B(n9099), .Z(n9062) );
  XOR U9077 ( .A(n9067), .B(n9066), .Z(n9055) );
  XNOR U9078 ( .A(n9100), .B(n9063), .Z(n9066) );
  XOR U9079 ( .A(n9101), .B(n9102), .Z(n9063) );
  AND U9080 ( .A(n9103), .B(n9104), .Z(n9102) );
  XOR U9081 ( .A(n9101), .B(n9105), .Z(n9103) );
  XNOR U9082 ( .A(n9106), .B(n9107), .Z(n9100) );
  NOR U9083 ( .A(n9108), .B(n9109), .Z(n9107) );
  XNOR U9084 ( .A(n9106), .B(n9110), .Z(n9108) );
  XOR U9085 ( .A(n9111), .B(n9112), .Z(n9067) );
  NOR U9086 ( .A(n9113), .B(n9114), .Z(n9112) );
  XNOR U9087 ( .A(n9111), .B(n9115), .Z(n9113) );
  XNOR U9088 ( .A(n9005), .B(n9072), .Z(n9074) );
  XOR U9089 ( .A(n9116), .B(n9117), .Z(n9005) );
  AND U9090 ( .A(n219), .B(n9118), .Z(n9117) );
  XOR U9091 ( .A(n9119), .B(n9116), .Z(n9118) );
  AND U9092 ( .A(n9017), .B(n9020), .Z(n9072) );
  XOR U9093 ( .A(n9120), .B(n9099), .Z(n9020) );
  XNOR U9094 ( .A(p_input[1024]), .B(p_input[848]), .Z(n9099) );
  XOR U9095 ( .A(n9087), .B(n9086), .Z(n9120) );
  XNOR U9096 ( .A(n9121), .B(n9093), .Z(n9086) );
  XNOR U9097 ( .A(n9082), .B(n9081), .Z(n9093) );
  XOR U9098 ( .A(n9122), .B(n9078), .Z(n9081) );
  XOR U9099 ( .A(p_input[1034]), .B(p_input[858]), .Z(n9078) );
  XNOR U9100 ( .A(p_input[1035]), .B(p_input[859]), .Z(n9122) );
  XOR U9101 ( .A(p_input[1036]), .B(p_input[860]), .Z(n9082) );
  XNOR U9102 ( .A(n9092), .B(n9083), .Z(n9121) );
  XNOR U9103 ( .A(n3298), .B(p_input[849]), .Z(n9083) );
  XOR U9104 ( .A(n9123), .B(n9098), .Z(n9092) );
  XNOR U9105 ( .A(p_input[1039]), .B(p_input[863]), .Z(n9098) );
  XOR U9106 ( .A(n9089), .B(n9097), .Z(n9123) );
  XOR U9107 ( .A(n9124), .B(n9094), .Z(n9097) );
  XOR U9108 ( .A(p_input[1037]), .B(p_input[861]), .Z(n9094) );
  XNOR U9109 ( .A(p_input[1038]), .B(p_input[862]), .Z(n9124) );
  XOR U9110 ( .A(p_input[1033]), .B(p_input[857]), .Z(n9089) );
  XNOR U9111 ( .A(n9105), .B(n9104), .Z(n9087) );
  XNOR U9112 ( .A(n9125), .B(n9110), .Z(n9104) );
  XOR U9113 ( .A(p_input[1032]), .B(p_input[856]), .Z(n9110) );
  XOR U9114 ( .A(n9101), .B(n9109), .Z(n9125) );
  XOR U9115 ( .A(n9126), .B(n9106), .Z(n9109) );
  XOR U9116 ( .A(p_input[1030]), .B(p_input[854]), .Z(n9106) );
  XNOR U9117 ( .A(p_input[1031]), .B(p_input[855]), .Z(n9126) );
  XOR U9118 ( .A(p_input[1026]), .B(p_input[850]), .Z(n9101) );
  XNOR U9119 ( .A(n9115), .B(n9114), .Z(n9105) );
  XOR U9120 ( .A(n9127), .B(n9111), .Z(n9114) );
  XOR U9121 ( .A(p_input[1027]), .B(p_input[851]), .Z(n9111) );
  XNOR U9122 ( .A(p_input[1028]), .B(p_input[852]), .Z(n9127) );
  XOR U9123 ( .A(p_input[1029]), .B(p_input[853]), .Z(n9115) );
  XOR U9124 ( .A(n9128), .B(n9129), .Z(n9017) );
  AND U9125 ( .A(n219), .B(n9130), .Z(n9129) );
  XNOR U9126 ( .A(n9131), .B(n9128), .Z(n9130) );
  XNOR U9127 ( .A(n9132), .B(n9133), .Z(n219) );
  NOR U9128 ( .A(n9134), .B(n9135), .Z(n9133) );
  XOR U9129 ( .A(n9029), .B(n9132), .Z(n9135) );
  AND U9130 ( .A(n9136), .B(n9137), .Z(n9029) );
  NOR U9131 ( .A(n9132), .B(n9028), .Z(n9134) );
  AND U9132 ( .A(n9138), .B(n9139), .Z(n9028) );
  XOR U9133 ( .A(n9140), .B(n9141), .Z(n9132) );
  AND U9134 ( .A(n9142), .B(n9143), .Z(n9141) );
  XNOR U9135 ( .A(n9140), .B(n9138), .Z(n9143) );
  IV U9136 ( .A(n9044), .Z(n9138) );
  XOR U9137 ( .A(n9144), .B(n9145), .Z(n9044) );
  XOR U9138 ( .A(n9146), .B(n9139), .Z(n9145) );
  AND U9139 ( .A(n9071), .B(n9147), .Z(n9139) );
  AND U9140 ( .A(n9148), .B(n9149), .Z(n9146) );
  XOR U9141 ( .A(n9150), .B(n9144), .Z(n9148) );
  XNOR U9142 ( .A(n9041), .B(n9140), .Z(n9142) );
  XOR U9143 ( .A(n9151), .B(n9152), .Z(n9041) );
  AND U9144 ( .A(n223), .B(n9153), .Z(n9152) );
  XOR U9145 ( .A(n9154), .B(n9151), .Z(n9153) );
  XOR U9146 ( .A(n9155), .B(n9156), .Z(n9140) );
  AND U9147 ( .A(n9157), .B(n9158), .Z(n9156) );
  XNOR U9148 ( .A(n9155), .B(n9071), .Z(n9158) );
  XOR U9149 ( .A(n9159), .B(n9149), .Z(n9071) );
  XNOR U9150 ( .A(n9160), .B(n9144), .Z(n9149) );
  XOR U9151 ( .A(n9161), .B(n9162), .Z(n9144) );
  AND U9152 ( .A(n9163), .B(n9164), .Z(n9162) );
  XOR U9153 ( .A(n9165), .B(n9161), .Z(n9163) );
  XNOR U9154 ( .A(n9166), .B(n9167), .Z(n9160) );
  AND U9155 ( .A(n9168), .B(n9169), .Z(n9167) );
  XOR U9156 ( .A(n9166), .B(n9170), .Z(n9168) );
  XNOR U9157 ( .A(n9150), .B(n9147), .Z(n9159) );
  AND U9158 ( .A(n9171), .B(n9172), .Z(n9147) );
  XOR U9159 ( .A(n9173), .B(n9174), .Z(n9150) );
  AND U9160 ( .A(n9175), .B(n9176), .Z(n9174) );
  XOR U9161 ( .A(n9173), .B(n9177), .Z(n9175) );
  XNOR U9162 ( .A(n9068), .B(n9155), .Z(n9157) );
  XOR U9163 ( .A(n9178), .B(n9179), .Z(n9068) );
  AND U9164 ( .A(n223), .B(n9180), .Z(n9179) );
  XNOR U9165 ( .A(n9181), .B(n9178), .Z(n9180) );
  XOR U9166 ( .A(n9182), .B(n9183), .Z(n9155) );
  AND U9167 ( .A(n9184), .B(n9185), .Z(n9183) );
  XNOR U9168 ( .A(n9182), .B(n9171), .Z(n9185) );
  IV U9169 ( .A(n9119), .Z(n9171) );
  XNOR U9170 ( .A(n9186), .B(n9164), .Z(n9119) );
  XNOR U9171 ( .A(n9187), .B(n9170), .Z(n9164) );
  XOR U9172 ( .A(n9188), .B(n9189), .Z(n9170) );
  NOR U9173 ( .A(n9190), .B(n9191), .Z(n9189) );
  XNOR U9174 ( .A(n9188), .B(n9192), .Z(n9190) );
  XNOR U9175 ( .A(n9169), .B(n9161), .Z(n9187) );
  XOR U9176 ( .A(n9193), .B(n9194), .Z(n9161) );
  AND U9177 ( .A(n9195), .B(n9196), .Z(n9194) );
  XNOR U9178 ( .A(n9193), .B(n9197), .Z(n9195) );
  XNOR U9179 ( .A(n9198), .B(n9166), .Z(n9169) );
  XOR U9180 ( .A(n9199), .B(n9200), .Z(n9166) );
  AND U9181 ( .A(n9201), .B(n9202), .Z(n9200) );
  XOR U9182 ( .A(n9199), .B(n9203), .Z(n9201) );
  XNOR U9183 ( .A(n9204), .B(n9205), .Z(n9198) );
  NOR U9184 ( .A(n9206), .B(n9207), .Z(n9205) );
  XOR U9185 ( .A(n9204), .B(n9208), .Z(n9206) );
  XNOR U9186 ( .A(n9165), .B(n9172), .Z(n9186) );
  NOR U9187 ( .A(n9131), .B(n9209), .Z(n9172) );
  XOR U9188 ( .A(n9177), .B(n9176), .Z(n9165) );
  XNOR U9189 ( .A(n9210), .B(n9173), .Z(n9176) );
  XOR U9190 ( .A(n9211), .B(n9212), .Z(n9173) );
  AND U9191 ( .A(n9213), .B(n9214), .Z(n9212) );
  XOR U9192 ( .A(n9211), .B(n9215), .Z(n9213) );
  XNOR U9193 ( .A(n9216), .B(n9217), .Z(n9210) );
  NOR U9194 ( .A(n9218), .B(n9219), .Z(n9217) );
  XNOR U9195 ( .A(n9216), .B(n9220), .Z(n9218) );
  XOR U9196 ( .A(n9221), .B(n9222), .Z(n9177) );
  NOR U9197 ( .A(n9223), .B(n9224), .Z(n9222) );
  XNOR U9198 ( .A(n9221), .B(n9225), .Z(n9223) );
  XNOR U9199 ( .A(n9116), .B(n9182), .Z(n9184) );
  XOR U9200 ( .A(n9226), .B(n9227), .Z(n9116) );
  AND U9201 ( .A(n223), .B(n9228), .Z(n9227) );
  XOR U9202 ( .A(n9229), .B(n9226), .Z(n9228) );
  AND U9203 ( .A(n9128), .B(n9131), .Z(n9182) );
  XOR U9204 ( .A(n9230), .B(n9209), .Z(n9131) );
  XNOR U9205 ( .A(p_input[1024]), .B(p_input[864]), .Z(n9209) );
  XOR U9206 ( .A(n9197), .B(n9196), .Z(n9230) );
  XNOR U9207 ( .A(n9231), .B(n9203), .Z(n9196) );
  XNOR U9208 ( .A(n9192), .B(n9191), .Z(n9203) );
  XOR U9209 ( .A(n9232), .B(n9188), .Z(n9191) );
  XOR U9210 ( .A(p_input[1034]), .B(p_input[874]), .Z(n9188) );
  XNOR U9211 ( .A(p_input[1035]), .B(p_input[875]), .Z(n9232) );
  XOR U9212 ( .A(p_input[1036]), .B(p_input[876]), .Z(n9192) );
  XNOR U9213 ( .A(n9202), .B(n9193), .Z(n9231) );
  XNOR U9214 ( .A(n3298), .B(p_input[865]), .Z(n9193) );
  XOR U9215 ( .A(n9233), .B(n9208), .Z(n9202) );
  XNOR U9216 ( .A(p_input[1039]), .B(p_input[879]), .Z(n9208) );
  XOR U9217 ( .A(n9199), .B(n9207), .Z(n9233) );
  XOR U9218 ( .A(n9234), .B(n9204), .Z(n9207) );
  XOR U9219 ( .A(p_input[1037]), .B(p_input[877]), .Z(n9204) );
  XNOR U9220 ( .A(p_input[1038]), .B(p_input[878]), .Z(n9234) );
  XOR U9221 ( .A(p_input[1033]), .B(p_input[873]), .Z(n9199) );
  XNOR U9222 ( .A(n9215), .B(n9214), .Z(n9197) );
  XNOR U9223 ( .A(n9235), .B(n9220), .Z(n9214) );
  XOR U9224 ( .A(p_input[1032]), .B(p_input[872]), .Z(n9220) );
  XOR U9225 ( .A(n9211), .B(n9219), .Z(n9235) );
  XOR U9226 ( .A(n9236), .B(n9216), .Z(n9219) );
  XOR U9227 ( .A(p_input[1030]), .B(p_input[870]), .Z(n9216) );
  XNOR U9228 ( .A(p_input[1031]), .B(p_input[871]), .Z(n9236) );
  XOR U9229 ( .A(p_input[1026]), .B(p_input[866]), .Z(n9211) );
  XNOR U9230 ( .A(n9225), .B(n9224), .Z(n9215) );
  XOR U9231 ( .A(n9237), .B(n9221), .Z(n9224) );
  XOR U9232 ( .A(p_input[1027]), .B(p_input[867]), .Z(n9221) );
  XNOR U9233 ( .A(p_input[1028]), .B(p_input[868]), .Z(n9237) );
  XOR U9234 ( .A(p_input[1029]), .B(p_input[869]), .Z(n9225) );
  XOR U9235 ( .A(n9238), .B(n9239), .Z(n9128) );
  AND U9236 ( .A(n223), .B(n9240), .Z(n9239) );
  XNOR U9237 ( .A(n9241), .B(n9238), .Z(n9240) );
  XNOR U9238 ( .A(n9242), .B(n9243), .Z(n223) );
  NOR U9239 ( .A(n9244), .B(n9245), .Z(n9243) );
  XOR U9240 ( .A(n9137), .B(n9242), .Z(n9245) );
  AND U9241 ( .A(n9246), .B(n9247), .Z(n9137) );
  NOR U9242 ( .A(n9242), .B(n9136), .Z(n9244) );
  AND U9243 ( .A(n9248), .B(n9249), .Z(n9136) );
  XOR U9244 ( .A(n9250), .B(n9251), .Z(n9242) );
  AND U9245 ( .A(n9252), .B(n9253), .Z(n9251) );
  XNOR U9246 ( .A(n9250), .B(n9248), .Z(n9253) );
  IV U9247 ( .A(n9154), .Z(n9248) );
  XOR U9248 ( .A(n9254), .B(n9255), .Z(n9154) );
  XOR U9249 ( .A(n9256), .B(n9249), .Z(n9255) );
  AND U9250 ( .A(n9181), .B(n9257), .Z(n9249) );
  AND U9251 ( .A(n9258), .B(n9259), .Z(n9256) );
  XOR U9252 ( .A(n9260), .B(n9254), .Z(n9258) );
  XNOR U9253 ( .A(n9151), .B(n9250), .Z(n9252) );
  XOR U9254 ( .A(n9261), .B(n9262), .Z(n9151) );
  AND U9255 ( .A(n227), .B(n9263), .Z(n9262) );
  XOR U9256 ( .A(n9264), .B(n9261), .Z(n9263) );
  XOR U9257 ( .A(n9265), .B(n9266), .Z(n9250) );
  AND U9258 ( .A(n9267), .B(n9268), .Z(n9266) );
  XNOR U9259 ( .A(n9265), .B(n9181), .Z(n9268) );
  XOR U9260 ( .A(n9269), .B(n9259), .Z(n9181) );
  XNOR U9261 ( .A(n9270), .B(n9254), .Z(n9259) );
  XOR U9262 ( .A(n9271), .B(n9272), .Z(n9254) );
  AND U9263 ( .A(n9273), .B(n9274), .Z(n9272) );
  XOR U9264 ( .A(n9275), .B(n9271), .Z(n9273) );
  XNOR U9265 ( .A(n9276), .B(n9277), .Z(n9270) );
  AND U9266 ( .A(n9278), .B(n9279), .Z(n9277) );
  XOR U9267 ( .A(n9276), .B(n9280), .Z(n9278) );
  XNOR U9268 ( .A(n9260), .B(n9257), .Z(n9269) );
  AND U9269 ( .A(n9281), .B(n9282), .Z(n9257) );
  XOR U9270 ( .A(n9283), .B(n9284), .Z(n9260) );
  AND U9271 ( .A(n9285), .B(n9286), .Z(n9284) );
  XOR U9272 ( .A(n9283), .B(n9287), .Z(n9285) );
  XNOR U9273 ( .A(n9178), .B(n9265), .Z(n9267) );
  XOR U9274 ( .A(n9288), .B(n9289), .Z(n9178) );
  AND U9275 ( .A(n227), .B(n9290), .Z(n9289) );
  XNOR U9276 ( .A(n9291), .B(n9288), .Z(n9290) );
  XOR U9277 ( .A(n9292), .B(n9293), .Z(n9265) );
  AND U9278 ( .A(n9294), .B(n9295), .Z(n9293) );
  XNOR U9279 ( .A(n9292), .B(n9281), .Z(n9295) );
  IV U9280 ( .A(n9229), .Z(n9281) );
  XNOR U9281 ( .A(n9296), .B(n9274), .Z(n9229) );
  XNOR U9282 ( .A(n9297), .B(n9280), .Z(n9274) );
  XOR U9283 ( .A(n9298), .B(n9299), .Z(n9280) );
  NOR U9284 ( .A(n9300), .B(n9301), .Z(n9299) );
  XNOR U9285 ( .A(n9298), .B(n9302), .Z(n9300) );
  XNOR U9286 ( .A(n9279), .B(n9271), .Z(n9297) );
  XOR U9287 ( .A(n9303), .B(n9304), .Z(n9271) );
  AND U9288 ( .A(n9305), .B(n9306), .Z(n9304) );
  XNOR U9289 ( .A(n9303), .B(n9307), .Z(n9305) );
  XNOR U9290 ( .A(n9308), .B(n9276), .Z(n9279) );
  XOR U9291 ( .A(n9309), .B(n9310), .Z(n9276) );
  AND U9292 ( .A(n9311), .B(n9312), .Z(n9310) );
  XOR U9293 ( .A(n9309), .B(n9313), .Z(n9311) );
  XNOR U9294 ( .A(n9314), .B(n9315), .Z(n9308) );
  NOR U9295 ( .A(n9316), .B(n9317), .Z(n9315) );
  XOR U9296 ( .A(n9314), .B(n9318), .Z(n9316) );
  XNOR U9297 ( .A(n9275), .B(n9282), .Z(n9296) );
  NOR U9298 ( .A(n9241), .B(n9319), .Z(n9282) );
  XOR U9299 ( .A(n9287), .B(n9286), .Z(n9275) );
  XNOR U9300 ( .A(n9320), .B(n9283), .Z(n9286) );
  XOR U9301 ( .A(n9321), .B(n9322), .Z(n9283) );
  AND U9302 ( .A(n9323), .B(n9324), .Z(n9322) );
  XOR U9303 ( .A(n9321), .B(n9325), .Z(n9323) );
  XNOR U9304 ( .A(n9326), .B(n9327), .Z(n9320) );
  NOR U9305 ( .A(n9328), .B(n9329), .Z(n9327) );
  XNOR U9306 ( .A(n9326), .B(n9330), .Z(n9328) );
  XOR U9307 ( .A(n9331), .B(n9332), .Z(n9287) );
  NOR U9308 ( .A(n9333), .B(n9334), .Z(n9332) );
  XNOR U9309 ( .A(n9331), .B(n9335), .Z(n9333) );
  XNOR U9310 ( .A(n9226), .B(n9292), .Z(n9294) );
  XOR U9311 ( .A(n9336), .B(n9337), .Z(n9226) );
  AND U9312 ( .A(n227), .B(n9338), .Z(n9337) );
  XOR U9313 ( .A(n9339), .B(n9336), .Z(n9338) );
  AND U9314 ( .A(n9238), .B(n9241), .Z(n9292) );
  XOR U9315 ( .A(n9340), .B(n9319), .Z(n9241) );
  XNOR U9316 ( .A(p_input[1024]), .B(p_input[880]), .Z(n9319) );
  XOR U9317 ( .A(n9307), .B(n9306), .Z(n9340) );
  XNOR U9318 ( .A(n9341), .B(n9313), .Z(n9306) );
  XNOR U9319 ( .A(n9302), .B(n9301), .Z(n9313) );
  XOR U9320 ( .A(n9342), .B(n9298), .Z(n9301) );
  XOR U9321 ( .A(p_input[1034]), .B(p_input[890]), .Z(n9298) );
  XNOR U9322 ( .A(p_input[1035]), .B(p_input[891]), .Z(n9342) );
  XOR U9323 ( .A(p_input[1036]), .B(p_input[892]), .Z(n9302) );
  XNOR U9324 ( .A(n9312), .B(n9303), .Z(n9341) );
  XNOR U9325 ( .A(n3298), .B(p_input[881]), .Z(n9303) );
  XOR U9326 ( .A(n9343), .B(n9318), .Z(n9312) );
  XNOR U9327 ( .A(p_input[1039]), .B(p_input[895]), .Z(n9318) );
  XOR U9328 ( .A(n9309), .B(n9317), .Z(n9343) );
  XOR U9329 ( .A(n9344), .B(n9314), .Z(n9317) );
  XOR U9330 ( .A(p_input[1037]), .B(p_input[893]), .Z(n9314) );
  XNOR U9331 ( .A(p_input[1038]), .B(p_input[894]), .Z(n9344) );
  XOR U9332 ( .A(p_input[1033]), .B(p_input[889]), .Z(n9309) );
  XNOR U9333 ( .A(n9325), .B(n9324), .Z(n9307) );
  XNOR U9334 ( .A(n9345), .B(n9330), .Z(n9324) );
  XOR U9335 ( .A(p_input[1032]), .B(p_input[888]), .Z(n9330) );
  XOR U9336 ( .A(n9321), .B(n9329), .Z(n9345) );
  XOR U9337 ( .A(n9346), .B(n9326), .Z(n9329) );
  XOR U9338 ( .A(p_input[1030]), .B(p_input[886]), .Z(n9326) );
  XNOR U9339 ( .A(p_input[1031]), .B(p_input[887]), .Z(n9346) );
  XOR U9340 ( .A(p_input[1026]), .B(p_input[882]), .Z(n9321) );
  XNOR U9341 ( .A(n9335), .B(n9334), .Z(n9325) );
  XOR U9342 ( .A(n9347), .B(n9331), .Z(n9334) );
  XOR U9343 ( .A(p_input[1027]), .B(p_input[883]), .Z(n9331) );
  XNOR U9344 ( .A(p_input[1028]), .B(p_input[884]), .Z(n9347) );
  XOR U9345 ( .A(p_input[1029]), .B(p_input[885]), .Z(n9335) );
  XOR U9346 ( .A(n9348), .B(n9349), .Z(n9238) );
  AND U9347 ( .A(n227), .B(n9350), .Z(n9349) );
  XNOR U9348 ( .A(n9351), .B(n9348), .Z(n9350) );
  XNOR U9349 ( .A(n9352), .B(n9353), .Z(n227) );
  NOR U9350 ( .A(n9354), .B(n9355), .Z(n9353) );
  XOR U9351 ( .A(n9247), .B(n9352), .Z(n9355) );
  AND U9352 ( .A(n9356), .B(n9357), .Z(n9247) );
  NOR U9353 ( .A(n9352), .B(n9246), .Z(n9354) );
  AND U9354 ( .A(n9358), .B(n9359), .Z(n9246) );
  XOR U9355 ( .A(n9360), .B(n9361), .Z(n9352) );
  AND U9356 ( .A(n9362), .B(n9363), .Z(n9361) );
  XNOR U9357 ( .A(n9360), .B(n9358), .Z(n9363) );
  IV U9358 ( .A(n9264), .Z(n9358) );
  XOR U9359 ( .A(n9364), .B(n9365), .Z(n9264) );
  XOR U9360 ( .A(n9366), .B(n9359), .Z(n9365) );
  AND U9361 ( .A(n9291), .B(n9367), .Z(n9359) );
  AND U9362 ( .A(n9368), .B(n9369), .Z(n9366) );
  XOR U9363 ( .A(n9370), .B(n9364), .Z(n9368) );
  XNOR U9364 ( .A(n9261), .B(n9360), .Z(n9362) );
  XOR U9365 ( .A(n9371), .B(n9372), .Z(n9261) );
  AND U9366 ( .A(n231), .B(n9373), .Z(n9372) );
  XOR U9367 ( .A(n9374), .B(n9371), .Z(n9373) );
  XOR U9368 ( .A(n9375), .B(n9376), .Z(n9360) );
  AND U9369 ( .A(n9377), .B(n9378), .Z(n9376) );
  XNOR U9370 ( .A(n9375), .B(n9291), .Z(n9378) );
  XOR U9371 ( .A(n9379), .B(n9369), .Z(n9291) );
  XNOR U9372 ( .A(n9380), .B(n9364), .Z(n9369) );
  XOR U9373 ( .A(n9381), .B(n9382), .Z(n9364) );
  AND U9374 ( .A(n9383), .B(n9384), .Z(n9382) );
  XOR U9375 ( .A(n9385), .B(n9381), .Z(n9383) );
  XNOR U9376 ( .A(n9386), .B(n9387), .Z(n9380) );
  AND U9377 ( .A(n9388), .B(n9389), .Z(n9387) );
  XOR U9378 ( .A(n9386), .B(n9390), .Z(n9388) );
  XNOR U9379 ( .A(n9370), .B(n9367), .Z(n9379) );
  AND U9380 ( .A(n9391), .B(n9392), .Z(n9367) );
  XOR U9381 ( .A(n9393), .B(n9394), .Z(n9370) );
  AND U9382 ( .A(n9395), .B(n9396), .Z(n9394) );
  XOR U9383 ( .A(n9393), .B(n9397), .Z(n9395) );
  XNOR U9384 ( .A(n9288), .B(n9375), .Z(n9377) );
  XOR U9385 ( .A(n9398), .B(n9399), .Z(n9288) );
  AND U9386 ( .A(n231), .B(n9400), .Z(n9399) );
  XNOR U9387 ( .A(n9401), .B(n9398), .Z(n9400) );
  XOR U9388 ( .A(n9402), .B(n9403), .Z(n9375) );
  AND U9389 ( .A(n9404), .B(n9405), .Z(n9403) );
  XNOR U9390 ( .A(n9402), .B(n9391), .Z(n9405) );
  IV U9391 ( .A(n9339), .Z(n9391) );
  XNOR U9392 ( .A(n9406), .B(n9384), .Z(n9339) );
  XNOR U9393 ( .A(n9407), .B(n9390), .Z(n9384) );
  XOR U9394 ( .A(n9408), .B(n9409), .Z(n9390) );
  NOR U9395 ( .A(n9410), .B(n9411), .Z(n9409) );
  XNOR U9396 ( .A(n9408), .B(n9412), .Z(n9410) );
  XNOR U9397 ( .A(n9389), .B(n9381), .Z(n9407) );
  XOR U9398 ( .A(n9413), .B(n9414), .Z(n9381) );
  AND U9399 ( .A(n9415), .B(n9416), .Z(n9414) );
  XNOR U9400 ( .A(n9413), .B(n9417), .Z(n9415) );
  XNOR U9401 ( .A(n9418), .B(n9386), .Z(n9389) );
  XOR U9402 ( .A(n9419), .B(n9420), .Z(n9386) );
  AND U9403 ( .A(n9421), .B(n9422), .Z(n9420) );
  XOR U9404 ( .A(n9419), .B(n9423), .Z(n9421) );
  XNOR U9405 ( .A(n9424), .B(n9425), .Z(n9418) );
  NOR U9406 ( .A(n9426), .B(n9427), .Z(n9425) );
  XOR U9407 ( .A(n9424), .B(n9428), .Z(n9426) );
  XNOR U9408 ( .A(n9385), .B(n9392), .Z(n9406) );
  NOR U9409 ( .A(n9351), .B(n9429), .Z(n9392) );
  XOR U9410 ( .A(n9397), .B(n9396), .Z(n9385) );
  XNOR U9411 ( .A(n9430), .B(n9393), .Z(n9396) );
  XOR U9412 ( .A(n9431), .B(n9432), .Z(n9393) );
  AND U9413 ( .A(n9433), .B(n9434), .Z(n9432) );
  XOR U9414 ( .A(n9431), .B(n9435), .Z(n9433) );
  XNOR U9415 ( .A(n9436), .B(n9437), .Z(n9430) );
  NOR U9416 ( .A(n9438), .B(n9439), .Z(n9437) );
  XNOR U9417 ( .A(n9436), .B(n9440), .Z(n9438) );
  XOR U9418 ( .A(n9441), .B(n9442), .Z(n9397) );
  NOR U9419 ( .A(n9443), .B(n9444), .Z(n9442) );
  XNOR U9420 ( .A(n9441), .B(n9445), .Z(n9443) );
  XNOR U9421 ( .A(n9336), .B(n9402), .Z(n9404) );
  XOR U9422 ( .A(n9446), .B(n9447), .Z(n9336) );
  AND U9423 ( .A(n231), .B(n9448), .Z(n9447) );
  XOR U9424 ( .A(n9449), .B(n9446), .Z(n9448) );
  AND U9425 ( .A(n9348), .B(n9351), .Z(n9402) );
  XOR U9426 ( .A(n9450), .B(n9429), .Z(n9351) );
  XNOR U9427 ( .A(p_input[1024]), .B(p_input[896]), .Z(n9429) );
  XOR U9428 ( .A(n9417), .B(n9416), .Z(n9450) );
  XNOR U9429 ( .A(n9451), .B(n9423), .Z(n9416) );
  XNOR U9430 ( .A(n9412), .B(n9411), .Z(n9423) );
  XOR U9431 ( .A(n9452), .B(n9408), .Z(n9411) );
  XOR U9432 ( .A(p_input[1034]), .B(p_input[906]), .Z(n9408) );
  XNOR U9433 ( .A(p_input[1035]), .B(p_input[907]), .Z(n9452) );
  XOR U9434 ( .A(p_input[1036]), .B(p_input[908]), .Z(n9412) );
  XNOR U9435 ( .A(n9422), .B(n9413), .Z(n9451) );
  XNOR U9436 ( .A(n3298), .B(p_input[897]), .Z(n9413) );
  XOR U9437 ( .A(n9453), .B(n9428), .Z(n9422) );
  XNOR U9438 ( .A(p_input[1039]), .B(p_input[911]), .Z(n9428) );
  XOR U9439 ( .A(n9419), .B(n9427), .Z(n9453) );
  XOR U9440 ( .A(n9454), .B(n9424), .Z(n9427) );
  XOR U9441 ( .A(p_input[1037]), .B(p_input[909]), .Z(n9424) );
  XNOR U9442 ( .A(p_input[1038]), .B(p_input[910]), .Z(n9454) );
  XOR U9443 ( .A(p_input[1033]), .B(p_input[905]), .Z(n9419) );
  XNOR U9444 ( .A(n9435), .B(n9434), .Z(n9417) );
  XNOR U9445 ( .A(n9455), .B(n9440), .Z(n9434) );
  XOR U9446 ( .A(p_input[1032]), .B(p_input[904]), .Z(n9440) );
  XOR U9447 ( .A(n9431), .B(n9439), .Z(n9455) );
  XOR U9448 ( .A(n9456), .B(n9436), .Z(n9439) );
  XOR U9449 ( .A(p_input[1030]), .B(p_input[902]), .Z(n9436) );
  XNOR U9450 ( .A(p_input[1031]), .B(p_input[903]), .Z(n9456) );
  XOR U9451 ( .A(p_input[1026]), .B(p_input[898]), .Z(n9431) );
  XNOR U9452 ( .A(n9445), .B(n9444), .Z(n9435) );
  XOR U9453 ( .A(n9457), .B(n9441), .Z(n9444) );
  XOR U9454 ( .A(p_input[1027]), .B(p_input[899]), .Z(n9441) );
  XNOR U9455 ( .A(p_input[1028]), .B(p_input[900]), .Z(n9457) );
  XOR U9456 ( .A(p_input[1029]), .B(p_input[901]), .Z(n9445) );
  XOR U9457 ( .A(n9458), .B(n9459), .Z(n9348) );
  AND U9458 ( .A(n231), .B(n9460), .Z(n9459) );
  XNOR U9459 ( .A(n9461), .B(n9458), .Z(n9460) );
  XNOR U9460 ( .A(n9462), .B(n9463), .Z(n231) );
  NOR U9461 ( .A(n9464), .B(n9465), .Z(n9463) );
  XOR U9462 ( .A(n9357), .B(n9462), .Z(n9465) );
  AND U9463 ( .A(n9466), .B(n9467), .Z(n9357) );
  NOR U9464 ( .A(n9462), .B(n9356), .Z(n9464) );
  AND U9465 ( .A(n9468), .B(n9469), .Z(n9356) );
  XOR U9466 ( .A(n9470), .B(n9471), .Z(n9462) );
  AND U9467 ( .A(n9472), .B(n9473), .Z(n9471) );
  XNOR U9468 ( .A(n9470), .B(n9468), .Z(n9473) );
  IV U9469 ( .A(n9374), .Z(n9468) );
  XOR U9470 ( .A(n9474), .B(n9475), .Z(n9374) );
  XOR U9471 ( .A(n9476), .B(n9469), .Z(n9475) );
  AND U9472 ( .A(n9401), .B(n9477), .Z(n9469) );
  AND U9473 ( .A(n9478), .B(n9479), .Z(n9476) );
  XOR U9474 ( .A(n9480), .B(n9474), .Z(n9478) );
  XNOR U9475 ( .A(n9371), .B(n9470), .Z(n9472) );
  XOR U9476 ( .A(n9481), .B(n9482), .Z(n9371) );
  AND U9477 ( .A(n235), .B(n9483), .Z(n9482) );
  XOR U9478 ( .A(n9484), .B(n9481), .Z(n9483) );
  XOR U9479 ( .A(n9485), .B(n9486), .Z(n9470) );
  AND U9480 ( .A(n9487), .B(n9488), .Z(n9486) );
  XNOR U9481 ( .A(n9485), .B(n9401), .Z(n9488) );
  XOR U9482 ( .A(n9489), .B(n9479), .Z(n9401) );
  XNOR U9483 ( .A(n9490), .B(n9474), .Z(n9479) );
  XOR U9484 ( .A(n9491), .B(n9492), .Z(n9474) );
  AND U9485 ( .A(n9493), .B(n9494), .Z(n9492) );
  XOR U9486 ( .A(n9495), .B(n9491), .Z(n9493) );
  XNOR U9487 ( .A(n9496), .B(n9497), .Z(n9490) );
  AND U9488 ( .A(n9498), .B(n9499), .Z(n9497) );
  XOR U9489 ( .A(n9496), .B(n9500), .Z(n9498) );
  XNOR U9490 ( .A(n9480), .B(n9477), .Z(n9489) );
  AND U9491 ( .A(n9501), .B(n9502), .Z(n9477) );
  XOR U9492 ( .A(n9503), .B(n9504), .Z(n9480) );
  AND U9493 ( .A(n9505), .B(n9506), .Z(n9504) );
  XOR U9494 ( .A(n9503), .B(n9507), .Z(n9505) );
  XNOR U9495 ( .A(n9398), .B(n9485), .Z(n9487) );
  XOR U9496 ( .A(n9508), .B(n9509), .Z(n9398) );
  AND U9497 ( .A(n235), .B(n9510), .Z(n9509) );
  XNOR U9498 ( .A(n9511), .B(n9508), .Z(n9510) );
  XOR U9499 ( .A(n9512), .B(n9513), .Z(n9485) );
  AND U9500 ( .A(n9514), .B(n9515), .Z(n9513) );
  XNOR U9501 ( .A(n9512), .B(n9501), .Z(n9515) );
  IV U9502 ( .A(n9449), .Z(n9501) );
  XNOR U9503 ( .A(n9516), .B(n9494), .Z(n9449) );
  XNOR U9504 ( .A(n9517), .B(n9500), .Z(n9494) );
  XOR U9505 ( .A(n9518), .B(n9519), .Z(n9500) );
  NOR U9506 ( .A(n9520), .B(n9521), .Z(n9519) );
  XNOR U9507 ( .A(n9518), .B(n9522), .Z(n9520) );
  XNOR U9508 ( .A(n9499), .B(n9491), .Z(n9517) );
  XOR U9509 ( .A(n9523), .B(n9524), .Z(n9491) );
  AND U9510 ( .A(n9525), .B(n9526), .Z(n9524) );
  XNOR U9511 ( .A(n9523), .B(n9527), .Z(n9525) );
  XNOR U9512 ( .A(n9528), .B(n9496), .Z(n9499) );
  XOR U9513 ( .A(n9529), .B(n9530), .Z(n9496) );
  AND U9514 ( .A(n9531), .B(n9532), .Z(n9530) );
  XOR U9515 ( .A(n9529), .B(n9533), .Z(n9531) );
  XNOR U9516 ( .A(n9534), .B(n9535), .Z(n9528) );
  NOR U9517 ( .A(n9536), .B(n9537), .Z(n9535) );
  XOR U9518 ( .A(n9534), .B(n9538), .Z(n9536) );
  XNOR U9519 ( .A(n9495), .B(n9502), .Z(n9516) );
  NOR U9520 ( .A(n9461), .B(n9539), .Z(n9502) );
  XOR U9521 ( .A(n9507), .B(n9506), .Z(n9495) );
  XNOR U9522 ( .A(n9540), .B(n9503), .Z(n9506) );
  XOR U9523 ( .A(n9541), .B(n9542), .Z(n9503) );
  AND U9524 ( .A(n9543), .B(n9544), .Z(n9542) );
  XOR U9525 ( .A(n9541), .B(n9545), .Z(n9543) );
  XNOR U9526 ( .A(n9546), .B(n9547), .Z(n9540) );
  NOR U9527 ( .A(n9548), .B(n9549), .Z(n9547) );
  XNOR U9528 ( .A(n9546), .B(n9550), .Z(n9548) );
  XOR U9529 ( .A(n9551), .B(n9552), .Z(n9507) );
  NOR U9530 ( .A(n9553), .B(n9554), .Z(n9552) );
  XNOR U9531 ( .A(n9551), .B(n9555), .Z(n9553) );
  XNOR U9532 ( .A(n9446), .B(n9512), .Z(n9514) );
  XOR U9533 ( .A(n9556), .B(n9557), .Z(n9446) );
  AND U9534 ( .A(n235), .B(n9558), .Z(n9557) );
  XOR U9535 ( .A(n9559), .B(n9556), .Z(n9558) );
  AND U9536 ( .A(n9458), .B(n9461), .Z(n9512) );
  XOR U9537 ( .A(n9560), .B(n9539), .Z(n9461) );
  XNOR U9538 ( .A(p_input[1024]), .B(p_input[912]), .Z(n9539) );
  XOR U9539 ( .A(n9527), .B(n9526), .Z(n9560) );
  XNOR U9540 ( .A(n9561), .B(n9533), .Z(n9526) );
  XNOR U9541 ( .A(n9522), .B(n9521), .Z(n9533) );
  XOR U9542 ( .A(n9562), .B(n9518), .Z(n9521) );
  XOR U9543 ( .A(p_input[1034]), .B(p_input[922]), .Z(n9518) );
  XNOR U9544 ( .A(p_input[1035]), .B(p_input[923]), .Z(n9562) );
  XOR U9545 ( .A(p_input[1036]), .B(p_input[924]), .Z(n9522) );
  XNOR U9546 ( .A(n9532), .B(n9523), .Z(n9561) );
  XNOR U9547 ( .A(n3298), .B(p_input[913]), .Z(n9523) );
  XOR U9548 ( .A(n9563), .B(n9538), .Z(n9532) );
  XNOR U9549 ( .A(p_input[1039]), .B(p_input[927]), .Z(n9538) );
  XOR U9550 ( .A(n9529), .B(n9537), .Z(n9563) );
  XOR U9551 ( .A(n9564), .B(n9534), .Z(n9537) );
  XOR U9552 ( .A(p_input[1037]), .B(p_input[925]), .Z(n9534) );
  XNOR U9553 ( .A(p_input[1038]), .B(p_input[926]), .Z(n9564) );
  XOR U9554 ( .A(p_input[1033]), .B(p_input[921]), .Z(n9529) );
  XNOR U9555 ( .A(n9545), .B(n9544), .Z(n9527) );
  XNOR U9556 ( .A(n9565), .B(n9550), .Z(n9544) );
  XOR U9557 ( .A(p_input[1032]), .B(p_input[920]), .Z(n9550) );
  XOR U9558 ( .A(n9541), .B(n9549), .Z(n9565) );
  XOR U9559 ( .A(n9566), .B(n9546), .Z(n9549) );
  XOR U9560 ( .A(p_input[1030]), .B(p_input[918]), .Z(n9546) );
  XNOR U9561 ( .A(p_input[1031]), .B(p_input[919]), .Z(n9566) );
  XOR U9562 ( .A(p_input[1026]), .B(p_input[914]), .Z(n9541) );
  XNOR U9563 ( .A(n9555), .B(n9554), .Z(n9545) );
  XOR U9564 ( .A(n9567), .B(n9551), .Z(n9554) );
  XOR U9565 ( .A(p_input[1027]), .B(p_input[915]), .Z(n9551) );
  XNOR U9566 ( .A(p_input[1028]), .B(p_input[916]), .Z(n9567) );
  XOR U9567 ( .A(p_input[1029]), .B(p_input[917]), .Z(n9555) );
  XOR U9568 ( .A(n9568), .B(n9569), .Z(n9458) );
  AND U9569 ( .A(n235), .B(n9570), .Z(n9569) );
  XNOR U9570 ( .A(n9571), .B(n9568), .Z(n9570) );
  XNOR U9571 ( .A(n9572), .B(n9573), .Z(n235) );
  NOR U9572 ( .A(n9574), .B(n9575), .Z(n9573) );
  XOR U9573 ( .A(n9467), .B(n9572), .Z(n9575) );
  AND U9574 ( .A(n9576), .B(n9577), .Z(n9467) );
  NOR U9575 ( .A(n9572), .B(n9466), .Z(n9574) );
  AND U9576 ( .A(n9578), .B(n9579), .Z(n9466) );
  XOR U9577 ( .A(n9580), .B(n9581), .Z(n9572) );
  AND U9578 ( .A(n9582), .B(n9583), .Z(n9581) );
  XNOR U9579 ( .A(n9580), .B(n9578), .Z(n9583) );
  IV U9580 ( .A(n9484), .Z(n9578) );
  XOR U9581 ( .A(n9584), .B(n9585), .Z(n9484) );
  XOR U9582 ( .A(n9586), .B(n9579), .Z(n9585) );
  AND U9583 ( .A(n9511), .B(n9587), .Z(n9579) );
  AND U9584 ( .A(n9588), .B(n9589), .Z(n9586) );
  XOR U9585 ( .A(n9590), .B(n9584), .Z(n9588) );
  XNOR U9586 ( .A(n9481), .B(n9580), .Z(n9582) );
  XOR U9587 ( .A(n9591), .B(n9592), .Z(n9481) );
  AND U9588 ( .A(n239), .B(n9593), .Z(n9592) );
  XOR U9589 ( .A(n9594), .B(n9591), .Z(n9593) );
  XOR U9590 ( .A(n9595), .B(n9596), .Z(n9580) );
  AND U9591 ( .A(n9597), .B(n9598), .Z(n9596) );
  XNOR U9592 ( .A(n9595), .B(n9511), .Z(n9598) );
  XOR U9593 ( .A(n9599), .B(n9589), .Z(n9511) );
  XNOR U9594 ( .A(n9600), .B(n9584), .Z(n9589) );
  XOR U9595 ( .A(n9601), .B(n9602), .Z(n9584) );
  AND U9596 ( .A(n9603), .B(n9604), .Z(n9602) );
  XOR U9597 ( .A(n9605), .B(n9601), .Z(n9603) );
  XNOR U9598 ( .A(n9606), .B(n9607), .Z(n9600) );
  AND U9599 ( .A(n9608), .B(n9609), .Z(n9607) );
  XOR U9600 ( .A(n9606), .B(n9610), .Z(n9608) );
  XNOR U9601 ( .A(n9590), .B(n9587), .Z(n9599) );
  AND U9602 ( .A(n9611), .B(n9612), .Z(n9587) );
  XOR U9603 ( .A(n9613), .B(n9614), .Z(n9590) );
  AND U9604 ( .A(n9615), .B(n9616), .Z(n9614) );
  XOR U9605 ( .A(n9613), .B(n9617), .Z(n9615) );
  XNOR U9606 ( .A(n9508), .B(n9595), .Z(n9597) );
  XOR U9607 ( .A(n9618), .B(n9619), .Z(n9508) );
  AND U9608 ( .A(n239), .B(n9620), .Z(n9619) );
  XNOR U9609 ( .A(n9621), .B(n9618), .Z(n9620) );
  XOR U9610 ( .A(n9622), .B(n9623), .Z(n9595) );
  AND U9611 ( .A(n9624), .B(n9625), .Z(n9623) );
  XNOR U9612 ( .A(n9622), .B(n9611), .Z(n9625) );
  IV U9613 ( .A(n9559), .Z(n9611) );
  XNOR U9614 ( .A(n9626), .B(n9604), .Z(n9559) );
  XNOR U9615 ( .A(n9627), .B(n9610), .Z(n9604) );
  XOR U9616 ( .A(n9628), .B(n9629), .Z(n9610) );
  NOR U9617 ( .A(n9630), .B(n9631), .Z(n9629) );
  XNOR U9618 ( .A(n9628), .B(n9632), .Z(n9630) );
  XNOR U9619 ( .A(n9609), .B(n9601), .Z(n9627) );
  XOR U9620 ( .A(n9633), .B(n9634), .Z(n9601) );
  AND U9621 ( .A(n9635), .B(n9636), .Z(n9634) );
  XNOR U9622 ( .A(n9633), .B(n9637), .Z(n9635) );
  XNOR U9623 ( .A(n9638), .B(n9606), .Z(n9609) );
  XOR U9624 ( .A(n9639), .B(n9640), .Z(n9606) );
  AND U9625 ( .A(n9641), .B(n9642), .Z(n9640) );
  XOR U9626 ( .A(n9639), .B(n9643), .Z(n9641) );
  XNOR U9627 ( .A(n9644), .B(n9645), .Z(n9638) );
  NOR U9628 ( .A(n9646), .B(n9647), .Z(n9645) );
  XOR U9629 ( .A(n9644), .B(n9648), .Z(n9646) );
  XNOR U9630 ( .A(n9605), .B(n9612), .Z(n9626) );
  NOR U9631 ( .A(n9571), .B(n9649), .Z(n9612) );
  XOR U9632 ( .A(n9617), .B(n9616), .Z(n9605) );
  XNOR U9633 ( .A(n9650), .B(n9613), .Z(n9616) );
  XOR U9634 ( .A(n9651), .B(n9652), .Z(n9613) );
  AND U9635 ( .A(n9653), .B(n9654), .Z(n9652) );
  XOR U9636 ( .A(n9651), .B(n9655), .Z(n9653) );
  XNOR U9637 ( .A(n9656), .B(n9657), .Z(n9650) );
  NOR U9638 ( .A(n9658), .B(n9659), .Z(n9657) );
  XNOR U9639 ( .A(n9656), .B(n9660), .Z(n9658) );
  XOR U9640 ( .A(n9661), .B(n9662), .Z(n9617) );
  NOR U9641 ( .A(n9663), .B(n9664), .Z(n9662) );
  XNOR U9642 ( .A(n9661), .B(n9665), .Z(n9663) );
  XNOR U9643 ( .A(n9556), .B(n9622), .Z(n9624) );
  XOR U9644 ( .A(n9666), .B(n9667), .Z(n9556) );
  AND U9645 ( .A(n239), .B(n9668), .Z(n9667) );
  XOR U9646 ( .A(n9669), .B(n9666), .Z(n9668) );
  AND U9647 ( .A(n9568), .B(n9571), .Z(n9622) );
  XOR U9648 ( .A(n9670), .B(n9649), .Z(n9571) );
  XNOR U9649 ( .A(p_input[1024]), .B(p_input[928]), .Z(n9649) );
  XOR U9650 ( .A(n9637), .B(n9636), .Z(n9670) );
  XNOR U9651 ( .A(n9671), .B(n9643), .Z(n9636) );
  XNOR U9652 ( .A(n9632), .B(n9631), .Z(n9643) );
  XOR U9653 ( .A(n9672), .B(n9628), .Z(n9631) );
  XOR U9654 ( .A(p_input[1034]), .B(p_input[938]), .Z(n9628) );
  XNOR U9655 ( .A(p_input[1035]), .B(p_input[939]), .Z(n9672) );
  XOR U9656 ( .A(p_input[1036]), .B(p_input[940]), .Z(n9632) );
  XNOR U9657 ( .A(n9642), .B(n9633), .Z(n9671) );
  XNOR U9658 ( .A(n3298), .B(p_input[929]), .Z(n9633) );
  XOR U9659 ( .A(n9673), .B(n9648), .Z(n9642) );
  XNOR U9660 ( .A(p_input[1039]), .B(p_input[943]), .Z(n9648) );
  XOR U9661 ( .A(n9639), .B(n9647), .Z(n9673) );
  XOR U9662 ( .A(n9674), .B(n9644), .Z(n9647) );
  XOR U9663 ( .A(p_input[1037]), .B(p_input[941]), .Z(n9644) );
  XNOR U9664 ( .A(p_input[1038]), .B(p_input[942]), .Z(n9674) );
  XOR U9665 ( .A(p_input[1033]), .B(p_input[937]), .Z(n9639) );
  XNOR U9666 ( .A(n9655), .B(n9654), .Z(n9637) );
  XNOR U9667 ( .A(n9675), .B(n9660), .Z(n9654) );
  XOR U9668 ( .A(p_input[1032]), .B(p_input[936]), .Z(n9660) );
  XOR U9669 ( .A(n9651), .B(n9659), .Z(n9675) );
  XOR U9670 ( .A(n9676), .B(n9656), .Z(n9659) );
  XOR U9671 ( .A(p_input[1030]), .B(p_input[934]), .Z(n9656) );
  XNOR U9672 ( .A(p_input[1031]), .B(p_input[935]), .Z(n9676) );
  XOR U9673 ( .A(p_input[1026]), .B(p_input[930]), .Z(n9651) );
  XNOR U9674 ( .A(n9665), .B(n9664), .Z(n9655) );
  XOR U9675 ( .A(n9677), .B(n9661), .Z(n9664) );
  XOR U9676 ( .A(p_input[1027]), .B(p_input[931]), .Z(n9661) );
  XNOR U9677 ( .A(p_input[1028]), .B(p_input[932]), .Z(n9677) );
  XOR U9678 ( .A(p_input[1029]), .B(p_input[933]), .Z(n9665) );
  XOR U9679 ( .A(n9678), .B(n9679), .Z(n9568) );
  AND U9680 ( .A(n239), .B(n9680), .Z(n9679) );
  XNOR U9681 ( .A(n9681), .B(n9678), .Z(n9680) );
  XNOR U9682 ( .A(n9682), .B(n9683), .Z(n239) );
  NOR U9683 ( .A(n9684), .B(n9685), .Z(n9683) );
  XOR U9684 ( .A(n9577), .B(n9682), .Z(n9685) );
  AND U9685 ( .A(n9686), .B(n9687), .Z(n9577) );
  NOR U9686 ( .A(n9682), .B(n9576), .Z(n9684) );
  AND U9687 ( .A(n9688), .B(n9689), .Z(n9576) );
  XOR U9688 ( .A(n9690), .B(n9691), .Z(n9682) );
  AND U9689 ( .A(n9692), .B(n9693), .Z(n9691) );
  XNOR U9690 ( .A(n9690), .B(n9688), .Z(n9693) );
  IV U9691 ( .A(n9594), .Z(n9688) );
  XOR U9692 ( .A(n9694), .B(n9695), .Z(n9594) );
  XOR U9693 ( .A(n9696), .B(n9689), .Z(n9695) );
  AND U9694 ( .A(n9621), .B(n9697), .Z(n9689) );
  AND U9695 ( .A(n9698), .B(n9699), .Z(n9696) );
  XOR U9696 ( .A(n9700), .B(n9694), .Z(n9698) );
  XNOR U9697 ( .A(n9591), .B(n9690), .Z(n9692) );
  XOR U9698 ( .A(n9701), .B(n9702), .Z(n9591) );
  AND U9699 ( .A(n243), .B(n9703), .Z(n9702) );
  XOR U9700 ( .A(n9704), .B(n9701), .Z(n9703) );
  XOR U9701 ( .A(n9705), .B(n9706), .Z(n9690) );
  AND U9702 ( .A(n9707), .B(n9708), .Z(n9706) );
  XNOR U9703 ( .A(n9705), .B(n9621), .Z(n9708) );
  XOR U9704 ( .A(n9709), .B(n9699), .Z(n9621) );
  XNOR U9705 ( .A(n9710), .B(n9694), .Z(n9699) );
  XOR U9706 ( .A(n9711), .B(n9712), .Z(n9694) );
  AND U9707 ( .A(n9713), .B(n9714), .Z(n9712) );
  XOR U9708 ( .A(n9715), .B(n9711), .Z(n9713) );
  XNOR U9709 ( .A(n9716), .B(n9717), .Z(n9710) );
  AND U9710 ( .A(n9718), .B(n9719), .Z(n9717) );
  XOR U9711 ( .A(n9716), .B(n9720), .Z(n9718) );
  XNOR U9712 ( .A(n9700), .B(n9697), .Z(n9709) );
  AND U9713 ( .A(n9721), .B(n9722), .Z(n9697) );
  XOR U9714 ( .A(n9723), .B(n9724), .Z(n9700) );
  AND U9715 ( .A(n9725), .B(n9726), .Z(n9724) );
  XOR U9716 ( .A(n9723), .B(n9727), .Z(n9725) );
  XNOR U9717 ( .A(n9618), .B(n9705), .Z(n9707) );
  XOR U9718 ( .A(n9728), .B(n9729), .Z(n9618) );
  AND U9719 ( .A(n243), .B(n9730), .Z(n9729) );
  XNOR U9720 ( .A(n9731), .B(n9728), .Z(n9730) );
  XOR U9721 ( .A(n9732), .B(n9733), .Z(n9705) );
  AND U9722 ( .A(n9734), .B(n9735), .Z(n9733) );
  XNOR U9723 ( .A(n9732), .B(n9721), .Z(n9735) );
  IV U9724 ( .A(n9669), .Z(n9721) );
  XNOR U9725 ( .A(n9736), .B(n9714), .Z(n9669) );
  XNOR U9726 ( .A(n9737), .B(n9720), .Z(n9714) );
  XOR U9727 ( .A(n9738), .B(n9739), .Z(n9720) );
  NOR U9728 ( .A(n9740), .B(n9741), .Z(n9739) );
  XNOR U9729 ( .A(n9738), .B(n9742), .Z(n9740) );
  XNOR U9730 ( .A(n9719), .B(n9711), .Z(n9737) );
  XOR U9731 ( .A(n9743), .B(n9744), .Z(n9711) );
  AND U9732 ( .A(n9745), .B(n9746), .Z(n9744) );
  XNOR U9733 ( .A(n9743), .B(n9747), .Z(n9745) );
  XNOR U9734 ( .A(n9748), .B(n9716), .Z(n9719) );
  XOR U9735 ( .A(n9749), .B(n9750), .Z(n9716) );
  AND U9736 ( .A(n9751), .B(n9752), .Z(n9750) );
  XOR U9737 ( .A(n9749), .B(n9753), .Z(n9751) );
  XNOR U9738 ( .A(n9754), .B(n9755), .Z(n9748) );
  NOR U9739 ( .A(n9756), .B(n9757), .Z(n9755) );
  XOR U9740 ( .A(n9754), .B(n9758), .Z(n9756) );
  XNOR U9741 ( .A(n9715), .B(n9722), .Z(n9736) );
  NOR U9742 ( .A(n9681), .B(n9759), .Z(n9722) );
  XOR U9743 ( .A(n9727), .B(n9726), .Z(n9715) );
  XNOR U9744 ( .A(n9760), .B(n9723), .Z(n9726) );
  XOR U9745 ( .A(n9761), .B(n9762), .Z(n9723) );
  AND U9746 ( .A(n9763), .B(n9764), .Z(n9762) );
  XOR U9747 ( .A(n9761), .B(n9765), .Z(n9763) );
  XNOR U9748 ( .A(n9766), .B(n9767), .Z(n9760) );
  NOR U9749 ( .A(n9768), .B(n9769), .Z(n9767) );
  XNOR U9750 ( .A(n9766), .B(n9770), .Z(n9768) );
  XOR U9751 ( .A(n9771), .B(n9772), .Z(n9727) );
  NOR U9752 ( .A(n9773), .B(n9774), .Z(n9772) );
  XNOR U9753 ( .A(n9771), .B(n9775), .Z(n9773) );
  XNOR U9754 ( .A(n9666), .B(n9732), .Z(n9734) );
  XOR U9755 ( .A(n9776), .B(n9777), .Z(n9666) );
  AND U9756 ( .A(n243), .B(n9778), .Z(n9777) );
  XOR U9757 ( .A(n9779), .B(n9776), .Z(n9778) );
  AND U9758 ( .A(n9678), .B(n9681), .Z(n9732) );
  XOR U9759 ( .A(n9780), .B(n9759), .Z(n9681) );
  XNOR U9760 ( .A(p_input[1024]), .B(p_input[944]), .Z(n9759) );
  XOR U9761 ( .A(n9747), .B(n9746), .Z(n9780) );
  XNOR U9762 ( .A(n9781), .B(n9753), .Z(n9746) );
  XNOR U9763 ( .A(n9742), .B(n9741), .Z(n9753) );
  XOR U9764 ( .A(n9782), .B(n9738), .Z(n9741) );
  XOR U9765 ( .A(p_input[1034]), .B(p_input[954]), .Z(n9738) );
  XNOR U9766 ( .A(p_input[1035]), .B(p_input[955]), .Z(n9782) );
  XOR U9767 ( .A(p_input[1036]), .B(p_input[956]), .Z(n9742) );
  XNOR U9768 ( .A(n9752), .B(n9743), .Z(n9781) );
  XNOR U9769 ( .A(n3298), .B(p_input[945]), .Z(n9743) );
  XOR U9770 ( .A(n9783), .B(n9758), .Z(n9752) );
  XNOR U9771 ( .A(p_input[1039]), .B(p_input[959]), .Z(n9758) );
  XOR U9772 ( .A(n9749), .B(n9757), .Z(n9783) );
  XOR U9773 ( .A(n9784), .B(n9754), .Z(n9757) );
  XOR U9774 ( .A(p_input[1037]), .B(p_input[957]), .Z(n9754) );
  XNOR U9775 ( .A(p_input[1038]), .B(p_input[958]), .Z(n9784) );
  XOR U9776 ( .A(p_input[1033]), .B(p_input[953]), .Z(n9749) );
  XNOR U9777 ( .A(n9765), .B(n9764), .Z(n9747) );
  XNOR U9778 ( .A(n9785), .B(n9770), .Z(n9764) );
  XOR U9779 ( .A(p_input[1032]), .B(p_input[952]), .Z(n9770) );
  XOR U9780 ( .A(n9761), .B(n9769), .Z(n9785) );
  XOR U9781 ( .A(n9786), .B(n9766), .Z(n9769) );
  XOR U9782 ( .A(p_input[1030]), .B(p_input[950]), .Z(n9766) );
  XNOR U9783 ( .A(p_input[1031]), .B(p_input[951]), .Z(n9786) );
  XOR U9784 ( .A(p_input[1026]), .B(p_input[946]), .Z(n9761) );
  XNOR U9785 ( .A(n9775), .B(n9774), .Z(n9765) );
  XOR U9786 ( .A(n9787), .B(n9771), .Z(n9774) );
  XOR U9787 ( .A(p_input[1027]), .B(p_input[947]), .Z(n9771) );
  XNOR U9788 ( .A(p_input[1028]), .B(p_input[948]), .Z(n9787) );
  XOR U9789 ( .A(p_input[1029]), .B(p_input[949]), .Z(n9775) );
  XOR U9790 ( .A(n9788), .B(n9789), .Z(n9678) );
  AND U9791 ( .A(n243), .B(n9790), .Z(n9789) );
  XNOR U9792 ( .A(n9791), .B(n9788), .Z(n9790) );
  XNOR U9793 ( .A(n9792), .B(n9793), .Z(n243) );
  NOR U9794 ( .A(n9794), .B(n9795), .Z(n9793) );
  XOR U9795 ( .A(n9687), .B(n9792), .Z(n9795) );
  AND U9796 ( .A(n9796), .B(n9797), .Z(n9687) );
  NOR U9797 ( .A(n9792), .B(n9686), .Z(n9794) );
  AND U9798 ( .A(n9798), .B(n9799), .Z(n9686) );
  XOR U9799 ( .A(n9800), .B(n9801), .Z(n9792) );
  AND U9800 ( .A(n9802), .B(n9803), .Z(n9801) );
  XNOR U9801 ( .A(n9800), .B(n9798), .Z(n9803) );
  IV U9802 ( .A(n9704), .Z(n9798) );
  XOR U9803 ( .A(n9804), .B(n9805), .Z(n9704) );
  XOR U9804 ( .A(n9806), .B(n9799), .Z(n9805) );
  AND U9805 ( .A(n9731), .B(n9807), .Z(n9799) );
  AND U9806 ( .A(n9808), .B(n9809), .Z(n9806) );
  XOR U9807 ( .A(n9810), .B(n9804), .Z(n9808) );
  XNOR U9808 ( .A(n9701), .B(n9800), .Z(n9802) );
  XOR U9809 ( .A(n9811), .B(n9812), .Z(n9701) );
  AND U9810 ( .A(n247), .B(n9813), .Z(n9812) );
  XOR U9811 ( .A(n9814), .B(n9811), .Z(n9813) );
  XOR U9812 ( .A(n9815), .B(n9816), .Z(n9800) );
  AND U9813 ( .A(n9817), .B(n9818), .Z(n9816) );
  XNOR U9814 ( .A(n9815), .B(n9731), .Z(n9818) );
  XOR U9815 ( .A(n9819), .B(n9809), .Z(n9731) );
  XNOR U9816 ( .A(n9820), .B(n9804), .Z(n9809) );
  XOR U9817 ( .A(n9821), .B(n9822), .Z(n9804) );
  AND U9818 ( .A(n9823), .B(n9824), .Z(n9822) );
  XOR U9819 ( .A(n9825), .B(n9821), .Z(n9823) );
  XNOR U9820 ( .A(n9826), .B(n9827), .Z(n9820) );
  AND U9821 ( .A(n9828), .B(n9829), .Z(n9827) );
  XOR U9822 ( .A(n9826), .B(n9830), .Z(n9828) );
  XNOR U9823 ( .A(n9810), .B(n9807), .Z(n9819) );
  AND U9824 ( .A(n9831), .B(n9832), .Z(n9807) );
  XOR U9825 ( .A(n9833), .B(n9834), .Z(n9810) );
  AND U9826 ( .A(n9835), .B(n9836), .Z(n9834) );
  XOR U9827 ( .A(n9833), .B(n9837), .Z(n9835) );
  XNOR U9828 ( .A(n9728), .B(n9815), .Z(n9817) );
  XOR U9829 ( .A(n9838), .B(n9839), .Z(n9728) );
  AND U9830 ( .A(n247), .B(n9840), .Z(n9839) );
  XNOR U9831 ( .A(n9841), .B(n9838), .Z(n9840) );
  XOR U9832 ( .A(n9842), .B(n9843), .Z(n9815) );
  AND U9833 ( .A(n9844), .B(n9845), .Z(n9843) );
  XNOR U9834 ( .A(n9842), .B(n9831), .Z(n9845) );
  IV U9835 ( .A(n9779), .Z(n9831) );
  XNOR U9836 ( .A(n9846), .B(n9824), .Z(n9779) );
  XNOR U9837 ( .A(n9847), .B(n9830), .Z(n9824) );
  XOR U9838 ( .A(n9848), .B(n9849), .Z(n9830) );
  NOR U9839 ( .A(n9850), .B(n9851), .Z(n9849) );
  XNOR U9840 ( .A(n9848), .B(n9852), .Z(n9850) );
  XNOR U9841 ( .A(n9829), .B(n9821), .Z(n9847) );
  XOR U9842 ( .A(n9853), .B(n9854), .Z(n9821) );
  AND U9843 ( .A(n9855), .B(n9856), .Z(n9854) );
  XNOR U9844 ( .A(n9853), .B(n9857), .Z(n9855) );
  XNOR U9845 ( .A(n9858), .B(n9826), .Z(n9829) );
  XOR U9846 ( .A(n9859), .B(n9860), .Z(n9826) );
  AND U9847 ( .A(n9861), .B(n9862), .Z(n9860) );
  XOR U9848 ( .A(n9859), .B(n9863), .Z(n9861) );
  XNOR U9849 ( .A(n9864), .B(n9865), .Z(n9858) );
  NOR U9850 ( .A(n9866), .B(n9867), .Z(n9865) );
  XOR U9851 ( .A(n9864), .B(n9868), .Z(n9866) );
  XNOR U9852 ( .A(n9825), .B(n9832), .Z(n9846) );
  NOR U9853 ( .A(n9791), .B(n9869), .Z(n9832) );
  XOR U9854 ( .A(n9837), .B(n9836), .Z(n9825) );
  XNOR U9855 ( .A(n9870), .B(n9833), .Z(n9836) );
  XOR U9856 ( .A(n9871), .B(n9872), .Z(n9833) );
  AND U9857 ( .A(n9873), .B(n9874), .Z(n9872) );
  XOR U9858 ( .A(n9871), .B(n9875), .Z(n9873) );
  XNOR U9859 ( .A(n9876), .B(n9877), .Z(n9870) );
  NOR U9860 ( .A(n9878), .B(n9879), .Z(n9877) );
  XNOR U9861 ( .A(n9876), .B(n9880), .Z(n9878) );
  XOR U9862 ( .A(n9881), .B(n9882), .Z(n9837) );
  NOR U9863 ( .A(n9883), .B(n9884), .Z(n9882) );
  XNOR U9864 ( .A(n9881), .B(n9885), .Z(n9883) );
  XNOR U9865 ( .A(n9776), .B(n9842), .Z(n9844) );
  XOR U9866 ( .A(n9886), .B(n9887), .Z(n9776) );
  AND U9867 ( .A(n247), .B(n9888), .Z(n9887) );
  XOR U9868 ( .A(n9889), .B(n9886), .Z(n9888) );
  AND U9869 ( .A(n9788), .B(n9791), .Z(n9842) );
  XOR U9870 ( .A(n9890), .B(n9869), .Z(n9791) );
  XNOR U9871 ( .A(p_input[1024]), .B(p_input[960]), .Z(n9869) );
  XOR U9872 ( .A(n9857), .B(n9856), .Z(n9890) );
  XNOR U9873 ( .A(n9891), .B(n9863), .Z(n9856) );
  XNOR U9874 ( .A(n9852), .B(n9851), .Z(n9863) );
  XOR U9875 ( .A(n9892), .B(n9848), .Z(n9851) );
  XOR U9876 ( .A(p_input[1034]), .B(p_input[970]), .Z(n9848) );
  XNOR U9877 ( .A(p_input[1035]), .B(p_input[971]), .Z(n9892) );
  XOR U9878 ( .A(p_input[1036]), .B(p_input[972]), .Z(n9852) );
  XNOR U9879 ( .A(n9862), .B(n9853), .Z(n9891) );
  XNOR U9880 ( .A(n3298), .B(p_input[961]), .Z(n9853) );
  XOR U9881 ( .A(n9893), .B(n9868), .Z(n9862) );
  XNOR U9882 ( .A(p_input[1039]), .B(p_input[975]), .Z(n9868) );
  XOR U9883 ( .A(n9859), .B(n9867), .Z(n9893) );
  XOR U9884 ( .A(n9894), .B(n9864), .Z(n9867) );
  XOR U9885 ( .A(p_input[1037]), .B(p_input[973]), .Z(n9864) );
  XNOR U9886 ( .A(p_input[1038]), .B(p_input[974]), .Z(n9894) );
  XOR U9887 ( .A(p_input[1033]), .B(p_input[969]), .Z(n9859) );
  XNOR U9888 ( .A(n9875), .B(n9874), .Z(n9857) );
  XNOR U9889 ( .A(n9895), .B(n9880), .Z(n9874) );
  XOR U9890 ( .A(p_input[1032]), .B(p_input[968]), .Z(n9880) );
  XOR U9891 ( .A(n9871), .B(n9879), .Z(n9895) );
  XOR U9892 ( .A(n9896), .B(n9876), .Z(n9879) );
  XOR U9893 ( .A(p_input[1030]), .B(p_input[966]), .Z(n9876) );
  XNOR U9894 ( .A(p_input[1031]), .B(p_input[967]), .Z(n9896) );
  XOR U9895 ( .A(p_input[1026]), .B(p_input[962]), .Z(n9871) );
  XNOR U9896 ( .A(n9885), .B(n9884), .Z(n9875) );
  XOR U9897 ( .A(n9897), .B(n9881), .Z(n9884) );
  XOR U9898 ( .A(p_input[1027]), .B(p_input[963]), .Z(n9881) );
  XNOR U9899 ( .A(p_input[1028]), .B(p_input[964]), .Z(n9897) );
  XOR U9900 ( .A(p_input[1029]), .B(p_input[965]), .Z(n9885) );
  XOR U9901 ( .A(n9898), .B(n9899), .Z(n9788) );
  AND U9902 ( .A(n247), .B(n9900), .Z(n9899) );
  XNOR U9903 ( .A(n9901), .B(n9898), .Z(n9900) );
  XNOR U9904 ( .A(n9902), .B(n9903), .Z(n247) );
  NOR U9905 ( .A(n9904), .B(n9905), .Z(n9903) );
  XOR U9906 ( .A(n9797), .B(n9902), .Z(n9905) );
  AND U9907 ( .A(n9906), .B(n9907), .Z(n9797) );
  NOR U9908 ( .A(n9902), .B(n9796), .Z(n9904) );
  AND U9909 ( .A(n9908), .B(n9909), .Z(n9796) );
  XOR U9910 ( .A(n9910), .B(n9911), .Z(n9902) );
  AND U9911 ( .A(n9912), .B(n9913), .Z(n9911) );
  XNOR U9912 ( .A(n9910), .B(n9908), .Z(n9913) );
  IV U9913 ( .A(n9814), .Z(n9908) );
  XOR U9914 ( .A(n9914), .B(n9915), .Z(n9814) );
  XOR U9915 ( .A(n9916), .B(n9909), .Z(n9915) );
  AND U9916 ( .A(n9841), .B(n9917), .Z(n9909) );
  AND U9917 ( .A(n9918), .B(n9919), .Z(n9916) );
  XOR U9918 ( .A(n9920), .B(n9914), .Z(n9918) );
  XNOR U9919 ( .A(n9811), .B(n9910), .Z(n9912) );
  XNOR U9920 ( .A(n9921), .B(n9922), .Z(n9811) );
  AND U9921 ( .A(n250), .B(n9923), .Z(n9922) );
  XNOR U9922 ( .A(n9924), .B(n9921), .Z(n9923) );
  XOR U9923 ( .A(n9925), .B(n9926), .Z(n9910) );
  AND U9924 ( .A(n9927), .B(n9928), .Z(n9926) );
  XNOR U9925 ( .A(n9925), .B(n9841), .Z(n9928) );
  XOR U9926 ( .A(n9929), .B(n9919), .Z(n9841) );
  XNOR U9927 ( .A(n9930), .B(n9914), .Z(n9919) );
  XOR U9928 ( .A(n9931), .B(n9932), .Z(n9914) );
  AND U9929 ( .A(n9933), .B(n9934), .Z(n9932) );
  XOR U9930 ( .A(n9935), .B(n9931), .Z(n9933) );
  XNOR U9931 ( .A(n9936), .B(n9937), .Z(n9930) );
  AND U9932 ( .A(n9938), .B(n9939), .Z(n9937) );
  XOR U9933 ( .A(n9936), .B(n9940), .Z(n9938) );
  XNOR U9934 ( .A(n9920), .B(n9917), .Z(n9929) );
  AND U9935 ( .A(n9941), .B(n9942), .Z(n9917) );
  XOR U9936 ( .A(n9943), .B(n9944), .Z(n9920) );
  AND U9937 ( .A(n9945), .B(n9946), .Z(n9944) );
  XOR U9938 ( .A(n9943), .B(n9947), .Z(n9945) );
  XNOR U9939 ( .A(n9838), .B(n9925), .Z(n9927) );
  XNOR U9940 ( .A(n9948), .B(n9949), .Z(n9838) );
  AND U9941 ( .A(n250), .B(n9950), .Z(n9949) );
  XOR U9942 ( .A(n9951), .B(n9948), .Z(n9950) );
  XOR U9943 ( .A(n9952), .B(n9953), .Z(n9925) );
  AND U9944 ( .A(n9954), .B(n9955), .Z(n9953) );
  XNOR U9945 ( .A(n9952), .B(n9941), .Z(n9955) );
  IV U9946 ( .A(n9889), .Z(n9941) );
  XNOR U9947 ( .A(n9956), .B(n9934), .Z(n9889) );
  XNOR U9948 ( .A(n9957), .B(n9940), .Z(n9934) );
  XOR U9949 ( .A(n9958), .B(n9959), .Z(n9940) );
  NOR U9950 ( .A(n9960), .B(n9961), .Z(n9959) );
  XNOR U9951 ( .A(n9958), .B(n9962), .Z(n9960) );
  XNOR U9952 ( .A(n9939), .B(n9931), .Z(n9957) );
  XOR U9953 ( .A(n9963), .B(n9964), .Z(n9931) );
  AND U9954 ( .A(n9965), .B(n9966), .Z(n9964) );
  XNOR U9955 ( .A(n9963), .B(n9967), .Z(n9965) );
  XNOR U9956 ( .A(n9968), .B(n9936), .Z(n9939) );
  XOR U9957 ( .A(n9969), .B(n9970), .Z(n9936) );
  AND U9958 ( .A(n9971), .B(n9972), .Z(n9970) );
  XOR U9959 ( .A(n9969), .B(n9973), .Z(n9971) );
  XNOR U9960 ( .A(n9974), .B(n9975), .Z(n9968) );
  NOR U9961 ( .A(n9976), .B(n9977), .Z(n9975) );
  XOR U9962 ( .A(n9974), .B(n9978), .Z(n9976) );
  XNOR U9963 ( .A(n9935), .B(n9942), .Z(n9956) );
  NOR U9964 ( .A(n9901), .B(n9979), .Z(n9942) );
  XOR U9965 ( .A(n9947), .B(n9946), .Z(n9935) );
  XNOR U9966 ( .A(n9980), .B(n9943), .Z(n9946) );
  XOR U9967 ( .A(n9981), .B(n9982), .Z(n9943) );
  AND U9968 ( .A(n9983), .B(n9984), .Z(n9982) );
  XOR U9969 ( .A(n9981), .B(n9985), .Z(n9983) );
  XNOR U9970 ( .A(n9986), .B(n9987), .Z(n9980) );
  NOR U9971 ( .A(n9988), .B(n9989), .Z(n9987) );
  XNOR U9972 ( .A(n9986), .B(n9990), .Z(n9988) );
  XOR U9973 ( .A(n9991), .B(n9992), .Z(n9947) );
  NOR U9974 ( .A(n9993), .B(n9994), .Z(n9992) );
  XNOR U9975 ( .A(n9991), .B(n9995), .Z(n9993) );
  XNOR U9976 ( .A(n9886), .B(n9952), .Z(n9954) );
  XNOR U9977 ( .A(n9996), .B(n9997), .Z(n9886) );
  AND U9978 ( .A(n250), .B(n9998), .Z(n9997) );
  XNOR U9979 ( .A(n9999), .B(n9996), .Z(n9998) );
  AND U9980 ( .A(n9898), .B(n9901), .Z(n9952) );
  XOR U9981 ( .A(n10000), .B(n9979), .Z(n9901) );
  XNOR U9982 ( .A(p_input[1024]), .B(p_input[976]), .Z(n9979) );
  XOR U9983 ( .A(n9967), .B(n9966), .Z(n10000) );
  XNOR U9984 ( .A(n10001), .B(n9973), .Z(n9966) );
  XNOR U9985 ( .A(n9962), .B(n9961), .Z(n9973) );
  XOR U9986 ( .A(n10002), .B(n9958), .Z(n9961) );
  XOR U9987 ( .A(p_input[1034]), .B(p_input[986]), .Z(n9958) );
  XNOR U9988 ( .A(p_input[1035]), .B(p_input[987]), .Z(n10002) );
  XOR U9989 ( .A(p_input[1036]), .B(p_input[988]), .Z(n9962) );
  XNOR U9990 ( .A(n9972), .B(n9963), .Z(n10001) );
  XNOR U9991 ( .A(n3298), .B(p_input[977]), .Z(n9963) );
  XOR U9992 ( .A(n10003), .B(n9978), .Z(n9972) );
  XNOR U9993 ( .A(p_input[1039]), .B(p_input[991]), .Z(n9978) );
  XOR U9994 ( .A(n9969), .B(n9977), .Z(n10003) );
  XOR U9995 ( .A(n10004), .B(n9974), .Z(n9977) );
  XOR U9996 ( .A(p_input[1037]), .B(p_input[989]), .Z(n9974) );
  XNOR U9997 ( .A(p_input[1038]), .B(p_input[990]), .Z(n10004) );
  XOR U9998 ( .A(p_input[1033]), .B(p_input[985]), .Z(n9969) );
  XNOR U9999 ( .A(n9985), .B(n9984), .Z(n9967) );
  XNOR U10000 ( .A(n10005), .B(n9990), .Z(n9984) );
  XOR U10001 ( .A(p_input[1032]), .B(p_input[984]), .Z(n9990) );
  XOR U10002 ( .A(n9981), .B(n9989), .Z(n10005) );
  XOR U10003 ( .A(n10006), .B(n9986), .Z(n9989) );
  XOR U10004 ( .A(p_input[1030]), .B(p_input[982]), .Z(n9986) );
  XNOR U10005 ( .A(p_input[1031]), .B(p_input[983]), .Z(n10006) );
  XOR U10006 ( .A(p_input[1026]), .B(p_input[978]), .Z(n9981) );
  XNOR U10007 ( .A(n9995), .B(n9994), .Z(n9985) );
  XOR U10008 ( .A(n10007), .B(n9991), .Z(n9994) );
  XOR U10009 ( .A(p_input[1027]), .B(p_input[979]), .Z(n9991) );
  XNOR U10010 ( .A(p_input[1028]), .B(p_input[980]), .Z(n10007) );
  XOR U10011 ( .A(p_input[1029]), .B(p_input[981]), .Z(n9995) );
  XOR U10012 ( .A(n10008), .B(n10009), .Z(n9898) );
  AND U10013 ( .A(n250), .B(n10010), .Z(n10009) );
  XNOR U10014 ( .A(n10011), .B(n10008), .Z(n10010) );
  XNOR U10015 ( .A(n10012), .B(n10013), .Z(n250) );
  NOR U10016 ( .A(n10014), .B(n10015), .Z(n10013) );
  XOR U10017 ( .A(n9907), .B(n10012), .Z(n10015) );
  AND U10018 ( .A(n9921), .B(n10016), .Z(n9907) );
  NOR U10019 ( .A(n10012), .B(n9906), .Z(n10014) );
  AND U10020 ( .A(n10017), .B(n10018), .Z(n9906) );
  XOR U10021 ( .A(n10019), .B(n10020), .Z(n10012) );
  AND U10022 ( .A(n10021), .B(n10022), .Z(n10020) );
  XNOR U10023 ( .A(n10019), .B(n10017), .Z(n10022) );
  IV U10024 ( .A(n9924), .Z(n10017) );
  XOR U10025 ( .A(n10023), .B(n10024), .Z(n9924) );
  XOR U10026 ( .A(n10025), .B(n10018), .Z(n10024) );
  AND U10027 ( .A(n9951), .B(n10026), .Z(n10018) );
  AND U10028 ( .A(n10027), .B(n10028), .Z(n10025) );
  XOR U10029 ( .A(n10029), .B(n10023), .Z(n10027) );
  XNOR U10030 ( .A(n10030), .B(n10019), .Z(n10021) );
  IV U10031 ( .A(n9921), .Z(n10030) );
  XNOR U10032 ( .A(n10031), .B(n10032), .Z(n9921) );
  XOR U10033 ( .A(n10033), .B(n10016), .Z(n10032) );
  AND U10034 ( .A(n9948), .B(n10034), .Z(n10016) );
  AND U10035 ( .A(n10035), .B(n10036), .Z(n10033) );
  XNOR U10036 ( .A(n10031), .B(n10037), .Z(n10035) );
  XOR U10037 ( .A(n10038), .B(n10039), .Z(n10019) );
  AND U10038 ( .A(n10040), .B(n10041), .Z(n10039) );
  XNOR U10039 ( .A(n10038), .B(n9951), .Z(n10041) );
  XOR U10040 ( .A(n10042), .B(n10028), .Z(n9951) );
  XNOR U10041 ( .A(n10043), .B(n10023), .Z(n10028) );
  XOR U10042 ( .A(n10044), .B(n10045), .Z(n10023) );
  AND U10043 ( .A(n10046), .B(n10047), .Z(n10045) );
  XOR U10044 ( .A(n10048), .B(n10044), .Z(n10046) );
  XNOR U10045 ( .A(n10049), .B(n10050), .Z(n10043) );
  AND U10046 ( .A(n10051), .B(n10052), .Z(n10050) );
  XOR U10047 ( .A(n10049), .B(n10053), .Z(n10051) );
  XNOR U10048 ( .A(n10029), .B(n10026), .Z(n10042) );
  AND U10049 ( .A(n10054), .B(n10055), .Z(n10026) );
  XOR U10050 ( .A(n10056), .B(n10057), .Z(n10029) );
  AND U10051 ( .A(n10058), .B(n10059), .Z(n10057) );
  XOR U10052 ( .A(n10056), .B(n10060), .Z(n10058) );
  XOR U10053 ( .A(n9948), .B(n10038), .Z(n10040) );
  XNOR U10054 ( .A(n10061), .B(n10037), .Z(n9948) );
  XNOR U10055 ( .A(n10062), .B(n10063), .Z(n10037) );
  AND U10056 ( .A(n10064), .B(n10065), .Z(n10063) );
  XOR U10057 ( .A(n10062), .B(n10066), .Z(n10064) );
  XNOR U10058 ( .A(n10036), .B(n10034), .Z(n10061) );
  AND U10059 ( .A(n9996), .B(n10067), .Z(n10034) );
  XNOR U10060 ( .A(n10068), .B(n10031), .Z(n10036) );
  XOR U10061 ( .A(n10069), .B(n10070), .Z(n10031) );
  AND U10062 ( .A(n10071), .B(n10072), .Z(n10070) );
  XOR U10063 ( .A(n10069), .B(n10073), .Z(n10071) );
  XNOR U10064 ( .A(n10074), .B(n10075), .Z(n10068) );
  AND U10065 ( .A(n10076), .B(n10077), .Z(n10075) );
  XNOR U10066 ( .A(n10074), .B(n10078), .Z(n10076) );
  XOR U10067 ( .A(n10079), .B(n10080), .Z(n10038) );
  AND U10068 ( .A(n10081), .B(n10082), .Z(n10080) );
  XNOR U10069 ( .A(n10079), .B(n10054), .Z(n10082) );
  IV U10070 ( .A(n9999), .Z(n10054) );
  XNOR U10071 ( .A(n10083), .B(n10047), .Z(n9999) );
  XNOR U10072 ( .A(n10084), .B(n10053), .Z(n10047) );
  XOR U10073 ( .A(n10085), .B(n10086), .Z(n10053) );
  NOR U10074 ( .A(n10087), .B(n10088), .Z(n10086) );
  XNOR U10075 ( .A(n10085), .B(n10089), .Z(n10087) );
  XNOR U10076 ( .A(n10052), .B(n10044), .Z(n10084) );
  XOR U10077 ( .A(n10090), .B(n10091), .Z(n10044) );
  AND U10078 ( .A(n10092), .B(n10093), .Z(n10091) );
  XOR U10079 ( .A(n10090), .B(n10094), .Z(n10092) );
  XNOR U10080 ( .A(n10095), .B(n10049), .Z(n10052) );
  XOR U10081 ( .A(n10096), .B(n10097), .Z(n10049) );
  NOR U10082 ( .A(n10098), .B(n10099), .Z(n10097) );
  XNOR U10083 ( .A(n10096), .B(n10100), .Z(n10098) );
  XNOR U10084 ( .A(n10101), .B(n10102), .Z(n10095) );
  NOR U10085 ( .A(n10103), .B(n10104), .Z(n10102) );
  XNOR U10086 ( .A(n10101), .B(n10105), .Z(n10103) );
  XNOR U10087 ( .A(n10048), .B(n10055), .Z(n10083) );
  NOR U10088 ( .A(n10011), .B(n10106), .Z(n10055) );
  XOR U10089 ( .A(n10060), .B(n10059), .Z(n10048) );
  XNOR U10090 ( .A(n10107), .B(n10056), .Z(n10059) );
  XOR U10091 ( .A(n10108), .B(n10109), .Z(n10056) );
  NOR U10092 ( .A(n10110), .B(n10111), .Z(n10109) );
  XNOR U10093 ( .A(n10108), .B(n10112), .Z(n10110) );
  XNOR U10094 ( .A(n10113), .B(n10114), .Z(n10107) );
  NOR U10095 ( .A(n10115), .B(n10116), .Z(n10114) );
  XNOR U10096 ( .A(n10113), .B(n10117), .Z(n10115) );
  XOR U10097 ( .A(n10118), .B(n10119), .Z(n10060) );
  NOR U10098 ( .A(n10120), .B(n10121), .Z(n10119) );
  XNOR U10099 ( .A(n10118), .B(n10122), .Z(n10120) );
  XNOR U10100 ( .A(n10123), .B(n10079), .Z(n10081) );
  IV U10101 ( .A(n9996), .Z(n10123) );
  XOR U10102 ( .A(n10124), .B(n10073), .Z(n9996) );
  XOR U10103 ( .A(n10066), .B(n10065), .Z(n10073) );
  XNOR U10104 ( .A(n10125), .B(n10062), .Z(n10065) );
  XOR U10105 ( .A(n10126), .B(n10127), .Z(n10062) );
  AND U10106 ( .A(n10128), .B(n10129), .Z(n10127) );
  XNOR U10107 ( .A(n10130), .B(n10131), .Z(n10128) );
  IV U10108 ( .A(n10126), .Z(n10130) );
  XNOR U10109 ( .A(n10132), .B(n10133), .Z(n10125) );
  NOR U10110 ( .A(n10134), .B(n10135), .Z(n10133) );
  XNOR U10111 ( .A(n10132), .B(n10136), .Z(n10134) );
  XOR U10112 ( .A(n10137), .B(n10138), .Z(n10066) );
  AND U10113 ( .A(n10139), .B(n10140), .Z(n10138) );
  XOR U10114 ( .A(n10137), .B(n10141), .Z(n10139) );
  XNOR U10115 ( .A(n10072), .B(n10067), .Z(n10124) );
  AND U10116 ( .A(n10008), .B(n10142), .Z(n10067) );
  XOR U10117 ( .A(n10143), .B(n10078), .Z(n10072) );
  XNOR U10118 ( .A(n10144), .B(n10145), .Z(n10078) );
  NOR U10119 ( .A(n10146), .B(n10147), .Z(n10145) );
  XNOR U10120 ( .A(n10144), .B(n10148), .Z(n10146) );
  XNOR U10121 ( .A(n10077), .B(n10069), .Z(n10143) );
  XOR U10122 ( .A(n10149), .B(n10150), .Z(n10069) );
  AND U10123 ( .A(n10151), .B(n10152), .Z(n10150) );
  XOR U10124 ( .A(n10149), .B(n10153), .Z(n10151) );
  XNOR U10125 ( .A(n10154), .B(n10074), .Z(n10077) );
  XOR U10126 ( .A(n10155), .B(n10156), .Z(n10074) );
  AND U10127 ( .A(n10157), .B(n10158), .Z(n10156) );
  XOR U10128 ( .A(n10155), .B(n10159), .Z(n10157) );
  XNOR U10129 ( .A(n10160), .B(n10161), .Z(n10154) );
  NOR U10130 ( .A(n10162), .B(n10163), .Z(n10161) );
  XOR U10131 ( .A(n10160), .B(n10164), .Z(n10162) );
  AND U10132 ( .A(n10008), .B(n10011), .Z(n10079) );
  XOR U10133 ( .A(n10165), .B(n10106), .Z(n10011) );
  XNOR U10134 ( .A(p_input[1024]), .B(p_input[992]), .Z(n10106) );
  XNOR U10135 ( .A(n10094), .B(n10093), .Z(n10165) );
  XNOR U10136 ( .A(n10166), .B(n10100), .Z(n10093) );
  XNOR U10137 ( .A(n10089), .B(n10088), .Z(n10100) );
  XOR U10138 ( .A(n10167), .B(n10085), .Z(n10088) );
  XOR U10139 ( .A(p_input[1002]), .B(p_input[1034]), .Z(n10085) );
  XNOR U10140 ( .A(p_input[1003]), .B(p_input[1035]), .Z(n10167) );
  XOR U10141 ( .A(p_input[1004]), .B(p_input[1036]), .Z(n10089) );
  XOR U10142 ( .A(n10099), .B(n10090), .Z(n10166) );
  XNOR U10143 ( .A(n3298), .B(p_input[993]), .Z(n10090) );
  IV U10144 ( .A(p_input[1025]), .Z(n3298) );
  XOR U10145 ( .A(n10168), .B(n10105), .Z(n10099) );
  XOR U10146 ( .A(p_input[1007]), .B(p_input[1039]), .Z(n10105) );
  XOR U10147 ( .A(n10096), .B(n10104), .Z(n10168) );
  XOR U10148 ( .A(n10169), .B(n10101), .Z(n10104) );
  XOR U10149 ( .A(p_input[1005]), .B(p_input[1037]), .Z(n10101) );
  XNOR U10150 ( .A(p_input[1006]), .B(p_input[1038]), .Z(n10169) );
  XOR U10151 ( .A(p_input[1001]), .B(p_input[1033]), .Z(n10096) );
  XNOR U10152 ( .A(n10112), .B(n10111), .Z(n10094) );
  XOR U10153 ( .A(n10170), .B(n10117), .Z(n10111) );
  XOR U10154 ( .A(p_input[1000]), .B(p_input[1032]), .Z(n10117) );
  XOR U10155 ( .A(n10108), .B(n10116), .Z(n10170) );
  XOR U10156 ( .A(n10171), .B(n10113), .Z(n10116) );
  XOR U10157 ( .A(p_input[1030]), .B(p_input[998]), .Z(n10113) );
  XNOR U10158 ( .A(p_input[1031]), .B(p_input[999]), .Z(n10171) );
  XOR U10159 ( .A(p_input[1026]), .B(p_input[994]), .Z(n10108) );
  XNOR U10160 ( .A(n10122), .B(n10121), .Z(n10112) );
  XOR U10161 ( .A(n10172), .B(n10118), .Z(n10121) );
  XOR U10162 ( .A(p_input[1027]), .B(p_input[995]), .Z(n10118) );
  XNOR U10163 ( .A(p_input[1028]), .B(p_input[996]), .Z(n10172) );
  XOR U10164 ( .A(p_input[1029]), .B(p_input[997]), .Z(n10122) );
  XOR U10165 ( .A(n10173), .B(n10153), .Z(n10008) );
  XOR U10166 ( .A(n10131), .B(n10129), .Z(n10153) );
  XNOR U10167 ( .A(n10174), .B(n10136), .Z(n10129) );
  XOR U10168 ( .A(\knn_comb_/min_val_out[0][8] ), .B(p_input[1032]), .Z(n10136) );
  XOR U10169 ( .A(n10126), .B(n10135), .Z(n10174) );
  XOR U10170 ( .A(n10175), .B(n10132), .Z(n10135) );
  XOR U10171 ( .A(\knn_comb_/min_val_out[0][6] ), .B(p_input[1030]), .Z(n10132) );
  XNOR U10172 ( .A(\knn_comb_/min_val_out[0][7] ), .B(p_input[1031]), .Z(
        n10175) );
  XOR U10173 ( .A(\knn_comb_/min_val_out[0][2] ), .B(p_input[1026]), .Z(n10126) );
  XOR U10174 ( .A(n10141), .B(n10140), .Z(n10131) );
  XNOR U10175 ( .A(n10176), .B(n10137), .Z(n10140) );
  XOR U10176 ( .A(\knn_comb_/min_val_out[0][3] ), .B(p_input[1027]), .Z(n10137) );
  XOR U10177 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n3864), .Z(n10176) );
  IV U10178 ( .A(p_input[1028]), .Z(n3864) );
  XOR U10179 ( .A(\knn_comb_/min_val_out[0][5] ), .B(p_input[1029]), .Z(n10141) );
  XNOR U10180 ( .A(n10152), .B(n10142), .Z(n10173) );
  XOR U10181 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[1024]), .Z(n10142) );
  XNOR U10182 ( .A(n10177), .B(n10159), .Z(n10152) );
  XNOR U10183 ( .A(n10148), .B(n10147), .Z(n10159) );
  XOR U10184 ( .A(n10178), .B(n10144), .Z(n10147) );
  XOR U10185 ( .A(\knn_comb_/min_val_out[0][10] ), .B(p_input[1034]), .Z(
        n10144) );
  XNOR U10186 ( .A(\knn_comb_/min_val_out[0][11] ), .B(p_input[1035]), .Z(
        n10178) );
  XOR U10187 ( .A(\knn_comb_/min_val_out[0][12] ), .B(p_input[1036]), .Z(
        n10148) );
  XNOR U10188 ( .A(n10158), .B(n10149), .Z(n10177) );
  XOR U10189 ( .A(\knn_comb_/min_val_out[0][1] ), .B(p_input[1025]), .Z(n10149) );
  XOR U10190 ( .A(n10179), .B(n10164), .Z(n10158) );
  XNOR U10191 ( .A(\knn_comb_/min_val_out[0][15] ), .B(p_input[1039]), .Z(
        n10164) );
  XOR U10192 ( .A(n10155), .B(n10163), .Z(n10179) );
  XOR U10193 ( .A(n10180), .B(n10160), .Z(n10163) );
  XOR U10194 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[1037]), .Z(
        n10160) );
  XNOR U10195 ( .A(\knn_comb_/min_val_out[0][14] ), .B(p_input[1038]), .Z(
        n10180) );
  XOR U10196 ( .A(\knn_comb_/min_val_out[0][9] ), .B(p_input[1033]), .Z(n10155) );
endmodule

