
module psi_BMR_b1000_n10 ( p_input, o );
  input [9999:0] p_input;
  output [999:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000;

  AND U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(n3), .B(n4), .Z(n2) );
  AND U3 ( .A(n5), .B(p_input[3009]), .Z(n4) );
  AND U4 ( .A(p_input[2009]), .B(p_input[1009]), .Z(n5) );
  AND U5 ( .A(p_input[5009]), .B(p_input[4009]), .Z(n3) );
  AND U6 ( .A(n6), .B(n7), .Z(n1) );
  AND U7 ( .A(n8), .B(p_input[8009]), .Z(n7) );
  AND U8 ( .A(p_input[7009]), .B(p_input[6009]), .Z(n8) );
  AND U9 ( .A(p_input[9]), .B(p_input[9009]), .Z(n6) );
  AND U10 ( .A(n9), .B(n10), .Z(o[99]) );
  AND U11 ( .A(n11), .B(n12), .Z(n10) );
  AND U12 ( .A(n13), .B(p_input[3099]), .Z(n12) );
  AND U13 ( .A(p_input[2099]), .B(p_input[1099]), .Z(n13) );
  AND U14 ( .A(p_input[5099]), .B(p_input[4099]), .Z(n11) );
  AND U15 ( .A(n14), .B(n15), .Z(n9) );
  AND U16 ( .A(n16), .B(p_input[8099]), .Z(n15) );
  AND U17 ( .A(p_input[7099]), .B(p_input[6099]), .Z(n16) );
  AND U18 ( .A(p_input[99]), .B(p_input[9099]), .Z(n14) );
  AND U19 ( .A(n17), .B(n18), .Z(o[999]) );
  AND U20 ( .A(n19), .B(n20), .Z(n18) );
  AND U21 ( .A(n21), .B(p_input[3999]), .Z(n20) );
  AND U22 ( .A(p_input[2999]), .B(p_input[1999]), .Z(n21) );
  AND U23 ( .A(p_input[5999]), .B(p_input[4999]), .Z(n19) );
  AND U24 ( .A(n22), .B(n23), .Z(n17) );
  AND U25 ( .A(n24), .B(p_input[8999]), .Z(n23) );
  AND U26 ( .A(p_input[7999]), .B(p_input[6999]), .Z(n24) );
  AND U27 ( .A(p_input[999]), .B(p_input[9999]), .Z(n22) );
  AND U28 ( .A(n25), .B(n26), .Z(o[998]) );
  AND U29 ( .A(n27), .B(n28), .Z(n26) );
  AND U30 ( .A(n29), .B(p_input[3998]), .Z(n28) );
  AND U31 ( .A(p_input[2998]), .B(p_input[1998]), .Z(n29) );
  AND U32 ( .A(p_input[5998]), .B(p_input[4998]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n25) );
  AND U34 ( .A(n32), .B(p_input[8998]), .Z(n31) );
  AND U35 ( .A(p_input[7998]), .B(p_input[6998]), .Z(n32) );
  AND U36 ( .A(p_input[9998]), .B(p_input[998]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(o[997]) );
  AND U38 ( .A(n35), .B(n36), .Z(n34) );
  AND U39 ( .A(n37), .B(p_input[3997]), .Z(n36) );
  AND U40 ( .A(p_input[2997]), .B(p_input[1997]), .Z(n37) );
  AND U41 ( .A(p_input[5997]), .B(p_input[4997]), .Z(n35) );
  AND U42 ( .A(n38), .B(n39), .Z(n33) );
  AND U43 ( .A(n40), .B(p_input[8997]), .Z(n39) );
  AND U44 ( .A(p_input[7997]), .B(p_input[6997]), .Z(n40) );
  AND U45 ( .A(p_input[9997]), .B(p_input[997]), .Z(n38) );
  AND U46 ( .A(n41), .B(n42), .Z(o[996]) );
  AND U47 ( .A(n43), .B(n44), .Z(n42) );
  AND U48 ( .A(n45), .B(p_input[3996]), .Z(n44) );
  AND U49 ( .A(p_input[2996]), .B(p_input[1996]), .Z(n45) );
  AND U50 ( .A(p_input[5996]), .B(p_input[4996]), .Z(n43) );
  AND U51 ( .A(n46), .B(n47), .Z(n41) );
  AND U52 ( .A(n48), .B(p_input[8996]), .Z(n47) );
  AND U53 ( .A(p_input[7996]), .B(p_input[6996]), .Z(n48) );
  AND U54 ( .A(p_input[9996]), .B(p_input[996]), .Z(n46) );
  AND U55 ( .A(n49), .B(n50), .Z(o[995]) );
  AND U56 ( .A(n51), .B(n52), .Z(n50) );
  AND U57 ( .A(n53), .B(p_input[3995]), .Z(n52) );
  AND U58 ( .A(p_input[2995]), .B(p_input[1995]), .Z(n53) );
  AND U59 ( .A(p_input[5995]), .B(p_input[4995]), .Z(n51) );
  AND U60 ( .A(n54), .B(n55), .Z(n49) );
  AND U61 ( .A(n56), .B(p_input[8995]), .Z(n55) );
  AND U62 ( .A(p_input[7995]), .B(p_input[6995]), .Z(n56) );
  AND U63 ( .A(p_input[9995]), .B(p_input[995]), .Z(n54) );
  AND U64 ( .A(n57), .B(n58), .Z(o[994]) );
  AND U65 ( .A(n59), .B(n60), .Z(n58) );
  AND U66 ( .A(n61), .B(p_input[3994]), .Z(n60) );
  AND U67 ( .A(p_input[2994]), .B(p_input[1994]), .Z(n61) );
  AND U68 ( .A(p_input[5994]), .B(p_input[4994]), .Z(n59) );
  AND U69 ( .A(n62), .B(n63), .Z(n57) );
  AND U70 ( .A(n64), .B(p_input[8994]), .Z(n63) );
  AND U71 ( .A(p_input[7994]), .B(p_input[6994]), .Z(n64) );
  AND U72 ( .A(p_input[9994]), .B(p_input[994]), .Z(n62) );
  AND U73 ( .A(n65), .B(n66), .Z(o[993]) );
  AND U74 ( .A(n67), .B(n68), .Z(n66) );
  AND U75 ( .A(n69), .B(p_input[3993]), .Z(n68) );
  AND U76 ( .A(p_input[2993]), .B(p_input[1993]), .Z(n69) );
  AND U77 ( .A(p_input[5993]), .B(p_input[4993]), .Z(n67) );
  AND U78 ( .A(n70), .B(n71), .Z(n65) );
  AND U79 ( .A(n72), .B(p_input[8993]), .Z(n71) );
  AND U80 ( .A(p_input[7993]), .B(p_input[6993]), .Z(n72) );
  AND U81 ( .A(p_input[9993]), .B(p_input[993]), .Z(n70) );
  AND U82 ( .A(n73), .B(n74), .Z(o[992]) );
  AND U83 ( .A(n75), .B(n76), .Z(n74) );
  AND U84 ( .A(n77), .B(p_input[3992]), .Z(n76) );
  AND U85 ( .A(p_input[2992]), .B(p_input[1992]), .Z(n77) );
  AND U86 ( .A(p_input[5992]), .B(p_input[4992]), .Z(n75) );
  AND U87 ( .A(n78), .B(n79), .Z(n73) );
  AND U88 ( .A(n80), .B(p_input[8992]), .Z(n79) );
  AND U89 ( .A(p_input[7992]), .B(p_input[6992]), .Z(n80) );
  AND U90 ( .A(p_input[9992]), .B(p_input[992]), .Z(n78) );
  AND U91 ( .A(n81), .B(n82), .Z(o[991]) );
  AND U92 ( .A(n83), .B(n84), .Z(n82) );
  AND U93 ( .A(n85), .B(p_input[3991]), .Z(n84) );
  AND U94 ( .A(p_input[2991]), .B(p_input[1991]), .Z(n85) );
  AND U95 ( .A(p_input[5991]), .B(p_input[4991]), .Z(n83) );
  AND U96 ( .A(n86), .B(n87), .Z(n81) );
  AND U97 ( .A(n88), .B(p_input[8991]), .Z(n87) );
  AND U98 ( .A(p_input[7991]), .B(p_input[6991]), .Z(n88) );
  AND U99 ( .A(p_input[9991]), .B(p_input[991]), .Z(n86) );
  AND U100 ( .A(n89), .B(n90), .Z(o[990]) );
  AND U101 ( .A(n91), .B(n92), .Z(n90) );
  AND U102 ( .A(n93), .B(p_input[3990]), .Z(n92) );
  AND U103 ( .A(p_input[2990]), .B(p_input[1990]), .Z(n93) );
  AND U104 ( .A(p_input[5990]), .B(p_input[4990]), .Z(n91) );
  AND U105 ( .A(n94), .B(n95), .Z(n89) );
  AND U106 ( .A(n96), .B(p_input[8990]), .Z(n95) );
  AND U107 ( .A(p_input[7990]), .B(p_input[6990]), .Z(n96) );
  AND U108 ( .A(p_input[9990]), .B(p_input[990]), .Z(n94) );
  AND U109 ( .A(n97), .B(n98), .Z(o[98]) );
  AND U110 ( .A(n99), .B(n100), .Z(n98) );
  AND U111 ( .A(n101), .B(p_input[3098]), .Z(n100) );
  AND U112 ( .A(p_input[2098]), .B(p_input[1098]), .Z(n101) );
  AND U113 ( .A(p_input[5098]), .B(p_input[4098]), .Z(n99) );
  AND U114 ( .A(n102), .B(n103), .Z(n97) );
  AND U115 ( .A(n104), .B(p_input[8098]), .Z(n103) );
  AND U116 ( .A(p_input[7098]), .B(p_input[6098]), .Z(n104) );
  AND U117 ( .A(p_input[98]), .B(p_input[9098]), .Z(n102) );
  AND U118 ( .A(n105), .B(n106), .Z(o[989]) );
  AND U119 ( .A(n107), .B(n108), .Z(n106) );
  AND U120 ( .A(n109), .B(p_input[3989]), .Z(n108) );
  AND U121 ( .A(p_input[2989]), .B(p_input[1989]), .Z(n109) );
  AND U122 ( .A(p_input[5989]), .B(p_input[4989]), .Z(n107) );
  AND U123 ( .A(n110), .B(n111), .Z(n105) );
  AND U124 ( .A(n112), .B(p_input[8989]), .Z(n111) );
  AND U125 ( .A(p_input[7989]), .B(p_input[6989]), .Z(n112) );
  AND U126 ( .A(p_input[9989]), .B(p_input[989]), .Z(n110) );
  AND U127 ( .A(n113), .B(n114), .Z(o[988]) );
  AND U128 ( .A(n115), .B(n116), .Z(n114) );
  AND U129 ( .A(n117), .B(p_input[3988]), .Z(n116) );
  AND U130 ( .A(p_input[2988]), .B(p_input[1988]), .Z(n117) );
  AND U131 ( .A(p_input[5988]), .B(p_input[4988]), .Z(n115) );
  AND U132 ( .A(n118), .B(n119), .Z(n113) );
  AND U133 ( .A(n120), .B(p_input[8988]), .Z(n119) );
  AND U134 ( .A(p_input[7988]), .B(p_input[6988]), .Z(n120) );
  AND U135 ( .A(p_input[9988]), .B(p_input[988]), .Z(n118) );
  AND U136 ( .A(n121), .B(n122), .Z(o[987]) );
  AND U137 ( .A(n123), .B(n124), .Z(n122) );
  AND U138 ( .A(n125), .B(p_input[3987]), .Z(n124) );
  AND U139 ( .A(p_input[2987]), .B(p_input[1987]), .Z(n125) );
  AND U140 ( .A(p_input[5987]), .B(p_input[4987]), .Z(n123) );
  AND U141 ( .A(n126), .B(n127), .Z(n121) );
  AND U142 ( .A(n128), .B(p_input[8987]), .Z(n127) );
  AND U143 ( .A(p_input[7987]), .B(p_input[6987]), .Z(n128) );
  AND U144 ( .A(p_input[9987]), .B(p_input[987]), .Z(n126) );
  AND U145 ( .A(n129), .B(n130), .Z(o[986]) );
  AND U146 ( .A(n131), .B(n132), .Z(n130) );
  AND U147 ( .A(n133), .B(p_input[3986]), .Z(n132) );
  AND U148 ( .A(p_input[2986]), .B(p_input[1986]), .Z(n133) );
  AND U149 ( .A(p_input[5986]), .B(p_input[4986]), .Z(n131) );
  AND U150 ( .A(n134), .B(n135), .Z(n129) );
  AND U151 ( .A(n136), .B(p_input[8986]), .Z(n135) );
  AND U152 ( .A(p_input[7986]), .B(p_input[6986]), .Z(n136) );
  AND U153 ( .A(p_input[9986]), .B(p_input[986]), .Z(n134) );
  AND U154 ( .A(n137), .B(n138), .Z(o[985]) );
  AND U155 ( .A(n139), .B(n140), .Z(n138) );
  AND U156 ( .A(n141), .B(p_input[3985]), .Z(n140) );
  AND U157 ( .A(p_input[2985]), .B(p_input[1985]), .Z(n141) );
  AND U158 ( .A(p_input[5985]), .B(p_input[4985]), .Z(n139) );
  AND U159 ( .A(n142), .B(n143), .Z(n137) );
  AND U160 ( .A(n144), .B(p_input[8985]), .Z(n143) );
  AND U161 ( .A(p_input[7985]), .B(p_input[6985]), .Z(n144) );
  AND U162 ( .A(p_input[9985]), .B(p_input[985]), .Z(n142) );
  AND U163 ( .A(n145), .B(n146), .Z(o[984]) );
  AND U164 ( .A(n147), .B(n148), .Z(n146) );
  AND U165 ( .A(n149), .B(p_input[3984]), .Z(n148) );
  AND U166 ( .A(p_input[2984]), .B(p_input[1984]), .Z(n149) );
  AND U167 ( .A(p_input[5984]), .B(p_input[4984]), .Z(n147) );
  AND U168 ( .A(n150), .B(n151), .Z(n145) );
  AND U169 ( .A(n152), .B(p_input[8984]), .Z(n151) );
  AND U170 ( .A(p_input[7984]), .B(p_input[6984]), .Z(n152) );
  AND U171 ( .A(p_input[9984]), .B(p_input[984]), .Z(n150) );
  AND U172 ( .A(n153), .B(n154), .Z(o[983]) );
  AND U173 ( .A(n155), .B(n156), .Z(n154) );
  AND U174 ( .A(n157), .B(p_input[3983]), .Z(n156) );
  AND U175 ( .A(p_input[2983]), .B(p_input[1983]), .Z(n157) );
  AND U176 ( .A(p_input[5983]), .B(p_input[4983]), .Z(n155) );
  AND U177 ( .A(n158), .B(n159), .Z(n153) );
  AND U178 ( .A(n160), .B(p_input[8983]), .Z(n159) );
  AND U179 ( .A(p_input[7983]), .B(p_input[6983]), .Z(n160) );
  AND U180 ( .A(p_input[9983]), .B(p_input[983]), .Z(n158) );
  AND U181 ( .A(n161), .B(n162), .Z(o[982]) );
  AND U182 ( .A(n163), .B(n164), .Z(n162) );
  AND U183 ( .A(n165), .B(p_input[3982]), .Z(n164) );
  AND U184 ( .A(p_input[2982]), .B(p_input[1982]), .Z(n165) );
  AND U185 ( .A(p_input[5982]), .B(p_input[4982]), .Z(n163) );
  AND U186 ( .A(n166), .B(n167), .Z(n161) );
  AND U187 ( .A(n168), .B(p_input[8982]), .Z(n167) );
  AND U188 ( .A(p_input[7982]), .B(p_input[6982]), .Z(n168) );
  AND U189 ( .A(p_input[9982]), .B(p_input[982]), .Z(n166) );
  AND U190 ( .A(n169), .B(n170), .Z(o[981]) );
  AND U191 ( .A(n171), .B(n172), .Z(n170) );
  AND U192 ( .A(n173), .B(p_input[3981]), .Z(n172) );
  AND U193 ( .A(p_input[2981]), .B(p_input[1981]), .Z(n173) );
  AND U194 ( .A(p_input[5981]), .B(p_input[4981]), .Z(n171) );
  AND U195 ( .A(n174), .B(n175), .Z(n169) );
  AND U196 ( .A(n176), .B(p_input[8981]), .Z(n175) );
  AND U197 ( .A(p_input[7981]), .B(p_input[6981]), .Z(n176) );
  AND U198 ( .A(p_input[9981]), .B(p_input[981]), .Z(n174) );
  AND U199 ( .A(n177), .B(n178), .Z(o[980]) );
  AND U200 ( .A(n179), .B(n180), .Z(n178) );
  AND U201 ( .A(n181), .B(p_input[3980]), .Z(n180) );
  AND U202 ( .A(p_input[2980]), .B(p_input[1980]), .Z(n181) );
  AND U203 ( .A(p_input[5980]), .B(p_input[4980]), .Z(n179) );
  AND U204 ( .A(n182), .B(n183), .Z(n177) );
  AND U205 ( .A(n184), .B(p_input[8980]), .Z(n183) );
  AND U206 ( .A(p_input[7980]), .B(p_input[6980]), .Z(n184) );
  AND U207 ( .A(p_input[9980]), .B(p_input[980]), .Z(n182) );
  AND U208 ( .A(n185), .B(n186), .Z(o[97]) );
  AND U209 ( .A(n187), .B(n188), .Z(n186) );
  AND U210 ( .A(n189), .B(p_input[3097]), .Z(n188) );
  AND U211 ( .A(p_input[2097]), .B(p_input[1097]), .Z(n189) );
  AND U212 ( .A(p_input[5097]), .B(p_input[4097]), .Z(n187) );
  AND U213 ( .A(n190), .B(n191), .Z(n185) );
  AND U214 ( .A(n192), .B(p_input[8097]), .Z(n191) );
  AND U215 ( .A(p_input[7097]), .B(p_input[6097]), .Z(n192) );
  AND U216 ( .A(p_input[97]), .B(p_input[9097]), .Z(n190) );
  AND U217 ( .A(n193), .B(n194), .Z(o[979]) );
  AND U218 ( .A(n195), .B(n196), .Z(n194) );
  AND U219 ( .A(n197), .B(p_input[3979]), .Z(n196) );
  AND U220 ( .A(p_input[2979]), .B(p_input[1979]), .Z(n197) );
  AND U221 ( .A(p_input[5979]), .B(p_input[4979]), .Z(n195) );
  AND U222 ( .A(n198), .B(n199), .Z(n193) );
  AND U223 ( .A(n200), .B(p_input[8979]), .Z(n199) );
  AND U224 ( .A(p_input[7979]), .B(p_input[6979]), .Z(n200) );
  AND U225 ( .A(p_input[9979]), .B(p_input[979]), .Z(n198) );
  AND U226 ( .A(n201), .B(n202), .Z(o[978]) );
  AND U227 ( .A(n203), .B(n204), .Z(n202) );
  AND U228 ( .A(n205), .B(p_input[3978]), .Z(n204) );
  AND U229 ( .A(p_input[2978]), .B(p_input[1978]), .Z(n205) );
  AND U230 ( .A(p_input[5978]), .B(p_input[4978]), .Z(n203) );
  AND U231 ( .A(n206), .B(n207), .Z(n201) );
  AND U232 ( .A(n208), .B(p_input[8978]), .Z(n207) );
  AND U233 ( .A(p_input[7978]), .B(p_input[6978]), .Z(n208) );
  AND U234 ( .A(p_input[9978]), .B(p_input[978]), .Z(n206) );
  AND U235 ( .A(n209), .B(n210), .Z(o[977]) );
  AND U236 ( .A(n211), .B(n212), .Z(n210) );
  AND U237 ( .A(n213), .B(p_input[3977]), .Z(n212) );
  AND U238 ( .A(p_input[2977]), .B(p_input[1977]), .Z(n213) );
  AND U239 ( .A(p_input[5977]), .B(p_input[4977]), .Z(n211) );
  AND U240 ( .A(n214), .B(n215), .Z(n209) );
  AND U241 ( .A(n216), .B(p_input[8977]), .Z(n215) );
  AND U242 ( .A(p_input[7977]), .B(p_input[6977]), .Z(n216) );
  AND U243 ( .A(p_input[9977]), .B(p_input[977]), .Z(n214) );
  AND U244 ( .A(n217), .B(n218), .Z(o[976]) );
  AND U245 ( .A(n219), .B(n220), .Z(n218) );
  AND U246 ( .A(n221), .B(p_input[3976]), .Z(n220) );
  AND U247 ( .A(p_input[2976]), .B(p_input[1976]), .Z(n221) );
  AND U248 ( .A(p_input[5976]), .B(p_input[4976]), .Z(n219) );
  AND U249 ( .A(n222), .B(n223), .Z(n217) );
  AND U250 ( .A(n224), .B(p_input[8976]), .Z(n223) );
  AND U251 ( .A(p_input[7976]), .B(p_input[6976]), .Z(n224) );
  AND U252 ( .A(p_input[9976]), .B(p_input[976]), .Z(n222) );
  AND U253 ( .A(n225), .B(n226), .Z(o[975]) );
  AND U254 ( .A(n227), .B(n228), .Z(n226) );
  AND U255 ( .A(n229), .B(p_input[3975]), .Z(n228) );
  AND U256 ( .A(p_input[2975]), .B(p_input[1975]), .Z(n229) );
  AND U257 ( .A(p_input[5975]), .B(p_input[4975]), .Z(n227) );
  AND U258 ( .A(n230), .B(n231), .Z(n225) );
  AND U259 ( .A(n232), .B(p_input[8975]), .Z(n231) );
  AND U260 ( .A(p_input[7975]), .B(p_input[6975]), .Z(n232) );
  AND U261 ( .A(p_input[9975]), .B(p_input[975]), .Z(n230) );
  AND U262 ( .A(n233), .B(n234), .Z(o[974]) );
  AND U263 ( .A(n235), .B(n236), .Z(n234) );
  AND U264 ( .A(n237), .B(p_input[3974]), .Z(n236) );
  AND U265 ( .A(p_input[2974]), .B(p_input[1974]), .Z(n237) );
  AND U266 ( .A(p_input[5974]), .B(p_input[4974]), .Z(n235) );
  AND U267 ( .A(n238), .B(n239), .Z(n233) );
  AND U268 ( .A(n240), .B(p_input[8974]), .Z(n239) );
  AND U269 ( .A(p_input[7974]), .B(p_input[6974]), .Z(n240) );
  AND U270 ( .A(p_input[9974]), .B(p_input[974]), .Z(n238) );
  AND U271 ( .A(n241), .B(n242), .Z(o[973]) );
  AND U272 ( .A(n243), .B(n244), .Z(n242) );
  AND U273 ( .A(n245), .B(p_input[3973]), .Z(n244) );
  AND U274 ( .A(p_input[2973]), .B(p_input[1973]), .Z(n245) );
  AND U275 ( .A(p_input[5973]), .B(p_input[4973]), .Z(n243) );
  AND U276 ( .A(n246), .B(n247), .Z(n241) );
  AND U277 ( .A(n248), .B(p_input[8973]), .Z(n247) );
  AND U278 ( .A(p_input[7973]), .B(p_input[6973]), .Z(n248) );
  AND U279 ( .A(p_input[9973]), .B(p_input[973]), .Z(n246) );
  AND U280 ( .A(n249), .B(n250), .Z(o[972]) );
  AND U281 ( .A(n251), .B(n252), .Z(n250) );
  AND U282 ( .A(n253), .B(p_input[3972]), .Z(n252) );
  AND U283 ( .A(p_input[2972]), .B(p_input[1972]), .Z(n253) );
  AND U284 ( .A(p_input[5972]), .B(p_input[4972]), .Z(n251) );
  AND U285 ( .A(n254), .B(n255), .Z(n249) );
  AND U286 ( .A(n256), .B(p_input[8972]), .Z(n255) );
  AND U287 ( .A(p_input[7972]), .B(p_input[6972]), .Z(n256) );
  AND U288 ( .A(p_input[9972]), .B(p_input[972]), .Z(n254) );
  AND U289 ( .A(n257), .B(n258), .Z(o[971]) );
  AND U290 ( .A(n259), .B(n260), .Z(n258) );
  AND U291 ( .A(n261), .B(p_input[3971]), .Z(n260) );
  AND U292 ( .A(p_input[2971]), .B(p_input[1971]), .Z(n261) );
  AND U293 ( .A(p_input[5971]), .B(p_input[4971]), .Z(n259) );
  AND U294 ( .A(n262), .B(n263), .Z(n257) );
  AND U295 ( .A(n264), .B(p_input[8971]), .Z(n263) );
  AND U296 ( .A(p_input[7971]), .B(p_input[6971]), .Z(n264) );
  AND U297 ( .A(p_input[9971]), .B(p_input[971]), .Z(n262) );
  AND U298 ( .A(n265), .B(n266), .Z(o[970]) );
  AND U299 ( .A(n267), .B(n268), .Z(n266) );
  AND U300 ( .A(n269), .B(p_input[3970]), .Z(n268) );
  AND U301 ( .A(p_input[2970]), .B(p_input[1970]), .Z(n269) );
  AND U302 ( .A(p_input[5970]), .B(p_input[4970]), .Z(n267) );
  AND U303 ( .A(n270), .B(n271), .Z(n265) );
  AND U304 ( .A(n272), .B(p_input[8970]), .Z(n271) );
  AND U305 ( .A(p_input[7970]), .B(p_input[6970]), .Z(n272) );
  AND U306 ( .A(p_input[9970]), .B(p_input[970]), .Z(n270) );
  AND U307 ( .A(n273), .B(n274), .Z(o[96]) );
  AND U308 ( .A(n275), .B(n276), .Z(n274) );
  AND U309 ( .A(n277), .B(p_input[3096]), .Z(n276) );
  AND U310 ( .A(p_input[2096]), .B(p_input[1096]), .Z(n277) );
  AND U311 ( .A(p_input[5096]), .B(p_input[4096]), .Z(n275) );
  AND U312 ( .A(n278), .B(n279), .Z(n273) );
  AND U313 ( .A(n280), .B(p_input[8096]), .Z(n279) );
  AND U314 ( .A(p_input[7096]), .B(p_input[6096]), .Z(n280) );
  AND U315 ( .A(p_input[96]), .B(p_input[9096]), .Z(n278) );
  AND U316 ( .A(n281), .B(n282), .Z(o[969]) );
  AND U317 ( .A(n283), .B(n284), .Z(n282) );
  AND U318 ( .A(n285), .B(p_input[3969]), .Z(n284) );
  AND U319 ( .A(p_input[2969]), .B(p_input[1969]), .Z(n285) );
  AND U320 ( .A(p_input[5969]), .B(p_input[4969]), .Z(n283) );
  AND U321 ( .A(n286), .B(n287), .Z(n281) );
  AND U322 ( .A(n288), .B(p_input[8969]), .Z(n287) );
  AND U323 ( .A(p_input[7969]), .B(p_input[6969]), .Z(n288) );
  AND U324 ( .A(p_input[9969]), .B(p_input[969]), .Z(n286) );
  AND U325 ( .A(n289), .B(n290), .Z(o[968]) );
  AND U326 ( .A(n291), .B(n292), .Z(n290) );
  AND U327 ( .A(n293), .B(p_input[3968]), .Z(n292) );
  AND U328 ( .A(p_input[2968]), .B(p_input[1968]), .Z(n293) );
  AND U329 ( .A(p_input[5968]), .B(p_input[4968]), .Z(n291) );
  AND U330 ( .A(n294), .B(n295), .Z(n289) );
  AND U331 ( .A(n296), .B(p_input[8968]), .Z(n295) );
  AND U332 ( .A(p_input[7968]), .B(p_input[6968]), .Z(n296) );
  AND U333 ( .A(p_input[9968]), .B(p_input[968]), .Z(n294) );
  AND U334 ( .A(n297), .B(n298), .Z(o[967]) );
  AND U335 ( .A(n299), .B(n300), .Z(n298) );
  AND U336 ( .A(n301), .B(p_input[3967]), .Z(n300) );
  AND U337 ( .A(p_input[2967]), .B(p_input[1967]), .Z(n301) );
  AND U338 ( .A(p_input[5967]), .B(p_input[4967]), .Z(n299) );
  AND U339 ( .A(n302), .B(n303), .Z(n297) );
  AND U340 ( .A(n304), .B(p_input[8967]), .Z(n303) );
  AND U341 ( .A(p_input[7967]), .B(p_input[6967]), .Z(n304) );
  AND U342 ( .A(p_input[9967]), .B(p_input[967]), .Z(n302) );
  AND U343 ( .A(n305), .B(n306), .Z(o[966]) );
  AND U344 ( .A(n307), .B(n308), .Z(n306) );
  AND U345 ( .A(n309), .B(p_input[3966]), .Z(n308) );
  AND U346 ( .A(p_input[2966]), .B(p_input[1966]), .Z(n309) );
  AND U347 ( .A(p_input[5966]), .B(p_input[4966]), .Z(n307) );
  AND U348 ( .A(n310), .B(n311), .Z(n305) );
  AND U349 ( .A(n312), .B(p_input[8966]), .Z(n311) );
  AND U350 ( .A(p_input[7966]), .B(p_input[6966]), .Z(n312) );
  AND U351 ( .A(p_input[9966]), .B(p_input[966]), .Z(n310) );
  AND U352 ( .A(n313), .B(n314), .Z(o[965]) );
  AND U353 ( .A(n315), .B(n316), .Z(n314) );
  AND U354 ( .A(n317), .B(p_input[3965]), .Z(n316) );
  AND U355 ( .A(p_input[2965]), .B(p_input[1965]), .Z(n317) );
  AND U356 ( .A(p_input[5965]), .B(p_input[4965]), .Z(n315) );
  AND U357 ( .A(n318), .B(n319), .Z(n313) );
  AND U358 ( .A(n320), .B(p_input[8965]), .Z(n319) );
  AND U359 ( .A(p_input[7965]), .B(p_input[6965]), .Z(n320) );
  AND U360 ( .A(p_input[9965]), .B(p_input[965]), .Z(n318) );
  AND U361 ( .A(n321), .B(n322), .Z(o[964]) );
  AND U362 ( .A(n323), .B(n324), .Z(n322) );
  AND U363 ( .A(n325), .B(p_input[3964]), .Z(n324) );
  AND U364 ( .A(p_input[2964]), .B(p_input[1964]), .Z(n325) );
  AND U365 ( .A(p_input[5964]), .B(p_input[4964]), .Z(n323) );
  AND U366 ( .A(n326), .B(n327), .Z(n321) );
  AND U367 ( .A(n328), .B(p_input[8964]), .Z(n327) );
  AND U368 ( .A(p_input[7964]), .B(p_input[6964]), .Z(n328) );
  AND U369 ( .A(p_input[9964]), .B(p_input[964]), .Z(n326) );
  AND U370 ( .A(n329), .B(n330), .Z(o[963]) );
  AND U371 ( .A(n331), .B(n332), .Z(n330) );
  AND U372 ( .A(n333), .B(p_input[3963]), .Z(n332) );
  AND U373 ( .A(p_input[2963]), .B(p_input[1963]), .Z(n333) );
  AND U374 ( .A(p_input[5963]), .B(p_input[4963]), .Z(n331) );
  AND U375 ( .A(n334), .B(n335), .Z(n329) );
  AND U376 ( .A(n336), .B(p_input[8963]), .Z(n335) );
  AND U377 ( .A(p_input[7963]), .B(p_input[6963]), .Z(n336) );
  AND U378 ( .A(p_input[9963]), .B(p_input[963]), .Z(n334) );
  AND U379 ( .A(n337), .B(n338), .Z(o[962]) );
  AND U380 ( .A(n339), .B(n340), .Z(n338) );
  AND U381 ( .A(n341), .B(p_input[3962]), .Z(n340) );
  AND U382 ( .A(p_input[2962]), .B(p_input[1962]), .Z(n341) );
  AND U383 ( .A(p_input[5962]), .B(p_input[4962]), .Z(n339) );
  AND U384 ( .A(n342), .B(n343), .Z(n337) );
  AND U385 ( .A(n344), .B(p_input[8962]), .Z(n343) );
  AND U386 ( .A(p_input[7962]), .B(p_input[6962]), .Z(n344) );
  AND U387 ( .A(p_input[9962]), .B(p_input[962]), .Z(n342) );
  AND U388 ( .A(n345), .B(n346), .Z(o[961]) );
  AND U389 ( .A(n347), .B(n348), .Z(n346) );
  AND U390 ( .A(n349), .B(p_input[3961]), .Z(n348) );
  AND U391 ( .A(p_input[2961]), .B(p_input[1961]), .Z(n349) );
  AND U392 ( .A(p_input[5961]), .B(p_input[4961]), .Z(n347) );
  AND U393 ( .A(n350), .B(n351), .Z(n345) );
  AND U394 ( .A(n352), .B(p_input[8961]), .Z(n351) );
  AND U395 ( .A(p_input[7961]), .B(p_input[6961]), .Z(n352) );
  AND U396 ( .A(p_input[9961]), .B(p_input[961]), .Z(n350) );
  AND U397 ( .A(n353), .B(n354), .Z(o[960]) );
  AND U398 ( .A(n355), .B(n356), .Z(n354) );
  AND U399 ( .A(n357), .B(p_input[3960]), .Z(n356) );
  AND U400 ( .A(p_input[2960]), .B(p_input[1960]), .Z(n357) );
  AND U401 ( .A(p_input[5960]), .B(p_input[4960]), .Z(n355) );
  AND U402 ( .A(n358), .B(n359), .Z(n353) );
  AND U403 ( .A(n360), .B(p_input[8960]), .Z(n359) );
  AND U404 ( .A(p_input[7960]), .B(p_input[6960]), .Z(n360) );
  AND U405 ( .A(p_input[9960]), .B(p_input[960]), .Z(n358) );
  AND U406 ( .A(n361), .B(n362), .Z(o[95]) );
  AND U407 ( .A(n363), .B(n364), .Z(n362) );
  AND U408 ( .A(n365), .B(p_input[3095]), .Z(n364) );
  AND U409 ( .A(p_input[2095]), .B(p_input[1095]), .Z(n365) );
  AND U410 ( .A(p_input[5095]), .B(p_input[4095]), .Z(n363) );
  AND U411 ( .A(n366), .B(n367), .Z(n361) );
  AND U412 ( .A(n368), .B(p_input[8095]), .Z(n367) );
  AND U413 ( .A(p_input[7095]), .B(p_input[6095]), .Z(n368) );
  AND U414 ( .A(p_input[95]), .B(p_input[9095]), .Z(n366) );
  AND U415 ( .A(n369), .B(n370), .Z(o[959]) );
  AND U416 ( .A(n371), .B(n372), .Z(n370) );
  AND U417 ( .A(n373), .B(p_input[3959]), .Z(n372) );
  AND U418 ( .A(p_input[2959]), .B(p_input[1959]), .Z(n373) );
  AND U419 ( .A(p_input[5959]), .B(p_input[4959]), .Z(n371) );
  AND U420 ( .A(n374), .B(n375), .Z(n369) );
  AND U421 ( .A(n376), .B(p_input[8959]), .Z(n375) );
  AND U422 ( .A(p_input[7959]), .B(p_input[6959]), .Z(n376) );
  AND U423 ( .A(p_input[9959]), .B(p_input[959]), .Z(n374) );
  AND U424 ( .A(n377), .B(n378), .Z(o[958]) );
  AND U425 ( .A(n379), .B(n380), .Z(n378) );
  AND U426 ( .A(n381), .B(p_input[3958]), .Z(n380) );
  AND U427 ( .A(p_input[2958]), .B(p_input[1958]), .Z(n381) );
  AND U428 ( .A(p_input[5958]), .B(p_input[4958]), .Z(n379) );
  AND U429 ( .A(n382), .B(n383), .Z(n377) );
  AND U430 ( .A(n384), .B(p_input[8958]), .Z(n383) );
  AND U431 ( .A(p_input[7958]), .B(p_input[6958]), .Z(n384) );
  AND U432 ( .A(p_input[9958]), .B(p_input[958]), .Z(n382) );
  AND U433 ( .A(n385), .B(n386), .Z(o[957]) );
  AND U434 ( .A(n387), .B(n388), .Z(n386) );
  AND U435 ( .A(n389), .B(p_input[3957]), .Z(n388) );
  AND U436 ( .A(p_input[2957]), .B(p_input[1957]), .Z(n389) );
  AND U437 ( .A(p_input[5957]), .B(p_input[4957]), .Z(n387) );
  AND U438 ( .A(n390), .B(n391), .Z(n385) );
  AND U439 ( .A(n392), .B(p_input[8957]), .Z(n391) );
  AND U440 ( .A(p_input[7957]), .B(p_input[6957]), .Z(n392) );
  AND U441 ( .A(p_input[9957]), .B(p_input[957]), .Z(n390) );
  AND U442 ( .A(n393), .B(n394), .Z(o[956]) );
  AND U443 ( .A(n395), .B(n396), .Z(n394) );
  AND U444 ( .A(n397), .B(p_input[3956]), .Z(n396) );
  AND U445 ( .A(p_input[2956]), .B(p_input[1956]), .Z(n397) );
  AND U446 ( .A(p_input[5956]), .B(p_input[4956]), .Z(n395) );
  AND U447 ( .A(n398), .B(n399), .Z(n393) );
  AND U448 ( .A(n400), .B(p_input[8956]), .Z(n399) );
  AND U449 ( .A(p_input[7956]), .B(p_input[6956]), .Z(n400) );
  AND U450 ( .A(p_input[9956]), .B(p_input[956]), .Z(n398) );
  AND U451 ( .A(n401), .B(n402), .Z(o[955]) );
  AND U452 ( .A(n403), .B(n404), .Z(n402) );
  AND U453 ( .A(n405), .B(p_input[3955]), .Z(n404) );
  AND U454 ( .A(p_input[2955]), .B(p_input[1955]), .Z(n405) );
  AND U455 ( .A(p_input[5955]), .B(p_input[4955]), .Z(n403) );
  AND U456 ( .A(n406), .B(n407), .Z(n401) );
  AND U457 ( .A(n408), .B(p_input[8955]), .Z(n407) );
  AND U458 ( .A(p_input[7955]), .B(p_input[6955]), .Z(n408) );
  AND U459 ( .A(p_input[9955]), .B(p_input[955]), .Z(n406) );
  AND U460 ( .A(n409), .B(n410), .Z(o[954]) );
  AND U461 ( .A(n411), .B(n412), .Z(n410) );
  AND U462 ( .A(n413), .B(p_input[3954]), .Z(n412) );
  AND U463 ( .A(p_input[2954]), .B(p_input[1954]), .Z(n413) );
  AND U464 ( .A(p_input[5954]), .B(p_input[4954]), .Z(n411) );
  AND U465 ( .A(n414), .B(n415), .Z(n409) );
  AND U466 ( .A(n416), .B(p_input[8954]), .Z(n415) );
  AND U467 ( .A(p_input[7954]), .B(p_input[6954]), .Z(n416) );
  AND U468 ( .A(p_input[9954]), .B(p_input[954]), .Z(n414) );
  AND U469 ( .A(n417), .B(n418), .Z(o[953]) );
  AND U470 ( .A(n419), .B(n420), .Z(n418) );
  AND U471 ( .A(n421), .B(p_input[3953]), .Z(n420) );
  AND U472 ( .A(p_input[2953]), .B(p_input[1953]), .Z(n421) );
  AND U473 ( .A(p_input[5953]), .B(p_input[4953]), .Z(n419) );
  AND U474 ( .A(n422), .B(n423), .Z(n417) );
  AND U475 ( .A(n424), .B(p_input[8953]), .Z(n423) );
  AND U476 ( .A(p_input[7953]), .B(p_input[6953]), .Z(n424) );
  AND U477 ( .A(p_input[9953]), .B(p_input[953]), .Z(n422) );
  AND U478 ( .A(n425), .B(n426), .Z(o[952]) );
  AND U479 ( .A(n427), .B(n428), .Z(n426) );
  AND U480 ( .A(n429), .B(p_input[3952]), .Z(n428) );
  AND U481 ( .A(p_input[2952]), .B(p_input[1952]), .Z(n429) );
  AND U482 ( .A(p_input[5952]), .B(p_input[4952]), .Z(n427) );
  AND U483 ( .A(n430), .B(n431), .Z(n425) );
  AND U484 ( .A(n432), .B(p_input[8952]), .Z(n431) );
  AND U485 ( .A(p_input[7952]), .B(p_input[6952]), .Z(n432) );
  AND U486 ( .A(p_input[9952]), .B(p_input[952]), .Z(n430) );
  AND U487 ( .A(n433), .B(n434), .Z(o[951]) );
  AND U488 ( .A(n435), .B(n436), .Z(n434) );
  AND U489 ( .A(n437), .B(p_input[3951]), .Z(n436) );
  AND U490 ( .A(p_input[2951]), .B(p_input[1951]), .Z(n437) );
  AND U491 ( .A(p_input[5951]), .B(p_input[4951]), .Z(n435) );
  AND U492 ( .A(n438), .B(n439), .Z(n433) );
  AND U493 ( .A(n440), .B(p_input[8951]), .Z(n439) );
  AND U494 ( .A(p_input[7951]), .B(p_input[6951]), .Z(n440) );
  AND U495 ( .A(p_input[9951]), .B(p_input[951]), .Z(n438) );
  AND U496 ( .A(n441), .B(n442), .Z(o[950]) );
  AND U497 ( .A(n443), .B(n444), .Z(n442) );
  AND U498 ( .A(n445), .B(p_input[3950]), .Z(n444) );
  AND U499 ( .A(p_input[2950]), .B(p_input[1950]), .Z(n445) );
  AND U500 ( .A(p_input[5950]), .B(p_input[4950]), .Z(n443) );
  AND U501 ( .A(n446), .B(n447), .Z(n441) );
  AND U502 ( .A(n448), .B(p_input[8950]), .Z(n447) );
  AND U503 ( .A(p_input[7950]), .B(p_input[6950]), .Z(n448) );
  AND U504 ( .A(p_input[9950]), .B(p_input[950]), .Z(n446) );
  AND U505 ( .A(n449), .B(n450), .Z(o[94]) );
  AND U506 ( .A(n451), .B(n452), .Z(n450) );
  AND U507 ( .A(n453), .B(p_input[3094]), .Z(n452) );
  AND U508 ( .A(p_input[2094]), .B(p_input[1094]), .Z(n453) );
  AND U509 ( .A(p_input[5094]), .B(p_input[4094]), .Z(n451) );
  AND U510 ( .A(n454), .B(n455), .Z(n449) );
  AND U511 ( .A(n456), .B(p_input[8094]), .Z(n455) );
  AND U512 ( .A(p_input[7094]), .B(p_input[6094]), .Z(n456) );
  AND U513 ( .A(p_input[94]), .B(p_input[9094]), .Z(n454) );
  AND U514 ( .A(n457), .B(n458), .Z(o[949]) );
  AND U515 ( .A(n459), .B(n460), .Z(n458) );
  AND U516 ( .A(n461), .B(p_input[3949]), .Z(n460) );
  AND U517 ( .A(p_input[2949]), .B(p_input[1949]), .Z(n461) );
  AND U518 ( .A(p_input[5949]), .B(p_input[4949]), .Z(n459) );
  AND U519 ( .A(n462), .B(n463), .Z(n457) );
  AND U520 ( .A(n464), .B(p_input[8949]), .Z(n463) );
  AND U521 ( .A(p_input[7949]), .B(p_input[6949]), .Z(n464) );
  AND U522 ( .A(p_input[9949]), .B(p_input[949]), .Z(n462) );
  AND U523 ( .A(n465), .B(n466), .Z(o[948]) );
  AND U524 ( .A(n467), .B(n468), .Z(n466) );
  AND U525 ( .A(n469), .B(p_input[3948]), .Z(n468) );
  AND U526 ( .A(p_input[2948]), .B(p_input[1948]), .Z(n469) );
  AND U527 ( .A(p_input[5948]), .B(p_input[4948]), .Z(n467) );
  AND U528 ( .A(n470), .B(n471), .Z(n465) );
  AND U529 ( .A(n472), .B(p_input[8948]), .Z(n471) );
  AND U530 ( .A(p_input[7948]), .B(p_input[6948]), .Z(n472) );
  AND U531 ( .A(p_input[9948]), .B(p_input[948]), .Z(n470) );
  AND U532 ( .A(n473), .B(n474), .Z(o[947]) );
  AND U533 ( .A(n475), .B(n476), .Z(n474) );
  AND U534 ( .A(n477), .B(p_input[3947]), .Z(n476) );
  AND U535 ( .A(p_input[2947]), .B(p_input[1947]), .Z(n477) );
  AND U536 ( .A(p_input[5947]), .B(p_input[4947]), .Z(n475) );
  AND U537 ( .A(n478), .B(n479), .Z(n473) );
  AND U538 ( .A(n480), .B(p_input[8947]), .Z(n479) );
  AND U539 ( .A(p_input[7947]), .B(p_input[6947]), .Z(n480) );
  AND U540 ( .A(p_input[9947]), .B(p_input[947]), .Z(n478) );
  AND U541 ( .A(n481), .B(n482), .Z(o[946]) );
  AND U542 ( .A(n483), .B(n484), .Z(n482) );
  AND U543 ( .A(n485), .B(p_input[3946]), .Z(n484) );
  AND U544 ( .A(p_input[2946]), .B(p_input[1946]), .Z(n485) );
  AND U545 ( .A(p_input[5946]), .B(p_input[4946]), .Z(n483) );
  AND U546 ( .A(n486), .B(n487), .Z(n481) );
  AND U547 ( .A(n488), .B(p_input[8946]), .Z(n487) );
  AND U548 ( .A(p_input[7946]), .B(p_input[6946]), .Z(n488) );
  AND U549 ( .A(p_input[9946]), .B(p_input[946]), .Z(n486) );
  AND U550 ( .A(n489), .B(n490), .Z(o[945]) );
  AND U551 ( .A(n491), .B(n492), .Z(n490) );
  AND U552 ( .A(n493), .B(p_input[3945]), .Z(n492) );
  AND U553 ( .A(p_input[2945]), .B(p_input[1945]), .Z(n493) );
  AND U554 ( .A(p_input[5945]), .B(p_input[4945]), .Z(n491) );
  AND U555 ( .A(n494), .B(n495), .Z(n489) );
  AND U556 ( .A(n496), .B(p_input[8945]), .Z(n495) );
  AND U557 ( .A(p_input[7945]), .B(p_input[6945]), .Z(n496) );
  AND U558 ( .A(p_input[9945]), .B(p_input[945]), .Z(n494) );
  AND U559 ( .A(n497), .B(n498), .Z(o[944]) );
  AND U560 ( .A(n499), .B(n500), .Z(n498) );
  AND U561 ( .A(n501), .B(p_input[3944]), .Z(n500) );
  AND U562 ( .A(p_input[2944]), .B(p_input[1944]), .Z(n501) );
  AND U563 ( .A(p_input[5944]), .B(p_input[4944]), .Z(n499) );
  AND U564 ( .A(n502), .B(n503), .Z(n497) );
  AND U565 ( .A(n504), .B(p_input[8944]), .Z(n503) );
  AND U566 ( .A(p_input[7944]), .B(p_input[6944]), .Z(n504) );
  AND U567 ( .A(p_input[9944]), .B(p_input[944]), .Z(n502) );
  AND U568 ( .A(n505), .B(n506), .Z(o[943]) );
  AND U569 ( .A(n507), .B(n508), .Z(n506) );
  AND U570 ( .A(n509), .B(p_input[3943]), .Z(n508) );
  AND U571 ( .A(p_input[2943]), .B(p_input[1943]), .Z(n509) );
  AND U572 ( .A(p_input[5943]), .B(p_input[4943]), .Z(n507) );
  AND U573 ( .A(n510), .B(n511), .Z(n505) );
  AND U574 ( .A(n512), .B(p_input[8943]), .Z(n511) );
  AND U575 ( .A(p_input[7943]), .B(p_input[6943]), .Z(n512) );
  AND U576 ( .A(p_input[9943]), .B(p_input[943]), .Z(n510) );
  AND U577 ( .A(n513), .B(n514), .Z(o[942]) );
  AND U578 ( .A(n515), .B(n516), .Z(n514) );
  AND U579 ( .A(n517), .B(p_input[3942]), .Z(n516) );
  AND U580 ( .A(p_input[2942]), .B(p_input[1942]), .Z(n517) );
  AND U581 ( .A(p_input[5942]), .B(p_input[4942]), .Z(n515) );
  AND U582 ( .A(n518), .B(n519), .Z(n513) );
  AND U583 ( .A(n520), .B(p_input[8942]), .Z(n519) );
  AND U584 ( .A(p_input[7942]), .B(p_input[6942]), .Z(n520) );
  AND U585 ( .A(p_input[9942]), .B(p_input[942]), .Z(n518) );
  AND U586 ( .A(n521), .B(n522), .Z(o[941]) );
  AND U587 ( .A(n523), .B(n524), .Z(n522) );
  AND U588 ( .A(n525), .B(p_input[3941]), .Z(n524) );
  AND U589 ( .A(p_input[2941]), .B(p_input[1941]), .Z(n525) );
  AND U590 ( .A(p_input[5941]), .B(p_input[4941]), .Z(n523) );
  AND U591 ( .A(n526), .B(n527), .Z(n521) );
  AND U592 ( .A(n528), .B(p_input[8941]), .Z(n527) );
  AND U593 ( .A(p_input[7941]), .B(p_input[6941]), .Z(n528) );
  AND U594 ( .A(p_input[9941]), .B(p_input[941]), .Z(n526) );
  AND U595 ( .A(n529), .B(n530), .Z(o[940]) );
  AND U596 ( .A(n531), .B(n532), .Z(n530) );
  AND U597 ( .A(n533), .B(p_input[3940]), .Z(n532) );
  AND U598 ( .A(p_input[2940]), .B(p_input[1940]), .Z(n533) );
  AND U599 ( .A(p_input[5940]), .B(p_input[4940]), .Z(n531) );
  AND U600 ( .A(n534), .B(n535), .Z(n529) );
  AND U601 ( .A(n536), .B(p_input[8940]), .Z(n535) );
  AND U602 ( .A(p_input[7940]), .B(p_input[6940]), .Z(n536) );
  AND U603 ( .A(p_input[9940]), .B(p_input[940]), .Z(n534) );
  AND U604 ( .A(n537), .B(n538), .Z(o[93]) );
  AND U605 ( .A(n539), .B(n540), .Z(n538) );
  AND U606 ( .A(n541), .B(p_input[3093]), .Z(n540) );
  AND U607 ( .A(p_input[2093]), .B(p_input[1093]), .Z(n541) );
  AND U608 ( .A(p_input[5093]), .B(p_input[4093]), .Z(n539) );
  AND U609 ( .A(n542), .B(n543), .Z(n537) );
  AND U610 ( .A(n544), .B(p_input[8093]), .Z(n543) );
  AND U611 ( .A(p_input[7093]), .B(p_input[6093]), .Z(n544) );
  AND U612 ( .A(p_input[93]), .B(p_input[9093]), .Z(n542) );
  AND U613 ( .A(n545), .B(n546), .Z(o[939]) );
  AND U614 ( .A(n547), .B(n548), .Z(n546) );
  AND U615 ( .A(n549), .B(p_input[3939]), .Z(n548) );
  AND U616 ( .A(p_input[2939]), .B(p_input[1939]), .Z(n549) );
  AND U617 ( .A(p_input[5939]), .B(p_input[4939]), .Z(n547) );
  AND U618 ( .A(n550), .B(n551), .Z(n545) );
  AND U619 ( .A(n552), .B(p_input[8939]), .Z(n551) );
  AND U620 ( .A(p_input[7939]), .B(p_input[6939]), .Z(n552) );
  AND U621 ( .A(p_input[9939]), .B(p_input[939]), .Z(n550) );
  AND U622 ( .A(n553), .B(n554), .Z(o[938]) );
  AND U623 ( .A(n555), .B(n556), .Z(n554) );
  AND U624 ( .A(n557), .B(p_input[3938]), .Z(n556) );
  AND U625 ( .A(p_input[2938]), .B(p_input[1938]), .Z(n557) );
  AND U626 ( .A(p_input[5938]), .B(p_input[4938]), .Z(n555) );
  AND U627 ( .A(n558), .B(n559), .Z(n553) );
  AND U628 ( .A(n560), .B(p_input[8938]), .Z(n559) );
  AND U629 ( .A(p_input[7938]), .B(p_input[6938]), .Z(n560) );
  AND U630 ( .A(p_input[9938]), .B(p_input[938]), .Z(n558) );
  AND U631 ( .A(n561), .B(n562), .Z(o[937]) );
  AND U632 ( .A(n563), .B(n564), .Z(n562) );
  AND U633 ( .A(n565), .B(p_input[3937]), .Z(n564) );
  AND U634 ( .A(p_input[2937]), .B(p_input[1937]), .Z(n565) );
  AND U635 ( .A(p_input[5937]), .B(p_input[4937]), .Z(n563) );
  AND U636 ( .A(n566), .B(n567), .Z(n561) );
  AND U637 ( .A(n568), .B(p_input[8937]), .Z(n567) );
  AND U638 ( .A(p_input[7937]), .B(p_input[6937]), .Z(n568) );
  AND U639 ( .A(p_input[9937]), .B(p_input[937]), .Z(n566) );
  AND U640 ( .A(n569), .B(n570), .Z(o[936]) );
  AND U641 ( .A(n571), .B(n572), .Z(n570) );
  AND U642 ( .A(n573), .B(p_input[3936]), .Z(n572) );
  AND U643 ( .A(p_input[2936]), .B(p_input[1936]), .Z(n573) );
  AND U644 ( .A(p_input[5936]), .B(p_input[4936]), .Z(n571) );
  AND U645 ( .A(n574), .B(n575), .Z(n569) );
  AND U646 ( .A(n576), .B(p_input[8936]), .Z(n575) );
  AND U647 ( .A(p_input[7936]), .B(p_input[6936]), .Z(n576) );
  AND U648 ( .A(p_input[9936]), .B(p_input[936]), .Z(n574) );
  AND U649 ( .A(n577), .B(n578), .Z(o[935]) );
  AND U650 ( .A(n579), .B(n580), .Z(n578) );
  AND U651 ( .A(n581), .B(p_input[3935]), .Z(n580) );
  AND U652 ( .A(p_input[2935]), .B(p_input[1935]), .Z(n581) );
  AND U653 ( .A(p_input[5935]), .B(p_input[4935]), .Z(n579) );
  AND U654 ( .A(n582), .B(n583), .Z(n577) );
  AND U655 ( .A(n584), .B(p_input[8935]), .Z(n583) );
  AND U656 ( .A(p_input[7935]), .B(p_input[6935]), .Z(n584) );
  AND U657 ( .A(p_input[9935]), .B(p_input[935]), .Z(n582) );
  AND U658 ( .A(n585), .B(n586), .Z(o[934]) );
  AND U659 ( .A(n587), .B(n588), .Z(n586) );
  AND U660 ( .A(n589), .B(p_input[3934]), .Z(n588) );
  AND U661 ( .A(p_input[2934]), .B(p_input[1934]), .Z(n589) );
  AND U662 ( .A(p_input[5934]), .B(p_input[4934]), .Z(n587) );
  AND U663 ( .A(n590), .B(n591), .Z(n585) );
  AND U664 ( .A(n592), .B(p_input[8934]), .Z(n591) );
  AND U665 ( .A(p_input[7934]), .B(p_input[6934]), .Z(n592) );
  AND U666 ( .A(p_input[9934]), .B(p_input[934]), .Z(n590) );
  AND U667 ( .A(n593), .B(n594), .Z(o[933]) );
  AND U668 ( .A(n595), .B(n596), .Z(n594) );
  AND U669 ( .A(n597), .B(p_input[3933]), .Z(n596) );
  AND U670 ( .A(p_input[2933]), .B(p_input[1933]), .Z(n597) );
  AND U671 ( .A(p_input[5933]), .B(p_input[4933]), .Z(n595) );
  AND U672 ( .A(n598), .B(n599), .Z(n593) );
  AND U673 ( .A(n600), .B(p_input[8933]), .Z(n599) );
  AND U674 ( .A(p_input[7933]), .B(p_input[6933]), .Z(n600) );
  AND U675 ( .A(p_input[9933]), .B(p_input[933]), .Z(n598) );
  AND U676 ( .A(n601), .B(n602), .Z(o[932]) );
  AND U677 ( .A(n603), .B(n604), .Z(n602) );
  AND U678 ( .A(n605), .B(p_input[3932]), .Z(n604) );
  AND U679 ( .A(p_input[2932]), .B(p_input[1932]), .Z(n605) );
  AND U680 ( .A(p_input[5932]), .B(p_input[4932]), .Z(n603) );
  AND U681 ( .A(n606), .B(n607), .Z(n601) );
  AND U682 ( .A(n608), .B(p_input[8932]), .Z(n607) );
  AND U683 ( .A(p_input[7932]), .B(p_input[6932]), .Z(n608) );
  AND U684 ( .A(p_input[9932]), .B(p_input[932]), .Z(n606) );
  AND U685 ( .A(n609), .B(n610), .Z(o[931]) );
  AND U686 ( .A(n611), .B(n612), .Z(n610) );
  AND U687 ( .A(n613), .B(p_input[3931]), .Z(n612) );
  AND U688 ( .A(p_input[2931]), .B(p_input[1931]), .Z(n613) );
  AND U689 ( .A(p_input[5931]), .B(p_input[4931]), .Z(n611) );
  AND U690 ( .A(n614), .B(n615), .Z(n609) );
  AND U691 ( .A(n616), .B(p_input[8931]), .Z(n615) );
  AND U692 ( .A(p_input[7931]), .B(p_input[6931]), .Z(n616) );
  AND U693 ( .A(p_input[9931]), .B(p_input[931]), .Z(n614) );
  AND U694 ( .A(n617), .B(n618), .Z(o[930]) );
  AND U695 ( .A(n619), .B(n620), .Z(n618) );
  AND U696 ( .A(n621), .B(p_input[3930]), .Z(n620) );
  AND U697 ( .A(p_input[2930]), .B(p_input[1930]), .Z(n621) );
  AND U698 ( .A(p_input[5930]), .B(p_input[4930]), .Z(n619) );
  AND U699 ( .A(n622), .B(n623), .Z(n617) );
  AND U700 ( .A(n624), .B(p_input[8930]), .Z(n623) );
  AND U701 ( .A(p_input[7930]), .B(p_input[6930]), .Z(n624) );
  AND U702 ( .A(p_input[9930]), .B(p_input[930]), .Z(n622) );
  AND U703 ( .A(n625), .B(n626), .Z(o[92]) );
  AND U704 ( .A(n627), .B(n628), .Z(n626) );
  AND U705 ( .A(n629), .B(p_input[3092]), .Z(n628) );
  AND U706 ( .A(p_input[2092]), .B(p_input[1092]), .Z(n629) );
  AND U707 ( .A(p_input[5092]), .B(p_input[4092]), .Z(n627) );
  AND U708 ( .A(n630), .B(n631), .Z(n625) );
  AND U709 ( .A(n632), .B(p_input[8092]), .Z(n631) );
  AND U710 ( .A(p_input[7092]), .B(p_input[6092]), .Z(n632) );
  AND U711 ( .A(p_input[92]), .B(p_input[9092]), .Z(n630) );
  AND U712 ( .A(n633), .B(n634), .Z(o[929]) );
  AND U713 ( .A(n635), .B(n636), .Z(n634) );
  AND U714 ( .A(n637), .B(p_input[3929]), .Z(n636) );
  AND U715 ( .A(p_input[2929]), .B(p_input[1929]), .Z(n637) );
  AND U716 ( .A(p_input[5929]), .B(p_input[4929]), .Z(n635) );
  AND U717 ( .A(n638), .B(n639), .Z(n633) );
  AND U718 ( .A(n640), .B(p_input[8929]), .Z(n639) );
  AND U719 ( .A(p_input[7929]), .B(p_input[6929]), .Z(n640) );
  AND U720 ( .A(p_input[9929]), .B(p_input[929]), .Z(n638) );
  AND U721 ( .A(n641), .B(n642), .Z(o[928]) );
  AND U722 ( .A(n643), .B(n644), .Z(n642) );
  AND U723 ( .A(n645), .B(p_input[3928]), .Z(n644) );
  AND U724 ( .A(p_input[2928]), .B(p_input[1928]), .Z(n645) );
  AND U725 ( .A(p_input[5928]), .B(p_input[4928]), .Z(n643) );
  AND U726 ( .A(n646), .B(n647), .Z(n641) );
  AND U727 ( .A(n648), .B(p_input[8928]), .Z(n647) );
  AND U728 ( .A(p_input[7928]), .B(p_input[6928]), .Z(n648) );
  AND U729 ( .A(p_input[9928]), .B(p_input[928]), .Z(n646) );
  AND U730 ( .A(n649), .B(n650), .Z(o[927]) );
  AND U731 ( .A(n651), .B(n652), .Z(n650) );
  AND U732 ( .A(n653), .B(p_input[3927]), .Z(n652) );
  AND U733 ( .A(p_input[2927]), .B(p_input[1927]), .Z(n653) );
  AND U734 ( .A(p_input[5927]), .B(p_input[4927]), .Z(n651) );
  AND U735 ( .A(n654), .B(n655), .Z(n649) );
  AND U736 ( .A(n656), .B(p_input[8927]), .Z(n655) );
  AND U737 ( .A(p_input[7927]), .B(p_input[6927]), .Z(n656) );
  AND U738 ( .A(p_input[9927]), .B(p_input[927]), .Z(n654) );
  AND U739 ( .A(n657), .B(n658), .Z(o[926]) );
  AND U740 ( .A(n659), .B(n660), .Z(n658) );
  AND U741 ( .A(n661), .B(p_input[3926]), .Z(n660) );
  AND U742 ( .A(p_input[2926]), .B(p_input[1926]), .Z(n661) );
  AND U743 ( .A(p_input[5926]), .B(p_input[4926]), .Z(n659) );
  AND U744 ( .A(n662), .B(n663), .Z(n657) );
  AND U745 ( .A(n664), .B(p_input[8926]), .Z(n663) );
  AND U746 ( .A(p_input[7926]), .B(p_input[6926]), .Z(n664) );
  AND U747 ( .A(p_input[9926]), .B(p_input[926]), .Z(n662) );
  AND U748 ( .A(n665), .B(n666), .Z(o[925]) );
  AND U749 ( .A(n667), .B(n668), .Z(n666) );
  AND U750 ( .A(n669), .B(p_input[3925]), .Z(n668) );
  AND U751 ( .A(p_input[2925]), .B(p_input[1925]), .Z(n669) );
  AND U752 ( .A(p_input[5925]), .B(p_input[4925]), .Z(n667) );
  AND U753 ( .A(n670), .B(n671), .Z(n665) );
  AND U754 ( .A(n672), .B(p_input[8925]), .Z(n671) );
  AND U755 ( .A(p_input[7925]), .B(p_input[6925]), .Z(n672) );
  AND U756 ( .A(p_input[9925]), .B(p_input[925]), .Z(n670) );
  AND U757 ( .A(n673), .B(n674), .Z(o[924]) );
  AND U758 ( .A(n675), .B(n676), .Z(n674) );
  AND U759 ( .A(n677), .B(p_input[3924]), .Z(n676) );
  AND U760 ( .A(p_input[2924]), .B(p_input[1924]), .Z(n677) );
  AND U761 ( .A(p_input[5924]), .B(p_input[4924]), .Z(n675) );
  AND U762 ( .A(n678), .B(n679), .Z(n673) );
  AND U763 ( .A(n680), .B(p_input[8924]), .Z(n679) );
  AND U764 ( .A(p_input[7924]), .B(p_input[6924]), .Z(n680) );
  AND U765 ( .A(p_input[9924]), .B(p_input[924]), .Z(n678) );
  AND U766 ( .A(n681), .B(n682), .Z(o[923]) );
  AND U767 ( .A(n683), .B(n684), .Z(n682) );
  AND U768 ( .A(n685), .B(p_input[3923]), .Z(n684) );
  AND U769 ( .A(p_input[2923]), .B(p_input[1923]), .Z(n685) );
  AND U770 ( .A(p_input[5923]), .B(p_input[4923]), .Z(n683) );
  AND U771 ( .A(n686), .B(n687), .Z(n681) );
  AND U772 ( .A(n688), .B(p_input[8923]), .Z(n687) );
  AND U773 ( .A(p_input[7923]), .B(p_input[6923]), .Z(n688) );
  AND U774 ( .A(p_input[9923]), .B(p_input[923]), .Z(n686) );
  AND U775 ( .A(n689), .B(n690), .Z(o[922]) );
  AND U776 ( .A(n691), .B(n692), .Z(n690) );
  AND U777 ( .A(n693), .B(p_input[3922]), .Z(n692) );
  AND U778 ( .A(p_input[2922]), .B(p_input[1922]), .Z(n693) );
  AND U779 ( .A(p_input[5922]), .B(p_input[4922]), .Z(n691) );
  AND U780 ( .A(n694), .B(n695), .Z(n689) );
  AND U781 ( .A(n696), .B(p_input[8922]), .Z(n695) );
  AND U782 ( .A(p_input[7922]), .B(p_input[6922]), .Z(n696) );
  AND U783 ( .A(p_input[9922]), .B(p_input[922]), .Z(n694) );
  AND U784 ( .A(n697), .B(n698), .Z(o[921]) );
  AND U785 ( .A(n699), .B(n700), .Z(n698) );
  AND U786 ( .A(n701), .B(p_input[3921]), .Z(n700) );
  AND U787 ( .A(p_input[2921]), .B(p_input[1921]), .Z(n701) );
  AND U788 ( .A(p_input[5921]), .B(p_input[4921]), .Z(n699) );
  AND U789 ( .A(n702), .B(n703), .Z(n697) );
  AND U790 ( .A(n704), .B(p_input[8921]), .Z(n703) );
  AND U791 ( .A(p_input[7921]), .B(p_input[6921]), .Z(n704) );
  AND U792 ( .A(p_input[9921]), .B(p_input[921]), .Z(n702) );
  AND U793 ( .A(n705), .B(n706), .Z(o[920]) );
  AND U794 ( .A(n707), .B(n708), .Z(n706) );
  AND U795 ( .A(n709), .B(p_input[3920]), .Z(n708) );
  AND U796 ( .A(p_input[2920]), .B(p_input[1920]), .Z(n709) );
  AND U797 ( .A(p_input[5920]), .B(p_input[4920]), .Z(n707) );
  AND U798 ( .A(n710), .B(n711), .Z(n705) );
  AND U799 ( .A(n712), .B(p_input[8920]), .Z(n711) );
  AND U800 ( .A(p_input[7920]), .B(p_input[6920]), .Z(n712) );
  AND U801 ( .A(p_input[9920]), .B(p_input[920]), .Z(n710) );
  AND U802 ( .A(n713), .B(n714), .Z(o[91]) );
  AND U803 ( .A(n715), .B(n716), .Z(n714) );
  AND U804 ( .A(n717), .B(p_input[3091]), .Z(n716) );
  AND U805 ( .A(p_input[2091]), .B(p_input[1091]), .Z(n717) );
  AND U806 ( .A(p_input[5091]), .B(p_input[4091]), .Z(n715) );
  AND U807 ( .A(n718), .B(n719), .Z(n713) );
  AND U808 ( .A(n720), .B(p_input[8091]), .Z(n719) );
  AND U809 ( .A(p_input[7091]), .B(p_input[6091]), .Z(n720) );
  AND U810 ( .A(p_input[91]), .B(p_input[9091]), .Z(n718) );
  AND U811 ( .A(n721), .B(n722), .Z(o[919]) );
  AND U812 ( .A(n723), .B(n724), .Z(n722) );
  AND U813 ( .A(n725), .B(p_input[3919]), .Z(n724) );
  AND U814 ( .A(p_input[2919]), .B(p_input[1919]), .Z(n725) );
  AND U815 ( .A(p_input[5919]), .B(p_input[4919]), .Z(n723) );
  AND U816 ( .A(n726), .B(n727), .Z(n721) );
  AND U817 ( .A(n728), .B(p_input[8919]), .Z(n727) );
  AND U818 ( .A(p_input[7919]), .B(p_input[6919]), .Z(n728) );
  AND U819 ( .A(p_input[9919]), .B(p_input[919]), .Z(n726) );
  AND U820 ( .A(n729), .B(n730), .Z(o[918]) );
  AND U821 ( .A(n731), .B(n732), .Z(n730) );
  AND U822 ( .A(n733), .B(p_input[3918]), .Z(n732) );
  AND U823 ( .A(p_input[2918]), .B(p_input[1918]), .Z(n733) );
  AND U824 ( .A(p_input[5918]), .B(p_input[4918]), .Z(n731) );
  AND U825 ( .A(n734), .B(n735), .Z(n729) );
  AND U826 ( .A(n736), .B(p_input[8918]), .Z(n735) );
  AND U827 ( .A(p_input[7918]), .B(p_input[6918]), .Z(n736) );
  AND U828 ( .A(p_input[9918]), .B(p_input[918]), .Z(n734) );
  AND U829 ( .A(n737), .B(n738), .Z(o[917]) );
  AND U830 ( .A(n739), .B(n740), .Z(n738) );
  AND U831 ( .A(n741), .B(p_input[3917]), .Z(n740) );
  AND U832 ( .A(p_input[2917]), .B(p_input[1917]), .Z(n741) );
  AND U833 ( .A(p_input[5917]), .B(p_input[4917]), .Z(n739) );
  AND U834 ( .A(n742), .B(n743), .Z(n737) );
  AND U835 ( .A(n744), .B(p_input[8917]), .Z(n743) );
  AND U836 ( .A(p_input[7917]), .B(p_input[6917]), .Z(n744) );
  AND U837 ( .A(p_input[9917]), .B(p_input[917]), .Z(n742) );
  AND U838 ( .A(n745), .B(n746), .Z(o[916]) );
  AND U839 ( .A(n747), .B(n748), .Z(n746) );
  AND U840 ( .A(n749), .B(p_input[3916]), .Z(n748) );
  AND U841 ( .A(p_input[2916]), .B(p_input[1916]), .Z(n749) );
  AND U842 ( .A(p_input[5916]), .B(p_input[4916]), .Z(n747) );
  AND U843 ( .A(n750), .B(n751), .Z(n745) );
  AND U844 ( .A(n752), .B(p_input[8916]), .Z(n751) );
  AND U845 ( .A(p_input[7916]), .B(p_input[6916]), .Z(n752) );
  AND U846 ( .A(p_input[9916]), .B(p_input[916]), .Z(n750) );
  AND U847 ( .A(n753), .B(n754), .Z(o[915]) );
  AND U848 ( .A(n755), .B(n756), .Z(n754) );
  AND U849 ( .A(n757), .B(p_input[3915]), .Z(n756) );
  AND U850 ( .A(p_input[2915]), .B(p_input[1915]), .Z(n757) );
  AND U851 ( .A(p_input[5915]), .B(p_input[4915]), .Z(n755) );
  AND U852 ( .A(n758), .B(n759), .Z(n753) );
  AND U853 ( .A(n760), .B(p_input[8915]), .Z(n759) );
  AND U854 ( .A(p_input[7915]), .B(p_input[6915]), .Z(n760) );
  AND U855 ( .A(p_input[9915]), .B(p_input[915]), .Z(n758) );
  AND U856 ( .A(n761), .B(n762), .Z(o[914]) );
  AND U857 ( .A(n763), .B(n764), .Z(n762) );
  AND U858 ( .A(n765), .B(p_input[3914]), .Z(n764) );
  AND U859 ( .A(p_input[2914]), .B(p_input[1914]), .Z(n765) );
  AND U860 ( .A(p_input[5914]), .B(p_input[4914]), .Z(n763) );
  AND U861 ( .A(n766), .B(n767), .Z(n761) );
  AND U862 ( .A(n768), .B(p_input[8914]), .Z(n767) );
  AND U863 ( .A(p_input[7914]), .B(p_input[6914]), .Z(n768) );
  AND U864 ( .A(p_input[9914]), .B(p_input[914]), .Z(n766) );
  AND U865 ( .A(n769), .B(n770), .Z(o[913]) );
  AND U866 ( .A(n771), .B(n772), .Z(n770) );
  AND U867 ( .A(n773), .B(p_input[3913]), .Z(n772) );
  AND U868 ( .A(p_input[2913]), .B(p_input[1913]), .Z(n773) );
  AND U869 ( .A(p_input[5913]), .B(p_input[4913]), .Z(n771) );
  AND U870 ( .A(n774), .B(n775), .Z(n769) );
  AND U871 ( .A(n776), .B(p_input[8913]), .Z(n775) );
  AND U872 ( .A(p_input[7913]), .B(p_input[6913]), .Z(n776) );
  AND U873 ( .A(p_input[9913]), .B(p_input[913]), .Z(n774) );
  AND U874 ( .A(n777), .B(n778), .Z(o[912]) );
  AND U875 ( .A(n779), .B(n780), .Z(n778) );
  AND U876 ( .A(n781), .B(p_input[3912]), .Z(n780) );
  AND U877 ( .A(p_input[2912]), .B(p_input[1912]), .Z(n781) );
  AND U878 ( .A(p_input[5912]), .B(p_input[4912]), .Z(n779) );
  AND U879 ( .A(n782), .B(n783), .Z(n777) );
  AND U880 ( .A(n784), .B(p_input[8912]), .Z(n783) );
  AND U881 ( .A(p_input[7912]), .B(p_input[6912]), .Z(n784) );
  AND U882 ( .A(p_input[9912]), .B(p_input[912]), .Z(n782) );
  AND U883 ( .A(n785), .B(n786), .Z(o[911]) );
  AND U884 ( .A(n787), .B(n788), .Z(n786) );
  AND U885 ( .A(n789), .B(p_input[3911]), .Z(n788) );
  AND U886 ( .A(p_input[2911]), .B(p_input[1911]), .Z(n789) );
  AND U887 ( .A(p_input[5911]), .B(p_input[4911]), .Z(n787) );
  AND U888 ( .A(n790), .B(n791), .Z(n785) );
  AND U889 ( .A(n792), .B(p_input[8911]), .Z(n791) );
  AND U890 ( .A(p_input[7911]), .B(p_input[6911]), .Z(n792) );
  AND U891 ( .A(p_input[9911]), .B(p_input[911]), .Z(n790) );
  AND U892 ( .A(n793), .B(n794), .Z(o[910]) );
  AND U893 ( .A(n795), .B(n796), .Z(n794) );
  AND U894 ( .A(n797), .B(p_input[3910]), .Z(n796) );
  AND U895 ( .A(p_input[2910]), .B(p_input[1910]), .Z(n797) );
  AND U896 ( .A(p_input[5910]), .B(p_input[4910]), .Z(n795) );
  AND U897 ( .A(n798), .B(n799), .Z(n793) );
  AND U898 ( .A(n800), .B(p_input[8910]), .Z(n799) );
  AND U899 ( .A(p_input[7910]), .B(p_input[6910]), .Z(n800) );
  AND U900 ( .A(p_input[9910]), .B(p_input[910]), .Z(n798) );
  AND U901 ( .A(n801), .B(n802), .Z(o[90]) );
  AND U902 ( .A(n803), .B(n804), .Z(n802) );
  AND U903 ( .A(n805), .B(p_input[3090]), .Z(n804) );
  AND U904 ( .A(p_input[2090]), .B(p_input[1090]), .Z(n805) );
  AND U905 ( .A(p_input[5090]), .B(p_input[4090]), .Z(n803) );
  AND U906 ( .A(n806), .B(n807), .Z(n801) );
  AND U907 ( .A(n808), .B(p_input[8090]), .Z(n807) );
  AND U908 ( .A(p_input[7090]), .B(p_input[6090]), .Z(n808) );
  AND U909 ( .A(p_input[90]), .B(p_input[9090]), .Z(n806) );
  AND U910 ( .A(n809), .B(n810), .Z(o[909]) );
  AND U911 ( .A(n811), .B(n812), .Z(n810) );
  AND U912 ( .A(n813), .B(p_input[3909]), .Z(n812) );
  AND U913 ( .A(p_input[2909]), .B(p_input[1909]), .Z(n813) );
  AND U914 ( .A(p_input[5909]), .B(p_input[4909]), .Z(n811) );
  AND U915 ( .A(n814), .B(n815), .Z(n809) );
  AND U916 ( .A(n816), .B(p_input[8909]), .Z(n815) );
  AND U917 ( .A(p_input[7909]), .B(p_input[6909]), .Z(n816) );
  AND U918 ( .A(p_input[9909]), .B(p_input[909]), .Z(n814) );
  AND U919 ( .A(n817), .B(n818), .Z(o[908]) );
  AND U920 ( .A(n819), .B(n820), .Z(n818) );
  AND U921 ( .A(n821), .B(p_input[3908]), .Z(n820) );
  AND U922 ( .A(p_input[2908]), .B(p_input[1908]), .Z(n821) );
  AND U923 ( .A(p_input[5908]), .B(p_input[4908]), .Z(n819) );
  AND U924 ( .A(n822), .B(n823), .Z(n817) );
  AND U925 ( .A(n824), .B(p_input[8908]), .Z(n823) );
  AND U926 ( .A(p_input[7908]), .B(p_input[6908]), .Z(n824) );
  AND U927 ( .A(p_input[9908]), .B(p_input[908]), .Z(n822) );
  AND U928 ( .A(n825), .B(n826), .Z(o[907]) );
  AND U929 ( .A(n827), .B(n828), .Z(n826) );
  AND U930 ( .A(n829), .B(p_input[3907]), .Z(n828) );
  AND U931 ( .A(p_input[2907]), .B(p_input[1907]), .Z(n829) );
  AND U932 ( .A(p_input[5907]), .B(p_input[4907]), .Z(n827) );
  AND U933 ( .A(n830), .B(n831), .Z(n825) );
  AND U934 ( .A(n832), .B(p_input[8907]), .Z(n831) );
  AND U935 ( .A(p_input[7907]), .B(p_input[6907]), .Z(n832) );
  AND U936 ( .A(p_input[9907]), .B(p_input[907]), .Z(n830) );
  AND U937 ( .A(n833), .B(n834), .Z(o[906]) );
  AND U938 ( .A(n835), .B(n836), .Z(n834) );
  AND U939 ( .A(n837), .B(p_input[3906]), .Z(n836) );
  AND U940 ( .A(p_input[2906]), .B(p_input[1906]), .Z(n837) );
  AND U941 ( .A(p_input[5906]), .B(p_input[4906]), .Z(n835) );
  AND U942 ( .A(n838), .B(n839), .Z(n833) );
  AND U943 ( .A(n840), .B(p_input[8906]), .Z(n839) );
  AND U944 ( .A(p_input[7906]), .B(p_input[6906]), .Z(n840) );
  AND U945 ( .A(p_input[9906]), .B(p_input[906]), .Z(n838) );
  AND U946 ( .A(n841), .B(n842), .Z(o[905]) );
  AND U947 ( .A(n843), .B(n844), .Z(n842) );
  AND U948 ( .A(n845), .B(p_input[3905]), .Z(n844) );
  AND U949 ( .A(p_input[2905]), .B(p_input[1905]), .Z(n845) );
  AND U950 ( .A(p_input[5905]), .B(p_input[4905]), .Z(n843) );
  AND U951 ( .A(n846), .B(n847), .Z(n841) );
  AND U952 ( .A(n848), .B(p_input[8905]), .Z(n847) );
  AND U953 ( .A(p_input[7905]), .B(p_input[6905]), .Z(n848) );
  AND U954 ( .A(p_input[9905]), .B(p_input[905]), .Z(n846) );
  AND U955 ( .A(n849), .B(n850), .Z(o[904]) );
  AND U956 ( .A(n851), .B(n852), .Z(n850) );
  AND U957 ( .A(n853), .B(p_input[3904]), .Z(n852) );
  AND U958 ( .A(p_input[2904]), .B(p_input[1904]), .Z(n853) );
  AND U959 ( .A(p_input[5904]), .B(p_input[4904]), .Z(n851) );
  AND U960 ( .A(n854), .B(n855), .Z(n849) );
  AND U961 ( .A(n856), .B(p_input[8904]), .Z(n855) );
  AND U962 ( .A(p_input[7904]), .B(p_input[6904]), .Z(n856) );
  AND U963 ( .A(p_input[9904]), .B(p_input[904]), .Z(n854) );
  AND U964 ( .A(n857), .B(n858), .Z(o[903]) );
  AND U965 ( .A(n859), .B(n860), .Z(n858) );
  AND U966 ( .A(n861), .B(p_input[3903]), .Z(n860) );
  AND U967 ( .A(p_input[2903]), .B(p_input[1903]), .Z(n861) );
  AND U968 ( .A(p_input[5903]), .B(p_input[4903]), .Z(n859) );
  AND U969 ( .A(n862), .B(n863), .Z(n857) );
  AND U970 ( .A(n864), .B(p_input[8903]), .Z(n863) );
  AND U971 ( .A(p_input[7903]), .B(p_input[6903]), .Z(n864) );
  AND U972 ( .A(p_input[9903]), .B(p_input[903]), .Z(n862) );
  AND U973 ( .A(n865), .B(n866), .Z(o[902]) );
  AND U974 ( .A(n867), .B(n868), .Z(n866) );
  AND U975 ( .A(n869), .B(p_input[3902]), .Z(n868) );
  AND U976 ( .A(p_input[2902]), .B(p_input[1902]), .Z(n869) );
  AND U977 ( .A(p_input[5902]), .B(p_input[4902]), .Z(n867) );
  AND U978 ( .A(n870), .B(n871), .Z(n865) );
  AND U979 ( .A(n872), .B(p_input[8902]), .Z(n871) );
  AND U980 ( .A(p_input[7902]), .B(p_input[6902]), .Z(n872) );
  AND U981 ( .A(p_input[9902]), .B(p_input[902]), .Z(n870) );
  AND U982 ( .A(n873), .B(n874), .Z(o[901]) );
  AND U983 ( .A(n875), .B(n876), .Z(n874) );
  AND U984 ( .A(n877), .B(p_input[3901]), .Z(n876) );
  AND U985 ( .A(p_input[2901]), .B(p_input[1901]), .Z(n877) );
  AND U986 ( .A(p_input[5901]), .B(p_input[4901]), .Z(n875) );
  AND U987 ( .A(n878), .B(n879), .Z(n873) );
  AND U988 ( .A(n880), .B(p_input[8901]), .Z(n879) );
  AND U989 ( .A(p_input[7901]), .B(p_input[6901]), .Z(n880) );
  AND U990 ( .A(p_input[9901]), .B(p_input[901]), .Z(n878) );
  AND U991 ( .A(n881), .B(n882), .Z(o[900]) );
  AND U992 ( .A(n883), .B(n884), .Z(n882) );
  AND U993 ( .A(n885), .B(p_input[3900]), .Z(n884) );
  AND U994 ( .A(p_input[2900]), .B(p_input[1900]), .Z(n885) );
  AND U995 ( .A(p_input[5900]), .B(p_input[4900]), .Z(n883) );
  AND U996 ( .A(n886), .B(n887), .Z(n881) );
  AND U997 ( .A(n888), .B(p_input[8900]), .Z(n887) );
  AND U998 ( .A(p_input[7900]), .B(p_input[6900]), .Z(n888) );
  AND U999 ( .A(p_input[9900]), .B(p_input[900]), .Z(n886) );
  AND U1000 ( .A(n889), .B(n890), .Z(o[8]) );
  AND U1001 ( .A(n891), .B(n892), .Z(n890) );
  AND U1002 ( .A(n893), .B(p_input[3008]), .Z(n892) );
  AND U1003 ( .A(p_input[2008]), .B(p_input[1008]), .Z(n893) );
  AND U1004 ( .A(p_input[5008]), .B(p_input[4008]), .Z(n891) );
  AND U1005 ( .A(n894), .B(n895), .Z(n889) );
  AND U1006 ( .A(n896), .B(p_input[8008]), .Z(n895) );
  AND U1007 ( .A(p_input[7008]), .B(p_input[6008]), .Z(n896) );
  AND U1008 ( .A(p_input[9008]), .B(p_input[8]), .Z(n894) );
  AND U1009 ( .A(n897), .B(n898), .Z(o[89]) );
  AND U1010 ( .A(n899), .B(n900), .Z(n898) );
  AND U1011 ( .A(n901), .B(p_input[3089]), .Z(n900) );
  AND U1012 ( .A(p_input[2089]), .B(p_input[1089]), .Z(n901) );
  AND U1013 ( .A(p_input[5089]), .B(p_input[4089]), .Z(n899) );
  AND U1014 ( .A(n902), .B(n903), .Z(n897) );
  AND U1015 ( .A(n904), .B(p_input[8089]), .Z(n903) );
  AND U1016 ( .A(p_input[7089]), .B(p_input[6089]), .Z(n904) );
  AND U1017 ( .A(p_input[9089]), .B(p_input[89]), .Z(n902) );
  AND U1018 ( .A(n905), .B(n906), .Z(o[899]) );
  AND U1019 ( .A(n907), .B(n908), .Z(n906) );
  AND U1020 ( .A(n909), .B(p_input[3899]), .Z(n908) );
  AND U1021 ( .A(p_input[2899]), .B(p_input[1899]), .Z(n909) );
  AND U1022 ( .A(p_input[5899]), .B(p_input[4899]), .Z(n907) );
  AND U1023 ( .A(n910), .B(n911), .Z(n905) );
  AND U1024 ( .A(n912), .B(p_input[8899]), .Z(n911) );
  AND U1025 ( .A(p_input[7899]), .B(p_input[6899]), .Z(n912) );
  AND U1026 ( .A(p_input[9899]), .B(p_input[899]), .Z(n910) );
  AND U1027 ( .A(n913), .B(n914), .Z(o[898]) );
  AND U1028 ( .A(n915), .B(n916), .Z(n914) );
  AND U1029 ( .A(n917), .B(p_input[3898]), .Z(n916) );
  AND U1030 ( .A(p_input[2898]), .B(p_input[1898]), .Z(n917) );
  AND U1031 ( .A(p_input[5898]), .B(p_input[4898]), .Z(n915) );
  AND U1032 ( .A(n918), .B(n919), .Z(n913) );
  AND U1033 ( .A(n920), .B(p_input[8898]), .Z(n919) );
  AND U1034 ( .A(p_input[7898]), .B(p_input[6898]), .Z(n920) );
  AND U1035 ( .A(p_input[9898]), .B(p_input[898]), .Z(n918) );
  AND U1036 ( .A(n921), .B(n922), .Z(o[897]) );
  AND U1037 ( .A(n923), .B(n924), .Z(n922) );
  AND U1038 ( .A(n925), .B(p_input[3897]), .Z(n924) );
  AND U1039 ( .A(p_input[2897]), .B(p_input[1897]), .Z(n925) );
  AND U1040 ( .A(p_input[5897]), .B(p_input[4897]), .Z(n923) );
  AND U1041 ( .A(n926), .B(n927), .Z(n921) );
  AND U1042 ( .A(n928), .B(p_input[8897]), .Z(n927) );
  AND U1043 ( .A(p_input[7897]), .B(p_input[6897]), .Z(n928) );
  AND U1044 ( .A(p_input[9897]), .B(p_input[897]), .Z(n926) );
  AND U1045 ( .A(n929), .B(n930), .Z(o[896]) );
  AND U1046 ( .A(n931), .B(n932), .Z(n930) );
  AND U1047 ( .A(n933), .B(p_input[3896]), .Z(n932) );
  AND U1048 ( .A(p_input[2896]), .B(p_input[1896]), .Z(n933) );
  AND U1049 ( .A(p_input[5896]), .B(p_input[4896]), .Z(n931) );
  AND U1050 ( .A(n934), .B(n935), .Z(n929) );
  AND U1051 ( .A(n936), .B(p_input[8896]), .Z(n935) );
  AND U1052 ( .A(p_input[7896]), .B(p_input[6896]), .Z(n936) );
  AND U1053 ( .A(p_input[9896]), .B(p_input[896]), .Z(n934) );
  AND U1054 ( .A(n937), .B(n938), .Z(o[895]) );
  AND U1055 ( .A(n939), .B(n940), .Z(n938) );
  AND U1056 ( .A(n941), .B(p_input[3895]), .Z(n940) );
  AND U1057 ( .A(p_input[2895]), .B(p_input[1895]), .Z(n941) );
  AND U1058 ( .A(p_input[5895]), .B(p_input[4895]), .Z(n939) );
  AND U1059 ( .A(n942), .B(n943), .Z(n937) );
  AND U1060 ( .A(n944), .B(p_input[8895]), .Z(n943) );
  AND U1061 ( .A(p_input[7895]), .B(p_input[6895]), .Z(n944) );
  AND U1062 ( .A(p_input[9895]), .B(p_input[895]), .Z(n942) );
  AND U1063 ( .A(n945), .B(n946), .Z(o[894]) );
  AND U1064 ( .A(n947), .B(n948), .Z(n946) );
  AND U1065 ( .A(n949), .B(p_input[3894]), .Z(n948) );
  AND U1066 ( .A(p_input[2894]), .B(p_input[1894]), .Z(n949) );
  AND U1067 ( .A(p_input[5894]), .B(p_input[4894]), .Z(n947) );
  AND U1068 ( .A(n950), .B(n951), .Z(n945) );
  AND U1069 ( .A(n952), .B(p_input[8894]), .Z(n951) );
  AND U1070 ( .A(p_input[7894]), .B(p_input[6894]), .Z(n952) );
  AND U1071 ( .A(p_input[9894]), .B(p_input[894]), .Z(n950) );
  AND U1072 ( .A(n953), .B(n954), .Z(o[893]) );
  AND U1073 ( .A(n955), .B(n956), .Z(n954) );
  AND U1074 ( .A(n957), .B(p_input[3893]), .Z(n956) );
  AND U1075 ( .A(p_input[2893]), .B(p_input[1893]), .Z(n957) );
  AND U1076 ( .A(p_input[5893]), .B(p_input[4893]), .Z(n955) );
  AND U1077 ( .A(n958), .B(n959), .Z(n953) );
  AND U1078 ( .A(n960), .B(p_input[8893]), .Z(n959) );
  AND U1079 ( .A(p_input[7893]), .B(p_input[6893]), .Z(n960) );
  AND U1080 ( .A(p_input[9893]), .B(p_input[893]), .Z(n958) );
  AND U1081 ( .A(n961), .B(n962), .Z(o[892]) );
  AND U1082 ( .A(n963), .B(n964), .Z(n962) );
  AND U1083 ( .A(n965), .B(p_input[3892]), .Z(n964) );
  AND U1084 ( .A(p_input[2892]), .B(p_input[1892]), .Z(n965) );
  AND U1085 ( .A(p_input[5892]), .B(p_input[4892]), .Z(n963) );
  AND U1086 ( .A(n966), .B(n967), .Z(n961) );
  AND U1087 ( .A(n968), .B(p_input[8892]), .Z(n967) );
  AND U1088 ( .A(p_input[7892]), .B(p_input[6892]), .Z(n968) );
  AND U1089 ( .A(p_input[9892]), .B(p_input[892]), .Z(n966) );
  AND U1090 ( .A(n969), .B(n970), .Z(o[891]) );
  AND U1091 ( .A(n971), .B(n972), .Z(n970) );
  AND U1092 ( .A(n973), .B(p_input[3891]), .Z(n972) );
  AND U1093 ( .A(p_input[2891]), .B(p_input[1891]), .Z(n973) );
  AND U1094 ( .A(p_input[5891]), .B(p_input[4891]), .Z(n971) );
  AND U1095 ( .A(n974), .B(n975), .Z(n969) );
  AND U1096 ( .A(n976), .B(p_input[8891]), .Z(n975) );
  AND U1097 ( .A(p_input[7891]), .B(p_input[6891]), .Z(n976) );
  AND U1098 ( .A(p_input[9891]), .B(p_input[891]), .Z(n974) );
  AND U1099 ( .A(n977), .B(n978), .Z(o[890]) );
  AND U1100 ( .A(n979), .B(n980), .Z(n978) );
  AND U1101 ( .A(n981), .B(p_input[3890]), .Z(n980) );
  AND U1102 ( .A(p_input[2890]), .B(p_input[1890]), .Z(n981) );
  AND U1103 ( .A(p_input[5890]), .B(p_input[4890]), .Z(n979) );
  AND U1104 ( .A(n982), .B(n983), .Z(n977) );
  AND U1105 ( .A(n984), .B(p_input[8890]), .Z(n983) );
  AND U1106 ( .A(p_input[7890]), .B(p_input[6890]), .Z(n984) );
  AND U1107 ( .A(p_input[9890]), .B(p_input[890]), .Z(n982) );
  AND U1108 ( .A(n985), .B(n986), .Z(o[88]) );
  AND U1109 ( .A(n987), .B(n988), .Z(n986) );
  AND U1110 ( .A(n989), .B(p_input[3088]), .Z(n988) );
  AND U1111 ( .A(p_input[2088]), .B(p_input[1088]), .Z(n989) );
  AND U1112 ( .A(p_input[5088]), .B(p_input[4088]), .Z(n987) );
  AND U1113 ( .A(n990), .B(n991), .Z(n985) );
  AND U1114 ( .A(n992), .B(p_input[8088]), .Z(n991) );
  AND U1115 ( .A(p_input[7088]), .B(p_input[6088]), .Z(n992) );
  AND U1116 ( .A(p_input[9088]), .B(p_input[88]), .Z(n990) );
  AND U1117 ( .A(n993), .B(n994), .Z(o[889]) );
  AND U1118 ( .A(n995), .B(n996), .Z(n994) );
  AND U1119 ( .A(n997), .B(p_input[3889]), .Z(n996) );
  AND U1120 ( .A(p_input[2889]), .B(p_input[1889]), .Z(n997) );
  AND U1121 ( .A(p_input[5889]), .B(p_input[4889]), .Z(n995) );
  AND U1122 ( .A(n998), .B(n999), .Z(n993) );
  AND U1123 ( .A(n1000), .B(p_input[8889]), .Z(n999) );
  AND U1124 ( .A(p_input[7889]), .B(p_input[6889]), .Z(n1000) );
  AND U1125 ( .A(p_input[9889]), .B(p_input[889]), .Z(n998) );
  AND U1126 ( .A(n1001), .B(n1002), .Z(o[888]) );
  AND U1127 ( .A(n1003), .B(n1004), .Z(n1002) );
  AND U1128 ( .A(n1005), .B(p_input[3888]), .Z(n1004) );
  AND U1129 ( .A(p_input[2888]), .B(p_input[1888]), .Z(n1005) );
  AND U1130 ( .A(p_input[5888]), .B(p_input[4888]), .Z(n1003) );
  AND U1131 ( .A(n1006), .B(n1007), .Z(n1001) );
  AND U1132 ( .A(n1008), .B(p_input[8888]), .Z(n1007) );
  AND U1133 ( .A(p_input[7888]), .B(p_input[6888]), .Z(n1008) );
  AND U1134 ( .A(p_input[9888]), .B(p_input[888]), .Z(n1006) );
  AND U1135 ( .A(n1009), .B(n1010), .Z(o[887]) );
  AND U1136 ( .A(n1011), .B(n1012), .Z(n1010) );
  AND U1137 ( .A(n1013), .B(p_input[3887]), .Z(n1012) );
  AND U1138 ( .A(p_input[2887]), .B(p_input[1887]), .Z(n1013) );
  AND U1139 ( .A(p_input[5887]), .B(p_input[4887]), .Z(n1011) );
  AND U1140 ( .A(n1014), .B(n1015), .Z(n1009) );
  AND U1141 ( .A(n1016), .B(p_input[887]), .Z(n1015) );
  AND U1142 ( .A(p_input[7887]), .B(p_input[6887]), .Z(n1016) );
  AND U1143 ( .A(p_input[9887]), .B(p_input[8887]), .Z(n1014) );
  AND U1144 ( .A(n1017), .B(n1018), .Z(o[886]) );
  AND U1145 ( .A(n1019), .B(n1020), .Z(n1018) );
  AND U1146 ( .A(n1021), .B(p_input[3886]), .Z(n1020) );
  AND U1147 ( .A(p_input[2886]), .B(p_input[1886]), .Z(n1021) );
  AND U1148 ( .A(p_input[5886]), .B(p_input[4886]), .Z(n1019) );
  AND U1149 ( .A(n1022), .B(n1023), .Z(n1017) );
  AND U1150 ( .A(n1024), .B(p_input[886]), .Z(n1023) );
  AND U1151 ( .A(p_input[7886]), .B(p_input[6886]), .Z(n1024) );
  AND U1152 ( .A(p_input[9886]), .B(p_input[8886]), .Z(n1022) );
  AND U1153 ( .A(n1025), .B(n1026), .Z(o[885]) );
  AND U1154 ( .A(n1027), .B(n1028), .Z(n1026) );
  AND U1155 ( .A(n1029), .B(p_input[3885]), .Z(n1028) );
  AND U1156 ( .A(p_input[2885]), .B(p_input[1885]), .Z(n1029) );
  AND U1157 ( .A(p_input[5885]), .B(p_input[4885]), .Z(n1027) );
  AND U1158 ( .A(n1030), .B(n1031), .Z(n1025) );
  AND U1159 ( .A(n1032), .B(p_input[885]), .Z(n1031) );
  AND U1160 ( .A(p_input[7885]), .B(p_input[6885]), .Z(n1032) );
  AND U1161 ( .A(p_input[9885]), .B(p_input[8885]), .Z(n1030) );
  AND U1162 ( .A(n1033), .B(n1034), .Z(o[884]) );
  AND U1163 ( .A(n1035), .B(n1036), .Z(n1034) );
  AND U1164 ( .A(n1037), .B(p_input[3884]), .Z(n1036) );
  AND U1165 ( .A(p_input[2884]), .B(p_input[1884]), .Z(n1037) );
  AND U1166 ( .A(p_input[5884]), .B(p_input[4884]), .Z(n1035) );
  AND U1167 ( .A(n1038), .B(n1039), .Z(n1033) );
  AND U1168 ( .A(n1040), .B(p_input[884]), .Z(n1039) );
  AND U1169 ( .A(p_input[7884]), .B(p_input[6884]), .Z(n1040) );
  AND U1170 ( .A(p_input[9884]), .B(p_input[8884]), .Z(n1038) );
  AND U1171 ( .A(n1041), .B(n1042), .Z(o[883]) );
  AND U1172 ( .A(n1043), .B(n1044), .Z(n1042) );
  AND U1173 ( .A(n1045), .B(p_input[3883]), .Z(n1044) );
  AND U1174 ( .A(p_input[2883]), .B(p_input[1883]), .Z(n1045) );
  AND U1175 ( .A(p_input[5883]), .B(p_input[4883]), .Z(n1043) );
  AND U1176 ( .A(n1046), .B(n1047), .Z(n1041) );
  AND U1177 ( .A(n1048), .B(p_input[883]), .Z(n1047) );
  AND U1178 ( .A(p_input[7883]), .B(p_input[6883]), .Z(n1048) );
  AND U1179 ( .A(p_input[9883]), .B(p_input[8883]), .Z(n1046) );
  AND U1180 ( .A(n1049), .B(n1050), .Z(o[882]) );
  AND U1181 ( .A(n1051), .B(n1052), .Z(n1050) );
  AND U1182 ( .A(n1053), .B(p_input[3882]), .Z(n1052) );
  AND U1183 ( .A(p_input[2882]), .B(p_input[1882]), .Z(n1053) );
  AND U1184 ( .A(p_input[5882]), .B(p_input[4882]), .Z(n1051) );
  AND U1185 ( .A(n1054), .B(n1055), .Z(n1049) );
  AND U1186 ( .A(n1056), .B(p_input[882]), .Z(n1055) );
  AND U1187 ( .A(p_input[7882]), .B(p_input[6882]), .Z(n1056) );
  AND U1188 ( .A(p_input[9882]), .B(p_input[8882]), .Z(n1054) );
  AND U1189 ( .A(n1057), .B(n1058), .Z(o[881]) );
  AND U1190 ( .A(n1059), .B(n1060), .Z(n1058) );
  AND U1191 ( .A(n1061), .B(p_input[3881]), .Z(n1060) );
  AND U1192 ( .A(p_input[2881]), .B(p_input[1881]), .Z(n1061) );
  AND U1193 ( .A(p_input[5881]), .B(p_input[4881]), .Z(n1059) );
  AND U1194 ( .A(n1062), .B(n1063), .Z(n1057) );
  AND U1195 ( .A(n1064), .B(p_input[881]), .Z(n1063) );
  AND U1196 ( .A(p_input[7881]), .B(p_input[6881]), .Z(n1064) );
  AND U1197 ( .A(p_input[9881]), .B(p_input[8881]), .Z(n1062) );
  AND U1198 ( .A(n1065), .B(n1066), .Z(o[880]) );
  AND U1199 ( .A(n1067), .B(n1068), .Z(n1066) );
  AND U1200 ( .A(n1069), .B(p_input[3880]), .Z(n1068) );
  AND U1201 ( .A(p_input[2880]), .B(p_input[1880]), .Z(n1069) );
  AND U1202 ( .A(p_input[5880]), .B(p_input[4880]), .Z(n1067) );
  AND U1203 ( .A(n1070), .B(n1071), .Z(n1065) );
  AND U1204 ( .A(n1072), .B(p_input[880]), .Z(n1071) );
  AND U1205 ( .A(p_input[7880]), .B(p_input[6880]), .Z(n1072) );
  AND U1206 ( .A(p_input[9880]), .B(p_input[8880]), .Z(n1070) );
  AND U1207 ( .A(n1073), .B(n1074), .Z(o[87]) );
  AND U1208 ( .A(n1075), .B(n1076), .Z(n1074) );
  AND U1209 ( .A(n1077), .B(p_input[3087]), .Z(n1076) );
  AND U1210 ( .A(p_input[2087]), .B(p_input[1087]), .Z(n1077) );
  AND U1211 ( .A(p_input[5087]), .B(p_input[4087]), .Z(n1075) );
  AND U1212 ( .A(n1078), .B(n1079), .Z(n1073) );
  AND U1213 ( .A(n1080), .B(p_input[8087]), .Z(n1079) );
  AND U1214 ( .A(p_input[7087]), .B(p_input[6087]), .Z(n1080) );
  AND U1215 ( .A(p_input[9087]), .B(p_input[87]), .Z(n1078) );
  AND U1216 ( .A(n1081), .B(n1082), .Z(o[879]) );
  AND U1217 ( .A(n1083), .B(n1084), .Z(n1082) );
  AND U1218 ( .A(n1085), .B(p_input[3879]), .Z(n1084) );
  AND U1219 ( .A(p_input[2879]), .B(p_input[1879]), .Z(n1085) );
  AND U1220 ( .A(p_input[5879]), .B(p_input[4879]), .Z(n1083) );
  AND U1221 ( .A(n1086), .B(n1087), .Z(n1081) );
  AND U1222 ( .A(n1088), .B(p_input[879]), .Z(n1087) );
  AND U1223 ( .A(p_input[7879]), .B(p_input[6879]), .Z(n1088) );
  AND U1224 ( .A(p_input[9879]), .B(p_input[8879]), .Z(n1086) );
  AND U1225 ( .A(n1089), .B(n1090), .Z(o[878]) );
  AND U1226 ( .A(n1091), .B(n1092), .Z(n1090) );
  AND U1227 ( .A(n1093), .B(p_input[3878]), .Z(n1092) );
  AND U1228 ( .A(p_input[2878]), .B(p_input[1878]), .Z(n1093) );
  AND U1229 ( .A(p_input[5878]), .B(p_input[4878]), .Z(n1091) );
  AND U1230 ( .A(n1094), .B(n1095), .Z(n1089) );
  AND U1231 ( .A(n1096), .B(p_input[878]), .Z(n1095) );
  AND U1232 ( .A(p_input[7878]), .B(p_input[6878]), .Z(n1096) );
  AND U1233 ( .A(p_input[9878]), .B(p_input[8878]), .Z(n1094) );
  AND U1234 ( .A(n1097), .B(n1098), .Z(o[877]) );
  AND U1235 ( .A(n1099), .B(n1100), .Z(n1098) );
  AND U1236 ( .A(n1101), .B(p_input[3877]), .Z(n1100) );
  AND U1237 ( .A(p_input[2877]), .B(p_input[1877]), .Z(n1101) );
  AND U1238 ( .A(p_input[5877]), .B(p_input[4877]), .Z(n1099) );
  AND U1239 ( .A(n1102), .B(n1103), .Z(n1097) );
  AND U1240 ( .A(n1104), .B(p_input[877]), .Z(n1103) );
  AND U1241 ( .A(p_input[7877]), .B(p_input[6877]), .Z(n1104) );
  AND U1242 ( .A(p_input[9877]), .B(p_input[8877]), .Z(n1102) );
  AND U1243 ( .A(n1105), .B(n1106), .Z(o[876]) );
  AND U1244 ( .A(n1107), .B(n1108), .Z(n1106) );
  AND U1245 ( .A(n1109), .B(p_input[3876]), .Z(n1108) );
  AND U1246 ( .A(p_input[2876]), .B(p_input[1876]), .Z(n1109) );
  AND U1247 ( .A(p_input[5876]), .B(p_input[4876]), .Z(n1107) );
  AND U1248 ( .A(n1110), .B(n1111), .Z(n1105) );
  AND U1249 ( .A(n1112), .B(p_input[876]), .Z(n1111) );
  AND U1250 ( .A(p_input[7876]), .B(p_input[6876]), .Z(n1112) );
  AND U1251 ( .A(p_input[9876]), .B(p_input[8876]), .Z(n1110) );
  AND U1252 ( .A(n1113), .B(n1114), .Z(o[875]) );
  AND U1253 ( .A(n1115), .B(n1116), .Z(n1114) );
  AND U1254 ( .A(n1117), .B(p_input[3875]), .Z(n1116) );
  AND U1255 ( .A(p_input[2875]), .B(p_input[1875]), .Z(n1117) );
  AND U1256 ( .A(p_input[5875]), .B(p_input[4875]), .Z(n1115) );
  AND U1257 ( .A(n1118), .B(n1119), .Z(n1113) );
  AND U1258 ( .A(n1120), .B(p_input[875]), .Z(n1119) );
  AND U1259 ( .A(p_input[7875]), .B(p_input[6875]), .Z(n1120) );
  AND U1260 ( .A(p_input[9875]), .B(p_input[8875]), .Z(n1118) );
  AND U1261 ( .A(n1121), .B(n1122), .Z(o[874]) );
  AND U1262 ( .A(n1123), .B(n1124), .Z(n1122) );
  AND U1263 ( .A(n1125), .B(p_input[3874]), .Z(n1124) );
  AND U1264 ( .A(p_input[2874]), .B(p_input[1874]), .Z(n1125) );
  AND U1265 ( .A(p_input[5874]), .B(p_input[4874]), .Z(n1123) );
  AND U1266 ( .A(n1126), .B(n1127), .Z(n1121) );
  AND U1267 ( .A(n1128), .B(p_input[874]), .Z(n1127) );
  AND U1268 ( .A(p_input[7874]), .B(p_input[6874]), .Z(n1128) );
  AND U1269 ( .A(p_input[9874]), .B(p_input[8874]), .Z(n1126) );
  AND U1270 ( .A(n1129), .B(n1130), .Z(o[873]) );
  AND U1271 ( .A(n1131), .B(n1132), .Z(n1130) );
  AND U1272 ( .A(n1133), .B(p_input[3873]), .Z(n1132) );
  AND U1273 ( .A(p_input[2873]), .B(p_input[1873]), .Z(n1133) );
  AND U1274 ( .A(p_input[5873]), .B(p_input[4873]), .Z(n1131) );
  AND U1275 ( .A(n1134), .B(n1135), .Z(n1129) );
  AND U1276 ( .A(n1136), .B(p_input[873]), .Z(n1135) );
  AND U1277 ( .A(p_input[7873]), .B(p_input[6873]), .Z(n1136) );
  AND U1278 ( .A(p_input[9873]), .B(p_input[8873]), .Z(n1134) );
  AND U1279 ( .A(n1137), .B(n1138), .Z(o[872]) );
  AND U1280 ( .A(n1139), .B(n1140), .Z(n1138) );
  AND U1281 ( .A(n1141), .B(p_input[3872]), .Z(n1140) );
  AND U1282 ( .A(p_input[2872]), .B(p_input[1872]), .Z(n1141) );
  AND U1283 ( .A(p_input[5872]), .B(p_input[4872]), .Z(n1139) );
  AND U1284 ( .A(n1142), .B(n1143), .Z(n1137) );
  AND U1285 ( .A(n1144), .B(p_input[872]), .Z(n1143) );
  AND U1286 ( .A(p_input[7872]), .B(p_input[6872]), .Z(n1144) );
  AND U1287 ( .A(p_input[9872]), .B(p_input[8872]), .Z(n1142) );
  AND U1288 ( .A(n1145), .B(n1146), .Z(o[871]) );
  AND U1289 ( .A(n1147), .B(n1148), .Z(n1146) );
  AND U1290 ( .A(n1149), .B(p_input[3871]), .Z(n1148) );
  AND U1291 ( .A(p_input[2871]), .B(p_input[1871]), .Z(n1149) );
  AND U1292 ( .A(p_input[5871]), .B(p_input[4871]), .Z(n1147) );
  AND U1293 ( .A(n1150), .B(n1151), .Z(n1145) );
  AND U1294 ( .A(n1152), .B(p_input[871]), .Z(n1151) );
  AND U1295 ( .A(p_input[7871]), .B(p_input[6871]), .Z(n1152) );
  AND U1296 ( .A(p_input[9871]), .B(p_input[8871]), .Z(n1150) );
  AND U1297 ( .A(n1153), .B(n1154), .Z(o[870]) );
  AND U1298 ( .A(n1155), .B(n1156), .Z(n1154) );
  AND U1299 ( .A(n1157), .B(p_input[3870]), .Z(n1156) );
  AND U1300 ( .A(p_input[2870]), .B(p_input[1870]), .Z(n1157) );
  AND U1301 ( .A(p_input[5870]), .B(p_input[4870]), .Z(n1155) );
  AND U1302 ( .A(n1158), .B(n1159), .Z(n1153) );
  AND U1303 ( .A(n1160), .B(p_input[870]), .Z(n1159) );
  AND U1304 ( .A(p_input[7870]), .B(p_input[6870]), .Z(n1160) );
  AND U1305 ( .A(p_input[9870]), .B(p_input[8870]), .Z(n1158) );
  AND U1306 ( .A(n1161), .B(n1162), .Z(o[86]) );
  AND U1307 ( .A(n1163), .B(n1164), .Z(n1162) );
  AND U1308 ( .A(n1165), .B(p_input[3086]), .Z(n1164) );
  AND U1309 ( .A(p_input[2086]), .B(p_input[1086]), .Z(n1165) );
  AND U1310 ( .A(p_input[5086]), .B(p_input[4086]), .Z(n1163) );
  AND U1311 ( .A(n1166), .B(n1167), .Z(n1161) );
  AND U1312 ( .A(n1168), .B(p_input[8086]), .Z(n1167) );
  AND U1313 ( .A(p_input[7086]), .B(p_input[6086]), .Z(n1168) );
  AND U1314 ( .A(p_input[9086]), .B(p_input[86]), .Z(n1166) );
  AND U1315 ( .A(n1169), .B(n1170), .Z(o[869]) );
  AND U1316 ( .A(n1171), .B(n1172), .Z(n1170) );
  AND U1317 ( .A(n1173), .B(p_input[3869]), .Z(n1172) );
  AND U1318 ( .A(p_input[2869]), .B(p_input[1869]), .Z(n1173) );
  AND U1319 ( .A(p_input[5869]), .B(p_input[4869]), .Z(n1171) );
  AND U1320 ( .A(n1174), .B(n1175), .Z(n1169) );
  AND U1321 ( .A(n1176), .B(p_input[869]), .Z(n1175) );
  AND U1322 ( .A(p_input[7869]), .B(p_input[6869]), .Z(n1176) );
  AND U1323 ( .A(p_input[9869]), .B(p_input[8869]), .Z(n1174) );
  AND U1324 ( .A(n1177), .B(n1178), .Z(o[868]) );
  AND U1325 ( .A(n1179), .B(n1180), .Z(n1178) );
  AND U1326 ( .A(n1181), .B(p_input[3868]), .Z(n1180) );
  AND U1327 ( .A(p_input[2868]), .B(p_input[1868]), .Z(n1181) );
  AND U1328 ( .A(p_input[5868]), .B(p_input[4868]), .Z(n1179) );
  AND U1329 ( .A(n1182), .B(n1183), .Z(n1177) );
  AND U1330 ( .A(n1184), .B(p_input[868]), .Z(n1183) );
  AND U1331 ( .A(p_input[7868]), .B(p_input[6868]), .Z(n1184) );
  AND U1332 ( .A(p_input[9868]), .B(p_input[8868]), .Z(n1182) );
  AND U1333 ( .A(n1185), .B(n1186), .Z(o[867]) );
  AND U1334 ( .A(n1187), .B(n1188), .Z(n1186) );
  AND U1335 ( .A(n1189), .B(p_input[3867]), .Z(n1188) );
  AND U1336 ( .A(p_input[2867]), .B(p_input[1867]), .Z(n1189) );
  AND U1337 ( .A(p_input[5867]), .B(p_input[4867]), .Z(n1187) );
  AND U1338 ( .A(n1190), .B(n1191), .Z(n1185) );
  AND U1339 ( .A(n1192), .B(p_input[867]), .Z(n1191) );
  AND U1340 ( .A(p_input[7867]), .B(p_input[6867]), .Z(n1192) );
  AND U1341 ( .A(p_input[9867]), .B(p_input[8867]), .Z(n1190) );
  AND U1342 ( .A(n1193), .B(n1194), .Z(o[866]) );
  AND U1343 ( .A(n1195), .B(n1196), .Z(n1194) );
  AND U1344 ( .A(n1197), .B(p_input[3866]), .Z(n1196) );
  AND U1345 ( .A(p_input[2866]), .B(p_input[1866]), .Z(n1197) );
  AND U1346 ( .A(p_input[5866]), .B(p_input[4866]), .Z(n1195) );
  AND U1347 ( .A(n1198), .B(n1199), .Z(n1193) );
  AND U1348 ( .A(n1200), .B(p_input[866]), .Z(n1199) );
  AND U1349 ( .A(p_input[7866]), .B(p_input[6866]), .Z(n1200) );
  AND U1350 ( .A(p_input[9866]), .B(p_input[8866]), .Z(n1198) );
  AND U1351 ( .A(n1201), .B(n1202), .Z(o[865]) );
  AND U1352 ( .A(n1203), .B(n1204), .Z(n1202) );
  AND U1353 ( .A(n1205), .B(p_input[3865]), .Z(n1204) );
  AND U1354 ( .A(p_input[2865]), .B(p_input[1865]), .Z(n1205) );
  AND U1355 ( .A(p_input[5865]), .B(p_input[4865]), .Z(n1203) );
  AND U1356 ( .A(n1206), .B(n1207), .Z(n1201) );
  AND U1357 ( .A(n1208), .B(p_input[865]), .Z(n1207) );
  AND U1358 ( .A(p_input[7865]), .B(p_input[6865]), .Z(n1208) );
  AND U1359 ( .A(p_input[9865]), .B(p_input[8865]), .Z(n1206) );
  AND U1360 ( .A(n1209), .B(n1210), .Z(o[864]) );
  AND U1361 ( .A(n1211), .B(n1212), .Z(n1210) );
  AND U1362 ( .A(n1213), .B(p_input[3864]), .Z(n1212) );
  AND U1363 ( .A(p_input[2864]), .B(p_input[1864]), .Z(n1213) );
  AND U1364 ( .A(p_input[5864]), .B(p_input[4864]), .Z(n1211) );
  AND U1365 ( .A(n1214), .B(n1215), .Z(n1209) );
  AND U1366 ( .A(n1216), .B(p_input[864]), .Z(n1215) );
  AND U1367 ( .A(p_input[7864]), .B(p_input[6864]), .Z(n1216) );
  AND U1368 ( .A(p_input[9864]), .B(p_input[8864]), .Z(n1214) );
  AND U1369 ( .A(n1217), .B(n1218), .Z(o[863]) );
  AND U1370 ( .A(n1219), .B(n1220), .Z(n1218) );
  AND U1371 ( .A(n1221), .B(p_input[3863]), .Z(n1220) );
  AND U1372 ( .A(p_input[2863]), .B(p_input[1863]), .Z(n1221) );
  AND U1373 ( .A(p_input[5863]), .B(p_input[4863]), .Z(n1219) );
  AND U1374 ( .A(n1222), .B(n1223), .Z(n1217) );
  AND U1375 ( .A(n1224), .B(p_input[863]), .Z(n1223) );
  AND U1376 ( .A(p_input[7863]), .B(p_input[6863]), .Z(n1224) );
  AND U1377 ( .A(p_input[9863]), .B(p_input[8863]), .Z(n1222) );
  AND U1378 ( .A(n1225), .B(n1226), .Z(o[862]) );
  AND U1379 ( .A(n1227), .B(n1228), .Z(n1226) );
  AND U1380 ( .A(n1229), .B(p_input[3862]), .Z(n1228) );
  AND U1381 ( .A(p_input[2862]), .B(p_input[1862]), .Z(n1229) );
  AND U1382 ( .A(p_input[5862]), .B(p_input[4862]), .Z(n1227) );
  AND U1383 ( .A(n1230), .B(n1231), .Z(n1225) );
  AND U1384 ( .A(n1232), .B(p_input[862]), .Z(n1231) );
  AND U1385 ( .A(p_input[7862]), .B(p_input[6862]), .Z(n1232) );
  AND U1386 ( .A(p_input[9862]), .B(p_input[8862]), .Z(n1230) );
  AND U1387 ( .A(n1233), .B(n1234), .Z(o[861]) );
  AND U1388 ( .A(n1235), .B(n1236), .Z(n1234) );
  AND U1389 ( .A(n1237), .B(p_input[3861]), .Z(n1236) );
  AND U1390 ( .A(p_input[2861]), .B(p_input[1861]), .Z(n1237) );
  AND U1391 ( .A(p_input[5861]), .B(p_input[4861]), .Z(n1235) );
  AND U1392 ( .A(n1238), .B(n1239), .Z(n1233) );
  AND U1393 ( .A(n1240), .B(p_input[861]), .Z(n1239) );
  AND U1394 ( .A(p_input[7861]), .B(p_input[6861]), .Z(n1240) );
  AND U1395 ( .A(p_input[9861]), .B(p_input[8861]), .Z(n1238) );
  AND U1396 ( .A(n1241), .B(n1242), .Z(o[860]) );
  AND U1397 ( .A(n1243), .B(n1244), .Z(n1242) );
  AND U1398 ( .A(n1245), .B(p_input[3860]), .Z(n1244) );
  AND U1399 ( .A(p_input[2860]), .B(p_input[1860]), .Z(n1245) );
  AND U1400 ( .A(p_input[5860]), .B(p_input[4860]), .Z(n1243) );
  AND U1401 ( .A(n1246), .B(n1247), .Z(n1241) );
  AND U1402 ( .A(n1248), .B(p_input[860]), .Z(n1247) );
  AND U1403 ( .A(p_input[7860]), .B(p_input[6860]), .Z(n1248) );
  AND U1404 ( .A(p_input[9860]), .B(p_input[8860]), .Z(n1246) );
  AND U1405 ( .A(n1249), .B(n1250), .Z(o[85]) );
  AND U1406 ( .A(n1251), .B(n1252), .Z(n1250) );
  AND U1407 ( .A(n1253), .B(p_input[3085]), .Z(n1252) );
  AND U1408 ( .A(p_input[2085]), .B(p_input[1085]), .Z(n1253) );
  AND U1409 ( .A(p_input[5085]), .B(p_input[4085]), .Z(n1251) );
  AND U1410 ( .A(n1254), .B(n1255), .Z(n1249) );
  AND U1411 ( .A(n1256), .B(p_input[8085]), .Z(n1255) );
  AND U1412 ( .A(p_input[7085]), .B(p_input[6085]), .Z(n1256) );
  AND U1413 ( .A(p_input[9085]), .B(p_input[85]), .Z(n1254) );
  AND U1414 ( .A(n1257), .B(n1258), .Z(o[859]) );
  AND U1415 ( .A(n1259), .B(n1260), .Z(n1258) );
  AND U1416 ( .A(n1261), .B(p_input[3859]), .Z(n1260) );
  AND U1417 ( .A(p_input[2859]), .B(p_input[1859]), .Z(n1261) );
  AND U1418 ( .A(p_input[5859]), .B(p_input[4859]), .Z(n1259) );
  AND U1419 ( .A(n1262), .B(n1263), .Z(n1257) );
  AND U1420 ( .A(n1264), .B(p_input[859]), .Z(n1263) );
  AND U1421 ( .A(p_input[7859]), .B(p_input[6859]), .Z(n1264) );
  AND U1422 ( .A(p_input[9859]), .B(p_input[8859]), .Z(n1262) );
  AND U1423 ( .A(n1265), .B(n1266), .Z(o[858]) );
  AND U1424 ( .A(n1267), .B(n1268), .Z(n1266) );
  AND U1425 ( .A(n1269), .B(p_input[3858]), .Z(n1268) );
  AND U1426 ( .A(p_input[2858]), .B(p_input[1858]), .Z(n1269) );
  AND U1427 ( .A(p_input[5858]), .B(p_input[4858]), .Z(n1267) );
  AND U1428 ( .A(n1270), .B(n1271), .Z(n1265) );
  AND U1429 ( .A(n1272), .B(p_input[858]), .Z(n1271) );
  AND U1430 ( .A(p_input[7858]), .B(p_input[6858]), .Z(n1272) );
  AND U1431 ( .A(p_input[9858]), .B(p_input[8858]), .Z(n1270) );
  AND U1432 ( .A(n1273), .B(n1274), .Z(o[857]) );
  AND U1433 ( .A(n1275), .B(n1276), .Z(n1274) );
  AND U1434 ( .A(n1277), .B(p_input[3857]), .Z(n1276) );
  AND U1435 ( .A(p_input[2857]), .B(p_input[1857]), .Z(n1277) );
  AND U1436 ( .A(p_input[5857]), .B(p_input[4857]), .Z(n1275) );
  AND U1437 ( .A(n1278), .B(n1279), .Z(n1273) );
  AND U1438 ( .A(n1280), .B(p_input[857]), .Z(n1279) );
  AND U1439 ( .A(p_input[7857]), .B(p_input[6857]), .Z(n1280) );
  AND U1440 ( .A(p_input[9857]), .B(p_input[8857]), .Z(n1278) );
  AND U1441 ( .A(n1281), .B(n1282), .Z(o[856]) );
  AND U1442 ( .A(n1283), .B(n1284), .Z(n1282) );
  AND U1443 ( .A(n1285), .B(p_input[3856]), .Z(n1284) );
  AND U1444 ( .A(p_input[2856]), .B(p_input[1856]), .Z(n1285) );
  AND U1445 ( .A(p_input[5856]), .B(p_input[4856]), .Z(n1283) );
  AND U1446 ( .A(n1286), .B(n1287), .Z(n1281) );
  AND U1447 ( .A(n1288), .B(p_input[856]), .Z(n1287) );
  AND U1448 ( .A(p_input[7856]), .B(p_input[6856]), .Z(n1288) );
  AND U1449 ( .A(p_input[9856]), .B(p_input[8856]), .Z(n1286) );
  AND U1450 ( .A(n1289), .B(n1290), .Z(o[855]) );
  AND U1451 ( .A(n1291), .B(n1292), .Z(n1290) );
  AND U1452 ( .A(n1293), .B(p_input[3855]), .Z(n1292) );
  AND U1453 ( .A(p_input[2855]), .B(p_input[1855]), .Z(n1293) );
  AND U1454 ( .A(p_input[5855]), .B(p_input[4855]), .Z(n1291) );
  AND U1455 ( .A(n1294), .B(n1295), .Z(n1289) );
  AND U1456 ( .A(n1296), .B(p_input[855]), .Z(n1295) );
  AND U1457 ( .A(p_input[7855]), .B(p_input[6855]), .Z(n1296) );
  AND U1458 ( .A(p_input[9855]), .B(p_input[8855]), .Z(n1294) );
  AND U1459 ( .A(n1297), .B(n1298), .Z(o[854]) );
  AND U1460 ( .A(n1299), .B(n1300), .Z(n1298) );
  AND U1461 ( .A(n1301), .B(p_input[3854]), .Z(n1300) );
  AND U1462 ( .A(p_input[2854]), .B(p_input[1854]), .Z(n1301) );
  AND U1463 ( .A(p_input[5854]), .B(p_input[4854]), .Z(n1299) );
  AND U1464 ( .A(n1302), .B(n1303), .Z(n1297) );
  AND U1465 ( .A(n1304), .B(p_input[854]), .Z(n1303) );
  AND U1466 ( .A(p_input[7854]), .B(p_input[6854]), .Z(n1304) );
  AND U1467 ( .A(p_input[9854]), .B(p_input[8854]), .Z(n1302) );
  AND U1468 ( .A(n1305), .B(n1306), .Z(o[853]) );
  AND U1469 ( .A(n1307), .B(n1308), .Z(n1306) );
  AND U1470 ( .A(n1309), .B(p_input[3853]), .Z(n1308) );
  AND U1471 ( .A(p_input[2853]), .B(p_input[1853]), .Z(n1309) );
  AND U1472 ( .A(p_input[5853]), .B(p_input[4853]), .Z(n1307) );
  AND U1473 ( .A(n1310), .B(n1311), .Z(n1305) );
  AND U1474 ( .A(n1312), .B(p_input[853]), .Z(n1311) );
  AND U1475 ( .A(p_input[7853]), .B(p_input[6853]), .Z(n1312) );
  AND U1476 ( .A(p_input[9853]), .B(p_input[8853]), .Z(n1310) );
  AND U1477 ( .A(n1313), .B(n1314), .Z(o[852]) );
  AND U1478 ( .A(n1315), .B(n1316), .Z(n1314) );
  AND U1479 ( .A(n1317), .B(p_input[3852]), .Z(n1316) );
  AND U1480 ( .A(p_input[2852]), .B(p_input[1852]), .Z(n1317) );
  AND U1481 ( .A(p_input[5852]), .B(p_input[4852]), .Z(n1315) );
  AND U1482 ( .A(n1318), .B(n1319), .Z(n1313) );
  AND U1483 ( .A(n1320), .B(p_input[852]), .Z(n1319) );
  AND U1484 ( .A(p_input[7852]), .B(p_input[6852]), .Z(n1320) );
  AND U1485 ( .A(p_input[9852]), .B(p_input[8852]), .Z(n1318) );
  AND U1486 ( .A(n1321), .B(n1322), .Z(o[851]) );
  AND U1487 ( .A(n1323), .B(n1324), .Z(n1322) );
  AND U1488 ( .A(n1325), .B(p_input[3851]), .Z(n1324) );
  AND U1489 ( .A(p_input[2851]), .B(p_input[1851]), .Z(n1325) );
  AND U1490 ( .A(p_input[5851]), .B(p_input[4851]), .Z(n1323) );
  AND U1491 ( .A(n1326), .B(n1327), .Z(n1321) );
  AND U1492 ( .A(n1328), .B(p_input[851]), .Z(n1327) );
  AND U1493 ( .A(p_input[7851]), .B(p_input[6851]), .Z(n1328) );
  AND U1494 ( .A(p_input[9851]), .B(p_input[8851]), .Z(n1326) );
  AND U1495 ( .A(n1329), .B(n1330), .Z(o[850]) );
  AND U1496 ( .A(n1331), .B(n1332), .Z(n1330) );
  AND U1497 ( .A(n1333), .B(p_input[3850]), .Z(n1332) );
  AND U1498 ( .A(p_input[2850]), .B(p_input[1850]), .Z(n1333) );
  AND U1499 ( .A(p_input[5850]), .B(p_input[4850]), .Z(n1331) );
  AND U1500 ( .A(n1334), .B(n1335), .Z(n1329) );
  AND U1501 ( .A(n1336), .B(p_input[850]), .Z(n1335) );
  AND U1502 ( .A(p_input[7850]), .B(p_input[6850]), .Z(n1336) );
  AND U1503 ( .A(p_input[9850]), .B(p_input[8850]), .Z(n1334) );
  AND U1504 ( .A(n1337), .B(n1338), .Z(o[84]) );
  AND U1505 ( .A(n1339), .B(n1340), .Z(n1338) );
  AND U1506 ( .A(n1341), .B(p_input[3084]), .Z(n1340) );
  AND U1507 ( .A(p_input[2084]), .B(p_input[1084]), .Z(n1341) );
  AND U1508 ( .A(p_input[5084]), .B(p_input[4084]), .Z(n1339) );
  AND U1509 ( .A(n1342), .B(n1343), .Z(n1337) );
  AND U1510 ( .A(n1344), .B(p_input[8084]), .Z(n1343) );
  AND U1511 ( .A(p_input[7084]), .B(p_input[6084]), .Z(n1344) );
  AND U1512 ( .A(p_input[9084]), .B(p_input[84]), .Z(n1342) );
  AND U1513 ( .A(n1345), .B(n1346), .Z(o[849]) );
  AND U1514 ( .A(n1347), .B(n1348), .Z(n1346) );
  AND U1515 ( .A(n1349), .B(p_input[3849]), .Z(n1348) );
  AND U1516 ( .A(p_input[2849]), .B(p_input[1849]), .Z(n1349) );
  AND U1517 ( .A(p_input[5849]), .B(p_input[4849]), .Z(n1347) );
  AND U1518 ( .A(n1350), .B(n1351), .Z(n1345) );
  AND U1519 ( .A(n1352), .B(p_input[849]), .Z(n1351) );
  AND U1520 ( .A(p_input[7849]), .B(p_input[6849]), .Z(n1352) );
  AND U1521 ( .A(p_input[9849]), .B(p_input[8849]), .Z(n1350) );
  AND U1522 ( .A(n1353), .B(n1354), .Z(o[848]) );
  AND U1523 ( .A(n1355), .B(n1356), .Z(n1354) );
  AND U1524 ( .A(n1357), .B(p_input[3848]), .Z(n1356) );
  AND U1525 ( .A(p_input[2848]), .B(p_input[1848]), .Z(n1357) );
  AND U1526 ( .A(p_input[5848]), .B(p_input[4848]), .Z(n1355) );
  AND U1527 ( .A(n1358), .B(n1359), .Z(n1353) );
  AND U1528 ( .A(n1360), .B(p_input[848]), .Z(n1359) );
  AND U1529 ( .A(p_input[7848]), .B(p_input[6848]), .Z(n1360) );
  AND U1530 ( .A(p_input[9848]), .B(p_input[8848]), .Z(n1358) );
  AND U1531 ( .A(n1361), .B(n1362), .Z(o[847]) );
  AND U1532 ( .A(n1363), .B(n1364), .Z(n1362) );
  AND U1533 ( .A(n1365), .B(p_input[3847]), .Z(n1364) );
  AND U1534 ( .A(p_input[2847]), .B(p_input[1847]), .Z(n1365) );
  AND U1535 ( .A(p_input[5847]), .B(p_input[4847]), .Z(n1363) );
  AND U1536 ( .A(n1366), .B(n1367), .Z(n1361) );
  AND U1537 ( .A(n1368), .B(p_input[847]), .Z(n1367) );
  AND U1538 ( .A(p_input[7847]), .B(p_input[6847]), .Z(n1368) );
  AND U1539 ( .A(p_input[9847]), .B(p_input[8847]), .Z(n1366) );
  AND U1540 ( .A(n1369), .B(n1370), .Z(o[846]) );
  AND U1541 ( .A(n1371), .B(n1372), .Z(n1370) );
  AND U1542 ( .A(n1373), .B(p_input[3846]), .Z(n1372) );
  AND U1543 ( .A(p_input[2846]), .B(p_input[1846]), .Z(n1373) );
  AND U1544 ( .A(p_input[5846]), .B(p_input[4846]), .Z(n1371) );
  AND U1545 ( .A(n1374), .B(n1375), .Z(n1369) );
  AND U1546 ( .A(n1376), .B(p_input[846]), .Z(n1375) );
  AND U1547 ( .A(p_input[7846]), .B(p_input[6846]), .Z(n1376) );
  AND U1548 ( .A(p_input[9846]), .B(p_input[8846]), .Z(n1374) );
  AND U1549 ( .A(n1377), .B(n1378), .Z(o[845]) );
  AND U1550 ( .A(n1379), .B(n1380), .Z(n1378) );
  AND U1551 ( .A(n1381), .B(p_input[3845]), .Z(n1380) );
  AND U1552 ( .A(p_input[2845]), .B(p_input[1845]), .Z(n1381) );
  AND U1553 ( .A(p_input[5845]), .B(p_input[4845]), .Z(n1379) );
  AND U1554 ( .A(n1382), .B(n1383), .Z(n1377) );
  AND U1555 ( .A(n1384), .B(p_input[845]), .Z(n1383) );
  AND U1556 ( .A(p_input[7845]), .B(p_input[6845]), .Z(n1384) );
  AND U1557 ( .A(p_input[9845]), .B(p_input[8845]), .Z(n1382) );
  AND U1558 ( .A(n1385), .B(n1386), .Z(o[844]) );
  AND U1559 ( .A(n1387), .B(n1388), .Z(n1386) );
  AND U1560 ( .A(n1389), .B(p_input[3844]), .Z(n1388) );
  AND U1561 ( .A(p_input[2844]), .B(p_input[1844]), .Z(n1389) );
  AND U1562 ( .A(p_input[5844]), .B(p_input[4844]), .Z(n1387) );
  AND U1563 ( .A(n1390), .B(n1391), .Z(n1385) );
  AND U1564 ( .A(n1392), .B(p_input[844]), .Z(n1391) );
  AND U1565 ( .A(p_input[7844]), .B(p_input[6844]), .Z(n1392) );
  AND U1566 ( .A(p_input[9844]), .B(p_input[8844]), .Z(n1390) );
  AND U1567 ( .A(n1393), .B(n1394), .Z(o[843]) );
  AND U1568 ( .A(n1395), .B(n1396), .Z(n1394) );
  AND U1569 ( .A(n1397), .B(p_input[3843]), .Z(n1396) );
  AND U1570 ( .A(p_input[2843]), .B(p_input[1843]), .Z(n1397) );
  AND U1571 ( .A(p_input[5843]), .B(p_input[4843]), .Z(n1395) );
  AND U1572 ( .A(n1398), .B(n1399), .Z(n1393) );
  AND U1573 ( .A(n1400), .B(p_input[843]), .Z(n1399) );
  AND U1574 ( .A(p_input[7843]), .B(p_input[6843]), .Z(n1400) );
  AND U1575 ( .A(p_input[9843]), .B(p_input[8843]), .Z(n1398) );
  AND U1576 ( .A(n1401), .B(n1402), .Z(o[842]) );
  AND U1577 ( .A(n1403), .B(n1404), .Z(n1402) );
  AND U1578 ( .A(n1405), .B(p_input[3842]), .Z(n1404) );
  AND U1579 ( .A(p_input[2842]), .B(p_input[1842]), .Z(n1405) );
  AND U1580 ( .A(p_input[5842]), .B(p_input[4842]), .Z(n1403) );
  AND U1581 ( .A(n1406), .B(n1407), .Z(n1401) );
  AND U1582 ( .A(n1408), .B(p_input[842]), .Z(n1407) );
  AND U1583 ( .A(p_input[7842]), .B(p_input[6842]), .Z(n1408) );
  AND U1584 ( .A(p_input[9842]), .B(p_input[8842]), .Z(n1406) );
  AND U1585 ( .A(n1409), .B(n1410), .Z(o[841]) );
  AND U1586 ( .A(n1411), .B(n1412), .Z(n1410) );
  AND U1587 ( .A(n1413), .B(p_input[3841]), .Z(n1412) );
  AND U1588 ( .A(p_input[2841]), .B(p_input[1841]), .Z(n1413) );
  AND U1589 ( .A(p_input[5841]), .B(p_input[4841]), .Z(n1411) );
  AND U1590 ( .A(n1414), .B(n1415), .Z(n1409) );
  AND U1591 ( .A(n1416), .B(p_input[841]), .Z(n1415) );
  AND U1592 ( .A(p_input[7841]), .B(p_input[6841]), .Z(n1416) );
  AND U1593 ( .A(p_input[9841]), .B(p_input[8841]), .Z(n1414) );
  AND U1594 ( .A(n1417), .B(n1418), .Z(o[840]) );
  AND U1595 ( .A(n1419), .B(n1420), .Z(n1418) );
  AND U1596 ( .A(n1421), .B(p_input[3840]), .Z(n1420) );
  AND U1597 ( .A(p_input[2840]), .B(p_input[1840]), .Z(n1421) );
  AND U1598 ( .A(p_input[5840]), .B(p_input[4840]), .Z(n1419) );
  AND U1599 ( .A(n1422), .B(n1423), .Z(n1417) );
  AND U1600 ( .A(n1424), .B(p_input[840]), .Z(n1423) );
  AND U1601 ( .A(p_input[7840]), .B(p_input[6840]), .Z(n1424) );
  AND U1602 ( .A(p_input[9840]), .B(p_input[8840]), .Z(n1422) );
  AND U1603 ( .A(n1425), .B(n1426), .Z(o[83]) );
  AND U1604 ( .A(n1427), .B(n1428), .Z(n1426) );
  AND U1605 ( .A(n1429), .B(p_input[3083]), .Z(n1428) );
  AND U1606 ( .A(p_input[2083]), .B(p_input[1083]), .Z(n1429) );
  AND U1607 ( .A(p_input[5083]), .B(p_input[4083]), .Z(n1427) );
  AND U1608 ( .A(n1430), .B(n1431), .Z(n1425) );
  AND U1609 ( .A(n1432), .B(p_input[8083]), .Z(n1431) );
  AND U1610 ( .A(p_input[7083]), .B(p_input[6083]), .Z(n1432) );
  AND U1611 ( .A(p_input[9083]), .B(p_input[83]), .Z(n1430) );
  AND U1612 ( .A(n1433), .B(n1434), .Z(o[839]) );
  AND U1613 ( .A(n1435), .B(n1436), .Z(n1434) );
  AND U1614 ( .A(n1437), .B(p_input[3839]), .Z(n1436) );
  AND U1615 ( .A(p_input[2839]), .B(p_input[1839]), .Z(n1437) );
  AND U1616 ( .A(p_input[5839]), .B(p_input[4839]), .Z(n1435) );
  AND U1617 ( .A(n1438), .B(n1439), .Z(n1433) );
  AND U1618 ( .A(n1440), .B(p_input[839]), .Z(n1439) );
  AND U1619 ( .A(p_input[7839]), .B(p_input[6839]), .Z(n1440) );
  AND U1620 ( .A(p_input[9839]), .B(p_input[8839]), .Z(n1438) );
  AND U1621 ( .A(n1441), .B(n1442), .Z(o[838]) );
  AND U1622 ( .A(n1443), .B(n1444), .Z(n1442) );
  AND U1623 ( .A(n1445), .B(p_input[3838]), .Z(n1444) );
  AND U1624 ( .A(p_input[2838]), .B(p_input[1838]), .Z(n1445) );
  AND U1625 ( .A(p_input[5838]), .B(p_input[4838]), .Z(n1443) );
  AND U1626 ( .A(n1446), .B(n1447), .Z(n1441) );
  AND U1627 ( .A(n1448), .B(p_input[838]), .Z(n1447) );
  AND U1628 ( .A(p_input[7838]), .B(p_input[6838]), .Z(n1448) );
  AND U1629 ( .A(p_input[9838]), .B(p_input[8838]), .Z(n1446) );
  AND U1630 ( .A(n1449), .B(n1450), .Z(o[837]) );
  AND U1631 ( .A(n1451), .B(n1452), .Z(n1450) );
  AND U1632 ( .A(n1453), .B(p_input[3837]), .Z(n1452) );
  AND U1633 ( .A(p_input[2837]), .B(p_input[1837]), .Z(n1453) );
  AND U1634 ( .A(p_input[5837]), .B(p_input[4837]), .Z(n1451) );
  AND U1635 ( .A(n1454), .B(n1455), .Z(n1449) );
  AND U1636 ( .A(n1456), .B(p_input[837]), .Z(n1455) );
  AND U1637 ( .A(p_input[7837]), .B(p_input[6837]), .Z(n1456) );
  AND U1638 ( .A(p_input[9837]), .B(p_input[8837]), .Z(n1454) );
  AND U1639 ( .A(n1457), .B(n1458), .Z(o[836]) );
  AND U1640 ( .A(n1459), .B(n1460), .Z(n1458) );
  AND U1641 ( .A(n1461), .B(p_input[3836]), .Z(n1460) );
  AND U1642 ( .A(p_input[2836]), .B(p_input[1836]), .Z(n1461) );
  AND U1643 ( .A(p_input[5836]), .B(p_input[4836]), .Z(n1459) );
  AND U1644 ( .A(n1462), .B(n1463), .Z(n1457) );
  AND U1645 ( .A(n1464), .B(p_input[836]), .Z(n1463) );
  AND U1646 ( .A(p_input[7836]), .B(p_input[6836]), .Z(n1464) );
  AND U1647 ( .A(p_input[9836]), .B(p_input[8836]), .Z(n1462) );
  AND U1648 ( .A(n1465), .B(n1466), .Z(o[835]) );
  AND U1649 ( .A(n1467), .B(n1468), .Z(n1466) );
  AND U1650 ( .A(n1469), .B(p_input[3835]), .Z(n1468) );
  AND U1651 ( .A(p_input[2835]), .B(p_input[1835]), .Z(n1469) );
  AND U1652 ( .A(p_input[5835]), .B(p_input[4835]), .Z(n1467) );
  AND U1653 ( .A(n1470), .B(n1471), .Z(n1465) );
  AND U1654 ( .A(n1472), .B(p_input[835]), .Z(n1471) );
  AND U1655 ( .A(p_input[7835]), .B(p_input[6835]), .Z(n1472) );
  AND U1656 ( .A(p_input[9835]), .B(p_input[8835]), .Z(n1470) );
  AND U1657 ( .A(n1473), .B(n1474), .Z(o[834]) );
  AND U1658 ( .A(n1475), .B(n1476), .Z(n1474) );
  AND U1659 ( .A(n1477), .B(p_input[3834]), .Z(n1476) );
  AND U1660 ( .A(p_input[2834]), .B(p_input[1834]), .Z(n1477) );
  AND U1661 ( .A(p_input[5834]), .B(p_input[4834]), .Z(n1475) );
  AND U1662 ( .A(n1478), .B(n1479), .Z(n1473) );
  AND U1663 ( .A(n1480), .B(p_input[834]), .Z(n1479) );
  AND U1664 ( .A(p_input[7834]), .B(p_input[6834]), .Z(n1480) );
  AND U1665 ( .A(p_input[9834]), .B(p_input[8834]), .Z(n1478) );
  AND U1666 ( .A(n1481), .B(n1482), .Z(o[833]) );
  AND U1667 ( .A(n1483), .B(n1484), .Z(n1482) );
  AND U1668 ( .A(n1485), .B(p_input[3833]), .Z(n1484) );
  AND U1669 ( .A(p_input[2833]), .B(p_input[1833]), .Z(n1485) );
  AND U1670 ( .A(p_input[5833]), .B(p_input[4833]), .Z(n1483) );
  AND U1671 ( .A(n1486), .B(n1487), .Z(n1481) );
  AND U1672 ( .A(n1488), .B(p_input[833]), .Z(n1487) );
  AND U1673 ( .A(p_input[7833]), .B(p_input[6833]), .Z(n1488) );
  AND U1674 ( .A(p_input[9833]), .B(p_input[8833]), .Z(n1486) );
  AND U1675 ( .A(n1489), .B(n1490), .Z(o[832]) );
  AND U1676 ( .A(n1491), .B(n1492), .Z(n1490) );
  AND U1677 ( .A(n1493), .B(p_input[3832]), .Z(n1492) );
  AND U1678 ( .A(p_input[2832]), .B(p_input[1832]), .Z(n1493) );
  AND U1679 ( .A(p_input[5832]), .B(p_input[4832]), .Z(n1491) );
  AND U1680 ( .A(n1494), .B(n1495), .Z(n1489) );
  AND U1681 ( .A(n1496), .B(p_input[832]), .Z(n1495) );
  AND U1682 ( .A(p_input[7832]), .B(p_input[6832]), .Z(n1496) );
  AND U1683 ( .A(p_input[9832]), .B(p_input[8832]), .Z(n1494) );
  AND U1684 ( .A(n1497), .B(n1498), .Z(o[831]) );
  AND U1685 ( .A(n1499), .B(n1500), .Z(n1498) );
  AND U1686 ( .A(n1501), .B(p_input[3831]), .Z(n1500) );
  AND U1687 ( .A(p_input[2831]), .B(p_input[1831]), .Z(n1501) );
  AND U1688 ( .A(p_input[5831]), .B(p_input[4831]), .Z(n1499) );
  AND U1689 ( .A(n1502), .B(n1503), .Z(n1497) );
  AND U1690 ( .A(n1504), .B(p_input[831]), .Z(n1503) );
  AND U1691 ( .A(p_input[7831]), .B(p_input[6831]), .Z(n1504) );
  AND U1692 ( .A(p_input[9831]), .B(p_input[8831]), .Z(n1502) );
  AND U1693 ( .A(n1505), .B(n1506), .Z(o[830]) );
  AND U1694 ( .A(n1507), .B(n1508), .Z(n1506) );
  AND U1695 ( .A(n1509), .B(p_input[3830]), .Z(n1508) );
  AND U1696 ( .A(p_input[2830]), .B(p_input[1830]), .Z(n1509) );
  AND U1697 ( .A(p_input[5830]), .B(p_input[4830]), .Z(n1507) );
  AND U1698 ( .A(n1510), .B(n1511), .Z(n1505) );
  AND U1699 ( .A(n1512), .B(p_input[830]), .Z(n1511) );
  AND U1700 ( .A(p_input[7830]), .B(p_input[6830]), .Z(n1512) );
  AND U1701 ( .A(p_input[9830]), .B(p_input[8830]), .Z(n1510) );
  AND U1702 ( .A(n1513), .B(n1514), .Z(o[82]) );
  AND U1703 ( .A(n1515), .B(n1516), .Z(n1514) );
  AND U1704 ( .A(n1517), .B(p_input[3082]), .Z(n1516) );
  AND U1705 ( .A(p_input[2082]), .B(p_input[1082]), .Z(n1517) );
  AND U1706 ( .A(p_input[5082]), .B(p_input[4082]), .Z(n1515) );
  AND U1707 ( .A(n1518), .B(n1519), .Z(n1513) );
  AND U1708 ( .A(n1520), .B(p_input[8082]), .Z(n1519) );
  AND U1709 ( .A(p_input[7082]), .B(p_input[6082]), .Z(n1520) );
  AND U1710 ( .A(p_input[9082]), .B(p_input[82]), .Z(n1518) );
  AND U1711 ( .A(n1521), .B(n1522), .Z(o[829]) );
  AND U1712 ( .A(n1523), .B(n1524), .Z(n1522) );
  AND U1713 ( .A(n1525), .B(p_input[3829]), .Z(n1524) );
  AND U1714 ( .A(p_input[2829]), .B(p_input[1829]), .Z(n1525) );
  AND U1715 ( .A(p_input[5829]), .B(p_input[4829]), .Z(n1523) );
  AND U1716 ( .A(n1526), .B(n1527), .Z(n1521) );
  AND U1717 ( .A(n1528), .B(p_input[829]), .Z(n1527) );
  AND U1718 ( .A(p_input[7829]), .B(p_input[6829]), .Z(n1528) );
  AND U1719 ( .A(p_input[9829]), .B(p_input[8829]), .Z(n1526) );
  AND U1720 ( .A(n1529), .B(n1530), .Z(o[828]) );
  AND U1721 ( .A(n1531), .B(n1532), .Z(n1530) );
  AND U1722 ( .A(n1533), .B(p_input[3828]), .Z(n1532) );
  AND U1723 ( .A(p_input[2828]), .B(p_input[1828]), .Z(n1533) );
  AND U1724 ( .A(p_input[5828]), .B(p_input[4828]), .Z(n1531) );
  AND U1725 ( .A(n1534), .B(n1535), .Z(n1529) );
  AND U1726 ( .A(n1536), .B(p_input[828]), .Z(n1535) );
  AND U1727 ( .A(p_input[7828]), .B(p_input[6828]), .Z(n1536) );
  AND U1728 ( .A(p_input[9828]), .B(p_input[8828]), .Z(n1534) );
  AND U1729 ( .A(n1537), .B(n1538), .Z(o[827]) );
  AND U1730 ( .A(n1539), .B(n1540), .Z(n1538) );
  AND U1731 ( .A(n1541), .B(p_input[3827]), .Z(n1540) );
  AND U1732 ( .A(p_input[2827]), .B(p_input[1827]), .Z(n1541) );
  AND U1733 ( .A(p_input[5827]), .B(p_input[4827]), .Z(n1539) );
  AND U1734 ( .A(n1542), .B(n1543), .Z(n1537) );
  AND U1735 ( .A(n1544), .B(p_input[827]), .Z(n1543) );
  AND U1736 ( .A(p_input[7827]), .B(p_input[6827]), .Z(n1544) );
  AND U1737 ( .A(p_input[9827]), .B(p_input[8827]), .Z(n1542) );
  AND U1738 ( .A(n1545), .B(n1546), .Z(o[826]) );
  AND U1739 ( .A(n1547), .B(n1548), .Z(n1546) );
  AND U1740 ( .A(n1549), .B(p_input[3826]), .Z(n1548) );
  AND U1741 ( .A(p_input[2826]), .B(p_input[1826]), .Z(n1549) );
  AND U1742 ( .A(p_input[5826]), .B(p_input[4826]), .Z(n1547) );
  AND U1743 ( .A(n1550), .B(n1551), .Z(n1545) );
  AND U1744 ( .A(n1552), .B(p_input[826]), .Z(n1551) );
  AND U1745 ( .A(p_input[7826]), .B(p_input[6826]), .Z(n1552) );
  AND U1746 ( .A(p_input[9826]), .B(p_input[8826]), .Z(n1550) );
  AND U1747 ( .A(n1553), .B(n1554), .Z(o[825]) );
  AND U1748 ( .A(n1555), .B(n1556), .Z(n1554) );
  AND U1749 ( .A(n1557), .B(p_input[3825]), .Z(n1556) );
  AND U1750 ( .A(p_input[2825]), .B(p_input[1825]), .Z(n1557) );
  AND U1751 ( .A(p_input[5825]), .B(p_input[4825]), .Z(n1555) );
  AND U1752 ( .A(n1558), .B(n1559), .Z(n1553) );
  AND U1753 ( .A(n1560), .B(p_input[825]), .Z(n1559) );
  AND U1754 ( .A(p_input[7825]), .B(p_input[6825]), .Z(n1560) );
  AND U1755 ( .A(p_input[9825]), .B(p_input[8825]), .Z(n1558) );
  AND U1756 ( .A(n1561), .B(n1562), .Z(o[824]) );
  AND U1757 ( .A(n1563), .B(n1564), .Z(n1562) );
  AND U1758 ( .A(n1565), .B(p_input[3824]), .Z(n1564) );
  AND U1759 ( .A(p_input[2824]), .B(p_input[1824]), .Z(n1565) );
  AND U1760 ( .A(p_input[5824]), .B(p_input[4824]), .Z(n1563) );
  AND U1761 ( .A(n1566), .B(n1567), .Z(n1561) );
  AND U1762 ( .A(n1568), .B(p_input[824]), .Z(n1567) );
  AND U1763 ( .A(p_input[7824]), .B(p_input[6824]), .Z(n1568) );
  AND U1764 ( .A(p_input[9824]), .B(p_input[8824]), .Z(n1566) );
  AND U1765 ( .A(n1569), .B(n1570), .Z(o[823]) );
  AND U1766 ( .A(n1571), .B(n1572), .Z(n1570) );
  AND U1767 ( .A(n1573), .B(p_input[3823]), .Z(n1572) );
  AND U1768 ( .A(p_input[2823]), .B(p_input[1823]), .Z(n1573) );
  AND U1769 ( .A(p_input[5823]), .B(p_input[4823]), .Z(n1571) );
  AND U1770 ( .A(n1574), .B(n1575), .Z(n1569) );
  AND U1771 ( .A(n1576), .B(p_input[823]), .Z(n1575) );
  AND U1772 ( .A(p_input[7823]), .B(p_input[6823]), .Z(n1576) );
  AND U1773 ( .A(p_input[9823]), .B(p_input[8823]), .Z(n1574) );
  AND U1774 ( .A(n1577), .B(n1578), .Z(o[822]) );
  AND U1775 ( .A(n1579), .B(n1580), .Z(n1578) );
  AND U1776 ( .A(n1581), .B(p_input[3822]), .Z(n1580) );
  AND U1777 ( .A(p_input[2822]), .B(p_input[1822]), .Z(n1581) );
  AND U1778 ( .A(p_input[5822]), .B(p_input[4822]), .Z(n1579) );
  AND U1779 ( .A(n1582), .B(n1583), .Z(n1577) );
  AND U1780 ( .A(n1584), .B(p_input[822]), .Z(n1583) );
  AND U1781 ( .A(p_input[7822]), .B(p_input[6822]), .Z(n1584) );
  AND U1782 ( .A(p_input[9822]), .B(p_input[8822]), .Z(n1582) );
  AND U1783 ( .A(n1585), .B(n1586), .Z(o[821]) );
  AND U1784 ( .A(n1587), .B(n1588), .Z(n1586) );
  AND U1785 ( .A(n1589), .B(p_input[3821]), .Z(n1588) );
  AND U1786 ( .A(p_input[2821]), .B(p_input[1821]), .Z(n1589) );
  AND U1787 ( .A(p_input[5821]), .B(p_input[4821]), .Z(n1587) );
  AND U1788 ( .A(n1590), .B(n1591), .Z(n1585) );
  AND U1789 ( .A(n1592), .B(p_input[821]), .Z(n1591) );
  AND U1790 ( .A(p_input[7821]), .B(p_input[6821]), .Z(n1592) );
  AND U1791 ( .A(p_input[9821]), .B(p_input[8821]), .Z(n1590) );
  AND U1792 ( .A(n1593), .B(n1594), .Z(o[820]) );
  AND U1793 ( .A(n1595), .B(n1596), .Z(n1594) );
  AND U1794 ( .A(n1597), .B(p_input[3820]), .Z(n1596) );
  AND U1795 ( .A(p_input[2820]), .B(p_input[1820]), .Z(n1597) );
  AND U1796 ( .A(p_input[5820]), .B(p_input[4820]), .Z(n1595) );
  AND U1797 ( .A(n1598), .B(n1599), .Z(n1593) );
  AND U1798 ( .A(n1600), .B(p_input[820]), .Z(n1599) );
  AND U1799 ( .A(p_input[7820]), .B(p_input[6820]), .Z(n1600) );
  AND U1800 ( .A(p_input[9820]), .B(p_input[8820]), .Z(n1598) );
  AND U1801 ( .A(n1601), .B(n1602), .Z(o[81]) );
  AND U1802 ( .A(n1603), .B(n1604), .Z(n1602) );
  AND U1803 ( .A(n1605), .B(p_input[3081]), .Z(n1604) );
  AND U1804 ( .A(p_input[2081]), .B(p_input[1081]), .Z(n1605) );
  AND U1805 ( .A(p_input[5081]), .B(p_input[4081]), .Z(n1603) );
  AND U1806 ( .A(n1606), .B(n1607), .Z(n1601) );
  AND U1807 ( .A(n1608), .B(p_input[8081]), .Z(n1607) );
  AND U1808 ( .A(p_input[7081]), .B(p_input[6081]), .Z(n1608) );
  AND U1809 ( .A(p_input[9081]), .B(p_input[81]), .Z(n1606) );
  AND U1810 ( .A(n1609), .B(n1610), .Z(o[819]) );
  AND U1811 ( .A(n1611), .B(n1612), .Z(n1610) );
  AND U1812 ( .A(n1613), .B(p_input[3819]), .Z(n1612) );
  AND U1813 ( .A(p_input[2819]), .B(p_input[1819]), .Z(n1613) );
  AND U1814 ( .A(p_input[5819]), .B(p_input[4819]), .Z(n1611) );
  AND U1815 ( .A(n1614), .B(n1615), .Z(n1609) );
  AND U1816 ( .A(n1616), .B(p_input[819]), .Z(n1615) );
  AND U1817 ( .A(p_input[7819]), .B(p_input[6819]), .Z(n1616) );
  AND U1818 ( .A(p_input[9819]), .B(p_input[8819]), .Z(n1614) );
  AND U1819 ( .A(n1617), .B(n1618), .Z(o[818]) );
  AND U1820 ( .A(n1619), .B(n1620), .Z(n1618) );
  AND U1821 ( .A(n1621), .B(p_input[3818]), .Z(n1620) );
  AND U1822 ( .A(p_input[2818]), .B(p_input[1818]), .Z(n1621) );
  AND U1823 ( .A(p_input[5818]), .B(p_input[4818]), .Z(n1619) );
  AND U1824 ( .A(n1622), .B(n1623), .Z(n1617) );
  AND U1825 ( .A(n1624), .B(p_input[818]), .Z(n1623) );
  AND U1826 ( .A(p_input[7818]), .B(p_input[6818]), .Z(n1624) );
  AND U1827 ( .A(p_input[9818]), .B(p_input[8818]), .Z(n1622) );
  AND U1828 ( .A(n1625), .B(n1626), .Z(o[817]) );
  AND U1829 ( .A(n1627), .B(n1628), .Z(n1626) );
  AND U1830 ( .A(n1629), .B(p_input[3817]), .Z(n1628) );
  AND U1831 ( .A(p_input[2817]), .B(p_input[1817]), .Z(n1629) );
  AND U1832 ( .A(p_input[5817]), .B(p_input[4817]), .Z(n1627) );
  AND U1833 ( .A(n1630), .B(n1631), .Z(n1625) );
  AND U1834 ( .A(n1632), .B(p_input[817]), .Z(n1631) );
  AND U1835 ( .A(p_input[7817]), .B(p_input[6817]), .Z(n1632) );
  AND U1836 ( .A(p_input[9817]), .B(p_input[8817]), .Z(n1630) );
  AND U1837 ( .A(n1633), .B(n1634), .Z(o[816]) );
  AND U1838 ( .A(n1635), .B(n1636), .Z(n1634) );
  AND U1839 ( .A(n1637), .B(p_input[3816]), .Z(n1636) );
  AND U1840 ( .A(p_input[2816]), .B(p_input[1816]), .Z(n1637) );
  AND U1841 ( .A(p_input[5816]), .B(p_input[4816]), .Z(n1635) );
  AND U1842 ( .A(n1638), .B(n1639), .Z(n1633) );
  AND U1843 ( .A(n1640), .B(p_input[816]), .Z(n1639) );
  AND U1844 ( .A(p_input[7816]), .B(p_input[6816]), .Z(n1640) );
  AND U1845 ( .A(p_input[9816]), .B(p_input[8816]), .Z(n1638) );
  AND U1846 ( .A(n1641), .B(n1642), .Z(o[815]) );
  AND U1847 ( .A(n1643), .B(n1644), .Z(n1642) );
  AND U1848 ( .A(n1645), .B(p_input[3815]), .Z(n1644) );
  AND U1849 ( .A(p_input[2815]), .B(p_input[1815]), .Z(n1645) );
  AND U1850 ( .A(p_input[5815]), .B(p_input[4815]), .Z(n1643) );
  AND U1851 ( .A(n1646), .B(n1647), .Z(n1641) );
  AND U1852 ( .A(n1648), .B(p_input[815]), .Z(n1647) );
  AND U1853 ( .A(p_input[7815]), .B(p_input[6815]), .Z(n1648) );
  AND U1854 ( .A(p_input[9815]), .B(p_input[8815]), .Z(n1646) );
  AND U1855 ( .A(n1649), .B(n1650), .Z(o[814]) );
  AND U1856 ( .A(n1651), .B(n1652), .Z(n1650) );
  AND U1857 ( .A(n1653), .B(p_input[3814]), .Z(n1652) );
  AND U1858 ( .A(p_input[2814]), .B(p_input[1814]), .Z(n1653) );
  AND U1859 ( .A(p_input[5814]), .B(p_input[4814]), .Z(n1651) );
  AND U1860 ( .A(n1654), .B(n1655), .Z(n1649) );
  AND U1861 ( .A(n1656), .B(p_input[814]), .Z(n1655) );
  AND U1862 ( .A(p_input[7814]), .B(p_input[6814]), .Z(n1656) );
  AND U1863 ( .A(p_input[9814]), .B(p_input[8814]), .Z(n1654) );
  AND U1864 ( .A(n1657), .B(n1658), .Z(o[813]) );
  AND U1865 ( .A(n1659), .B(n1660), .Z(n1658) );
  AND U1866 ( .A(n1661), .B(p_input[3813]), .Z(n1660) );
  AND U1867 ( .A(p_input[2813]), .B(p_input[1813]), .Z(n1661) );
  AND U1868 ( .A(p_input[5813]), .B(p_input[4813]), .Z(n1659) );
  AND U1869 ( .A(n1662), .B(n1663), .Z(n1657) );
  AND U1870 ( .A(n1664), .B(p_input[813]), .Z(n1663) );
  AND U1871 ( .A(p_input[7813]), .B(p_input[6813]), .Z(n1664) );
  AND U1872 ( .A(p_input[9813]), .B(p_input[8813]), .Z(n1662) );
  AND U1873 ( .A(n1665), .B(n1666), .Z(o[812]) );
  AND U1874 ( .A(n1667), .B(n1668), .Z(n1666) );
  AND U1875 ( .A(n1669), .B(p_input[3812]), .Z(n1668) );
  AND U1876 ( .A(p_input[2812]), .B(p_input[1812]), .Z(n1669) );
  AND U1877 ( .A(p_input[5812]), .B(p_input[4812]), .Z(n1667) );
  AND U1878 ( .A(n1670), .B(n1671), .Z(n1665) );
  AND U1879 ( .A(n1672), .B(p_input[812]), .Z(n1671) );
  AND U1880 ( .A(p_input[7812]), .B(p_input[6812]), .Z(n1672) );
  AND U1881 ( .A(p_input[9812]), .B(p_input[8812]), .Z(n1670) );
  AND U1882 ( .A(n1673), .B(n1674), .Z(o[811]) );
  AND U1883 ( .A(n1675), .B(n1676), .Z(n1674) );
  AND U1884 ( .A(n1677), .B(p_input[3811]), .Z(n1676) );
  AND U1885 ( .A(p_input[2811]), .B(p_input[1811]), .Z(n1677) );
  AND U1886 ( .A(p_input[5811]), .B(p_input[4811]), .Z(n1675) );
  AND U1887 ( .A(n1678), .B(n1679), .Z(n1673) );
  AND U1888 ( .A(n1680), .B(p_input[811]), .Z(n1679) );
  AND U1889 ( .A(p_input[7811]), .B(p_input[6811]), .Z(n1680) );
  AND U1890 ( .A(p_input[9811]), .B(p_input[8811]), .Z(n1678) );
  AND U1891 ( .A(n1681), .B(n1682), .Z(o[810]) );
  AND U1892 ( .A(n1683), .B(n1684), .Z(n1682) );
  AND U1893 ( .A(n1685), .B(p_input[3810]), .Z(n1684) );
  AND U1894 ( .A(p_input[2810]), .B(p_input[1810]), .Z(n1685) );
  AND U1895 ( .A(p_input[5810]), .B(p_input[4810]), .Z(n1683) );
  AND U1896 ( .A(n1686), .B(n1687), .Z(n1681) );
  AND U1897 ( .A(n1688), .B(p_input[810]), .Z(n1687) );
  AND U1898 ( .A(p_input[7810]), .B(p_input[6810]), .Z(n1688) );
  AND U1899 ( .A(p_input[9810]), .B(p_input[8810]), .Z(n1686) );
  AND U1900 ( .A(n1689), .B(n1690), .Z(o[80]) );
  AND U1901 ( .A(n1691), .B(n1692), .Z(n1690) );
  AND U1902 ( .A(n1693), .B(p_input[3080]), .Z(n1692) );
  AND U1903 ( .A(p_input[2080]), .B(p_input[1080]), .Z(n1693) );
  AND U1904 ( .A(p_input[5080]), .B(p_input[4080]), .Z(n1691) );
  AND U1905 ( .A(n1694), .B(n1695), .Z(n1689) );
  AND U1906 ( .A(n1696), .B(p_input[8080]), .Z(n1695) );
  AND U1907 ( .A(p_input[7080]), .B(p_input[6080]), .Z(n1696) );
  AND U1908 ( .A(p_input[9080]), .B(p_input[80]), .Z(n1694) );
  AND U1909 ( .A(n1697), .B(n1698), .Z(o[809]) );
  AND U1910 ( .A(n1699), .B(n1700), .Z(n1698) );
  AND U1911 ( .A(n1701), .B(p_input[3809]), .Z(n1700) );
  AND U1912 ( .A(p_input[2809]), .B(p_input[1809]), .Z(n1701) );
  AND U1913 ( .A(p_input[5809]), .B(p_input[4809]), .Z(n1699) );
  AND U1914 ( .A(n1702), .B(n1703), .Z(n1697) );
  AND U1915 ( .A(n1704), .B(p_input[809]), .Z(n1703) );
  AND U1916 ( .A(p_input[7809]), .B(p_input[6809]), .Z(n1704) );
  AND U1917 ( .A(p_input[9809]), .B(p_input[8809]), .Z(n1702) );
  AND U1918 ( .A(n1705), .B(n1706), .Z(o[808]) );
  AND U1919 ( .A(n1707), .B(n1708), .Z(n1706) );
  AND U1920 ( .A(n1709), .B(p_input[3808]), .Z(n1708) );
  AND U1921 ( .A(p_input[2808]), .B(p_input[1808]), .Z(n1709) );
  AND U1922 ( .A(p_input[5808]), .B(p_input[4808]), .Z(n1707) );
  AND U1923 ( .A(n1710), .B(n1711), .Z(n1705) );
  AND U1924 ( .A(n1712), .B(p_input[808]), .Z(n1711) );
  AND U1925 ( .A(p_input[7808]), .B(p_input[6808]), .Z(n1712) );
  AND U1926 ( .A(p_input[9808]), .B(p_input[8808]), .Z(n1710) );
  AND U1927 ( .A(n1713), .B(n1714), .Z(o[807]) );
  AND U1928 ( .A(n1715), .B(n1716), .Z(n1714) );
  AND U1929 ( .A(n1717), .B(p_input[3807]), .Z(n1716) );
  AND U1930 ( .A(p_input[2807]), .B(p_input[1807]), .Z(n1717) );
  AND U1931 ( .A(p_input[5807]), .B(p_input[4807]), .Z(n1715) );
  AND U1932 ( .A(n1718), .B(n1719), .Z(n1713) );
  AND U1933 ( .A(n1720), .B(p_input[807]), .Z(n1719) );
  AND U1934 ( .A(p_input[7807]), .B(p_input[6807]), .Z(n1720) );
  AND U1935 ( .A(p_input[9807]), .B(p_input[8807]), .Z(n1718) );
  AND U1936 ( .A(n1721), .B(n1722), .Z(o[806]) );
  AND U1937 ( .A(n1723), .B(n1724), .Z(n1722) );
  AND U1938 ( .A(n1725), .B(p_input[3806]), .Z(n1724) );
  AND U1939 ( .A(p_input[2806]), .B(p_input[1806]), .Z(n1725) );
  AND U1940 ( .A(p_input[5806]), .B(p_input[4806]), .Z(n1723) );
  AND U1941 ( .A(n1726), .B(n1727), .Z(n1721) );
  AND U1942 ( .A(n1728), .B(p_input[806]), .Z(n1727) );
  AND U1943 ( .A(p_input[7806]), .B(p_input[6806]), .Z(n1728) );
  AND U1944 ( .A(p_input[9806]), .B(p_input[8806]), .Z(n1726) );
  AND U1945 ( .A(n1729), .B(n1730), .Z(o[805]) );
  AND U1946 ( .A(n1731), .B(n1732), .Z(n1730) );
  AND U1947 ( .A(n1733), .B(p_input[3805]), .Z(n1732) );
  AND U1948 ( .A(p_input[2805]), .B(p_input[1805]), .Z(n1733) );
  AND U1949 ( .A(p_input[5805]), .B(p_input[4805]), .Z(n1731) );
  AND U1950 ( .A(n1734), .B(n1735), .Z(n1729) );
  AND U1951 ( .A(n1736), .B(p_input[805]), .Z(n1735) );
  AND U1952 ( .A(p_input[7805]), .B(p_input[6805]), .Z(n1736) );
  AND U1953 ( .A(p_input[9805]), .B(p_input[8805]), .Z(n1734) );
  AND U1954 ( .A(n1737), .B(n1738), .Z(o[804]) );
  AND U1955 ( .A(n1739), .B(n1740), .Z(n1738) );
  AND U1956 ( .A(n1741), .B(p_input[3804]), .Z(n1740) );
  AND U1957 ( .A(p_input[2804]), .B(p_input[1804]), .Z(n1741) );
  AND U1958 ( .A(p_input[5804]), .B(p_input[4804]), .Z(n1739) );
  AND U1959 ( .A(n1742), .B(n1743), .Z(n1737) );
  AND U1960 ( .A(n1744), .B(p_input[804]), .Z(n1743) );
  AND U1961 ( .A(p_input[7804]), .B(p_input[6804]), .Z(n1744) );
  AND U1962 ( .A(p_input[9804]), .B(p_input[8804]), .Z(n1742) );
  AND U1963 ( .A(n1745), .B(n1746), .Z(o[803]) );
  AND U1964 ( .A(n1747), .B(n1748), .Z(n1746) );
  AND U1965 ( .A(n1749), .B(p_input[3803]), .Z(n1748) );
  AND U1966 ( .A(p_input[2803]), .B(p_input[1803]), .Z(n1749) );
  AND U1967 ( .A(p_input[5803]), .B(p_input[4803]), .Z(n1747) );
  AND U1968 ( .A(n1750), .B(n1751), .Z(n1745) );
  AND U1969 ( .A(n1752), .B(p_input[803]), .Z(n1751) );
  AND U1970 ( .A(p_input[7803]), .B(p_input[6803]), .Z(n1752) );
  AND U1971 ( .A(p_input[9803]), .B(p_input[8803]), .Z(n1750) );
  AND U1972 ( .A(n1753), .B(n1754), .Z(o[802]) );
  AND U1973 ( .A(n1755), .B(n1756), .Z(n1754) );
  AND U1974 ( .A(n1757), .B(p_input[3802]), .Z(n1756) );
  AND U1975 ( .A(p_input[2802]), .B(p_input[1802]), .Z(n1757) );
  AND U1976 ( .A(p_input[5802]), .B(p_input[4802]), .Z(n1755) );
  AND U1977 ( .A(n1758), .B(n1759), .Z(n1753) );
  AND U1978 ( .A(n1760), .B(p_input[802]), .Z(n1759) );
  AND U1979 ( .A(p_input[7802]), .B(p_input[6802]), .Z(n1760) );
  AND U1980 ( .A(p_input[9802]), .B(p_input[8802]), .Z(n1758) );
  AND U1981 ( .A(n1761), .B(n1762), .Z(o[801]) );
  AND U1982 ( .A(n1763), .B(n1764), .Z(n1762) );
  AND U1983 ( .A(n1765), .B(p_input[3801]), .Z(n1764) );
  AND U1984 ( .A(p_input[2801]), .B(p_input[1801]), .Z(n1765) );
  AND U1985 ( .A(p_input[5801]), .B(p_input[4801]), .Z(n1763) );
  AND U1986 ( .A(n1766), .B(n1767), .Z(n1761) );
  AND U1987 ( .A(n1768), .B(p_input[801]), .Z(n1767) );
  AND U1988 ( .A(p_input[7801]), .B(p_input[6801]), .Z(n1768) );
  AND U1989 ( .A(p_input[9801]), .B(p_input[8801]), .Z(n1766) );
  AND U1990 ( .A(n1769), .B(n1770), .Z(o[800]) );
  AND U1991 ( .A(n1771), .B(n1772), .Z(n1770) );
  AND U1992 ( .A(n1773), .B(p_input[3800]), .Z(n1772) );
  AND U1993 ( .A(p_input[2800]), .B(p_input[1800]), .Z(n1773) );
  AND U1994 ( .A(p_input[5800]), .B(p_input[4800]), .Z(n1771) );
  AND U1995 ( .A(n1774), .B(n1775), .Z(n1769) );
  AND U1996 ( .A(n1776), .B(p_input[800]), .Z(n1775) );
  AND U1997 ( .A(p_input[7800]), .B(p_input[6800]), .Z(n1776) );
  AND U1998 ( .A(p_input[9800]), .B(p_input[8800]), .Z(n1774) );
  AND U1999 ( .A(n1777), .B(n1778), .Z(o[7]) );
  AND U2000 ( .A(n1779), .B(n1780), .Z(n1778) );
  AND U2001 ( .A(n1781), .B(p_input[3007]), .Z(n1780) );
  AND U2002 ( .A(p_input[2007]), .B(p_input[1007]), .Z(n1781) );
  AND U2003 ( .A(p_input[5007]), .B(p_input[4007]), .Z(n1779) );
  AND U2004 ( .A(n1782), .B(n1783), .Z(n1777) );
  AND U2005 ( .A(n1784), .B(p_input[7]), .Z(n1783) );
  AND U2006 ( .A(p_input[7007]), .B(p_input[6007]), .Z(n1784) );
  AND U2007 ( .A(p_input[9007]), .B(p_input[8007]), .Z(n1782) );
  AND U2008 ( .A(n1785), .B(n1786), .Z(o[79]) );
  AND U2009 ( .A(n1787), .B(n1788), .Z(n1786) );
  AND U2010 ( .A(n1789), .B(p_input[3079]), .Z(n1788) );
  AND U2011 ( .A(p_input[2079]), .B(p_input[1079]), .Z(n1789) );
  AND U2012 ( .A(p_input[5079]), .B(p_input[4079]), .Z(n1787) );
  AND U2013 ( .A(n1790), .B(n1791), .Z(n1785) );
  AND U2014 ( .A(n1792), .B(p_input[79]), .Z(n1791) );
  AND U2015 ( .A(p_input[7079]), .B(p_input[6079]), .Z(n1792) );
  AND U2016 ( .A(p_input[9079]), .B(p_input[8079]), .Z(n1790) );
  AND U2017 ( .A(n1793), .B(n1794), .Z(o[799]) );
  AND U2018 ( .A(n1795), .B(n1796), .Z(n1794) );
  AND U2019 ( .A(n1797), .B(p_input[3799]), .Z(n1796) );
  AND U2020 ( .A(p_input[2799]), .B(p_input[1799]), .Z(n1797) );
  AND U2021 ( .A(p_input[5799]), .B(p_input[4799]), .Z(n1795) );
  AND U2022 ( .A(n1798), .B(n1799), .Z(n1793) );
  AND U2023 ( .A(n1800), .B(p_input[799]), .Z(n1799) );
  AND U2024 ( .A(p_input[7799]), .B(p_input[6799]), .Z(n1800) );
  AND U2025 ( .A(p_input[9799]), .B(p_input[8799]), .Z(n1798) );
  AND U2026 ( .A(n1801), .B(n1802), .Z(o[798]) );
  AND U2027 ( .A(n1803), .B(n1804), .Z(n1802) );
  AND U2028 ( .A(n1805), .B(p_input[3798]), .Z(n1804) );
  AND U2029 ( .A(p_input[2798]), .B(p_input[1798]), .Z(n1805) );
  AND U2030 ( .A(p_input[5798]), .B(p_input[4798]), .Z(n1803) );
  AND U2031 ( .A(n1806), .B(n1807), .Z(n1801) );
  AND U2032 ( .A(n1808), .B(p_input[798]), .Z(n1807) );
  AND U2033 ( .A(p_input[7798]), .B(p_input[6798]), .Z(n1808) );
  AND U2034 ( .A(p_input[9798]), .B(p_input[8798]), .Z(n1806) );
  AND U2035 ( .A(n1809), .B(n1810), .Z(o[797]) );
  AND U2036 ( .A(n1811), .B(n1812), .Z(n1810) );
  AND U2037 ( .A(n1813), .B(p_input[3797]), .Z(n1812) );
  AND U2038 ( .A(p_input[2797]), .B(p_input[1797]), .Z(n1813) );
  AND U2039 ( .A(p_input[5797]), .B(p_input[4797]), .Z(n1811) );
  AND U2040 ( .A(n1814), .B(n1815), .Z(n1809) );
  AND U2041 ( .A(n1816), .B(p_input[797]), .Z(n1815) );
  AND U2042 ( .A(p_input[7797]), .B(p_input[6797]), .Z(n1816) );
  AND U2043 ( .A(p_input[9797]), .B(p_input[8797]), .Z(n1814) );
  AND U2044 ( .A(n1817), .B(n1818), .Z(o[796]) );
  AND U2045 ( .A(n1819), .B(n1820), .Z(n1818) );
  AND U2046 ( .A(n1821), .B(p_input[3796]), .Z(n1820) );
  AND U2047 ( .A(p_input[2796]), .B(p_input[1796]), .Z(n1821) );
  AND U2048 ( .A(p_input[5796]), .B(p_input[4796]), .Z(n1819) );
  AND U2049 ( .A(n1822), .B(n1823), .Z(n1817) );
  AND U2050 ( .A(n1824), .B(p_input[796]), .Z(n1823) );
  AND U2051 ( .A(p_input[7796]), .B(p_input[6796]), .Z(n1824) );
  AND U2052 ( .A(p_input[9796]), .B(p_input[8796]), .Z(n1822) );
  AND U2053 ( .A(n1825), .B(n1826), .Z(o[795]) );
  AND U2054 ( .A(n1827), .B(n1828), .Z(n1826) );
  AND U2055 ( .A(n1829), .B(p_input[3795]), .Z(n1828) );
  AND U2056 ( .A(p_input[2795]), .B(p_input[1795]), .Z(n1829) );
  AND U2057 ( .A(p_input[5795]), .B(p_input[4795]), .Z(n1827) );
  AND U2058 ( .A(n1830), .B(n1831), .Z(n1825) );
  AND U2059 ( .A(n1832), .B(p_input[795]), .Z(n1831) );
  AND U2060 ( .A(p_input[7795]), .B(p_input[6795]), .Z(n1832) );
  AND U2061 ( .A(p_input[9795]), .B(p_input[8795]), .Z(n1830) );
  AND U2062 ( .A(n1833), .B(n1834), .Z(o[794]) );
  AND U2063 ( .A(n1835), .B(n1836), .Z(n1834) );
  AND U2064 ( .A(n1837), .B(p_input[3794]), .Z(n1836) );
  AND U2065 ( .A(p_input[2794]), .B(p_input[1794]), .Z(n1837) );
  AND U2066 ( .A(p_input[5794]), .B(p_input[4794]), .Z(n1835) );
  AND U2067 ( .A(n1838), .B(n1839), .Z(n1833) );
  AND U2068 ( .A(n1840), .B(p_input[794]), .Z(n1839) );
  AND U2069 ( .A(p_input[7794]), .B(p_input[6794]), .Z(n1840) );
  AND U2070 ( .A(p_input[9794]), .B(p_input[8794]), .Z(n1838) );
  AND U2071 ( .A(n1841), .B(n1842), .Z(o[793]) );
  AND U2072 ( .A(n1843), .B(n1844), .Z(n1842) );
  AND U2073 ( .A(n1845), .B(p_input[3793]), .Z(n1844) );
  AND U2074 ( .A(p_input[2793]), .B(p_input[1793]), .Z(n1845) );
  AND U2075 ( .A(p_input[5793]), .B(p_input[4793]), .Z(n1843) );
  AND U2076 ( .A(n1846), .B(n1847), .Z(n1841) );
  AND U2077 ( .A(n1848), .B(p_input[793]), .Z(n1847) );
  AND U2078 ( .A(p_input[7793]), .B(p_input[6793]), .Z(n1848) );
  AND U2079 ( .A(p_input[9793]), .B(p_input[8793]), .Z(n1846) );
  AND U2080 ( .A(n1849), .B(n1850), .Z(o[792]) );
  AND U2081 ( .A(n1851), .B(n1852), .Z(n1850) );
  AND U2082 ( .A(n1853), .B(p_input[3792]), .Z(n1852) );
  AND U2083 ( .A(p_input[2792]), .B(p_input[1792]), .Z(n1853) );
  AND U2084 ( .A(p_input[5792]), .B(p_input[4792]), .Z(n1851) );
  AND U2085 ( .A(n1854), .B(n1855), .Z(n1849) );
  AND U2086 ( .A(n1856), .B(p_input[792]), .Z(n1855) );
  AND U2087 ( .A(p_input[7792]), .B(p_input[6792]), .Z(n1856) );
  AND U2088 ( .A(p_input[9792]), .B(p_input[8792]), .Z(n1854) );
  AND U2089 ( .A(n1857), .B(n1858), .Z(o[791]) );
  AND U2090 ( .A(n1859), .B(n1860), .Z(n1858) );
  AND U2091 ( .A(n1861), .B(p_input[3791]), .Z(n1860) );
  AND U2092 ( .A(p_input[2791]), .B(p_input[1791]), .Z(n1861) );
  AND U2093 ( .A(p_input[5791]), .B(p_input[4791]), .Z(n1859) );
  AND U2094 ( .A(n1862), .B(n1863), .Z(n1857) );
  AND U2095 ( .A(n1864), .B(p_input[791]), .Z(n1863) );
  AND U2096 ( .A(p_input[7791]), .B(p_input[6791]), .Z(n1864) );
  AND U2097 ( .A(p_input[9791]), .B(p_input[8791]), .Z(n1862) );
  AND U2098 ( .A(n1865), .B(n1866), .Z(o[790]) );
  AND U2099 ( .A(n1867), .B(n1868), .Z(n1866) );
  AND U2100 ( .A(n1869), .B(p_input[3790]), .Z(n1868) );
  AND U2101 ( .A(p_input[2790]), .B(p_input[1790]), .Z(n1869) );
  AND U2102 ( .A(p_input[5790]), .B(p_input[4790]), .Z(n1867) );
  AND U2103 ( .A(n1870), .B(n1871), .Z(n1865) );
  AND U2104 ( .A(n1872), .B(p_input[790]), .Z(n1871) );
  AND U2105 ( .A(p_input[7790]), .B(p_input[6790]), .Z(n1872) );
  AND U2106 ( .A(p_input[9790]), .B(p_input[8790]), .Z(n1870) );
  AND U2107 ( .A(n1873), .B(n1874), .Z(o[78]) );
  AND U2108 ( .A(n1875), .B(n1876), .Z(n1874) );
  AND U2109 ( .A(n1877), .B(p_input[3078]), .Z(n1876) );
  AND U2110 ( .A(p_input[2078]), .B(p_input[1078]), .Z(n1877) );
  AND U2111 ( .A(p_input[5078]), .B(p_input[4078]), .Z(n1875) );
  AND U2112 ( .A(n1878), .B(n1879), .Z(n1873) );
  AND U2113 ( .A(n1880), .B(p_input[78]), .Z(n1879) );
  AND U2114 ( .A(p_input[7078]), .B(p_input[6078]), .Z(n1880) );
  AND U2115 ( .A(p_input[9078]), .B(p_input[8078]), .Z(n1878) );
  AND U2116 ( .A(n1881), .B(n1882), .Z(o[789]) );
  AND U2117 ( .A(n1883), .B(n1884), .Z(n1882) );
  AND U2118 ( .A(n1885), .B(p_input[3789]), .Z(n1884) );
  AND U2119 ( .A(p_input[2789]), .B(p_input[1789]), .Z(n1885) );
  AND U2120 ( .A(p_input[5789]), .B(p_input[4789]), .Z(n1883) );
  AND U2121 ( .A(n1886), .B(n1887), .Z(n1881) );
  AND U2122 ( .A(n1888), .B(p_input[789]), .Z(n1887) );
  AND U2123 ( .A(p_input[7789]), .B(p_input[6789]), .Z(n1888) );
  AND U2124 ( .A(p_input[9789]), .B(p_input[8789]), .Z(n1886) );
  AND U2125 ( .A(n1889), .B(n1890), .Z(o[788]) );
  AND U2126 ( .A(n1891), .B(n1892), .Z(n1890) );
  AND U2127 ( .A(n1893), .B(p_input[3788]), .Z(n1892) );
  AND U2128 ( .A(p_input[2788]), .B(p_input[1788]), .Z(n1893) );
  AND U2129 ( .A(p_input[5788]), .B(p_input[4788]), .Z(n1891) );
  AND U2130 ( .A(n1894), .B(n1895), .Z(n1889) );
  AND U2131 ( .A(n1896), .B(p_input[788]), .Z(n1895) );
  AND U2132 ( .A(p_input[7788]), .B(p_input[6788]), .Z(n1896) );
  AND U2133 ( .A(p_input[9788]), .B(p_input[8788]), .Z(n1894) );
  AND U2134 ( .A(n1897), .B(n1898), .Z(o[787]) );
  AND U2135 ( .A(n1899), .B(n1900), .Z(n1898) );
  AND U2136 ( .A(n1901), .B(p_input[3787]), .Z(n1900) );
  AND U2137 ( .A(p_input[2787]), .B(p_input[1787]), .Z(n1901) );
  AND U2138 ( .A(p_input[5787]), .B(p_input[4787]), .Z(n1899) );
  AND U2139 ( .A(n1902), .B(n1903), .Z(n1897) );
  AND U2140 ( .A(n1904), .B(p_input[787]), .Z(n1903) );
  AND U2141 ( .A(p_input[7787]), .B(p_input[6787]), .Z(n1904) );
  AND U2142 ( .A(p_input[9787]), .B(p_input[8787]), .Z(n1902) );
  AND U2143 ( .A(n1905), .B(n1906), .Z(o[786]) );
  AND U2144 ( .A(n1907), .B(n1908), .Z(n1906) );
  AND U2145 ( .A(n1909), .B(p_input[3786]), .Z(n1908) );
  AND U2146 ( .A(p_input[2786]), .B(p_input[1786]), .Z(n1909) );
  AND U2147 ( .A(p_input[5786]), .B(p_input[4786]), .Z(n1907) );
  AND U2148 ( .A(n1910), .B(n1911), .Z(n1905) );
  AND U2149 ( .A(n1912), .B(p_input[786]), .Z(n1911) );
  AND U2150 ( .A(p_input[7786]), .B(p_input[6786]), .Z(n1912) );
  AND U2151 ( .A(p_input[9786]), .B(p_input[8786]), .Z(n1910) );
  AND U2152 ( .A(n1913), .B(n1914), .Z(o[785]) );
  AND U2153 ( .A(n1915), .B(n1916), .Z(n1914) );
  AND U2154 ( .A(n1917), .B(p_input[3785]), .Z(n1916) );
  AND U2155 ( .A(p_input[2785]), .B(p_input[1785]), .Z(n1917) );
  AND U2156 ( .A(p_input[5785]), .B(p_input[4785]), .Z(n1915) );
  AND U2157 ( .A(n1918), .B(n1919), .Z(n1913) );
  AND U2158 ( .A(n1920), .B(p_input[785]), .Z(n1919) );
  AND U2159 ( .A(p_input[7785]), .B(p_input[6785]), .Z(n1920) );
  AND U2160 ( .A(p_input[9785]), .B(p_input[8785]), .Z(n1918) );
  AND U2161 ( .A(n1921), .B(n1922), .Z(o[784]) );
  AND U2162 ( .A(n1923), .B(n1924), .Z(n1922) );
  AND U2163 ( .A(n1925), .B(p_input[3784]), .Z(n1924) );
  AND U2164 ( .A(p_input[2784]), .B(p_input[1784]), .Z(n1925) );
  AND U2165 ( .A(p_input[5784]), .B(p_input[4784]), .Z(n1923) );
  AND U2166 ( .A(n1926), .B(n1927), .Z(n1921) );
  AND U2167 ( .A(n1928), .B(p_input[784]), .Z(n1927) );
  AND U2168 ( .A(p_input[7784]), .B(p_input[6784]), .Z(n1928) );
  AND U2169 ( .A(p_input[9784]), .B(p_input[8784]), .Z(n1926) );
  AND U2170 ( .A(n1929), .B(n1930), .Z(o[783]) );
  AND U2171 ( .A(n1931), .B(n1932), .Z(n1930) );
  AND U2172 ( .A(n1933), .B(p_input[3783]), .Z(n1932) );
  AND U2173 ( .A(p_input[2783]), .B(p_input[1783]), .Z(n1933) );
  AND U2174 ( .A(p_input[5783]), .B(p_input[4783]), .Z(n1931) );
  AND U2175 ( .A(n1934), .B(n1935), .Z(n1929) );
  AND U2176 ( .A(n1936), .B(p_input[783]), .Z(n1935) );
  AND U2177 ( .A(p_input[7783]), .B(p_input[6783]), .Z(n1936) );
  AND U2178 ( .A(p_input[9783]), .B(p_input[8783]), .Z(n1934) );
  AND U2179 ( .A(n1937), .B(n1938), .Z(o[782]) );
  AND U2180 ( .A(n1939), .B(n1940), .Z(n1938) );
  AND U2181 ( .A(n1941), .B(p_input[3782]), .Z(n1940) );
  AND U2182 ( .A(p_input[2782]), .B(p_input[1782]), .Z(n1941) );
  AND U2183 ( .A(p_input[5782]), .B(p_input[4782]), .Z(n1939) );
  AND U2184 ( .A(n1942), .B(n1943), .Z(n1937) );
  AND U2185 ( .A(n1944), .B(p_input[782]), .Z(n1943) );
  AND U2186 ( .A(p_input[7782]), .B(p_input[6782]), .Z(n1944) );
  AND U2187 ( .A(p_input[9782]), .B(p_input[8782]), .Z(n1942) );
  AND U2188 ( .A(n1945), .B(n1946), .Z(o[781]) );
  AND U2189 ( .A(n1947), .B(n1948), .Z(n1946) );
  AND U2190 ( .A(n1949), .B(p_input[3781]), .Z(n1948) );
  AND U2191 ( .A(p_input[2781]), .B(p_input[1781]), .Z(n1949) );
  AND U2192 ( .A(p_input[5781]), .B(p_input[4781]), .Z(n1947) );
  AND U2193 ( .A(n1950), .B(n1951), .Z(n1945) );
  AND U2194 ( .A(n1952), .B(p_input[781]), .Z(n1951) );
  AND U2195 ( .A(p_input[7781]), .B(p_input[6781]), .Z(n1952) );
  AND U2196 ( .A(p_input[9781]), .B(p_input[8781]), .Z(n1950) );
  AND U2197 ( .A(n1953), .B(n1954), .Z(o[780]) );
  AND U2198 ( .A(n1955), .B(n1956), .Z(n1954) );
  AND U2199 ( .A(n1957), .B(p_input[3780]), .Z(n1956) );
  AND U2200 ( .A(p_input[2780]), .B(p_input[1780]), .Z(n1957) );
  AND U2201 ( .A(p_input[5780]), .B(p_input[4780]), .Z(n1955) );
  AND U2202 ( .A(n1958), .B(n1959), .Z(n1953) );
  AND U2203 ( .A(n1960), .B(p_input[780]), .Z(n1959) );
  AND U2204 ( .A(p_input[7780]), .B(p_input[6780]), .Z(n1960) );
  AND U2205 ( .A(p_input[9780]), .B(p_input[8780]), .Z(n1958) );
  AND U2206 ( .A(n1961), .B(n1962), .Z(o[77]) );
  AND U2207 ( .A(n1963), .B(n1964), .Z(n1962) );
  AND U2208 ( .A(n1965), .B(p_input[3077]), .Z(n1964) );
  AND U2209 ( .A(p_input[2077]), .B(p_input[1077]), .Z(n1965) );
  AND U2210 ( .A(p_input[5077]), .B(p_input[4077]), .Z(n1963) );
  AND U2211 ( .A(n1966), .B(n1967), .Z(n1961) );
  AND U2212 ( .A(n1968), .B(p_input[77]), .Z(n1967) );
  AND U2213 ( .A(p_input[7077]), .B(p_input[6077]), .Z(n1968) );
  AND U2214 ( .A(p_input[9077]), .B(p_input[8077]), .Z(n1966) );
  AND U2215 ( .A(n1969), .B(n1970), .Z(o[779]) );
  AND U2216 ( .A(n1971), .B(n1972), .Z(n1970) );
  AND U2217 ( .A(n1973), .B(p_input[3779]), .Z(n1972) );
  AND U2218 ( .A(p_input[2779]), .B(p_input[1779]), .Z(n1973) );
  AND U2219 ( .A(p_input[5779]), .B(p_input[4779]), .Z(n1971) );
  AND U2220 ( .A(n1974), .B(n1975), .Z(n1969) );
  AND U2221 ( .A(n1976), .B(p_input[779]), .Z(n1975) );
  AND U2222 ( .A(p_input[7779]), .B(p_input[6779]), .Z(n1976) );
  AND U2223 ( .A(p_input[9779]), .B(p_input[8779]), .Z(n1974) );
  AND U2224 ( .A(n1977), .B(n1978), .Z(o[778]) );
  AND U2225 ( .A(n1979), .B(n1980), .Z(n1978) );
  AND U2226 ( .A(n1981), .B(p_input[3778]), .Z(n1980) );
  AND U2227 ( .A(p_input[2778]), .B(p_input[1778]), .Z(n1981) );
  AND U2228 ( .A(p_input[5778]), .B(p_input[4778]), .Z(n1979) );
  AND U2229 ( .A(n1982), .B(n1983), .Z(n1977) );
  AND U2230 ( .A(n1984), .B(p_input[778]), .Z(n1983) );
  AND U2231 ( .A(p_input[7778]), .B(p_input[6778]), .Z(n1984) );
  AND U2232 ( .A(p_input[9778]), .B(p_input[8778]), .Z(n1982) );
  AND U2233 ( .A(n1985), .B(n1986), .Z(o[777]) );
  AND U2234 ( .A(n1987), .B(n1988), .Z(n1986) );
  AND U2235 ( .A(n1989), .B(p_input[3777]), .Z(n1988) );
  AND U2236 ( .A(p_input[2777]), .B(p_input[1777]), .Z(n1989) );
  AND U2237 ( .A(p_input[5777]), .B(p_input[4777]), .Z(n1987) );
  AND U2238 ( .A(n1990), .B(n1991), .Z(n1985) );
  AND U2239 ( .A(n1992), .B(p_input[777]), .Z(n1991) );
  AND U2240 ( .A(p_input[7777]), .B(p_input[6777]), .Z(n1992) );
  AND U2241 ( .A(p_input[9777]), .B(p_input[8777]), .Z(n1990) );
  AND U2242 ( .A(n1993), .B(n1994), .Z(o[776]) );
  AND U2243 ( .A(n1995), .B(n1996), .Z(n1994) );
  AND U2244 ( .A(n1997), .B(p_input[3776]), .Z(n1996) );
  AND U2245 ( .A(p_input[2776]), .B(p_input[1776]), .Z(n1997) );
  AND U2246 ( .A(p_input[5776]), .B(p_input[4776]), .Z(n1995) );
  AND U2247 ( .A(n1998), .B(n1999), .Z(n1993) );
  AND U2248 ( .A(n2000), .B(p_input[7776]), .Z(n1999) );
  AND U2249 ( .A(p_input[776]), .B(p_input[6776]), .Z(n2000) );
  AND U2250 ( .A(p_input[9776]), .B(p_input[8776]), .Z(n1998) );
  AND U2251 ( .A(n2001), .B(n2002), .Z(o[775]) );
  AND U2252 ( .A(n2003), .B(n2004), .Z(n2002) );
  AND U2253 ( .A(n2005), .B(p_input[3775]), .Z(n2004) );
  AND U2254 ( .A(p_input[2775]), .B(p_input[1775]), .Z(n2005) );
  AND U2255 ( .A(p_input[5775]), .B(p_input[4775]), .Z(n2003) );
  AND U2256 ( .A(n2006), .B(n2007), .Z(n2001) );
  AND U2257 ( .A(n2008), .B(p_input[7775]), .Z(n2007) );
  AND U2258 ( .A(p_input[775]), .B(p_input[6775]), .Z(n2008) );
  AND U2259 ( .A(p_input[9775]), .B(p_input[8775]), .Z(n2006) );
  AND U2260 ( .A(n2009), .B(n2010), .Z(o[774]) );
  AND U2261 ( .A(n2011), .B(n2012), .Z(n2010) );
  AND U2262 ( .A(n2013), .B(p_input[3774]), .Z(n2012) );
  AND U2263 ( .A(p_input[2774]), .B(p_input[1774]), .Z(n2013) );
  AND U2264 ( .A(p_input[5774]), .B(p_input[4774]), .Z(n2011) );
  AND U2265 ( .A(n2014), .B(n2015), .Z(n2009) );
  AND U2266 ( .A(n2016), .B(p_input[7774]), .Z(n2015) );
  AND U2267 ( .A(p_input[774]), .B(p_input[6774]), .Z(n2016) );
  AND U2268 ( .A(p_input[9774]), .B(p_input[8774]), .Z(n2014) );
  AND U2269 ( .A(n2017), .B(n2018), .Z(o[773]) );
  AND U2270 ( .A(n2019), .B(n2020), .Z(n2018) );
  AND U2271 ( .A(n2021), .B(p_input[3773]), .Z(n2020) );
  AND U2272 ( .A(p_input[2773]), .B(p_input[1773]), .Z(n2021) );
  AND U2273 ( .A(p_input[5773]), .B(p_input[4773]), .Z(n2019) );
  AND U2274 ( .A(n2022), .B(n2023), .Z(n2017) );
  AND U2275 ( .A(n2024), .B(p_input[7773]), .Z(n2023) );
  AND U2276 ( .A(p_input[773]), .B(p_input[6773]), .Z(n2024) );
  AND U2277 ( .A(p_input[9773]), .B(p_input[8773]), .Z(n2022) );
  AND U2278 ( .A(n2025), .B(n2026), .Z(o[772]) );
  AND U2279 ( .A(n2027), .B(n2028), .Z(n2026) );
  AND U2280 ( .A(n2029), .B(p_input[3772]), .Z(n2028) );
  AND U2281 ( .A(p_input[2772]), .B(p_input[1772]), .Z(n2029) );
  AND U2282 ( .A(p_input[5772]), .B(p_input[4772]), .Z(n2027) );
  AND U2283 ( .A(n2030), .B(n2031), .Z(n2025) );
  AND U2284 ( .A(n2032), .B(p_input[7772]), .Z(n2031) );
  AND U2285 ( .A(p_input[772]), .B(p_input[6772]), .Z(n2032) );
  AND U2286 ( .A(p_input[9772]), .B(p_input[8772]), .Z(n2030) );
  AND U2287 ( .A(n2033), .B(n2034), .Z(o[771]) );
  AND U2288 ( .A(n2035), .B(n2036), .Z(n2034) );
  AND U2289 ( .A(n2037), .B(p_input[3771]), .Z(n2036) );
  AND U2290 ( .A(p_input[2771]), .B(p_input[1771]), .Z(n2037) );
  AND U2291 ( .A(p_input[5771]), .B(p_input[4771]), .Z(n2035) );
  AND U2292 ( .A(n2038), .B(n2039), .Z(n2033) );
  AND U2293 ( .A(n2040), .B(p_input[7771]), .Z(n2039) );
  AND U2294 ( .A(p_input[771]), .B(p_input[6771]), .Z(n2040) );
  AND U2295 ( .A(p_input[9771]), .B(p_input[8771]), .Z(n2038) );
  AND U2296 ( .A(n2041), .B(n2042), .Z(o[770]) );
  AND U2297 ( .A(n2043), .B(n2044), .Z(n2042) );
  AND U2298 ( .A(n2045), .B(p_input[3770]), .Z(n2044) );
  AND U2299 ( .A(p_input[2770]), .B(p_input[1770]), .Z(n2045) );
  AND U2300 ( .A(p_input[5770]), .B(p_input[4770]), .Z(n2043) );
  AND U2301 ( .A(n2046), .B(n2047), .Z(n2041) );
  AND U2302 ( .A(n2048), .B(p_input[7770]), .Z(n2047) );
  AND U2303 ( .A(p_input[770]), .B(p_input[6770]), .Z(n2048) );
  AND U2304 ( .A(p_input[9770]), .B(p_input[8770]), .Z(n2046) );
  AND U2305 ( .A(n2049), .B(n2050), .Z(o[76]) );
  AND U2306 ( .A(n2051), .B(n2052), .Z(n2050) );
  AND U2307 ( .A(n2053), .B(p_input[3076]), .Z(n2052) );
  AND U2308 ( .A(p_input[2076]), .B(p_input[1076]), .Z(n2053) );
  AND U2309 ( .A(p_input[5076]), .B(p_input[4076]), .Z(n2051) );
  AND U2310 ( .A(n2054), .B(n2055), .Z(n2049) );
  AND U2311 ( .A(n2056), .B(p_input[76]), .Z(n2055) );
  AND U2312 ( .A(p_input[7076]), .B(p_input[6076]), .Z(n2056) );
  AND U2313 ( .A(p_input[9076]), .B(p_input[8076]), .Z(n2054) );
  AND U2314 ( .A(n2057), .B(n2058), .Z(o[769]) );
  AND U2315 ( .A(n2059), .B(n2060), .Z(n2058) );
  AND U2316 ( .A(n2061), .B(p_input[3769]), .Z(n2060) );
  AND U2317 ( .A(p_input[2769]), .B(p_input[1769]), .Z(n2061) );
  AND U2318 ( .A(p_input[5769]), .B(p_input[4769]), .Z(n2059) );
  AND U2319 ( .A(n2062), .B(n2063), .Z(n2057) );
  AND U2320 ( .A(n2064), .B(p_input[7769]), .Z(n2063) );
  AND U2321 ( .A(p_input[769]), .B(p_input[6769]), .Z(n2064) );
  AND U2322 ( .A(p_input[9769]), .B(p_input[8769]), .Z(n2062) );
  AND U2323 ( .A(n2065), .B(n2066), .Z(o[768]) );
  AND U2324 ( .A(n2067), .B(n2068), .Z(n2066) );
  AND U2325 ( .A(n2069), .B(p_input[3768]), .Z(n2068) );
  AND U2326 ( .A(p_input[2768]), .B(p_input[1768]), .Z(n2069) );
  AND U2327 ( .A(p_input[5768]), .B(p_input[4768]), .Z(n2067) );
  AND U2328 ( .A(n2070), .B(n2071), .Z(n2065) );
  AND U2329 ( .A(n2072), .B(p_input[7768]), .Z(n2071) );
  AND U2330 ( .A(p_input[768]), .B(p_input[6768]), .Z(n2072) );
  AND U2331 ( .A(p_input[9768]), .B(p_input[8768]), .Z(n2070) );
  AND U2332 ( .A(n2073), .B(n2074), .Z(o[767]) );
  AND U2333 ( .A(n2075), .B(n2076), .Z(n2074) );
  AND U2334 ( .A(n2077), .B(p_input[3767]), .Z(n2076) );
  AND U2335 ( .A(p_input[2767]), .B(p_input[1767]), .Z(n2077) );
  AND U2336 ( .A(p_input[5767]), .B(p_input[4767]), .Z(n2075) );
  AND U2337 ( .A(n2078), .B(n2079), .Z(n2073) );
  AND U2338 ( .A(n2080), .B(p_input[7767]), .Z(n2079) );
  AND U2339 ( .A(p_input[767]), .B(p_input[6767]), .Z(n2080) );
  AND U2340 ( .A(p_input[9767]), .B(p_input[8767]), .Z(n2078) );
  AND U2341 ( .A(n2081), .B(n2082), .Z(o[766]) );
  AND U2342 ( .A(n2083), .B(n2084), .Z(n2082) );
  AND U2343 ( .A(n2085), .B(p_input[3766]), .Z(n2084) );
  AND U2344 ( .A(p_input[2766]), .B(p_input[1766]), .Z(n2085) );
  AND U2345 ( .A(p_input[5766]), .B(p_input[4766]), .Z(n2083) );
  AND U2346 ( .A(n2086), .B(n2087), .Z(n2081) );
  AND U2347 ( .A(n2088), .B(p_input[7766]), .Z(n2087) );
  AND U2348 ( .A(p_input[766]), .B(p_input[6766]), .Z(n2088) );
  AND U2349 ( .A(p_input[9766]), .B(p_input[8766]), .Z(n2086) );
  AND U2350 ( .A(n2089), .B(n2090), .Z(o[765]) );
  AND U2351 ( .A(n2091), .B(n2092), .Z(n2090) );
  AND U2352 ( .A(n2093), .B(p_input[3765]), .Z(n2092) );
  AND U2353 ( .A(p_input[2765]), .B(p_input[1765]), .Z(n2093) );
  AND U2354 ( .A(p_input[5765]), .B(p_input[4765]), .Z(n2091) );
  AND U2355 ( .A(n2094), .B(n2095), .Z(n2089) );
  AND U2356 ( .A(n2096), .B(p_input[7765]), .Z(n2095) );
  AND U2357 ( .A(p_input[765]), .B(p_input[6765]), .Z(n2096) );
  AND U2358 ( .A(p_input[9765]), .B(p_input[8765]), .Z(n2094) );
  AND U2359 ( .A(n2097), .B(n2098), .Z(o[764]) );
  AND U2360 ( .A(n2099), .B(n2100), .Z(n2098) );
  AND U2361 ( .A(n2101), .B(p_input[3764]), .Z(n2100) );
  AND U2362 ( .A(p_input[2764]), .B(p_input[1764]), .Z(n2101) );
  AND U2363 ( .A(p_input[5764]), .B(p_input[4764]), .Z(n2099) );
  AND U2364 ( .A(n2102), .B(n2103), .Z(n2097) );
  AND U2365 ( .A(n2104), .B(p_input[7764]), .Z(n2103) );
  AND U2366 ( .A(p_input[764]), .B(p_input[6764]), .Z(n2104) );
  AND U2367 ( .A(p_input[9764]), .B(p_input[8764]), .Z(n2102) );
  AND U2368 ( .A(n2105), .B(n2106), .Z(o[763]) );
  AND U2369 ( .A(n2107), .B(n2108), .Z(n2106) );
  AND U2370 ( .A(n2109), .B(p_input[3763]), .Z(n2108) );
  AND U2371 ( .A(p_input[2763]), .B(p_input[1763]), .Z(n2109) );
  AND U2372 ( .A(p_input[5763]), .B(p_input[4763]), .Z(n2107) );
  AND U2373 ( .A(n2110), .B(n2111), .Z(n2105) );
  AND U2374 ( .A(n2112), .B(p_input[7763]), .Z(n2111) );
  AND U2375 ( .A(p_input[763]), .B(p_input[6763]), .Z(n2112) );
  AND U2376 ( .A(p_input[9763]), .B(p_input[8763]), .Z(n2110) );
  AND U2377 ( .A(n2113), .B(n2114), .Z(o[762]) );
  AND U2378 ( .A(n2115), .B(n2116), .Z(n2114) );
  AND U2379 ( .A(n2117), .B(p_input[3762]), .Z(n2116) );
  AND U2380 ( .A(p_input[2762]), .B(p_input[1762]), .Z(n2117) );
  AND U2381 ( .A(p_input[5762]), .B(p_input[4762]), .Z(n2115) );
  AND U2382 ( .A(n2118), .B(n2119), .Z(n2113) );
  AND U2383 ( .A(n2120), .B(p_input[7762]), .Z(n2119) );
  AND U2384 ( .A(p_input[762]), .B(p_input[6762]), .Z(n2120) );
  AND U2385 ( .A(p_input[9762]), .B(p_input[8762]), .Z(n2118) );
  AND U2386 ( .A(n2121), .B(n2122), .Z(o[761]) );
  AND U2387 ( .A(n2123), .B(n2124), .Z(n2122) );
  AND U2388 ( .A(n2125), .B(p_input[3761]), .Z(n2124) );
  AND U2389 ( .A(p_input[2761]), .B(p_input[1761]), .Z(n2125) );
  AND U2390 ( .A(p_input[5761]), .B(p_input[4761]), .Z(n2123) );
  AND U2391 ( .A(n2126), .B(n2127), .Z(n2121) );
  AND U2392 ( .A(n2128), .B(p_input[7761]), .Z(n2127) );
  AND U2393 ( .A(p_input[761]), .B(p_input[6761]), .Z(n2128) );
  AND U2394 ( .A(p_input[9761]), .B(p_input[8761]), .Z(n2126) );
  AND U2395 ( .A(n2129), .B(n2130), .Z(o[760]) );
  AND U2396 ( .A(n2131), .B(n2132), .Z(n2130) );
  AND U2397 ( .A(n2133), .B(p_input[3760]), .Z(n2132) );
  AND U2398 ( .A(p_input[2760]), .B(p_input[1760]), .Z(n2133) );
  AND U2399 ( .A(p_input[5760]), .B(p_input[4760]), .Z(n2131) );
  AND U2400 ( .A(n2134), .B(n2135), .Z(n2129) );
  AND U2401 ( .A(n2136), .B(p_input[7760]), .Z(n2135) );
  AND U2402 ( .A(p_input[760]), .B(p_input[6760]), .Z(n2136) );
  AND U2403 ( .A(p_input[9760]), .B(p_input[8760]), .Z(n2134) );
  AND U2404 ( .A(n2137), .B(n2138), .Z(o[75]) );
  AND U2405 ( .A(n2139), .B(n2140), .Z(n2138) );
  AND U2406 ( .A(n2141), .B(p_input[3075]), .Z(n2140) );
  AND U2407 ( .A(p_input[2075]), .B(p_input[1075]), .Z(n2141) );
  AND U2408 ( .A(p_input[5075]), .B(p_input[4075]), .Z(n2139) );
  AND U2409 ( .A(n2142), .B(n2143), .Z(n2137) );
  AND U2410 ( .A(n2144), .B(p_input[75]), .Z(n2143) );
  AND U2411 ( .A(p_input[7075]), .B(p_input[6075]), .Z(n2144) );
  AND U2412 ( .A(p_input[9075]), .B(p_input[8075]), .Z(n2142) );
  AND U2413 ( .A(n2145), .B(n2146), .Z(o[759]) );
  AND U2414 ( .A(n2147), .B(n2148), .Z(n2146) );
  AND U2415 ( .A(n2149), .B(p_input[3759]), .Z(n2148) );
  AND U2416 ( .A(p_input[2759]), .B(p_input[1759]), .Z(n2149) );
  AND U2417 ( .A(p_input[5759]), .B(p_input[4759]), .Z(n2147) );
  AND U2418 ( .A(n2150), .B(n2151), .Z(n2145) );
  AND U2419 ( .A(n2152), .B(p_input[7759]), .Z(n2151) );
  AND U2420 ( .A(p_input[759]), .B(p_input[6759]), .Z(n2152) );
  AND U2421 ( .A(p_input[9759]), .B(p_input[8759]), .Z(n2150) );
  AND U2422 ( .A(n2153), .B(n2154), .Z(o[758]) );
  AND U2423 ( .A(n2155), .B(n2156), .Z(n2154) );
  AND U2424 ( .A(n2157), .B(p_input[3758]), .Z(n2156) );
  AND U2425 ( .A(p_input[2758]), .B(p_input[1758]), .Z(n2157) );
  AND U2426 ( .A(p_input[5758]), .B(p_input[4758]), .Z(n2155) );
  AND U2427 ( .A(n2158), .B(n2159), .Z(n2153) );
  AND U2428 ( .A(n2160), .B(p_input[7758]), .Z(n2159) );
  AND U2429 ( .A(p_input[758]), .B(p_input[6758]), .Z(n2160) );
  AND U2430 ( .A(p_input[9758]), .B(p_input[8758]), .Z(n2158) );
  AND U2431 ( .A(n2161), .B(n2162), .Z(o[757]) );
  AND U2432 ( .A(n2163), .B(n2164), .Z(n2162) );
  AND U2433 ( .A(n2165), .B(p_input[3757]), .Z(n2164) );
  AND U2434 ( .A(p_input[2757]), .B(p_input[1757]), .Z(n2165) );
  AND U2435 ( .A(p_input[5757]), .B(p_input[4757]), .Z(n2163) );
  AND U2436 ( .A(n2166), .B(n2167), .Z(n2161) );
  AND U2437 ( .A(n2168), .B(p_input[7757]), .Z(n2167) );
  AND U2438 ( .A(p_input[757]), .B(p_input[6757]), .Z(n2168) );
  AND U2439 ( .A(p_input[9757]), .B(p_input[8757]), .Z(n2166) );
  AND U2440 ( .A(n2169), .B(n2170), .Z(o[756]) );
  AND U2441 ( .A(n2171), .B(n2172), .Z(n2170) );
  AND U2442 ( .A(n2173), .B(p_input[3756]), .Z(n2172) );
  AND U2443 ( .A(p_input[2756]), .B(p_input[1756]), .Z(n2173) );
  AND U2444 ( .A(p_input[5756]), .B(p_input[4756]), .Z(n2171) );
  AND U2445 ( .A(n2174), .B(n2175), .Z(n2169) );
  AND U2446 ( .A(n2176), .B(p_input[7756]), .Z(n2175) );
  AND U2447 ( .A(p_input[756]), .B(p_input[6756]), .Z(n2176) );
  AND U2448 ( .A(p_input[9756]), .B(p_input[8756]), .Z(n2174) );
  AND U2449 ( .A(n2177), .B(n2178), .Z(o[755]) );
  AND U2450 ( .A(n2179), .B(n2180), .Z(n2178) );
  AND U2451 ( .A(n2181), .B(p_input[3755]), .Z(n2180) );
  AND U2452 ( .A(p_input[2755]), .B(p_input[1755]), .Z(n2181) );
  AND U2453 ( .A(p_input[5755]), .B(p_input[4755]), .Z(n2179) );
  AND U2454 ( .A(n2182), .B(n2183), .Z(n2177) );
  AND U2455 ( .A(n2184), .B(p_input[7755]), .Z(n2183) );
  AND U2456 ( .A(p_input[755]), .B(p_input[6755]), .Z(n2184) );
  AND U2457 ( .A(p_input[9755]), .B(p_input[8755]), .Z(n2182) );
  AND U2458 ( .A(n2185), .B(n2186), .Z(o[754]) );
  AND U2459 ( .A(n2187), .B(n2188), .Z(n2186) );
  AND U2460 ( .A(n2189), .B(p_input[3754]), .Z(n2188) );
  AND U2461 ( .A(p_input[2754]), .B(p_input[1754]), .Z(n2189) );
  AND U2462 ( .A(p_input[5754]), .B(p_input[4754]), .Z(n2187) );
  AND U2463 ( .A(n2190), .B(n2191), .Z(n2185) );
  AND U2464 ( .A(n2192), .B(p_input[7754]), .Z(n2191) );
  AND U2465 ( .A(p_input[754]), .B(p_input[6754]), .Z(n2192) );
  AND U2466 ( .A(p_input[9754]), .B(p_input[8754]), .Z(n2190) );
  AND U2467 ( .A(n2193), .B(n2194), .Z(o[753]) );
  AND U2468 ( .A(n2195), .B(n2196), .Z(n2194) );
  AND U2469 ( .A(n2197), .B(p_input[3753]), .Z(n2196) );
  AND U2470 ( .A(p_input[2753]), .B(p_input[1753]), .Z(n2197) );
  AND U2471 ( .A(p_input[5753]), .B(p_input[4753]), .Z(n2195) );
  AND U2472 ( .A(n2198), .B(n2199), .Z(n2193) );
  AND U2473 ( .A(n2200), .B(p_input[7753]), .Z(n2199) );
  AND U2474 ( .A(p_input[753]), .B(p_input[6753]), .Z(n2200) );
  AND U2475 ( .A(p_input[9753]), .B(p_input[8753]), .Z(n2198) );
  AND U2476 ( .A(n2201), .B(n2202), .Z(o[752]) );
  AND U2477 ( .A(n2203), .B(n2204), .Z(n2202) );
  AND U2478 ( .A(n2205), .B(p_input[3752]), .Z(n2204) );
  AND U2479 ( .A(p_input[2752]), .B(p_input[1752]), .Z(n2205) );
  AND U2480 ( .A(p_input[5752]), .B(p_input[4752]), .Z(n2203) );
  AND U2481 ( .A(n2206), .B(n2207), .Z(n2201) );
  AND U2482 ( .A(n2208), .B(p_input[7752]), .Z(n2207) );
  AND U2483 ( .A(p_input[752]), .B(p_input[6752]), .Z(n2208) );
  AND U2484 ( .A(p_input[9752]), .B(p_input[8752]), .Z(n2206) );
  AND U2485 ( .A(n2209), .B(n2210), .Z(o[751]) );
  AND U2486 ( .A(n2211), .B(n2212), .Z(n2210) );
  AND U2487 ( .A(n2213), .B(p_input[3751]), .Z(n2212) );
  AND U2488 ( .A(p_input[2751]), .B(p_input[1751]), .Z(n2213) );
  AND U2489 ( .A(p_input[5751]), .B(p_input[4751]), .Z(n2211) );
  AND U2490 ( .A(n2214), .B(n2215), .Z(n2209) );
  AND U2491 ( .A(n2216), .B(p_input[7751]), .Z(n2215) );
  AND U2492 ( .A(p_input[751]), .B(p_input[6751]), .Z(n2216) );
  AND U2493 ( .A(p_input[9751]), .B(p_input[8751]), .Z(n2214) );
  AND U2494 ( .A(n2217), .B(n2218), .Z(o[750]) );
  AND U2495 ( .A(n2219), .B(n2220), .Z(n2218) );
  AND U2496 ( .A(n2221), .B(p_input[3750]), .Z(n2220) );
  AND U2497 ( .A(p_input[2750]), .B(p_input[1750]), .Z(n2221) );
  AND U2498 ( .A(p_input[5750]), .B(p_input[4750]), .Z(n2219) );
  AND U2499 ( .A(n2222), .B(n2223), .Z(n2217) );
  AND U2500 ( .A(n2224), .B(p_input[7750]), .Z(n2223) );
  AND U2501 ( .A(p_input[750]), .B(p_input[6750]), .Z(n2224) );
  AND U2502 ( .A(p_input[9750]), .B(p_input[8750]), .Z(n2222) );
  AND U2503 ( .A(n2225), .B(n2226), .Z(o[74]) );
  AND U2504 ( .A(n2227), .B(n2228), .Z(n2226) );
  AND U2505 ( .A(n2229), .B(p_input[3074]), .Z(n2228) );
  AND U2506 ( .A(p_input[2074]), .B(p_input[1074]), .Z(n2229) );
  AND U2507 ( .A(p_input[5074]), .B(p_input[4074]), .Z(n2227) );
  AND U2508 ( .A(n2230), .B(n2231), .Z(n2225) );
  AND U2509 ( .A(n2232), .B(p_input[74]), .Z(n2231) );
  AND U2510 ( .A(p_input[7074]), .B(p_input[6074]), .Z(n2232) );
  AND U2511 ( .A(p_input[9074]), .B(p_input[8074]), .Z(n2230) );
  AND U2512 ( .A(n2233), .B(n2234), .Z(o[749]) );
  AND U2513 ( .A(n2235), .B(n2236), .Z(n2234) );
  AND U2514 ( .A(n2237), .B(p_input[3749]), .Z(n2236) );
  AND U2515 ( .A(p_input[2749]), .B(p_input[1749]), .Z(n2237) );
  AND U2516 ( .A(p_input[5749]), .B(p_input[4749]), .Z(n2235) );
  AND U2517 ( .A(n2238), .B(n2239), .Z(n2233) );
  AND U2518 ( .A(n2240), .B(p_input[7749]), .Z(n2239) );
  AND U2519 ( .A(p_input[749]), .B(p_input[6749]), .Z(n2240) );
  AND U2520 ( .A(p_input[9749]), .B(p_input[8749]), .Z(n2238) );
  AND U2521 ( .A(n2241), .B(n2242), .Z(o[748]) );
  AND U2522 ( .A(n2243), .B(n2244), .Z(n2242) );
  AND U2523 ( .A(n2245), .B(p_input[3748]), .Z(n2244) );
  AND U2524 ( .A(p_input[2748]), .B(p_input[1748]), .Z(n2245) );
  AND U2525 ( .A(p_input[5748]), .B(p_input[4748]), .Z(n2243) );
  AND U2526 ( .A(n2246), .B(n2247), .Z(n2241) );
  AND U2527 ( .A(n2248), .B(p_input[7748]), .Z(n2247) );
  AND U2528 ( .A(p_input[748]), .B(p_input[6748]), .Z(n2248) );
  AND U2529 ( .A(p_input[9748]), .B(p_input[8748]), .Z(n2246) );
  AND U2530 ( .A(n2249), .B(n2250), .Z(o[747]) );
  AND U2531 ( .A(n2251), .B(n2252), .Z(n2250) );
  AND U2532 ( .A(n2253), .B(p_input[3747]), .Z(n2252) );
  AND U2533 ( .A(p_input[2747]), .B(p_input[1747]), .Z(n2253) );
  AND U2534 ( .A(p_input[5747]), .B(p_input[4747]), .Z(n2251) );
  AND U2535 ( .A(n2254), .B(n2255), .Z(n2249) );
  AND U2536 ( .A(n2256), .B(p_input[7747]), .Z(n2255) );
  AND U2537 ( .A(p_input[747]), .B(p_input[6747]), .Z(n2256) );
  AND U2538 ( .A(p_input[9747]), .B(p_input[8747]), .Z(n2254) );
  AND U2539 ( .A(n2257), .B(n2258), .Z(o[746]) );
  AND U2540 ( .A(n2259), .B(n2260), .Z(n2258) );
  AND U2541 ( .A(n2261), .B(p_input[3746]), .Z(n2260) );
  AND U2542 ( .A(p_input[2746]), .B(p_input[1746]), .Z(n2261) );
  AND U2543 ( .A(p_input[5746]), .B(p_input[4746]), .Z(n2259) );
  AND U2544 ( .A(n2262), .B(n2263), .Z(n2257) );
  AND U2545 ( .A(n2264), .B(p_input[7746]), .Z(n2263) );
  AND U2546 ( .A(p_input[746]), .B(p_input[6746]), .Z(n2264) );
  AND U2547 ( .A(p_input[9746]), .B(p_input[8746]), .Z(n2262) );
  AND U2548 ( .A(n2265), .B(n2266), .Z(o[745]) );
  AND U2549 ( .A(n2267), .B(n2268), .Z(n2266) );
  AND U2550 ( .A(n2269), .B(p_input[3745]), .Z(n2268) );
  AND U2551 ( .A(p_input[2745]), .B(p_input[1745]), .Z(n2269) );
  AND U2552 ( .A(p_input[5745]), .B(p_input[4745]), .Z(n2267) );
  AND U2553 ( .A(n2270), .B(n2271), .Z(n2265) );
  AND U2554 ( .A(n2272), .B(p_input[7745]), .Z(n2271) );
  AND U2555 ( .A(p_input[745]), .B(p_input[6745]), .Z(n2272) );
  AND U2556 ( .A(p_input[9745]), .B(p_input[8745]), .Z(n2270) );
  AND U2557 ( .A(n2273), .B(n2274), .Z(o[744]) );
  AND U2558 ( .A(n2275), .B(n2276), .Z(n2274) );
  AND U2559 ( .A(n2277), .B(p_input[3744]), .Z(n2276) );
  AND U2560 ( .A(p_input[2744]), .B(p_input[1744]), .Z(n2277) );
  AND U2561 ( .A(p_input[5744]), .B(p_input[4744]), .Z(n2275) );
  AND U2562 ( .A(n2278), .B(n2279), .Z(n2273) );
  AND U2563 ( .A(n2280), .B(p_input[7744]), .Z(n2279) );
  AND U2564 ( .A(p_input[744]), .B(p_input[6744]), .Z(n2280) );
  AND U2565 ( .A(p_input[9744]), .B(p_input[8744]), .Z(n2278) );
  AND U2566 ( .A(n2281), .B(n2282), .Z(o[743]) );
  AND U2567 ( .A(n2283), .B(n2284), .Z(n2282) );
  AND U2568 ( .A(n2285), .B(p_input[3743]), .Z(n2284) );
  AND U2569 ( .A(p_input[2743]), .B(p_input[1743]), .Z(n2285) );
  AND U2570 ( .A(p_input[5743]), .B(p_input[4743]), .Z(n2283) );
  AND U2571 ( .A(n2286), .B(n2287), .Z(n2281) );
  AND U2572 ( .A(n2288), .B(p_input[7743]), .Z(n2287) );
  AND U2573 ( .A(p_input[743]), .B(p_input[6743]), .Z(n2288) );
  AND U2574 ( .A(p_input[9743]), .B(p_input[8743]), .Z(n2286) );
  AND U2575 ( .A(n2289), .B(n2290), .Z(o[742]) );
  AND U2576 ( .A(n2291), .B(n2292), .Z(n2290) );
  AND U2577 ( .A(n2293), .B(p_input[3742]), .Z(n2292) );
  AND U2578 ( .A(p_input[2742]), .B(p_input[1742]), .Z(n2293) );
  AND U2579 ( .A(p_input[5742]), .B(p_input[4742]), .Z(n2291) );
  AND U2580 ( .A(n2294), .B(n2295), .Z(n2289) );
  AND U2581 ( .A(n2296), .B(p_input[7742]), .Z(n2295) );
  AND U2582 ( .A(p_input[742]), .B(p_input[6742]), .Z(n2296) );
  AND U2583 ( .A(p_input[9742]), .B(p_input[8742]), .Z(n2294) );
  AND U2584 ( .A(n2297), .B(n2298), .Z(o[741]) );
  AND U2585 ( .A(n2299), .B(n2300), .Z(n2298) );
  AND U2586 ( .A(n2301), .B(p_input[3741]), .Z(n2300) );
  AND U2587 ( .A(p_input[2741]), .B(p_input[1741]), .Z(n2301) );
  AND U2588 ( .A(p_input[5741]), .B(p_input[4741]), .Z(n2299) );
  AND U2589 ( .A(n2302), .B(n2303), .Z(n2297) );
  AND U2590 ( .A(n2304), .B(p_input[7741]), .Z(n2303) );
  AND U2591 ( .A(p_input[741]), .B(p_input[6741]), .Z(n2304) );
  AND U2592 ( .A(p_input[9741]), .B(p_input[8741]), .Z(n2302) );
  AND U2593 ( .A(n2305), .B(n2306), .Z(o[740]) );
  AND U2594 ( .A(n2307), .B(n2308), .Z(n2306) );
  AND U2595 ( .A(n2309), .B(p_input[3740]), .Z(n2308) );
  AND U2596 ( .A(p_input[2740]), .B(p_input[1740]), .Z(n2309) );
  AND U2597 ( .A(p_input[5740]), .B(p_input[4740]), .Z(n2307) );
  AND U2598 ( .A(n2310), .B(n2311), .Z(n2305) );
  AND U2599 ( .A(n2312), .B(p_input[7740]), .Z(n2311) );
  AND U2600 ( .A(p_input[740]), .B(p_input[6740]), .Z(n2312) );
  AND U2601 ( .A(p_input[9740]), .B(p_input[8740]), .Z(n2310) );
  AND U2602 ( .A(n2313), .B(n2314), .Z(o[73]) );
  AND U2603 ( .A(n2315), .B(n2316), .Z(n2314) );
  AND U2604 ( .A(n2317), .B(p_input[3073]), .Z(n2316) );
  AND U2605 ( .A(p_input[2073]), .B(p_input[1073]), .Z(n2317) );
  AND U2606 ( .A(p_input[5073]), .B(p_input[4073]), .Z(n2315) );
  AND U2607 ( .A(n2318), .B(n2319), .Z(n2313) );
  AND U2608 ( .A(n2320), .B(p_input[73]), .Z(n2319) );
  AND U2609 ( .A(p_input[7073]), .B(p_input[6073]), .Z(n2320) );
  AND U2610 ( .A(p_input[9073]), .B(p_input[8073]), .Z(n2318) );
  AND U2611 ( .A(n2321), .B(n2322), .Z(o[739]) );
  AND U2612 ( .A(n2323), .B(n2324), .Z(n2322) );
  AND U2613 ( .A(n2325), .B(p_input[3739]), .Z(n2324) );
  AND U2614 ( .A(p_input[2739]), .B(p_input[1739]), .Z(n2325) );
  AND U2615 ( .A(p_input[5739]), .B(p_input[4739]), .Z(n2323) );
  AND U2616 ( .A(n2326), .B(n2327), .Z(n2321) );
  AND U2617 ( .A(n2328), .B(p_input[7739]), .Z(n2327) );
  AND U2618 ( .A(p_input[739]), .B(p_input[6739]), .Z(n2328) );
  AND U2619 ( .A(p_input[9739]), .B(p_input[8739]), .Z(n2326) );
  AND U2620 ( .A(n2329), .B(n2330), .Z(o[738]) );
  AND U2621 ( .A(n2331), .B(n2332), .Z(n2330) );
  AND U2622 ( .A(n2333), .B(p_input[3738]), .Z(n2332) );
  AND U2623 ( .A(p_input[2738]), .B(p_input[1738]), .Z(n2333) );
  AND U2624 ( .A(p_input[5738]), .B(p_input[4738]), .Z(n2331) );
  AND U2625 ( .A(n2334), .B(n2335), .Z(n2329) );
  AND U2626 ( .A(n2336), .B(p_input[7738]), .Z(n2335) );
  AND U2627 ( .A(p_input[738]), .B(p_input[6738]), .Z(n2336) );
  AND U2628 ( .A(p_input[9738]), .B(p_input[8738]), .Z(n2334) );
  AND U2629 ( .A(n2337), .B(n2338), .Z(o[737]) );
  AND U2630 ( .A(n2339), .B(n2340), .Z(n2338) );
  AND U2631 ( .A(n2341), .B(p_input[3737]), .Z(n2340) );
  AND U2632 ( .A(p_input[2737]), .B(p_input[1737]), .Z(n2341) );
  AND U2633 ( .A(p_input[5737]), .B(p_input[4737]), .Z(n2339) );
  AND U2634 ( .A(n2342), .B(n2343), .Z(n2337) );
  AND U2635 ( .A(n2344), .B(p_input[7737]), .Z(n2343) );
  AND U2636 ( .A(p_input[737]), .B(p_input[6737]), .Z(n2344) );
  AND U2637 ( .A(p_input[9737]), .B(p_input[8737]), .Z(n2342) );
  AND U2638 ( .A(n2345), .B(n2346), .Z(o[736]) );
  AND U2639 ( .A(n2347), .B(n2348), .Z(n2346) );
  AND U2640 ( .A(n2349), .B(p_input[3736]), .Z(n2348) );
  AND U2641 ( .A(p_input[2736]), .B(p_input[1736]), .Z(n2349) );
  AND U2642 ( .A(p_input[5736]), .B(p_input[4736]), .Z(n2347) );
  AND U2643 ( .A(n2350), .B(n2351), .Z(n2345) );
  AND U2644 ( .A(n2352), .B(p_input[7736]), .Z(n2351) );
  AND U2645 ( .A(p_input[736]), .B(p_input[6736]), .Z(n2352) );
  AND U2646 ( .A(p_input[9736]), .B(p_input[8736]), .Z(n2350) );
  AND U2647 ( .A(n2353), .B(n2354), .Z(o[735]) );
  AND U2648 ( .A(n2355), .B(n2356), .Z(n2354) );
  AND U2649 ( .A(n2357), .B(p_input[3735]), .Z(n2356) );
  AND U2650 ( .A(p_input[2735]), .B(p_input[1735]), .Z(n2357) );
  AND U2651 ( .A(p_input[5735]), .B(p_input[4735]), .Z(n2355) );
  AND U2652 ( .A(n2358), .B(n2359), .Z(n2353) );
  AND U2653 ( .A(n2360), .B(p_input[7735]), .Z(n2359) );
  AND U2654 ( .A(p_input[735]), .B(p_input[6735]), .Z(n2360) );
  AND U2655 ( .A(p_input[9735]), .B(p_input[8735]), .Z(n2358) );
  AND U2656 ( .A(n2361), .B(n2362), .Z(o[734]) );
  AND U2657 ( .A(n2363), .B(n2364), .Z(n2362) );
  AND U2658 ( .A(n2365), .B(p_input[3734]), .Z(n2364) );
  AND U2659 ( .A(p_input[2734]), .B(p_input[1734]), .Z(n2365) );
  AND U2660 ( .A(p_input[5734]), .B(p_input[4734]), .Z(n2363) );
  AND U2661 ( .A(n2366), .B(n2367), .Z(n2361) );
  AND U2662 ( .A(n2368), .B(p_input[7734]), .Z(n2367) );
  AND U2663 ( .A(p_input[734]), .B(p_input[6734]), .Z(n2368) );
  AND U2664 ( .A(p_input[9734]), .B(p_input[8734]), .Z(n2366) );
  AND U2665 ( .A(n2369), .B(n2370), .Z(o[733]) );
  AND U2666 ( .A(n2371), .B(n2372), .Z(n2370) );
  AND U2667 ( .A(n2373), .B(p_input[3733]), .Z(n2372) );
  AND U2668 ( .A(p_input[2733]), .B(p_input[1733]), .Z(n2373) );
  AND U2669 ( .A(p_input[5733]), .B(p_input[4733]), .Z(n2371) );
  AND U2670 ( .A(n2374), .B(n2375), .Z(n2369) );
  AND U2671 ( .A(n2376), .B(p_input[7733]), .Z(n2375) );
  AND U2672 ( .A(p_input[733]), .B(p_input[6733]), .Z(n2376) );
  AND U2673 ( .A(p_input[9733]), .B(p_input[8733]), .Z(n2374) );
  AND U2674 ( .A(n2377), .B(n2378), .Z(o[732]) );
  AND U2675 ( .A(n2379), .B(n2380), .Z(n2378) );
  AND U2676 ( .A(n2381), .B(p_input[3732]), .Z(n2380) );
  AND U2677 ( .A(p_input[2732]), .B(p_input[1732]), .Z(n2381) );
  AND U2678 ( .A(p_input[5732]), .B(p_input[4732]), .Z(n2379) );
  AND U2679 ( .A(n2382), .B(n2383), .Z(n2377) );
  AND U2680 ( .A(n2384), .B(p_input[7732]), .Z(n2383) );
  AND U2681 ( .A(p_input[732]), .B(p_input[6732]), .Z(n2384) );
  AND U2682 ( .A(p_input[9732]), .B(p_input[8732]), .Z(n2382) );
  AND U2683 ( .A(n2385), .B(n2386), .Z(o[731]) );
  AND U2684 ( .A(n2387), .B(n2388), .Z(n2386) );
  AND U2685 ( .A(n2389), .B(p_input[3731]), .Z(n2388) );
  AND U2686 ( .A(p_input[2731]), .B(p_input[1731]), .Z(n2389) );
  AND U2687 ( .A(p_input[5731]), .B(p_input[4731]), .Z(n2387) );
  AND U2688 ( .A(n2390), .B(n2391), .Z(n2385) );
  AND U2689 ( .A(n2392), .B(p_input[7731]), .Z(n2391) );
  AND U2690 ( .A(p_input[731]), .B(p_input[6731]), .Z(n2392) );
  AND U2691 ( .A(p_input[9731]), .B(p_input[8731]), .Z(n2390) );
  AND U2692 ( .A(n2393), .B(n2394), .Z(o[730]) );
  AND U2693 ( .A(n2395), .B(n2396), .Z(n2394) );
  AND U2694 ( .A(n2397), .B(p_input[3730]), .Z(n2396) );
  AND U2695 ( .A(p_input[2730]), .B(p_input[1730]), .Z(n2397) );
  AND U2696 ( .A(p_input[5730]), .B(p_input[4730]), .Z(n2395) );
  AND U2697 ( .A(n2398), .B(n2399), .Z(n2393) );
  AND U2698 ( .A(n2400), .B(p_input[7730]), .Z(n2399) );
  AND U2699 ( .A(p_input[730]), .B(p_input[6730]), .Z(n2400) );
  AND U2700 ( .A(p_input[9730]), .B(p_input[8730]), .Z(n2398) );
  AND U2701 ( .A(n2401), .B(n2402), .Z(o[72]) );
  AND U2702 ( .A(n2403), .B(n2404), .Z(n2402) );
  AND U2703 ( .A(n2405), .B(p_input[3072]), .Z(n2404) );
  AND U2704 ( .A(p_input[2072]), .B(p_input[1072]), .Z(n2405) );
  AND U2705 ( .A(p_input[5072]), .B(p_input[4072]), .Z(n2403) );
  AND U2706 ( .A(n2406), .B(n2407), .Z(n2401) );
  AND U2707 ( .A(n2408), .B(p_input[72]), .Z(n2407) );
  AND U2708 ( .A(p_input[7072]), .B(p_input[6072]), .Z(n2408) );
  AND U2709 ( .A(p_input[9072]), .B(p_input[8072]), .Z(n2406) );
  AND U2710 ( .A(n2409), .B(n2410), .Z(o[729]) );
  AND U2711 ( .A(n2411), .B(n2412), .Z(n2410) );
  AND U2712 ( .A(n2413), .B(p_input[3729]), .Z(n2412) );
  AND U2713 ( .A(p_input[2729]), .B(p_input[1729]), .Z(n2413) );
  AND U2714 ( .A(p_input[5729]), .B(p_input[4729]), .Z(n2411) );
  AND U2715 ( .A(n2414), .B(n2415), .Z(n2409) );
  AND U2716 ( .A(n2416), .B(p_input[7729]), .Z(n2415) );
  AND U2717 ( .A(p_input[729]), .B(p_input[6729]), .Z(n2416) );
  AND U2718 ( .A(p_input[9729]), .B(p_input[8729]), .Z(n2414) );
  AND U2719 ( .A(n2417), .B(n2418), .Z(o[728]) );
  AND U2720 ( .A(n2419), .B(n2420), .Z(n2418) );
  AND U2721 ( .A(n2421), .B(p_input[3728]), .Z(n2420) );
  AND U2722 ( .A(p_input[2728]), .B(p_input[1728]), .Z(n2421) );
  AND U2723 ( .A(p_input[5728]), .B(p_input[4728]), .Z(n2419) );
  AND U2724 ( .A(n2422), .B(n2423), .Z(n2417) );
  AND U2725 ( .A(n2424), .B(p_input[7728]), .Z(n2423) );
  AND U2726 ( .A(p_input[728]), .B(p_input[6728]), .Z(n2424) );
  AND U2727 ( .A(p_input[9728]), .B(p_input[8728]), .Z(n2422) );
  AND U2728 ( .A(n2425), .B(n2426), .Z(o[727]) );
  AND U2729 ( .A(n2427), .B(n2428), .Z(n2426) );
  AND U2730 ( .A(n2429), .B(p_input[3727]), .Z(n2428) );
  AND U2731 ( .A(p_input[2727]), .B(p_input[1727]), .Z(n2429) );
  AND U2732 ( .A(p_input[5727]), .B(p_input[4727]), .Z(n2427) );
  AND U2733 ( .A(n2430), .B(n2431), .Z(n2425) );
  AND U2734 ( .A(n2432), .B(p_input[7727]), .Z(n2431) );
  AND U2735 ( .A(p_input[727]), .B(p_input[6727]), .Z(n2432) );
  AND U2736 ( .A(p_input[9727]), .B(p_input[8727]), .Z(n2430) );
  AND U2737 ( .A(n2433), .B(n2434), .Z(o[726]) );
  AND U2738 ( .A(n2435), .B(n2436), .Z(n2434) );
  AND U2739 ( .A(n2437), .B(p_input[3726]), .Z(n2436) );
  AND U2740 ( .A(p_input[2726]), .B(p_input[1726]), .Z(n2437) );
  AND U2741 ( .A(p_input[5726]), .B(p_input[4726]), .Z(n2435) );
  AND U2742 ( .A(n2438), .B(n2439), .Z(n2433) );
  AND U2743 ( .A(n2440), .B(p_input[7726]), .Z(n2439) );
  AND U2744 ( .A(p_input[726]), .B(p_input[6726]), .Z(n2440) );
  AND U2745 ( .A(p_input[9726]), .B(p_input[8726]), .Z(n2438) );
  AND U2746 ( .A(n2441), .B(n2442), .Z(o[725]) );
  AND U2747 ( .A(n2443), .B(n2444), .Z(n2442) );
  AND U2748 ( .A(n2445), .B(p_input[3725]), .Z(n2444) );
  AND U2749 ( .A(p_input[2725]), .B(p_input[1725]), .Z(n2445) );
  AND U2750 ( .A(p_input[5725]), .B(p_input[4725]), .Z(n2443) );
  AND U2751 ( .A(n2446), .B(n2447), .Z(n2441) );
  AND U2752 ( .A(n2448), .B(p_input[7725]), .Z(n2447) );
  AND U2753 ( .A(p_input[725]), .B(p_input[6725]), .Z(n2448) );
  AND U2754 ( .A(p_input[9725]), .B(p_input[8725]), .Z(n2446) );
  AND U2755 ( .A(n2449), .B(n2450), .Z(o[724]) );
  AND U2756 ( .A(n2451), .B(n2452), .Z(n2450) );
  AND U2757 ( .A(n2453), .B(p_input[3724]), .Z(n2452) );
  AND U2758 ( .A(p_input[2724]), .B(p_input[1724]), .Z(n2453) );
  AND U2759 ( .A(p_input[5724]), .B(p_input[4724]), .Z(n2451) );
  AND U2760 ( .A(n2454), .B(n2455), .Z(n2449) );
  AND U2761 ( .A(n2456), .B(p_input[7724]), .Z(n2455) );
  AND U2762 ( .A(p_input[724]), .B(p_input[6724]), .Z(n2456) );
  AND U2763 ( .A(p_input[9724]), .B(p_input[8724]), .Z(n2454) );
  AND U2764 ( .A(n2457), .B(n2458), .Z(o[723]) );
  AND U2765 ( .A(n2459), .B(n2460), .Z(n2458) );
  AND U2766 ( .A(n2461), .B(p_input[3723]), .Z(n2460) );
  AND U2767 ( .A(p_input[2723]), .B(p_input[1723]), .Z(n2461) );
  AND U2768 ( .A(p_input[5723]), .B(p_input[4723]), .Z(n2459) );
  AND U2769 ( .A(n2462), .B(n2463), .Z(n2457) );
  AND U2770 ( .A(n2464), .B(p_input[7723]), .Z(n2463) );
  AND U2771 ( .A(p_input[723]), .B(p_input[6723]), .Z(n2464) );
  AND U2772 ( .A(p_input[9723]), .B(p_input[8723]), .Z(n2462) );
  AND U2773 ( .A(n2465), .B(n2466), .Z(o[722]) );
  AND U2774 ( .A(n2467), .B(n2468), .Z(n2466) );
  AND U2775 ( .A(n2469), .B(p_input[3722]), .Z(n2468) );
  AND U2776 ( .A(p_input[2722]), .B(p_input[1722]), .Z(n2469) );
  AND U2777 ( .A(p_input[5722]), .B(p_input[4722]), .Z(n2467) );
  AND U2778 ( .A(n2470), .B(n2471), .Z(n2465) );
  AND U2779 ( .A(n2472), .B(p_input[7722]), .Z(n2471) );
  AND U2780 ( .A(p_input[722]), .B(p_input[6722]), .Z(n2472) );
  AND U2781 ( .A(p_input[9722]), .B(p_input[8722]), .Z(n2470) );
  AND U2782 ( .A(n2473), .B(n2474), .Z(o[721]) );
  AND U2783 ( .A(n2475), .B(n2476), .Z(n2474) );
  AND U2784 ( .A(n2477), .B(p_input[3721]), .Z(n2476) );
  AND U2785 ( .A(p_input[2721]), .B(p_input[1721]), .Z(n2477) );
  AND U2786 ( .A(p_input[5721]), .B(p_input[4721]), .Z(n2475) );
  AND U2787 ( .A(n2478), .B(n2479), .Z(n2473) );
  AND U2788 ( .A(n2480), .B(p_input[7721]), .Z(n2479) );
  AND U2789 ( .A(p_input[721]), .B(p_input[6721]), .Z(n2480) );
  AND U2790 ( .A(p_input[9721]), .B(p_input[8721]), .Z(n2478) );
  AND U2791 ( .A(n2481), .B(n2482), .Z(o[720]) );
  AND U2792 ( .A(n2483), .B(n2484), .Z(n2482) );
  AND U2793 ( .A(n2485), .B(p_input[3720]), .Z(n2484) );
  AND U2794 ( .A(p_input[2720]), .B(p_input[1720]), .Z(n2485) );
  AND U2795 ( .A(p_input[5720]), .B(p_input[4720]), .Z(n2483) );
  AND U2796 ( .A(n2486), .B(n2487), .Z(n2481) );
  AND U2797 ( .A(n2488), .B(p_input[7720]), .Z(n2487) );
  AND U2798 ( .A(p_input[720]), .B(p_input[6720]), .Z(n2488) );
  AND U2799 ( .A(p_input[9720]), .B(p_input[8720]), .Z(n2486) );
  AND U2800 ( .A(n2489), .B(n2490), .Z(o[71]) );
  AND U2801 ( .A(n2491), .B(n2492), .Z(n2490) );
  AND U2802 ( .A(n2493), .B(p_input[3071]), .Z(n2492) );
  AND U2803 ( .A(p_input[2071]), .B(p_input[1071]), .Z(n2493) );
  AND U2804 ( .A(p_input[5071]), .B(p_input[4071]), .Z(n2491) );
  AND U2805 ( .A(n2494), .B(n2495), .Z(n2489) );
  AND U2806 ( .A(n2496), .B(p_input[71]), .Z(n2495) );
  AND U2807 ( .A(p_input[7071]), .B(p_input[6071]), .Z(n2496) );
  AND U2808 ( .A(p_input[9071]), .B(p_input[8071]), .Z(n2494) );
  AND U2809 ( .A(n2497), .B(n2498), .Z(o[719]) );
  AND U2810 ( .A(n2499), .B(n2500), .Z(n2498) );
  AND U2811 ( .A(n2501), .B(p_input[3719]), .Z(n2500) );
  AND U2812 ( .A(p_input[2719]), .B(p_input[1719]), .Z(n2501) );
  AND U2813 ( .A(p_input[5719]), .B(p_input[4719]), .Z(n2499) );
  AND U2814 ( .A(n2502), .B(n2503), .Z(n2497) );
  AND U2815 ( .A(n2504), .B(p_input[7719]), .Z(n2503) );
  AND U2816 ( .A(p_input[719]), .B(p_input[6719]), .Z(n2504) );
  AND U2817 ( .A(p_input[9719]), .B(p_input[8719]), .Z(n2502) );
  AND U2818 ( .A(n2505), .B(n2506), .Z(o[718]) );
  AND U2819 ( .A(n2507), .B(n2508), .Z(n2506) );
  AND U2820 ( .A(n2509), .B(p_input[3718]), .Z(n2508) );
  AND U2821 ( .A(p_input[2718]), .B(p_input[1718]), .Z(n2509) );
  AND U2822 ( .A(p_input[5718]), .B(p_input[4718]), .Z(n2507) );
  AND U2823 ( .A(n2510), .B(n2511), .Z(n2505) );
  AND U2824 ( .A(n2512), .B(p_input[7718]), .Z(n2511) );
  AND U2825 ( .A(p_input[718]), .B(p_input[6718]), .Z(n2512) );
  AND U2826 ( .A(p_input[9718]), .B(p_input[8718]), .Z(n2510) );
  AND U2827 ( .A(n2513), .B(n2514), .Z(o[717]) );
  AND U2828 ( .A(n2515), .B(n2516), .Z(n2514) );
  AND U2829 ( .A(n2517), .B(p_input[3717]), .Z(n2516) );
  AND U2830 ( .A(p_input[2717]), .B(p_input[1717]), .Z(n2517) );
  AND U2831 ( .A(p_input[5717]), .B(p_input[4717]), .Z(n2515) );
  AND U2832 ( .A(n2518), .B(n2519), .Z(n2513) );
  AND U2833 ( .A(n2520), .B(p_input[7717]), .Z(n2519) );
  AND U2834 ( .A(p_input[717]), .B(p_input[6717]), .Z(n2520) );
  AND U2835 ( .A(p_input[9717]), .B(p_input[8717]), .Z(n2518) );
  AND U2836 ( .A(n2521), .B(n2522), .Z(o[716]) );
  AND U2837 ( .A(n2523), .B(n2524), .Z(n2522) );
  AND U2838 ( .A(n2525), .B(p_input[3716]), .Z(n2524) );
  AND U2839 ( .A(p_input[2716]), .B(p_input[1716]), .Z(n2525) );
  AND U2840 ( .A(p_input[5716]), .B(p_input[4716]), .Z(n2523) );
  AND U2841 ( .A(n2526), .B(n2527), .Z(n2521) );
  AND U2842 ( .A(n2528), .B(p_input[7716]), .Z(n2527) );
  AND U2843 ( .A(p_input[716]), .B(p_input[6716]), .Z(n2528) );
  AND U2844 ( .A(p_input[9716]), .B(p_input[8716]), .Z(n2526) );
  AND U2845 ( .A(n2529), .B(n2530), .Z(o[715]) );
  AND U2846 ( .A(n2531), .B(n2532), .Z(n2530) );
  AND U2847 ( .A(n2533), .B(p_input[3715]), .Z(n2532) );
  AND U2848 ( .A(p_input[2715]), .B(p_input[1715]), .Z(n2533) );
  AND U2849 ( .A(p_input[5715]), .B(p_input[4715]), .Z(n2531) );
  AND U2850 ( .A(n2534), .B(n2535), .Z(n2529) );
  AND U2851 ( .A(n2536), .B(p_input[7715]), .Z(n2535) );
  AND U2852 ( .A(p_input[715]), .B(p_input[6715]), .Z(n2536) );
  AND U2853 ( .A(p_input[9715]), .B(p_input[8715]), .Z(n2534) );
  AND U2854 ( .A(n2537), .B(n2538), .Z(o[714]) );
  AND U2855 ( .A(n2539), .B(n2540), .Z(n2538) );
  AND U2856 ( .A(n2541), .B(p_input[3714]), .Z(n2540) );
  AND U2857 ( .A(p_input[2714]), .B(p_input[1714]), .Z(n2541) );
  AND U2858 ( .A(p_input[5714]), .B(p_input[4714]), .Z(n2539) );
  AND U2859 ( .A(n2542), .B(n2543), .Z(n2537) );
  AND U2860 ( .A(n2544), .B(p_input[7714]), .Z(n2543) );
  AND U2861 ( .A(p_input[714]), .B(p_input[6714]), .Z(n2544) );
  AND U2862 ( .A(p_input[9714]), .B(p_input[8714]), .Z(n2542) );
  AND U2863 ( .A(n2545), .B(n2546), .Z(o[713]) );
  AND U2864 ( .A(n2547), .B(n2548), .Z(n2546) );
  AND U2865 ( .A(n2549), .B(p_input[3713]), .Z(n2548) );
  AND U2866 ( .A(p_input[2713]), .B(p_input[1713]), .Z(n2549) );
  AND U2867 ( .A(p_input[5713]), .B(p_input[4713]), .Z(n2547) );
  AND U2868 ( .A(n2550), .B(n2551), .Z(n2545) );
  AND U2869 ( .A(n2552), .B(p_input[7713]), .Z(n2551) );
  AND U2870 ( .A(p_input[713]), .B(p_input[6713]), .Z(n2552) );
  AND U2871 ( .A(p_input[9713]), .B(p_input[8713]), .Z(n2550) );
  AND U2872 ( .A(n2553), .B(n2554), .Z(o[712]) );
  AND U2873 ( .A(n2555), .B(n2556), .Z(n2554) );
  AND U2874 ( .A(n2557), .B(p_input[3712]), .Z(n2556) );
  AND U2875 ( .A(p_input[2712]), .B(p_input[1712]), .Z(n2557) );
  AND U2876 ( .A(p_input[5712]), .B(p_input[4712]), .Z(n2555) );
  AND U2877 ( .A(n2558), .B(n2559), .Z(n2553) );
  AND U2878 ( .A(n2560), .B(p_input[7712]), .Z(n2559) );
  AND U2879 ( .A(p_input[712]), .B(p_input[6712]), .Z(n2560) );
  AND U2880 ( .A(p_input[9712]), .B(p_input[8712]), .Z(n2558) );
  AND U2881 ( .A(n2561), .B(n2562), .Z(o[711]) );
  AND U2882 ( .A(n2563), .B(n2564), .Z(n2562) );
  AND U2883 ( .A(n2565), .B(p_input[3711]), .Z(n2564) );
  AND U2884 ( .A(p_input[2711]), .B(p_input[1711]), .Z(n2565) );
  AND U2885 ( .A(p_input[5711]), .B(p_input[4711]), .Z(n2563) );
  AND U2886 ( .A(n2566), .B(n2567), .Z(n2561) );
  AND U2887 ( .A(n2568), .B(p_input[7711]), .Z(n2567) );
  AND U2888 ( .A(p_input[711]), .B(p_input[6711]), .Z(n2568) );
  AND U2889 ( .A(p_input[9711]), .B(p_input[8711]), .Z(n2566) );
  AND U2890 ( .A(n2569), .B(n2570), .Z(o[710]) );
  AND U2891 ( .A(n2571), .B(n2572), .Z(n2570) );
  AND U2892 ( .A(n2573), .B(p_input[3710]), .Z(n2572) );
  AND U2893 ( .A(p_input[2710]), .B(p_input[1710]), .Z(n2573) );
  AND U2894 ( .A(p_input[5710]), .B(p_input[4710]), .Z(n2571) );
  AND U2895 ( .A(n2574), .B(n2575), .Z(n2569) );
  AND U2896 ( .A(n2576), .B(p_input[7710]), .Z(n2575) );
  AND U2897 ( .A(p_input[710]), .B(p_input[6710]), .Z(n2576) );
  AND U2898 ( .A(p_input[9710]), .B(p_input[8710]), .Z(n2574) );
  AND U2899 ( .A(n2577), .B(n2578), .Z(o[70]) );
  AND U2900 ( .A(n2579), .B(n2580), .Z(n2578) );
  AND U2901 ( .A(n2581), .B(p_input[3070]), .Z(n2580) );
  AND U2902 ( .A(p_input[2070]), .B(p_input[1070]), .Z(n2581) );
  AND U2903 ( .A(p_input[5070]), .B(p_input[4070]), .Z(n2579) );
  AND U2904 ( .A(n2582), .B(n2583), .Z(n2577) );
  AND U2905 ( .A(n2584), .B(p_input[70]), .Z(n2583) );
  AND U2906 ( .A(p_input[7070]), .B(p_input[6070]), .Z(n2584) );
  AND U2907 ( .A(p_input[9070]), .B(p_input[8070]), .Z(n2582) );
  AND U2908 ( .A(n2585), .B(n2586), .Z(o[709]) );
  AND U2909 ( .A(n2587), .B(n2588), .Z(n2586) );
  AND U2910 ( .A(n2589), .B(p_input[3709]), .Z(n2588) );
  AND U2911 ( .A(p_input[2709]), .B(p_input[1709]), .Z(n2589) );
  AND U2912 ( .A(p_input[5709]), .B(p_input[4709]), .Z(n2587) );
  AND U2913 ( .A(n2590), .B(n2591), .Z(n2585) );
  AND U2914 ( .A(n2592), .B(p_input[7709]), .Z(n2591) );
  AND U2915 ( .A(p_input[709]), .B(p_input[6709]), .Z(n2592) );
  AND U2916 ( .A(p_input[9709]), .B(p_input[8709]), .Z(n2590) );
  AND U2917 ( .A(n2593), .B(n2594), .Z(o[708]) );
  AND U2918 ( .A(n2595), .B(n2596), .Z(n2594) );
  AND U2919 ( .A(n2597), .B(p_input[3708]), .Z(n2596) );
  AND U2920 ( .A(p_input[2708]), .B(p_input[1708]), .Z(n2597) );
  AND U2921 ( .A(p_input[5708]), .B(p_input[4708]), .Z(n2595) );
  AND U2922 ( .A(n2598), .B(n2599), .Z(n2593) );
  AND U2923 ( .A(n2600), .B(p_input[7708]), .Z(n2599) );
  AND U2924 ( .A(p_input[708]), .B(p_input[6708]), .Z(n2600) );
  AND U2925 ( .A(p_input[9708]), .B(p_input[8708]), .Z(n2598) );
  AND U2926 ( .A(n2601), .B(n2602), .Z(o[707]) );
  AND U2927 ( .A(n2603), .B(n2604), .Z(n2602) );
  AND U2928 ( .A(n2605), .B(p_input[3707]), .Z(n2604) );
  AND U2929 ( .A(p_input[2707]), .B(p_input[1707]), .Z(n2605) );
  AND U2930 ( .A(p_input[5707]), .B(p_input[4707]), .Z(n2603) );
  AND U2931 ( .A(n2606), .B(n2607), .Z(n2601) );
  AND U2932 ( .A(n2608), .B(p_input[7707]), .Z(n2607) );
  AND U2933 ( .A(p_input[707]), .B(p_input[6707]), .Z(n2608) );
  AND U2934 ( .A(p_input[9707]), .B(p_input[8707]), .Z(n2606) );
  AND U2935 ( .A(n2609), .B(n2610), .Z(o[706]) );
  AND U2936 ( .A(n2611), .B(n2612), .Z(n2610) );
  AND U2937 ( .A(n2613), .B(p_input[3706]), .Z(n2612) );
  AND U2938 ( .A(p_input[2706]), .B(p_input[1706]), .Z(n2613) );
  AND U2939 ( .A(p_input[5706]), .B(p_input[4706]), .Z(n2611) );
  AND U2940 ( .A(n2614), .B(n2615), .Z(n2609) );
  AND U2941 ( .A(n2616), .B(p_input[7706]), .Z(n2615) );
  AND U2942 ( .A(p_input[706]), .B(p_input[6706]), .Z(n2616) );
  AND U2943 ( .A(p_input[9706]), .B(p_input[8706]), .Z(n2614) );
  AND U2944 ( .A(n2617), .B(n2618), .Z(o[705]) );
  AND U2945 ( .A(n2619), .B(n2620), .Z(n2618) );
  AND U2946 ( .A(n2621), .B(p_input[3705]), .Z(n2620) );
  AND U2947 ( .A(p_input[2705]), .B(p_input[1705]), .Z(n2621) );
  AND U2948 ( .A(p_input[5705]), .B(p_input[4705]), .Z(n2619) );
  AND U2949 ( .A(n2622), .B(n2623), .Z(n2617) );
  AND U2950 ( .A(n2624), .B(p_input[7705]), .Z(n2623) );
  AND U2951 ( .A(p_input[705]), .B(p_input[6705]), .Z(n2624) );
  AND U2952 ( .A(p_input[9705]), .B(p_input[8705]), .Z(n2622) );
  AND U2953 ( .A(n2625), .B(n2626), .Z(o[704]) );
  AND U2954 ( .A(n2627), .B(n2628), .Z(n2626) );
  AND U2955 ( .A(n2629), .B(p_input[3704]), .Z(n2628) );
  AND U2956 ( .A(p_input[2704]), .B(p_input[1704]), .Z(n2629) );
  AND U2957 ( .A(p_input[5704]), .B(p_input[4704]), .Z(n2627) );
  AND U2958 ( .A(n2630), .B(n2631), .Z(n2625) );
  AND U2959 ( .A(n2632), .B(p_input[7704]), .Z(n2631) );
  AND U2960 ( .A(p_input[704]), .B(p_input[6704]), .Z(n2632) );
  AND U2961 ( .A(p_input[9704]), .B(p_input[8704]), .Z(n2630) );
  AND U2962 ( .A(n2633), .B(n2634), .Z(o[703]) );
  AND U2963 ( .A(n2635), .B(n2636), .Z(n2634) );
  AND U2964 ( .A(n2637), .B(p_input[3703]), .Z(n2636) );
  AND U2965 ( .A(p_input[2703]), .B(p_input[1703]), .Z(n2637) );
  AND U2966 ( .A(p_input[5703]), .B(p_input[4703]), .Z(n2635) );
  AND U2967 ( .A(n2638), .B(n2639), .Z(n2633) );
  AND U2968 ( .A(n2640), .B(p_input[7703]), .Z(n2639) );
  AND U2969 ( .A(p_input[703]), .B(p_input[6703]), .Z(n2640) );
  AND U2970 ( .A(p_input[9703]), .B(p_input[8703]), .Z(n2638) );
  AND U2971 ( .A(n2641), .B(n2642), .Z(o[702]) );
  AND U2972 ( .A(n2643), .B(n2644), .Z(n2642) );
  AND U2973 ( .A(n2645), .B(p_input[3702]), .Z(n2644) );
  AND U2974 ( .A(p_input[2702]), .B(p_input[1702]), .Z(n2645) );
  AND U2975 ( .A(p_input[5702]), .B(p_input[4702]), .Z(n2643) );
  AND U2976 ( .A(n2646), .B(n2647), .Z(n2641) );
  AND U2977 ( .A(n2648), .B(p_input[7702]), .Z(n2647) );
  AND U2978 ( .A(p_input[702]), .B(p_input[6702]), .Z(n2648) );
  AND U2979 ( .A(p_input[9702]), .B(p_input[8702]), .Z(n2646) );
  AND U2980 ( .A(n2649), .B(n2650), .Z(o[701]) );
  AND U2981 ( .A(n2651), .B(n2652), .Z(n2650) );
  AND U2982 ( .A(n2653), .B(p_input[3701]), .Z(n2652) );
  AND U2983 ( .A(p_input[2701]), .B(p_input[1701]), .Z(n2653) );
  AND U2984 ( .A(p_input[5701]), .B(p_input[4701]), .Z(n2651) );
  AND U2985 ( .A(n2654), .B(n2655), .Z(n2649) );
  AND U2986 ( .A(n2656), .B(p_input[7701]), .Z(n2655) );
  AND U2987 ( .A(p_input[701]), .B(p_input[6701]), .Z(n2656) );
  AND U2988 ( .A(p_input[9701]), .B(p_input[8701]), .Z(n2654) );
  AND U2989 ( .A(n2657), .B(n2658), .Z(o[700]) );
  AND U2990 ( .A(n2659), .B(n2660), .Z(n2658) );
  AND U2991 ( .A(n2661), .B(p_input[3700]), .Z(n2660) );
  AND U2992 ( .A(p_input[2700]), .B(p_input[1700]), .Z(n2661) );
  AND U2993 ( .A(p_input[5700]), .B(p_input[4700]), .Z(n2659) );
  AND U2994 ( .A(n2662), .B(n2663), .Z(n2657) );
  AND U2995 ( .A(n2664), .B(p_input[7700]), .Z(n2663) );
  AND U2996 ( .A(p_input[700]), .B(p_input[6700]), .Z(n2664) );
  AND U2997 ( .A(p_input[9700]), .B(p_input[8700]), .Z(n2662) );
  AND U2998 ( .A(n2665), .B(n2666), .Z(o[6]) );
  AND U2999 ( .A(n2667), .B(n2668), .Z(n2666) );
  AND U3000 ( .A(n2669), .B(p_input[3006]), .Z(n2668) );
  AND U3001 ( .A(p_input[2006]), .B(p_input[1006]), .Z(n2669) );
  AND U3002 ( .A(p_input[5006]), .B(p_input[4006]), .Z(n2667) );
  AND U3003 ( .A(n2670), .B(n2671), .Z(n2665) );
  AND U3004 ( .A(n2672), .B(p_input[7006]), .Z(n2671) );
  AND U3005 ( .A(p_input[6]), .B(p_input[6006]), .Z(n2672) );
  AND U3006 ( .A(p_input[9006]), .B(p_input[8006]), .Z(n2670) );
  AND U3007 ( .A(n2673), .B(n2674), .Z(o[69]) );
  AND U3008 ( .A(n2675), .B(n2676), .Z(n2674) );
  AND U3009 ( .A(n2677), .B(p_input[3069]), .Z(n2676) );
  AND U3010 ( .A(p_input[2069]), .B(p_input[1069]), .Z(n2677) );
  AND U3011 ( .A(p_input[5069]), .B(p_input[4069]), .Z(n2675) );
  AND U3012 ( .A(n2678), .B(n2679), .Z(n2673) );
  AND U3013 ( .A(n2680), .B(p_input[7069]), .Z(n2679) );
  AND U3014 ( .A(p_input[69]), .B(p_input[6069]), .Z(n2680) );
  AND U3015 ( .A(p_input[9069]), .B(p_input[8069]), .Z(n2678) );
  AND U3016 ( .A(n2681), .B(n2682), .Z(o[699]) );
  AND U3017 ( .A(n2683), .B(n2684), .Z(n2682) );
  AND U3018 ( .A(n2685), .B(p_input[3699]), .Z(n2684) );
  AND U3019 ( .A(p_input[2699]), .B(p_input[1699]), .Z(n2685) );
  AND U3020 ( .A(p_input[5699]), .B(p_input[4699]), .Z(n2683) );
  AND U3021 ( .A(n2686), .B(n2687), .Z(n2681) );
  AND U3022 ( .A(n2688), .B(p_input[7699]), .Z(n2687) );
  AND U3023 ( .A(p_input[699]), .B(p_input[6699]), .Z(n2688) );
  AND U3024 ( .A(p_input[9699]), .B(p_input[8699]), .Z(n2686) );
  AND U3025 ( .A(n2689), .B(n2690), .Z(o[698]) );
  AND U3026 ( .A(n2691), .B(n2692), .Z(n2690) );
  AND U3027 ( .A(n2693), .B(p_input[3698]), .Z(n2692) );
  AND U3028 ( .A(p_input[2698]), .B(p_input[1698]), .Z(n2693) );
  AND U3029 ( .A(p_input[5698]), .B(p_input[4698]), .Z(n2691) );
  AND U3030 ( .A(n2694), .B(n2695), .Z(n2689) );
  AND U3031 ( .A(n2696), .B(p_input[7698]), .Z(n2695) );
  AND U3032 ( .A(p_input[698]), .B(p_input[6698]), .Z(n2696) );
  AND U3033 ( .A(p_input[9698]), .B(p_input[8698]), .Z(n2694) );
  AND U3034 ( .A(n2697), .B(n2698), .Z(o[697]) );
  AND U3035 ( .A(n2699), .B(n2700), .Z(n2698) );
  AND U3036 ( .A(n2701), .B(p_input[3697]), .Z(n2700) );
  AND U3037 ( .A(p_input[2697]), .B(p_input[1697]), .Z(n2701) );
  AND U3038 ( .A(p_input[5697]), .B(p_input[4697]), .Z(n2699) );
  AND U3039 ( .A(n2702), .B(n2703), .Z(n2697) );
  AND U3040 ( .A(n2704), .B(p_input[7697]), .Z(n2703) );
  AND U3041 ( .A(p_input[697]), .B(p_input[6697]), .Z(n2704) );
  AND U3042 ( .A(p_input[9697]), .B(p_input[8697]), .Z(n2702) );
  AND U3043 ( .A(n2705), .B(n2706), .Z(o[696]) );
  AND U3044 ( .A(n2707), .B(n2708), .Z(n2706) );
  AND U3045 ( .A(n2709), .B(p_input[3696]), .Z(n2708) );
  AND U3046 ( .A(p_input[2696]), .B(p_input[1696]), .Z(n2709) );
  AND U3047 ( .A(p_input[5696]), .B(p_input[4696]), .Z(n2707) );
  AND U3048 ( .A(n2710), .B(n2711), .Z(n2705) );
  AND U3049 ( .A(n2712), .B(p_input[7696]), .Z(n2711) );
  AND U3050 ( .A(p_input[696]), .B(p_input[6696]), .Z(n2712) );
  AND U3051 ( .A(p_input[9696]), .B(p_input[8696]), .Z(n2710) );
  AND U3052 ( .A(n2713), .B(n2714), .Z(o[695]) );
  AND U3053 ( .A(n2715), .B(n2716), .Z(n2714) );
  AND U3054 ( .A(n2717), .B(p_input[3695]), .Z(n2716) );
  AND U3055 ( .A(p_input[2695]), .B(p_input[1695]), .Z(n2717) );
  AND U3056 ( .A(p_input[5695]), .B(p_input[4695]), .Z(n2715) );
  AND U3057 ( .A(n2718), .B(n2719), .Z(n2713) );
  AND U3058 ( .A(n2720), .B(p_input[7695]), .Z(n2719) );
  AND U3059 ( .A(p_input[695]), .B(p_input[6695]), .Z(n2720) );
  AND U3060 ( .A(p_input[9695]), .B(p_input[8695]), .Z(n2718) );
  AND U3061 ( .A(n2721), .B(n2722), .Z(o[694]) );
  AND U3062 ( .A(n2723), .B(n2724), .Z(n2722) );
  AND U3063 ( .A(n2725), .B(p_input[3694]), .Z(n2724) );
  AND U3064 ( .A(p_input[2694]), .B(p_input[1694]), .Z(n2725) );
  AND U3065 ( .A(p_input[5694]), .B(p_input[4694]), .Z(n2723) );
  AND U3066 ( .A(n2726), .B(n2727), .Z(n2721) );
  AND U3067 ( .A(n2728), .B(p_input[7694]), .Z(n2727) );
  AND U3068 ( .A(p_input[694]), .B(p_input[6694]), .Z(n2728) );
  AND U3069 ( .A(p_input[9694]), .B(p_input[8694]), .Z(n2726) );
  AND U3070 ( .A(n2729), .B(n2730), .Z(o[693]) );
  AND U3071 ( .A(n2731), .B(n2732), .Z(n2730) );
  AND U3072 ( .A(n2733), .B(p_input[3693]), .Z(n2732) );
  AND U3073 ( .A(p_input[2693]), .B(p_input[1693]), .Z(n2733) );
  AND U3074 ( .A(p_input[5693]), .B(p_input[4693]), .Z(n2731) );
  AND U3075 ( .A(n2734), .B(n2735), .Z(n2729) );
  AND U3076 ( .A(n2736), .B(p_input[7693]), .Z(n2735) );
  AND U3077 ( .A(p_input[693]), .B(p_input[6693]), .Z(n2736) );
  AND U3078 ( .A(p_input[9693]), .B(p_input[8693]), .Z(n2734) );
  AND U3079 ( .A(n2737), .B(n2738), .Z(o[692]) );
  AND U3080 ( .A(n2739), .B(n2740), .Z(n2738) );
  AND U3081 ( .A(n2741), .B(p_input[3692]), .Z(n2740) );
  AND U3082 ( .A(p_input[2692]), .B(p_input[1692]), .Z(n2741) );
  AND U3083 ( .A(p_input[5692]), .B(p_input[4692]), .Z(n2739) );
  AND U3084 ( .A(n2742), .B(n2743), .Z(n2737) );
  AND U3085 ( .A(n2744), .B(p_input[7692]), .Z(n2743) );
  AND U3086 ( .A(p_input[692]), .B(p_input[6692]), .Z(n2744) );
  AND U3087 ( .A(p_input[9692]), .B(p_input[8692]), .Z(n2742) );
  AND U3088 ( .A(n2745), .B(n2746), .Z(o[691]) );
  AND U3089 ( .A(n2747), .B(n2748), .Z(n2746) );
  AND U3090 ( .A(n2749), .B(p_input[3691]), .Z(n2748) );
  AND U3091 ( .A(p_input[2691]), .B(p_input[1691]), .Z(n2749) );
  AND U3092 ( .A(p_input[5691]), .B(p_input[4691]), .Z(n2747) );
  AND U3093 ( .A(n2750), .B(n2751), .Z(n2745) );
  AND U3094 ( .A(n2752), .B(p_input[7691]), .Z(n2751) );
  AND U3095 ( .A(p_input[691]), .B(p_input[6691]), .Z(n2752) );
  AND U3096 ( .A(p_input[9691]), .B(p_input[8691]), .Z(n2750) );
  AND U3097 ( .A(n2753), .B(n2754), .Z(o[690]) );
  AND U3098 ( .A(n2755), .B(n2756), .Z(n2754) );
  AND U3099 ( .A(n2757), .B(p_input[3690]), .Z(n2756) );
  AND U3100 ( .A(p_input[2690]), .B(p_input[1690]), .Z(n2757) );
  AND U3101 ( .A(p_input[5690]), .B(p_input[4690]), .Z(n2755) );
  AND U3102 ( .A(n2758), .B(n2759), .Z(n2753) );
  AND U3103 ( .A(n2760), .B(p_input[7690]), .Z(n2759) );
  AND U3104 ( .A(p_input[690]), .B(p_input[6690]), .Z(n2760) );
  AND U3105 ( .A(p_input[9690]), .B(p_input[8690]), .Z(n2758) );
  AND U3106 ( .A(n2761), .B(n2762), .Z(o[68]) );
  AND U3107 ( .A(n2763), .B(n2764), .Z(n2762) );
  AND U3108 ( .A(n2765), .B(p_input[3068]), .Z(n2764) );
  AND U3109 ( .A(p_input[2068]), .B(p_input[1068]), .Z(n2765) );
  AND U3110 ( .A(p_input[5068]), .B(p_input[4068]), .Z(n2763) );
  AND U3111 ( .A(n2766), .B(n2767), .Z(n2761) );
  AND U3112 ( .A(n2768), .B(p_input[7068]), .Z(n2767) );
  AND U3113 ( .A(p_input[68]), .B(p_input[6068]), .Z(n2768) );
  AND U3114 ( .A(p_input[9068]), .B(p_input[8068]), .Z(n2766) );
  AND U3115 ( .A(n2769), .B(n2770), .Z(o[689]) );
  AND U3116 ( .A(n2771), .B(n2772), .Z(n2770) );
  AND U3117 ( .A(n2773), .B(p_input[3689]), .Z(n2772) );
  AND U3118 ( .A(p_input[2689]), .B(p_input[1689]), .Z(n2773) );
  AND U3119 ( .A(p_input[5689]), .B(p_input[4689]), .Z(n2771) );
  AND U3120 ( .A(n2774), .B(n2775), .Z(n2769) );
  AND U3121 ( .A(n2776), .B(p_input[7689]), .Z(n2775) );
  AND U3122 ( .A(p_input[689]), .B(p_input[6689]), .Z(n2776) );
  AND U3123 ( .A(p_input[9689]), .B(p_input[8689]), .Z(n2774) );
  AND U3124 ( .A(n2777), .B(n2778), .Z(o[688]) );
  AND U3125 ( .A(n2779), .B(n2780), .Z(n2778) );
  AND U3126 ( .A(n2781), .B(p_input[3688]), .Z(n2780) );
  AND U3127 ( .A(p_input[2688]), .B(p_input[1688]), .Z(n2781) );
  AND U3128 ( .A(p_input[5688]), .B(p_input[4688]), .Z(n2779) );
  AND U3129 ( .A(n2782), .B(n2783), .Z(n2777) );
  AND U3130 ( .A(n2784), .B(p_input[7688]), .Z(n2783) );
  AND U3131 ( .A(p_input[688]), .B(p_input[6688]), .Z(n2784) );
  AND U3132 ( .A(p_input[9688]), .B(p_input[8688]), .Z(n2782) );
  AND U3133 ( .A(n2785), .B(n2786), .Z(o[687]) );
  AND U3134 ( .A(n2787), .B(n2788), .Z(n2786) );
  AND U3135 ( .A(n2789), .B(p_input[3687]), .Z(n2788) );
  AND U3136 ( .A(p_input[2687]), .B(p_input[1687]), .Z(n2789) );
  AND U3137 ( .A(p_input[5687]), .B(p_input[4687]), .Z(n2787) );
  AND U3138 ( .A(n2790), .B(n2791), .Z(n2785) );
  AND U3139 ( .A(n2792), .B(p_input[7687]), .Z(n2791) );
  AND U3140 ( .A(p_input[687]), .B(p_input[6687]), .Z(n2792) );
  AND U3141 ( .A(p_input[9687]), .B(p_input[8687]), .Z(n2790) );
  AND U3142 ( .A(n2793), .B(n2794), .Z(o[686]) );
  AND U3143 ( .A(n2795), .B(n2796), .Z(n2794) );
  AND U3144 ( .A(n2797), .B(p_input[3686]), .Z(n2796) );
  AND U3145 ( .A(p_input[2686]), .B(p_input[1686]), .Z(n2797) );
  AND U3146 ( .A(p_input[5686]), .B(p_input[4686]), .Z(n2795) );
  AND U3147 ( .A(n2798), .B(n2799), .Z(n2793) );
  AND U3148 ( .A(n2800), .B(p_input[7686]), .Z(n2799) );
  AND U3149 ( .A(p_input[686]), .B(p_input[6686]), .Z(n2800) );
  AND U3150 ( .A(p_input[9686]), .B(p_input[8686]), .Z(n2798) );
  AND U3151 ( .A(n2801), .B(n2802), .Z(o[685]) );
  AND U3152 ( .A(n2803), .B(n2804), .Z(n2802) );
  AND U3153 ( .A(n2805), .B(p_input[3685]), .Z(n2804) );
  AND U3154 ( .A(p_input[2685]), .B(p_input[1685]), .Z(n2805) );
  AND U3155 ( .A(p_input[5685]), .B(p_input[4685]), .Z(n2803) );
  AND U3156 ( .A(n2806), .B(n2807), .Z(n2801) );
  AND U3157 ( .A(n2808), .B(p_input[7685]), .Z(n2807) );
  AND U3158 ( .A(p_input[685]), .B(p_input[6685]), .Z(n2808) );
  AND U3159 ( .A(p_input[9685]), .B(p_input[8685]), .Z(n2806) );
  AND U3160 ( .A(n2809), .B(n2810), .Z(o[684]) );
  AND U3161 ( .A(n2811), .B(n2812), .Z(n2810) );
  AND U3162 ( .A(n2813), .B(p_input[3684]), .Z(n2812) );
  AND U3163 ( .A(p_input[2684]), .B(p_input[1684]), .Z(n2813) );
  AND U3164 ( .A(p_input[5684]), .B(p_input[4684]), .Z(n2811) );
  AND U3165 ( .A(n2814), .B(n2815), .Z(n2809) );
  AND U3166 ( .A(n2816), .B(p_input[7684]), .Z(n2815) );
  AND U3167 ( .A(p_input[684]), .B(p_input[6684]), .Z(n2816) );
  AND U3168 ( .A(p_input[9684]), .B(p_input[8684]), .Z(n2814) );
  AND U3169 ( .A(n2817), .B(n2818), .Z(o[683]) );
  AND U3170 ( .A(n2819), .B(n2820), .Z(n2818) );
  AND U3171 ( .A(n2821), .B(p_input[3683]), .Z(n2820) );
  AND U3172 ( .A(p_input[2683]), .B(p_input[1683]), .Z(n2821) );
  AND U3173 ( .A(p_input[5683]), .B(p_input[4683]), .Z(n2819) );
  AND U3174 ( .A(n2822), .B(n2823), .Z(n2817) );
  AND U3175 ( .A(n2824), .B(p_input[7683]), .Z(n2823) );
  AND U3176 ( .A(p_input[683]), .B(p_input[6683]), .Z(n2824) );
  AND U3177 ( .A(p_input[9683]), .B(p_input[8683]), .Z(n2822) );
  AND U3178 ( .A(n2825), .B(n2826), .Z(o[682]) );
  AND U3179 ( .A(n2827), .B(n2828), .Z(n2826) );
  AND U3180 ( .A(n2829), .B(p_input[3682]), .Z(n2828) );
  AND U3181 ( .A(p_input[2682]), .B(p_input[1682]), .Z(n2829) );
  AND U3182 ( .A(p_input[5682]), .B(p_input[4682]), .Z(n2827) );
  AND U3183 ( .A(n2830), .B(n2831), .Z(n2825) );
  AND U3184 ( .A(n2832), .B(p_input[7682]), .Z(n2831) );
  AND U3185 ( .A(p_input[682]), .B(p_input[6682]), .Z(n2832) );
  AND U3186 ( .A(p_input[9682]), .B(p_input[8682]), .Z(n2830) );
  AND U3187 ( .A(n2833), .B(n2834), .Z(o[681]) );
  AND U3188 ( .A(n2835), .B(n2836), .Z(n2834) );
  AND U3189 ( .A(n2837), .B(p_input[3681]), .Z(n2836) );
  AND U3190 ( .A(p_input[2681]), .B(p_input[1681]), .Z(n2837) );
  AND U3191 ( .A(p_input[5681]), .B(p_input[4681]), .Z(n2835) );
  AND U3192 ( .A(n2838), .B(n2839), .Z(n2833) );
  AND U3193 ( .A(n2840), .B(p_input[7681]), .Z(n2839) );
  AND U3194 ( .A(p_input[681]), .B(p_input[6681]), .Z(n2840) );
  AND U3195 ( .A(p_input[9681]), .B(p_input[8681]), .Z(n2838) );
  AND U3196 ( .A(n2841), .B(n2842), .Z(o[680]) );
  AND U3197 ( .A(n2843), .B(n2844), .Z(n2842) );
  AND U3198 ( .A(n2845), .B(p_input[3680]), .Z(n2844) );
  AND U3199 ( .A(p_input[2680]), .B(p_input[1680]), .Z(n2845) );
  AND U3200 ( .A(p_input[5680]), .B(p_input[4680]), .Z(n2843) );
  AND U3201 ( .A(n2846), .B(n2847), .Z(n2841) );
  AND U3202 ( .A(n2848), .B(p_input[7680]), .Z(n2847) );
  AND U3203 ( .A(p_input[680]), .B(p_input[6680]), .Z(n2848) );
  AND U3204 ( .A(p_input[9680]), .B(p_input[8680]), .Z(n2846) );
  AND U3205 ( .A(n2849), .B(n2850), .Z(o[67]) );
  AND U3206 ( .A(n2851), .B(n2852), .Z(n2850) );
  AND U3207 ( .A(n2853), .B(p_input[3067]), .Z(n2852) );
  AND U3208 ( .A(p_input[2067]), .B(p_input[1067]), .Z(n2853) );
  AND U3209 ( .A(p_input[5067]), .B(p_input[4067]), .Z(n2851) );
  AND U3210 ( .A(n2854), .B(n2855), .Z(n2849) );
  AND U3211 ( .A(n2856), .B(p_input[7067]), .Z(n2855) );
  AND U3212 ( .A(p_input[67]), .B(p_input[6067]), .Z(n2856) );
  AND U3213 ( .A(p_input[9067]), .B(p_input[8067]), .Z(n2854) );
  AND U3214 ( .A(n2857), .B(n2858), .Z(o[679]) );
  AND U3215 ( .A(n2859), .B(n2860), .Z(n2858) );
  AND U3216 ( .A(n2861), .B(p_input[3679]), .Z(n2860) );
  AND U3217 ( .A(p_input[2679]), .B(p_input[1679]), .Z(n2861) );
  AND U3218 ( .A(p_input[5679]), .B(p_input[4679]), .Z(n2859) );
  AND U3219 ( .A(n2862), .B(n2863), .Z(n2857) );
  AND U3220 ( .A(n2864), .B(p_input[7679]), .Z(n2863) );
  AND U3221 ( .A(p_input[679]), .B(p_input[6679]), .Z(n2864) );
  AND U3222 ( .A(p_input[9679]), .B(p_input[8679]), .Z(n2862) );
  AND U3223 ( .A(n2865), .B(n2866), .Z(o[678]) );
  AND U3224 ( .A(n2867), .B(n2868), .Z(n2866) );
  AND U3225 ( .A(n2869), .B(p_input[3678]), .Z(n2868) );
  AND U3226 ( .A(p_input[2678]), .B(p_input[1678]), .Z(n2869) );
  AND U3227 ( .A(p_input[5678]), .B(p_input[4678]), .Z(n2867) );
  AND U3228 ( .A(n2870), .B(n2871), .Z(n2865) );
  AND U3229 ( .A(n2872), .B(p_input[7678]), .Z(n2871) );
  AND U3230 ( .A(p_input[678]), .B(p_input[6678]), .Z(n2872) );
  AND U3231 ( .A(p_input[9678]), .B(p_input[8678]), .Z(n2870) );
  AND U3232 ( .A(n2873), .B(n2874), .Z(o[677]) );
  AND U3233 ( .A(n2875), .B(n2876), .Z(n2874) );
  AND U3234 ( .A(n2877), .B(p_input[3677]), .Z(n2876) );
  AND U3235 ( .A(p_input[2677]), .B(p_input[1677]), .Z(n2877) );
  AND U3236 ( .A(p_input[5677]), .B(p_input[4677]), .Z(n2875) );
  AND U3237 ( .A(n2878), .B(n2879), .Z(n2873) );
  AND U3238 ( .A(n2880), .B(p_input[7677]), .Z(n2879) );
  AND U3239 ( .A(p_input[677]), .B(p_input[6677]), .Z(n2880) );
  AND U3240 ( .A(p_input[9677]), .B(p_input[8677]), .Z(n2878) );
  AND U3241 ( .A(n2881), .B(n2882), .Z(o[676]) );
  AND U3242 ( .A(n2883), .B(n2884), .Z(n2882) );
  AND U3243 ( .A(n2885), .B(p_input[3676]), .Z(n2884) );
  AND U3244 ( .A(p_input[2676]), .B(p_input[1676]), .Z(n2885) );
  AND U3245 ( .A(p_input[5676]), .B(p_input[4676]), .Z(n2883) );
  AND U3246 ( .A(n2886), .B(n2887), .Z(n2881) );
  AND U3247 ( .A(n2888), .B(p_input[7676]), .Z(n2887) );
  AND U3248 ( .A(p_input[676]), .B(p_input[6676]), .Z(n2888) );
  AND U3249 ( .A(p_input[9676]), .B(p_input[8676]), .Z(n2886) );
  AND U3250 ( .A(n2889), .B(n2890), .Z(o[675]) );
  AND U3251 ( .A(n2891), .B(n2892), .Z(n2890) );
  AND U3252 ( .A(n2893), .B(p_input[3675]), .Z(n2892) );
  AND U3253 ( .A(p_input[2675]), .B(p_input[1675]), .Z(n2893) );
  AND U3254 ( .A(p_input[5675]), .B(p_input[4675]), .Z(n2891) );
  AND U3255 ( .A(n2894), .B(n2895), .Z(n2889) );
  AND U3256 ( .A(n2896), .B(p_input[7675]), .Z(n2895) );
  AND U3257 ( .A(p_input[675]), .B(p_input[6675]), .Z(n2896) );
  AND U3258 ( .A(p_input[9675]), .B(p_input[8675]), .Z(n2894) );
  AND U3259 ( .A(n2897), .B(n2898), .Z(o[674]) );
  AND U3260 ( .A(n2899), .B(n2900), .Z(n2898) );
  AND U3261 ( .A(n2901), .B(p_input[3674]), .Z(n2900) );
  AND U3262 ( .A(p_input[2674]), .B(p_input[1674]), .Z(n2901) );
  AND U3263 ( .A(p_input[5674]), .B(p_input[4674]), .Z(n2899) );
  AND U3264 ( .A(n2902), .B(n2903), .Z(n2897) );
  AND U3265 ( .A(n2904), .B(p_input[7674]), .Z(n2903) );
  AND U3266 ( .A(p_input[674]), .B(p_input[6674]), .Z(n2904) );
  AND U3267 ( .A(p_input[9674]), .B(p_input[8674]), .Z(n2902) );
  AND U3268 ( .A(n2905), .B(n2906), .Z(o[673]) );
  AND U3269 ( .A(n2907), .B(n2908), .Z(n2906) );
  AND U3270 ( .A(n2909), .B(p_input[3673]), .Z(n2908) );
  AND U3271 ( .A(p_input[2673]), .B(p_input[1673]), .Z(n2909) );
  AND U3272 ( .A(p_input[5673]), .B(p_input[4673]), .Z(n2907) );
  AND U3273 ( .A(n2910), .B(n2911), .Z(n2905) );
  AND U3274 ( .A(n2912), .B(p_input[7673]), .Z(n2911) );
  AND U3275 ( .A(p_input[673]), .B(p_input[6673]), .Z(n2912) );
  AND U3276 ( .A(p_input[9673]), .B(p_input[8673]), .Z(n2910) );
  AND U3277 ( .A(n2913), .B(n2914), .Z(o[672]) );
  AND U3278 ( .A(n2915), .B(n2916), .Z(n2914) );
  AND U3279 ( .A(n2917), .B(p_input[3672]), .Z(n2916) );
  AND U3280 ( .A(p_input[2672]), .B(p_input[1672]), .Z(n2917) );
  AND U3281 ( .A(p_input[5672]), .B(p_input[4672]), .Z(n2915) );
  AND U3282 ( .A(n2918), .B(n2919), .Z(n2913) );
  AND U3283 ( .A(n2920), .B(p_input[7672]), .Z(n2919) );
  AND U3284 ( .A(p_input[672]), .B(p_input[6672]), .Z(n2920) );
  AND U3285 ( .A(p_input[9672]), .B(p_input[8672]), .Z(n2918) );
  AND U3286 ( .A(n2921), .B(n2922), .Z(o[671]) );
  AND U3287 ( .A(n2923), .B(n2924), .Z(n2922) );
  AND U3288 ( .A(n2925), .B(p_input[3671]), .Z(n2924) );
  AND U3289 ( .A(p_input[2671]), .B(p_input[1671]), .Z(n2925) );
  AND U3290 ( .A(p_input[5671]), .B(p_input[4671]), .Z(n2923) );
  AND U3291 ( .A(n2926), .B(n2927), .Z(n2921) );
  AND U3292 ( .A(n2928), .B(p_input[7671]), .Z(n2927) );
  AND U3293 ( .A(p_input[671]), .B(p_input[6671]), .Z(n2928) );
  AND U3294 ( .A(p_input[9671]), .B(p_input[8671]), .Z(n2926) );
  AND U3295 ( .A(n2929), .B(n2930), .Z(o[670]) );
  AND U3296 ( .A(n2931), .B(n2932), .Z(n2930) );
  AND U3297 ( .A(n2933), .B(p_input[3670]), .Z(n2932) );
  AND U3298 ( .A(p_input[2670]), .B(p_input[1670]), .Z(n2933) );
  AND U3299 ( .A(p_input[5670]), .B(p_input[4670]), .Z(n2931) );
  AND U3300 ( .A(n2934), .B(n2935), .Z(n2929) );
  AND U3301 ( .A(n2936), .B(p_input[7670]), .Z(n2935) );
  AND U3302 ( .A(p_input[670]), .B(p_input[6670]), .Z(n2936) );
  AND U3303 ( .A(p_input[9670]), .B(p_input[8670]), .Z(n2934) );
  AND U3304 ( .A(n2937), .B(n2938), .Z(o[66]) );
  AND U3305 ( .A(n2939), .B(n2940), .Z(n2938) );
  AND U3306 ( .A(n2941), .B(p_input[3066]), .Z(n2940) );
  AND U3307 ( .A(p_input[2066]), .B(p_input[1066]), .Z(n2941) );
  AND U3308 ( .A(p_input[5066]), .B(p_input[4066]), .Z(n2939) );
  AND U3309 ( .A(n2942), .B(n2943), .Z(n2937) );
  AND U3310 ( .A(n2944), .B(p_input[7066]), .Z(n2943) );
  AND U3311 ( .A(p_input[66]), .B(p_input[6066]), .Z(n2944) );
  AND U3312 ( .A(p_input[9066]), .B(p_input[8066]), .Z(n2942) );
  AND U3313 ( .A(n2945), .B(n2946), .Z(o[669]) );
  AND U3314 ( .A(n2947), .B(n2948), .Z(n2946) );
  AND U3315 ( .A(n2949), .B(p_input[3669]), .Z(n2948) );
  AND U3316 ( .A(p_input[2669]), .B(p_input[1669]), .Z(n2949) );
  AND U3317 ( .A(p_input[5669]), .B(p_input[4669]), .Z(n2947) );
  AND U3318 ( .A(n2950), .B(n2951), .Z(n2945) );
  AND U3319 ( .A(n2952), .B(p_input[7669]), .Z(n2951) );
  AND U3320 ( .A(p_input[669]), .B(p_input[6669]), .Z(n2952) );
  AND U3321 ( .A(p_input[9669]), .B(p_input[8669]), .Z(n2950) );
  AND U3322 ( .A(n2953), .B(n2954), .Z(o[668]) );
  AND U3323 ( .A(n2955), .B(n2956), .Z(n2954) );
  AND U3324 ( .A(n2957), .B(p_input[3668]), .Z(n2956) );
  AND U3325 ( .A(p_input[2668]), .B(p_input[1668]), .Z(n2957) );
  AND U3326 ( .A(p_input[5668]), .B(p_input[4668]), .Z(n2955) );
  AND U3327 ( .A(n2958), .B(n2959), .Z(n2953) );
  AND U3328 ( .A(n2960), .B(p_input[7668]), .Z(n2959) );
  AND U3329 ( .A(p_input[668]), .B(p_input[6668]), .Z(n2960) );
  AND U3330 ( .A(p_input[9668]), .B(p_input[8668]), .Z(n2958) );
  AND U3331 ( .A(n2961), .B(n2962), .Z(o[667]) );
  AND U3332 ( .A(n2963), .B(n2964), .Z(n2962) );
  AND U3333 ( .A(n2965), .B(p_input[3667]), .Z(n2964) );
  AND U3334 ( .A(p_input[2667]), .B(p_input[1667]), .Z(n2965) );
  AND U3335 ( .A(p_input[5667]), .B(p_input[4667]), .Z(n2963) );
  AND U3336 ( .A(n2966), .B(n2967), .Z(n2961) );
  AND U3337 ( .A(n2968), .B(p_input[7667]), .Z(n2967) );
  AND U3338 ( .A(p_input[667]), .B(p_input[6667]), .Z(n2968) );
  AND U3339 ( .A(p_input[9667]), .B(p_input[8667]), .Z(n2966) );
  AND U3340 ( .A(n2969), .B(n2970), .Z(o[666]) );
  AND U3341 ( .A(n2971), .B(n2972), .Z(n2970) );
  AND U3342 ( .A(n2973), .B(p_input[3666]), .Z(n2972) );
  AND U3343 ( .A(p_input[2666]), .B(p_input[1666]), .Z(n2973) );
  AND U3344 ( .A(p_input[5666]), .B(p_input[4666]), .Z(n2971) );
  AND U3345 ( .A(n2974), .B(n2975), .Z(n2969) );
  AND U3346 ( .A(n2976), .B(p_input[7666]), .Z(n2975) );
  AND U3347 ( .A(p_input[666]), .B(p_input[6666]), .Z(n2976) );
  AND U3348 ( .A(p_input[9666]), .B(p_input[8666]), .Z(n2974) );
  AND U3349 ( .A(n2977), .B(n2978), .Z(o[665]) );
  AND U3350 ( .A(n2979), .B(n2980), .Z(n2978) );
  AND U3351 ( .A(n2981), .B(p_input[3665]), .Z(n2980) );
  AND U3352 ( .A(p_input[2665]), .B(p_input[1665]), .Z(n2981) );
  AND U3353 ( .A(p_input[5665]), .B(p_input[4665]), .Z(n2979) );
  AND U3354 ( .A(n2982), .B(n2983), .Z(n2977) );
  AND U3355 ( .A(n2984), .B(p_input[7665]), .Z(n2983) );
  AND U3356 ( .A(p_input[6665]), .B(p_input[665]), .Z(n2984) );
  AND U3357 ( .A(p_input[9665]), .B(p_input[8665]), .Z(n2982) );
  AND U3358 ( .A(n2985), .B(n2986), .Z(o[664]) );
  AND U3359 ( .A(n2987), .B(n2988), .Z(n2986) );
  AND U3360 ( .A(n2989), .B(p_input[3664]), .Z(n2988) );
  AND U3361 ( .A(p_input[2664]), .B(p_input[1664]), .Z(n2989) );
  AND U3362 ( .A(p_input[5664]), .B(p_input[4664]), .Z(n2987) );
  AND U3363 ( .A(n2990), .B(n2991), .Z(n2985) );
  AND U3364 ( .A(n2992), .B(p_input[7664]), .Z(n2991) );
  AND U3365 ( .A(p_input[6664]), .B(p_input[664]), .Z(n2992) );
  AND U3366 ( .A(p_input[9664]), .B(p_input[8664]), .Z(n2990) );
  AND U3367 ( .A(n2993), .B(n2994), .Z(o[663]) );
  AND U3368 ( .A(n2995), .B(n2996), .Z(n2994) );
  AND U3369 ( .A(n2997), .B(p_input[3663]), .Z(n2996) );
  AND U3370 ( .A(p_input[2663]), .B(p_input[1663]), .Z(n2997) );
  AND U3371 ( .A(p_input[5663]), .B(p_input[4663]), .Z(n2995) );
  AND U3372 ( .A(n2998), .B(n2999), .Z(n2993) );
  AND U3373 ( .A(n3000), .B(p_input[7663]), .Z(n2999) );
  AND U3374 ( .A(p_input[6663]), .B(p_input[663]), .Z(n3000) );
  AND U3375 ( .A(p_input[9663]), .B(p_input[8663]), .Z(n2998) );
  AND U3376 ( .A(n3001), .B(n3002), .Z(o[662]) );
  AND U3377 ( .A(n3003), .B(n3004), .Z(n3002) );
  AND U3378 ( .A(n3005), .B(p_input[3662]), .Z(n3004) );
  AND U3379 ( .A(p_input[2662]), .B(p_input[1662]), .Z(n3005) );
  AND U3380 ( .A(p_input[5662]), .B(p_input[4662]), .Z(n3003) );
  AND U3381 ( .A(n3006), .B(n3007), .Z(n3001) );
  AND U3382 ( .A(n3008), .B(p_input[7662]), .Z(n3007) );
  AND U3383 ( .A(p_input[6662]), .B(p_input[662]), .Z(n3008) );
  AND U3384 ( .A(p_input[9662]), .B(p_input[8662]), .Z(n3006) );
  AND U3385 ( .A(n3009), .B(n3010), .Z(o[661]) );
  AND U3386 ( .A(n3011), .B(n3012), .Z(n3010) );
  AND U3387 ( .A(n3013), .B(p_input[3661]), .Z(n3012) );
  AND U3388 ( .A(p_input[2661]), .B(p_input[1661]), .Z(n3013) );
  AND U3389 ( .A(p_input[5661]), .B(p_input[4661]), .Z(n3011) );
  AND U3390 ( .A(n3014), .B(n3015), .Z(n3009) );
  AND U3391 ( .A(n3016), .B(p_input[7661]), .Z(n3015) );
  AND U3392 ( .A(p_input[6661]), .B(p_input[661]), .Z(n3016) );
  AND U3393 ( .A(p_input[9661]), .B(p_input[8661]), .Z(n3014) );
  AND U3394 ( .A(n3017), .B(n3018), .Z(o[660]) );
  AND U3395 ( .A(n3019), .B(n3020), .Z(n3018) );
  AND U3396 ( .A(n3021), .B(p_input[3660]), .Z(n3020) );
  AND U3397 ( .A(p_input[2660]), .B(p_input[1660]), .Z(n3021) );
  AND U3398 ( .A(p_input[5660]), .B(p_input[4660]), .Z(n3019) );
  AND U3399 ( .A(n3022), .B(n3023), .Z(n3017) );
  AND U3400 ( .A(n3024), .B(p_input[7660]), .Z(n3023) );
  AND U3401 ( .A(p_input[6660]), .B(p_input[660]), .Z(n3024) );
  AND U3402 ( .A(p_input[9660]), .B(p_input[8660]), .Z(n3022) );
  AND U3403 ( .A(n3025), .B(n3026), .Z(o[65]) );
  AND U3404 ( .A(n3027), .B(n3028), .Z(n3026) );
  AND U3405 ( .A(n3029), .B(p_input[3065]), .Z(n3028) );
  AND U3406 ( .A(p_input[2065]), .B(p_input[1065]), .Z(n3029) );
  AND U3407 ( .A(p_input[5065]), .B(p_input[4065]), .Z(n3027) );
  AND U3408 ( .A(n3030), .B(n3031), .Z(n3025) );
  AND U3409 ( .A(n3032), .B(p_input[7065]), .Z(n3031) );
  AND U3410 ( .A(p_input[65]), .B(p_input[6065]), .Z(n3032) );
  AND U3411 ( .A(p_input[9065]), .B(p_input[8065]), .Z(n3030) );
  AND U3412 ( .A(n3033), .B(n3034), .Z(o[659]) );
  AND U3413 ( .A(n3035), .B(n3036), .Z(n3034) );
  AND U3414 ( .A(n3037), .B(p_input[3659]), .Z(n3036) );
  AND U3415 ( .A(p_input[2659]), .B(p_input[1659]), .Z(n3037) );
  AND U3416 ( .A(p_input[5659]), .B(p_input[4659]), .Z(n3035) );
  AND U3417 ( .A(n3038), .B(n3039), .Z(n3033) );
  AND U3418 ( .A(n3040), .B(p_input[7659]), .Z(n3039) );
  AND U3419 ( .A(p_input[6659]), .B(p_input[659]), .Z(n3040) );
  AND U3420 ( .A(p_input[9659]), .B(p_input[8659]), .Z(n3038) );
  AND U3421 ( .A(n3041), .B(n3042), .Z(o[658]) );
  AND U3422 ( .A(n3043), .B(n3044), .Z(n3042) );
  AND U3423 ( .A(n3045), .B(p_input[3658]), .Z(n3044) );
  AND U3424 ( .A(p_input[2658]), .B(p_input[1658]), .Z(n3045) );
  AND U3425 ( .A(p_input[5658]), .B(p_input[4658]), .Z(n3043) );
  AND U3426 ( .A(n3046), .B(n3047), .Z(n3041) );
  AND U3427 ( .A(n3048), .B(p_input[7658]), .Z(n3047) );
  AND U3428 ( .A(p_input[6658]), .B(p_input[658]), .Z(n3048) );
  AND U3429 ( .A(p_input[9658]), .B(p_input[8658]), .Z(n3046) );
  AND U3430 ( .A(n3049), .B(n3050), .Z(o[657]) );
  AND U3431 ( .A(n3051), .B(n3052), .Z(n3050) );
  AND U3432 ( .A(n3053), .B(p_input[3657]), .Z(n3052) );
  AND U3433 ( .A(p_input[2657]), .B(p_input[1657]), .Z(n3053) );
  AND U3434 ( .A(p_input[5657]), .B(p_input[4657]), .Z(n3051) );
  AND U3435 ( .A(n3054), .B(n3055), .Z(n3049) );
  AND U3436 ( .A(n3056), .B(p_input[7657]), .Z(n3055) );
  AND U3437 ( .A(p_input[6657]), .B(p_input[657]), .Z(n3056) );
  AND U3438 ( .A(p_input[9657]), .B(p_input[8657]), .Z(n3054) );
  AND U3439 ( .A(n3057), .B(n3058), .Z(o[656]) );
  AND U3440 ( .A(n3059), .B(n3060), .Z(n3058) );
  AND U3441 ( .A(n3061), .B(p_input[3656]), .Z(n3060) );
  AND U3442 ( .A(p_input[2656]), .B(p_input[1656]), .Z(n3061) );
  AND U3443 ( .A(p_input[5656]), .B(p_input[4656]), .Z(n3059) );
  AND U3444 ( .A(n3062), .B(n3063), .Z(n3057) );
  AND U3445 ( .A(n3064), .B(p_input[7656]), .Z(n3063) );
  AND U3446 ( .A(p_input[6656]), .B(p_input[656]), .Z(n3064) );
  AND U3447 ( .A(p_input[9656]), .B(p_input[8656]), .Z(n3062) );
  AND U3448 ( .A(n3065), .B(n3066), .Z(o[655]) );
  AND U3449 ( .A(n3067), .B(n3068), .Z(n3066) );
  AND U3450 ( .A(n3069), .B(p_input[3655]), .Z(n3068) );
  AND U3451 ( .A(p_input[2655]), .B(p_input[1655]), .Z(n3069) );
  AND U3452 ( .A(p_input[5655]), .B(p_input[4655]), .Z(n3067) );
  AND U3453 ( .A(n3070), .B(n3071), .Z(n3065) );
  AND U3454 ( .A(n3072), .B(p_input[7655]), .Z(n3071) );
  AND U3455 ( .A(p_input[6655]), .B(p_input[655]), .Z(n3072) );
  AND U3456 ( .A(p_input[9655]), .B(p_input[8655]), .Z(n3070) );
  AND U3457 ( .A(n3073), .B(n3074), .Z(o[654]) );
  AND U3458 ( .A(n3075), .B(n3076), .Z(n3074) );
  AND U3459 ( .A(n3077), .B(p_input[3654]), .Z(n3076) );
  AND U3460 ( .A(p_input[2654]), .B(p_input[1654]), .Z(n3077) );
  AND U3461 ( .A(p_input[5654]), .B(p_input[4654]), .Z(n3075) );
  AND U3462 ( .A(n3078), .B(n3079), .Z(n3073) );
  AND U3463 ( .A(n3080), .B(p_input[7654]), .Z(n3079) );
  AND U3464 ( .A(p_input[6654]), .B(p_input[654]), .Z(n3080) );
  AND U3465 ( .A(p_input[9654]), .B(p_input[8654]), .Z(n3078) );
  AND U3466 ( .A(n3081), .B(n3082), .Z(o[653]) );
  AND U3467 ( .A(n3083), .B(n3084), .Z(n3082) );
  AND U3468 ( .A(n3085), .B(p_input[3653]), .Z(n3084) );
  AND U3469 ( .A(p_input[2653]), .B(p_input[1653]), .Z(n3085) );
  AND U3470 ( .A(p_input[5653]), .B(p_input[4653]), .Z(n3083) );
  AND U3471 ( .A(n3086), .B(n3087), .Z(n3081) );
  AND U3472 ( .A(n3088), .B(p_input[7653]), .Z(n3087) );
  AND U3473 ( .A(p_input[6653]), .B(p_input[653]), .Z(n3088) );
  AND U3474 ( .A(p_input[9653]), .B(p_input[8653]), .Z(n3086) );
  AND U3475 ( .A(n3089), .B(n3090), .Z(o[652]) );
  AND U3476 ( .A(n3091), .B(n3092), .Z(n3090) );
  AND U3477 ( .A(n3093), .B(p_input[3652]), .Z(n3092) );
  AND U3478 ( .A(p_input[2652]), .B(p_input[1652]), .Z(n3093) );
  AND U3479 ( .A(p_input[5652]), .B(p_input[4652]), .Z(n3091) );
  AND U3480 ( .A(n3094), .B(n3095), .Z(n3089) );
  AND U3481 ( .A(n3096), .B(p_input[7652]), .Z(n3095) );
  AND U3482 ( .A(p_input[6652]), .B(p_input[652]), .Z(n3096) );
  AND U3483 ( .A(p_input[9652]), .B(p_input[8652]), .Z(n3094) );
  AND U3484 ( .A(n3097), .B(n3098), .Z(o[651]) );
  AND U3485 ( .A(n3099), .B(n3100), .Z(n3098) );
  AND U3486 ( .A(n3101), .B(p_input[3651]), .Z(n3100) );
  AND U3487 ( .A(p_input[2651]), .B(p_input[1651]), .Z(n3101) );
  AND U3488 ( .A(p_input[5651]), .B(p_input[4651]), .Z(n3099) );
  AND U3489 ( .A(n3102), .B(n3103), .Z(n3097) );
  AND U3490 ( .A(n3104), .B(p_input[7651]), .Z(n3103) );
  AND U3491 ( .A(p_input[6651]), .B(p_input[651]), .Z(n3104) );
  AND U3492 ( .A(p_input[9651]), .B(p_input[8651]), .Z(n3102) );
  AND U3493 ( .A(n3105), .B(n3106), .Z(o[650]) );
  AND U3494 ( .A(n3107), .B(n3108), .Z(n3106) );
  AND U3495 ( .A(n3109), .B(p_input[3650]), .Z(n3108) );
  AND U3496 ( .A(p_input[2650]), .B(p_input[1650]), .Z(n3109) );
  AND U3497 ( .A(p_input[5650]), .B(p_input[4650]), .Z(n3107) );
  AND U3498 ( .A(n3110), .B(n3111), .Z(n3105) );
  AND U3499 ( .A(n3112), .B(p_input[7650]), .Z(n3111) );
  AND U3500 ( .A(p_input[6650]), .B(p_input[650]), .Z(n3112) );
  AND U3501 ( .A(p_input[9650]), .B(p_input[8650]), .Z(n3110) );
  AND U3502 ( .A(n3113), .B(n3114), .Z(o[64]) );
  AND U3503 ( .A(n3115), .B(n3116), .Z(n3114) );
  AND U3504 ( .A(n3117), .B(p_input[3064]), .Z(n3116) );
  AND U3505 ( .A(p_input[2064]), .B(p_input[1064]), .Z(n3117) );
  AND U3506 ( .A(p_input[5064]), .B(p_input[4064]), .Z(n3115) );
  AND U3507 ( .A(n3118), .B(n3119), .Z(n3113) );
  AND U3508 ( .A(n3120), .B(p_input[7064]), .Z(n3119) );
  AND U3509 ( .A(p_input[64]), .B(p_input[6064]), .Z(n3120) );
  AND U3510 ( .A(p_input[9064]), .B(p_input[8064]), .Z(n3118) );
  AND U3511 ( .A(n3121), .B(n3122), .Z(o[649]) );
  AND U3512 ( .A(n3123), .B(n3124), .Z(n3122) );
  AND U3513 ( .A(n3125), .B(p_input[3649]), .Z(n3124) );
  AND U3514 ( .A(p_input[2649]), .B(p_input[1649]), .Z(n3125) );
  AND U3515 ( .A(p_input[5649]), .B(p_input[4649]), .Z(n3123) );
  AND U3516 ( .A(n3126), .B(n3127), .Z(n3121) );
  AND U3517 ( .A(n3128), .B(p_input[7649]), .Z(n3127) );
  AND U3518 ( .A(p_input[6649]), .B(p_input[649]), .Z(n3128) );
  AND U3519 ( .A(p_input[9649]), .B(p_input[8649]), .Z(n3126) );
  AND U3520 ( .A(n3129), .B(n3130), .Z(o[648]) );
  AND U3521 ( .A(n3131), .B(n3132), .Z(n3130) );
  AND U3522 ( .A(n3133), .B(p_input[3648]), .Z(n3132) );
  AND U3523 ( .A(p_input[2648]), .B(p_input[1648]), .Z(n3133) );
  AND U3524 ( .A(p_input[5648]), .B(p_input[4648]), .Z(n3131) );
  AND U3525 ( .A(n3134), .B(n3135), .Z(n3129) );
  AND U3526 ( .A(n3136), .B(p_input[7648]), .Z(n3135) );
  AND U3527 ( .A(p_input[6648]), .B(p_input[648]), .Z(n3136) );
  AND U3528 ( .A(p_input[9648]), .B(p_input[8648]), .Z(n3134) );
  AND U3529 ( .A(n3137), .B(n3138), .Z(o[647]) );
  AND U3530 ( .A(n3139), .B(n3140), .Z(n3138) );
  AND U3531 ( .A(n3141), .B(p_input[3647]), .Z(n3140) );
  AND U3532 ( .A(p_input[2647]), .B(p_input[1647]), .Z(n3141) );
  AND U3533 ( .A(p_input[5647]), .B(p_input[4647]), .Z(n3139) );
  AND U3534 ( .A(n3142), .B(n3143), .Z(n3137) );
  AND U3535 ( .A(n3144), .B(p_input[7647]), .Z(n3143) );
  AND U3536 ( .A(p_input[6647]), .B(p_input[647]), .Z(n3144) );
  AND U3537 ( .A(p_input[9647]), .B(p_input[8647]), .Z(n3142) );
  AND U3538 ( .A(n3145), .B(n3146), .Z(o[646]) );
  AND U3539 ( .A(n3147), .B(n3148), .Z(n3146) );
  AND U3540 ( .A(n3149), .B(p_input[3646]), .Z(n3148) );
  AND U3541 ( .A(p_input[2646]), .B(p_input[1646]), .Z(n3149) );
  AND U3542 ( .A(p_input[5646]), .B(p_input[4646]), .Z(n3147) );
  AND U3543 ( .A(n3150), .B(n3151), .Z(n3145) );
  AND U3544 ( .A(n3152), .B(p_input[7646]), .Z(n3151) );
  AND U3545 ( .A(p_input[6646]), .B(p_input[646]), .Z(n3152) );
  AND U3546 ( .A(p_input[9646]), .B(p_input[8646]), .Z(n3150) );
  AND U3547 ( .A(n3153), .B(n3154), .Z(o[645]) );
  AND U3548 ( .A(n3155), .B(n3156), .Z(n3154) );
  AND U3549 ( .A(n3157), .B(p_input[3645]), .Z(n3156) );
  AND U3550 ( .A(p_input[2645]), .B(p_input[1645]), .Z(n3157) );
  AND U3551 ( .A(p_input[5645]), .B(p_input[4645]), .Z(n3155) );
  AND U3552 ( .A(n3158), .B(n3159), .Z(n3153) );
  AND U3553 ( .A(n3160), .B(p_input[7645]), .Z(n3159) );
  AND U3554 ( .A(p_input[6645]), .B(p_input[645]), .Z(n3160) );
  AND U3555 ( .A(p_input[9645]), .B(p_input[8645]), .Z(n3158) );
  AND U3556 ( .A(n3161), .B(n3162), .Z(o[644]) );
  AND U3557 ( .A(n3163), .B(n3164), .Z(n3162) );
  AND U3558 ( .A(n3165), .B(p_input[3644]), .Z(n3164) );
  AND U3559 ( .A(p_input[2644]), .B(p_input[1644]), .Z(n3165) );
  AND U3560 ( .A(p_input[5644]), .B(p_input[4644]), .Z(n3163) );
  AND U3561 ( .A(n3166), .B(n3167), .Z(n3161) );
  AND U3562 ( .A(n3168), .B(p_input[7644]), .Z(n3167) );
  AND U3563 ( .A(p_input[6644]), .B(p_input[644]), .Z(n3168) );
  AND U3564 ( .A(p_input[9644]), .B(p_input[8644]), .Z(n3166) );
  AND U3565 ( .A(n3169), .B(n3170), .Z(o[643]) );
  AND U3566 ( .A(n3171), .B(n3172), .Z(n3170) );
  AND U3567 ( .A(n3173), .B(p_input[3643]), .Z(n3172) );
  AND U3568 ( .A(p_input[2643]), .B(p_input[1643]), .Z(n3173) );
  AND U3569 ( .A(p_input[5643]), .B(p_input[4643]), .Z(n3171) );
  AND U3570 ( .A(n3174), .B(n3175), .Z(n3169) );
  AND U3571 ( .A(n3176), .B(p_input[7643]), .Z(n3175) );
  AND U3572 ( .A(p_input[6643]), .B(p_input[643]), .Z(n3176) );
  AND U3573 ( .A(p_input[9643]), .B(p_input[8643]), .Z(n3174) );
  AND U3574 ( .A(n3177), .B(n3178), .Z(o[642]) );
  AND U3575 ( .A(n3179), .B(n3180), .Z(n3178) );
  AND U3576 ( .A(n3181), .B(p_input[3642]), .Z(n3180) );
  AND U3577 ( .A(p_input[2642]), .B(p_input[1642]), .Z(n3181) );
  AND U3578 ( .A(p_input[5642]), .B(p_input[4642]), .Z(n3179) );
  AND U3579 ( .A(n3182), .B(n3183), .Z(n3177) );
  AND U3580 ( .A(n3184), .B(p_input[7642]), .Z(n3183) );
  AND U3581 ( .A(p_input[6642]), .B(p_input[642]), .Z(n3184) );
  AND U3582 ( .A(p_input[9642]), .B(p_input[8642]), .Z(n3182) );
  AND U3583 ( .A(n3185), .B(n3186), .Z(o[641]) );
  AND U3584 ( .A(n3187), .B(n3188), .Z(n3186) );
  AND U3585 ( .A(n3189), .B(p_input[3641]), .Z(n3188) );
  AND U3586 ( .A(p_input[2641]), .B(p_input[1641]), .Z(n3189) );
  AND U3587 ( .A(p_input[5641]), .B(p_input[4641]), .Z(n3187) );
  AND U3588 ( .A(n3190), .B(n3191), .Z(n3185) );
  AND U3589 ( .A(n3192), .B(p_input[7641]), .Z(n3191) );
  AND U3590 ( .A(p_input[6641]), .B(p_input[641]), .Z(n3192) );
  AND U3591 ( .A(p_input[9641]), .B(p_input[8641]), .Z(n3190) );
  AND U3592 ( .A(n3193), .B(n3194), .Z(o[640]) );
  AND U3593 ( .A(n3195), .B(n3196), .Z(n3194) );
  AND U3594 ( .A(n3197), .B(p_input[3640]), .Z(n3196) );
  AND U3595 ( .A(p_input[2640]), .B(p_input[1640]), .Z(n3197) );
  AND U3596 ( .A(p_input[5640]), .B(p_input[4640]), .Z(n3195) );
  AND U3597 ( .A(n3198), .B(n3199), .Z(n3193) );
  AND U3598 ( .A(n3200), .B(p_input[7640]), .Z(n3199) );
  AND U3599 ( .A(p_input[6640]), .B(p_input[640]), .Z(n3200) );
  AND U3600 ( .A(p_input[9640]), .B(p_input[8640]), .Z(n3198) );
  AND U3601 ( .A(n3201), .B(n3202), .Z(o[63]) );
  AND U3602 ( .A(n3203), .B(n3204), .Z(n3202) );
  AND U3603 ( .A(n3205), .B(p_input[3063]), .Z(n3204) );
  AND U3604 ( .A(p_input[2063]), .B(p_input[1063]), .Z(n3205) );
  AND U3605 ( .A(p_input[5063]), .B(p_input[4063]), .Z(n3203) );
  AND U3606 ( .A(n3206), .B(n3207), .Z(n3201) );
  AND U3607 ( .A(n3208), .B(p_input[7063]), .Z(n3207) );
  AND U3608 ( .A(p_input[63]), .B(p_input[6063]), .Z(n3208) );
  AND U3609 ( .A(p_input[9063]), .B(p_input[8063]), .Z(n3206) );
  AND U3610 ( .A(n3209), .B(n3210), .Z(o[639]) );
  AND U3611 ( .A(n3211), .B(n3212), .Z(n3210) );
  AND U3612 ( .A(n3213), .B(p_input[3639]), .Z(n3212) );
  AND U3613 ( .A(p_input[2639]), .B(p_input[1639]), .Z(n3213) );
  AND U3614 ( .A(p_input[5639]), .B(p_input[4639]), .Z(n3211) );
  AND U3615 ( .A(n3214), .B(n3215), .Z(n3209) );
  AND U3616 ( .A(n3216), .B(p_input[7639]), .Z(n3215) );
  AND U3617 ( .A(p_input[6639]), .B(p_input[639]), .Z(n3216) );
  AND U3618 ( .A(p_input[9639]), .B(p_input[8639]), .Z(n3214) );
  AND U3619 ( .A(n3217), .B(n3218), .Z(o[638]) );
  AND U3620 ( .A(n3219), .B(n3220), .Z(n3218) );
  AND U3621 ( .A(n3221), .B(p_input[3638]), .Z(n3220) );
  AND U3622 ( .A(p_input[2638]), .B(p_input[1638]), .Z(n3221) );
  AND U3623 ( .A(p_input[5638]), .B(p_input[4638]), .Z(n3219) );
  AND U3624 ( .A(n3222), .B(n3223), .Z(n3217) );
  AND U3625 ( .A(n3224), .B(p_input[7638]), .Z(n3223) );
  AND U3626 ( .A(p_input[6638]), .B(p_input[638]), .Z(n3224) );
  AND U3627 ( .A(p_input[9638]), .B(p_input[8638]), .Z(n3222) );
  AND U3628 ( .A(n3225), .B(n3226), .Z(o[637]) );
  AND U3629 ( .A(n3227), .B(n3228), .Z(n3226) );
  AND U3630 ( .A(n3229), .B(p_input[3637]), .Z(n3228) );
  AND U3631 ( .A(p_input[2637]), .B(p_input[1637]), .Z(n3229) );
  AND U3632 ( .A(p_input[5637]), .B(p_input[4637]), .Z(n3227) );
  AND U3633 ( .A(n3230), .B(n3231), .Z(n3225) );
  AND U3634 ( .A(n3232), .B(p_input[7637]), .Z(n3231) );
  AND U3635 ( .A(p_input[6637]), .B(p_input[637]), .Z(n3232) );
  AND U3636 ( .A(p_input[9637]), .B(p_input[8637]), .Z(n3230) );
  AND U3637 ( .A(n3233), .B(n3234), .Z(o[636]) );
  AND U3638 ( .A(n3235), .B(n3236), .Z(n3234) );
  AND U3639 ( .A(n3237), .B(p_input[3636]), .Z(n3236) );
  AND U3640 ( .A(p_input[2636]), .B(p_input[1636]), .Z(n3237) );
  AND U3641 ( .A(p_input[5636]), .B(p_input[4636]), .Z(n3235) );
  AND U3642 ( .A(n3238), .B(n3239), .Z(n3233) );
  AND U3643 ( .A(n3240), .B(p_input[7636]), .Z(n3239) );
  AND U3644 ( .A(p_input[6636]), .B(p_input[636]), .Z(n3240) );
  AND U3645 ( .A(p_input[9636]), .B(p_input[8636]), .Z(n3238) );
  AND U3646 ( .A(n3241), .B(n3242), .Z(o[635]) );
  AND U3647 ( .A(n3243), .B(n3244), .Z(n3242) );
  AND U3648 ( .A(n3245), .B(p_input[3635]), .Z(n3244) );
  AND U3649 ( .A(p_input[2635]), .B(p_input[1635]), .Z(n3245) );
  AND U3650 ( .A(p_input[5635]), .B(p_input[4635]), .Z(n3243) );
  AND U3651 ( .A(n3246), .B(n3247), .Z(n3241) );
  AND U3652 ( .A(n3248), .B(p_input[7635]), .Z(n3247) );
  AND U3653 ( .A(p_input[6635]), .B(p_input[635]), .Z(n3248) );
  AND U3654 ( .A(p_input[9635]), .B(p_input[8635]), .Z(n3246) );
  AND U3655 ( .A(n3249), .B(n3250), .Z(o[634]) );
  AND U3656 ( .A(n3251), .B(n3252), .Z(n3250) );
  AND U3657 ( .A(n3253), .B(p_input[3634]), .Z(n3252) );
  AND U3658 ( .A(p_input[2634]), .B(p_input[1634]), .Z(n3253) );
  AND U3659 ( .A(p_input[5634]), .B(p_input[4634]), .Z(n3251) );
  AND U3660 ( .A(n3254), .B(n3255), .Z(n3249) );
  AND U3661 ( .A(n3256), .B(p_input[7634]), .Z(n3255) );
  AND U3662 ( .A(p_input[6634]), .B(p_input[634]), .Z(n3256) );
  AND U3663 ( .A(p_input[9634]), .B(p_input[8634]), .Z(n3254) );
  AND U3664 ( .A(n3257), .B(n3258), .Z(o[633]) );
  AND U3665 ( .A(n3259), .B(n3260), .Z(n3258) );
  AND U3666 ( .A(n3261), .B(p_input[3633]), .Z(n3260) );
  AND U3667 ( .A(p_input[2633]), .B(p_input[1633]), .Z(n3261) );
  AND U3668 ( .A(p_input[5633]), .B(p_input[4633]), .Z(n3259) );
  AND U3669 ( .A(n3262), .B(n3263), .Z(n3257) );
  AND U3670 ( .A(n3264), .B(p_input[7633]), .Z(n3263) );
  AND U3671 ( .A(p_input[6633]), .B(p_input[633]), .Z(n3264) );
  AND U3672 ( .A(p_input[9633]), .B(p_input[8633]), .Z(n3262) );
  AND U3673 ( .A(n3265), .B(n3266), .Z(o[632]) );
  AND U3674 ( .A(n3267), .B(n3268), .Z(n3266) );
  AND U3675 ( .A(n3269), .B(p_input[3632]), .Z(n3268) );
  AND U3676 ( .A(p_input[2632]), .B(p_input[1632]), .Z(n3269) );
  AND U3677 ( .A(p_input[5632]), .B(p_input[4632]), .Z(n3267) );
  AND U3678 ( .A(n3270), .B(n3271), .Z(n3265) );
  AND U3679 ( .A(n3272), .B(p_input[7632]), .Z(n3271) );
  AND U3680 ( .A(p_input[6632]), .B(p_input[632]), .Z(n3272) );
  AND U3681 ( .A(p_input[9632]), .B(p_input[8632]), .Z(n3270) );
  AND U3682 ( .A(n3273), .B(n3274), .Z(o[631]) );
  AND U3683 ( .A(n3275), .B(n3276), .Z(n3274) );
  AND U3684 ( .A(n3277), .B(p_input[3631]), .Z(n3276) );
  AND U3685 ( .A(p_input[2631]), .B(p_input[1631]), .Z(n3277) );
  AND U3686 ( .A(p_input[5631]), .B(p_input[4631]), .Z(n3275) );
  AND U3687 ( .A(n3278), .B(n3279), .Z(n3273) );
  AND U3688 ( .A(n3280), .B(p_input[7631]), .Z(n3279) );
  AND U3689 ( .A(p_input[6631]), .B(p_input[631]), .Z(n3280) );
  AND U3690 ( .A(p_input[9631]), .B(p_input[8631]), .Z(n3278) );
  AND U3691 ( .A(n3281), .B(n3282), .Z(o[630]) );
  AND U3692 ( .A(n3283), .B(n3284), .Z(n3282) );
  AND U3693 ( .A(n3285), .B(p_input[3630]), .Z(n3284) );
  AND U3694 ( .A(p_input[2630]), .B(p_input[1630]), .Z(n3285) );
  AND U3695 ( .A(p_input[5630]), .B(p_input[4630]), .Z(n3283) );
  AND U3696 ( .A(n3286), .B(n3287), .Z(n3281) );
  AND U3697 ( .A(n3288), .B(p_input[7630]), .Z(n3287) );
  AND U3698 ( .A(p_input[6630]), .B(p_input[630]), .Z(n3288) );
  AND U3699 ( .A(p_input[9630]), .B(p_input[8630]), .Z(n3286) );
  AND U3700 ( .A(n3289), .B(n3290), .Z(o[62]) );
  AND U3701 ( .A(n3291), .B(n3292), .Z(n3290) );
  AND U3702 ( .A(n3293), .B(p_input[3062]), .Z(n3292) );
  AND U3703 ( .A(p_input[2062]), .B(p_input[1062]), .Z(n3293) );
  AND U3704 ( .A(p_input[5062]), .B(p_input[4062]), .Z(n3291) );
  AND U3705 ( .A(n3294), .B(n3295), .Z(n3289) );
  AND U3706 ( .A(n3296), .B(p_input[7062]), .Z(n3295) );
  AND U3707 ( .A(p_input[62]), .B(p_input[6062]), .Z(n3296) );
  AND U3708 ( .A(p_input[9062]), .B(p_input[8062]), .Z(n3294) );
  AND U3709 ( .A(n3297), .B(n3298), .Z(o[629]) );
  AND U3710 ( .A(n3299), .B(n3300), .Z(n3298) );
  AND U3711 ( .A(n3301), .B(p_input[3629]), .Z(n3300) );
  AND U3712 ( .A(p_input[2629]), .B(p_input[1629]), .Z(n3301) );
  AND U3713 ( .A(p_input[5629]), .B(p_input[4629]), .Z(n3299) );
  AND U3714 ( .A(n3302), .B(n3303), .Z(n3297) );
  AND U3715 ( .A(n3304), .B(p_input[7629]), .Z(n3303) );
  AND U3716 ( .A(p_input[6629]), .B(p_input[629]), .Z(n3304) );
  AND U3717 ( .A(p_input[9629]), .B(p_input[8629]), .Z(n3302) );
  AND U3718 ( .A(n3305), .B(n3306), .Z(o[628]) );
  AND U3719 ( .A(n3307), .B(n3308), .Z(n3306) );
  AND U3720 ( .A(n3309), .B(p_input[3628]), .Z(n3308) );
  AND U3721 ( .A(p_input[2628]), .B(p_input[1628]), .Z(n3309) );
  AND U3722 ( .A(p_input[5628]), .B(p_input[4628]), .Z(n3307) );
  AND U3723 ( .A(n3310), .B(n3311), .Z(n3305) );
  AND U3724 ( .A(n3312), .B(p_input[7628]), .Z(n3311) );
  AND U3725 ( .A(p_input[6628]), .B(p_input[628]), .Z(n3312) );
  AND U3726 ( .A(p_input[9628]), .B(p_input[8628]), .Z(n3310) );
  AND U3727 ( .A(n3313), .B(n3314), .Z(o[627]) );
  AND U3728 ( .A(n3315), .B(n3316), .Z(n3314) );
  AND U3729 ( .A(n3317), .B(p_input[3627]), .Z(n3316) );
  AND U3730 ( .A(p_input[2627]), .B(p_input[1627]), .Z(n3317) );
  AND U3731 ( .A(p_input[5627]), .B(p_input[4627]), .Z(n3315) );
  AND U3732 ( .A(n3318), .B(n3319), .Z(n3313) );
  AND U3733 ( .A(n3320), .B(p_input[7627]), .Z(n3319) );
  AND U3734 ( .A(p_input[6627]), .B(p_input[627]), .Z(n3320) );
  AND U3735 ( .A(p_input[9627]), .B(p_input[8627]), .Z(n3318) );
  AND U3736 ( .A(n3321), .B(n3322), .Z(o[626]) );
  AND U3737 ( .A(n3323), .B(n3324), .Z(n3322) );
  AND U3738 ( .A(n3325), .B(p_input[3626]), .Z(n3324) );
  AND U3739 ( .A(p_input[2626]), .B(p_input[1626]), .Z(n3325) );
  AND U3740 ( .A(p_input[5626]), .B(p_input[4626]), .Z(n3323) );
  AND U3741 ( .A(n3326), .B(n3327), .Z(n3321) );
  AND U3742 ( .A(n3328), .B(p_input[7626]), .Z(n3327) );
  AND U3743 ( .A(p_input[6626]), .B(p_input[626]), .Z(n3328) );
  AND U3744 ( .A(p_input[9626]), .B(p_input[8626]), .Z(n3326) );
  AND U3745 ( .A(n3329), .B(n3330), .Z(o[625]) );
  AND U3746 ( .A(n3331), .B(n3332), .Z(n3330) );
  AND U3747 ( .A(n3333), .B(p_input[3625]), .Z(n3332) );
  AND U3748 ( .A(p_input[2625]), .B(p_input[1625]), .Z(n3333) );
  AND U3749 ( .A(p_input[5625]), .B(p_input[4625]), .Z(n3331) );
  AND U3750 ( .A(n3334), .B(n3335), .Z(n3329) );
  AND U3751 ( .A(n3336), .B(p_input[7625]), .Z(n3335) );
  AND U3752 ( .A(p_input[6625]), .B(p_input[625]), .Z(n3336) );
  AND U3753 ( .A(p_input[9625]), .B(p_input[8625]), .Z(n3334) );
  AND U3754 ( .A(n3337), .B(n3338), .Z(o[624]) );
  AND U3755 ( .A(n3339), .B(n3340), .Z(n3338) );
  AND U3756 ( .A(n3341), .B(p_input[3624]), .Z(n3340) );
  AND U3757 ( .A(p_input[2624]), .B(p_input[1624]), .Z(n3341) );
  AND U3758 ( .A(p_input[5624]), .B(p_input[4624]), .Z(n3339) );
  AND U3759 ( .A(n3342), .B(n3343), .Z(n3337) );
  AND U3760 ( .A(n3344), .B(p_input[7624]), .Z(n3343) );
  AND U3761 ( .A(p_input[6624]), .B(p_input[624]), .Z(n3344) );
  AND U3762 ( .A(p_input[9624]), .B(p_input[8624]), .Z(n3342) );
  AND U3763 ( .A(n3345), .B(n3346), .Z(o[623]) );
  AND U3764 ( .A(n3347), .B(n3348), .Z(n3346) );
  AND U3765 ( .A(n3349), .B(p_input[3623]), .Z(n3348) );
  AND U3766 ( .A(p_input[2623]), .B(p_input[1623]), .Z(n3349) );
  AND U3767 ( .A(p_input[5623]), .B(p_input[4623]), .Z(n3347) );
  AND U3768 ( .A(n3350), .B(n3351), .Z(n3345) );
  AND U3769 ( .A(n3352), .B(p_input[7623]), .Z(n3351) );
  AND U3770 ( .A(p_input[6623]), .B(p_input[623]), .Z(n3352) );
  AND U3771 ( .A(p_input[9623]), .B(p_input[8623]), .Z(n3350) );
  AND U3772 ( .A(n3353), .B(n3354), .Z(o[622]) );
  AND U3773 ( .A(n3355), .B(n3356), .Z(n3354) );
  AND U3774 ( .A(n3357), .B(p_input[3622]), .Z(n3356) );
  AND U3775 ( .A(p_input[2622]), .B(p_input[1622]), .Z(n3357) );
  AND U3776 ( .A(p_input[5622]), .B(p_input[4622]), .Z(n3355) );
  AND U3777 ( .A(n3358), .B(n3359), .Z(n3353) );
  AND U3778 ( .A(n3360), .B(p_input[7622]), .Z(n3359) );
  AND U3779 ( .A(p_input[6622]), .B(p_input[622]), .Z(n3360) );
  AND U3780 ( .A(p_input[9622]), .B(p_input[8622]), .Z(n3358) );
  AND U3781 ( .A(n3361), .B(n3362), .Z(o[621]) );
  AND U3782 ( .A(n3363), .B(n3364), .Z(n3362) );
  AND U3783 ( .A(n3365), .B(p_input[3621]), .Z(n3364) );
  AND U3784 ( .A(p_input[2621]), .B(p_input[1621]), .Z(n3365) );
  AND U3785 ( .A(p_input[5621]), .B(p_input[4621]), .Z(n3363) );
  AND U3786 ( .A(n3366), .B(n3367), .Z(n3361) );
  AND U3787 ( .A(n3368), .B(p_input[7621]), .Z(n3367) );
  AND U3788 ( .A(p_input[6621]), .B(p_input[621]), .Z(n3368) );
  AND U3789 ( .A(p_input[9621]), .B(p_input[8621]), .Z(n3366) );
  AND U3790 ( .A(n3369), .B(n3370), .Z(o[620]) );
  AND U3791 ( .A(n3371), .B(n3372), .Z(n3370) );
  AND U3792 ( .A(n3373), .B(p_input[3620]), .Z(n3372) );
  AND U3793 ( .A(p_input[2620]), .B(p_input[1620]), .Z(n3373) );
  AND U3794 ( .A(p_input[5620]), .B(p_input[4620]), .Z(n3371) );
  AND U3795 ( .A(n3374), .B(n3375), .Z(n3369) );
  AND U3796 ( .A(n3376), .B(p_input[7620]), .Z(n3375) );
  AND U3797 ( .A(p_input[6620]), .B(p_input[620]), .Z(n3376) );
  AND U3798 ( .A(p_input[9620]), .B(p_input[8620]), .Z(n3374) );
  AND U3799 ( .A(n3377), .B(n3378), .Z(o[61]) );
  AND U3800 ( .A(n3379), .B(n3380), .Z(n3378) );
  AND U3801 ( .A(n3381), .B(p_input[3061]), .Z(n3380) );
  AND U3802 ( .A(p_input[2061]), .B(p_input[1061]), .Z(n3381) );
  AND U3803 ( .A(p_input[5061]), .B(p_input[4061]), .Z(n3379) );
  AND U3804 ( .A(n3382), .B(n3383), .Z(n3377) );
  AND U3805 ( .A(n3384), .B(p_input[7061]), .Z(n3383) );
  AND U3806 ( .A(p_input[61]), .B(p_input[6061]), .Z(n3384) );
  AND U3807 ( .A(p_input[9061]), .B(p_input[8061]), .Z(n3382) );
  AND U3808 ( .A(n3385), .B(n3386), .Z(o[619]) );
  AND U3809 ( .A(n3387), .B(n3388), .Z(n3386) );
  AND U3810 ( .A(n3389), .B(p_input[3619]), .Z(n3388) );
  AND U3811 ( .A(p_input[2619]), .B(p_input[1619]), .Z(n3389) );
  AND U3812 ( .A(p_input[5619]), .B(p_input[4619]), .Z(n3387) );
  AND U3813 ( .A(n3390), .B(n3391), .Z(n3385) );
  AND U3814 ( .A(n3392), .B(p_input[7619]), .Z(n3391) );
  AND U3815 ( .A(p_input[6619]), .B(p_input[619]), .Z(n3392) );
  AND U3816 ( .A(p_input[9619]), .B(p_input[8619]), .Z(n3390) );
  AND U3817 ( .A(n3393), .B(n3394), .Z(o[618]) );
  AND U3818 ( .A(n3395), .B(n3396), .Z(n3394) );
  AND U3819 ( .A(n3397), .B(p_input[3618]), .Z(n3396) );
  AND U3820 ( .A(p_input[2618]), .B(p_input[1618]), .Z(n3397) );
  AND U3821 ( .A(p_input[5618]), .B(p_input[4618]), .Z(n3395) );
  AND U3822 ( .A(n3398), .B(n3399), .Z(n3393) );
  AND U3823 ( .A(n3400), .B(p_input[7618]), .Z(n3399) );
  AND U3824 ( .A(p_input[6618]), .B(p_input[618]), .Z(n3400) );
  AND U3825 ( .A(p_input[9618]), .B(p_input[8618]), .Z(n3398) );
  AND U3826 ( .A(n3401), .B(n3402), .Z(o[617]) );
  AND U3827 ( .A(n3403), .B(n3404), .Z(n3402) );
  AND U3828 ( .A(n3405), .B(p_input[3617]), .Z(n3404) );
  AND U3829 ( .A(p_input[2617]), .B(p_input[1617]), .Z(n3405) );
  AND U3830 ( .A(p_input[5617]), .B(p_input[4617]), .Z(n3403) );
  AND U3831 ( .A(n3406), .B(n3407), .Z(n3401) );
  AND U3832 ( .A(n3408), .B(p_input[7617]), .Z(n3407) );
  AND U3833 ( .A(p_input[6617]), .B(p_input[617]), .Z(n3408) );
  AND U3834 ( .A(p_input[9617]), .B(p_input[8617]), .Z(n3406) );
  AND U3835 ( .A(n3409), .B(n3410), .Z(o[616]) );
  AND U3836 ( .A(n3411), .B(n3412), .Z(n3410) );
  AND U3837 ( .A(n3413), .B(p_input[3616]), .Z(n3412) );
  AND U3838 ( .A(p_input[2616]), .B(p_input[1616]), .Z(n3413) );
  AND U3839 ( .A(p_input[5616]), .B(p_input[4616]), .Z(n3411) );
  AND U3840 ( .A(n3414), .B(n3415), .Z(n3409) );
  AND U3841 ( .A(n3416), .B(p_input[7616]), .Z(n3415) );
  AND U3842 ( .A(p_input[6616]), .B(p_input[616]), .Z(n3416) );
  AND U3843 ( .A(p_input[9616]), .B(p_input[8616]), .Z(n3414) );
  AND U3844 ( .A(n3417), .B(n3418), .Z(o[615]) );
  AND U3845 ( .A(n3419), .B(n3420), .Z(n3418) );
  AND U3846 ( .A(n3421), .B(p_input[3615]), .Z(n3420) );
  AND U3847 ( .A(p_input[2615]), .B(p_input[1615]), .Z(n3421) );
  AND U3848 ( .A(p_input[5615]), .B(p_input[4615]), .Z(n3419) );
  AND U3849 ( .A(n3422), .B(n3423), .Z(n3417) );
  AND U3850 ( .A(n3424), .B(p_input[7615]), .Z(n3423) );
  AND U3851 ( .A(p_input[6615]), .B(p_input[615]), .Z(n3424) );
  AND U3852 ( .A(p_input[9615]), .B(p_input[8615]), .Z(n3422) );
  AND U3853 ( .A(n3425), .B(n3426), .Z(o[614]) );
  AND U3854 ( .A(n3427), .B(n3428), .Z(n3426) );
  AND U3855 ( .A(n3429), .B(p_input[3614]), .Z(n3428) );
  AND U3856 ( .A(p_input[2614]), .B(p_input[1614]), .Z(n3429) );
  AND U3857 ( .A(p_input[5614]), .B(p_input[4614]), .Z(n3427) );
  AND U3858 ( .A(n3430), .B(n3431), .Z(n3425) );
  AND U3859 ( .A(n3432), .B(p_input[7614]), .Z(n3431) );
  AND U3860 ( .A(p_input[6614]), .B(p_input[614]), .Z(n3432) );
  AND U3861 ( .A(p_input[9614]), .B(p_input[8614]), .Z(n3430) );
  AND U3862 ( .A(n3433), .B(n3434), .Z(o[613]) );
  AND U3863 ( .A(n3435), .B(n3436), .Z(n3434) );
  AND U3864 ( .A(n3437), .B(p_input[3613]), .Z(n3436) );
  AND U3865 ( .A(p_input[2613]), .B(p_input[1613]), .Z(n3437) );
  AND U3866 ( .A(p_input[5613]), .B(p_input[4613]), .Z(n3435) );
  AND U3867 ( .A(n3438), .B(n3439), .Z(n3433) );
  AND U3868 ( .A(n3440), .B(p_input[7613]), .Z(n3439) );
  AND U3869 ( .A(p_input[6613]), .B(p_input[613]), .Z(n3440) );
  AND U3870 ( .A(p_input[9613]), .B(p_input[8613]), .Z(n3438) );
  AND U3871 ( .A(n3441), .B(n3442), .Z(o[612]) );
  AND U3872 ( .A(n3443), .B(n3444), .Z(n3442) );
  AND U3873 ( .A(n3445), .B(p_input[3612]), .Z(n3444) );
  AND U3874 ( .A(p_input[2612]), .B(p_input[1612]), .Z(n3445) );
  AND U3875 ( .A(p_input[5612]), .B(p_input[4612]), .Z(n3443) );
  AND U3876 ( .A(n3446), .B(n3447), .Z(n3441) );
  AND U3877 ( .A(n3448), .B(p_input[7612]), .Z(n3447) );
  AND U3878 ( .A(p_input[6612]), .B(p_input[612]), .Z(n3448) );
  AND U3879 ( .A(p_input[9612]), .B(p_input[8612]), .Z(n3446) );
  AND U3880 ( .A(n3449), .B(n3450), .Z(o[611]) );
  AND U3881 ( .A(n3451), .B(n3452), .Z(n3450) );
  AND U3882 ( .A(n3453), .B(p_input[3611]), .Z(n3452) );
  AND U3883 ( .A(p_input[2611]), .B(p_input[1611]), .Z(n3453) );
  AND U3884 ( .A(p_input[5611]), .B(p_input[4611]), .Z(n3451) );
  AND U3885 ( .A(n3454), .B(n3455), .Z(n3449) );
  AND U3886 ( .A(n3456), .B(p_input[7611]), .Z(n3455) );
  AND U3887 ( .A(p_input[6611]), .B(p_input[611]), .Z(n3456) );
  AND U3888 ( .A(p_input[9611]), .B(p_input[8611]), .Z(n3454) );
  AND U3889 ( .A(n3457), .B(n3458), .Z(o[610]) );
  AND U3890 ( .A(n3459), .B(n3460), .Z(n3458) );
  AND U3891 ( .A(n3461), .B(p_input[3610]), .Z(n3460) );
  AND U3892 ( .A(p_input[2610]), .B(p_input[1610]), .Z(n3461) );
  AND U3893 ( .A(p_input[5610]), .B(p_input[4610]), .Z(n3459) );
  AND U3894 ( .A(n3462), .B(n3463), .Z(n3457) );
  AND U3895 ( .A(n3464), .B(p_input[7610]), .Z(n3463) );
  AND U3896 ( .A(p_input[6610]), .B(p_input[610]), .Z(n3464) );
  AND U3897 ( .A(p_input[9610]), .B(p_input[8610]), .Z(n3462) );
  AND U3898 ( .A(n3465), .B(n3466), .Z(o[60]) );
  AND U3899 ( .A(n3467), .B(n3468), .Z(n3466) );
  AND U3900 ( .A(n3469), .B(p_input[3060]), .Z(n3468) );
  AND U3901 ( .A(p_input[2060]), .B(p_input[1060]), .Z(n3469) );
  AND U3902 ( .A(p_input[5060]), .B(p_input[4060]), .Z(n3467) );
  AND U3903 ( .A(n3470), .B(n3471), .Z(n3465) );
  AND U3904 ( .A(n3472), .B(p_input[7060]), .Z(n3471) );
  AND U3905 ( .A(p_input[60]), .B(p_input[6060]), .Z(n3472) );
  AND U3906 ( .A(p_input[9060]), .B(p_input[8060]), .Z(n3470) );
  AND U3907 ( .A(n3473), .B(n3474), .Z(o[609]) );
  AND U3908 ( .A(n3475), .B(n3476), .Z(n3474) );
  AND U3909 ( .A(n3477), .B(p_input[3609]), .Z(n3476) );
  AND U3910 ( .A(p_input[2609]), .B(p_input[1609]), .Z(n3477) );
  AND U3911 ( .A(p_input[5609]), .B(p_input[4609]), .Z(n3475) );
  AND U3912 ( .A(n3478), .B(n3479), .Z(n3473) );
  AND U3913 ( .A(n3480), .B(p_input[7609]), .Z(n3479) );
  AND U3914 ( .A(p_input[6609]), .B(p_input[609]), .Z(n3480) );
  AND U3915 ( .A(p_input[9609]), .B(p_input[8609]), .Z(n3478) );
  AND U3916 ( .A(n3481), .B(n3482), .Z(o[608]) );
  AND U3917 ( .A(n3483), .B(n3484), .Z(n3482) );
  AND U3918 ( .A(n3485), .B(p_input[3608]), .Z(n3484) );
  AND U3919 ( .A(p_input[2608]), .B(p_input[1608]), .Z(n3485) );
  AND U3920 ( .A(p_input[5608]), .B(p_input[4608]), .Z(n3483) );
  AND U3921 ( .A(n3486), .B(n3487), .Z(n3481) );
  AND U3922 ( .A(n3488), .B(p_input[7608]), .Z(n3487) );
  AND U3923 ( .A(p_input[6608]), .B(p_input[608]), .Z(n3488) );
  AND U3924 ( .A(p_input[9608]), .B(p_input[8608]), .Z(n3486) );
  AND U3925 ( .A(n3489), .B(n3490), .Z(o[607]) );
  AND U3926 ( .A(n3491), .B(n3492), .Z(n3490) );
  AND U3927 ( .A(n3493), .B(p_input[3607]), .Z(n3492) );
  AND U3928 ( .A(p_input[2607]), .B(p_input[1607]), .Z(n3493) );
  AND U3929 ( .A(p_input[5607]), .B(p_input[4607]), .Z(n3491) );
  AND U3930 ( .A(n3494), .B(n3495), .Z(n3489) );
  AND U3931 ( .A(n3496), .B(p_input[7607]), .Z(n3495) );
  AND U3932 ( .A(p_input[6607]), .B(p_input[607]), .Z(n3496) );
  AND U3933 ( .A(p_input[9607]), .B(p_input[8607]), .Z(n3494) );
  AND U3934 ( .A(n3497), .B(n3498), .Z(o[606]) );
  AND U3935 ( .A(n3499), .B(n3500), .Z(n3498) );
  AND U3936 ( .A(n3501), .B(p_input[3606]), .Z(n3500) );
  AND U3937 ( .A(p_input[2606]), .B(p_input[1606]), .Z(n3501) );
  AND U3938 ( .A(p_input[5606]), .B(p_input[4606]), .Z(n3499) );
  AND U3939 ( .A(n3502), .B(n3503), .Z(n3497) );
  AND U3940 ( .A(n3504), .B(p_input[7606]), .Z(n3503) );
  AND U3941 ( .A(p_input[6606]), .B(p_input[606]), .Z(n3504) );
  AND U3942 ( .A(p_input[9606]), .B(p_input[8606]), .Z(n3502) );
  AND U3943 ( .A(n3505), .B(n3506), .Z(o[605]) );
  AND U3944 ( .A(n3507), .B(n3508), .Z(n3506) );
  AND U3945 ( .A(n3509), .B(p_input[3605]), .Z(n3508) );
  AND U3946 ( .A(p_input[2605]), .B(p_input[1605]), .Z(n3509) );
  AND U3947 ( .A(p_input[5605]), .B(p_input[4605]), .Z(n3507) );
  AND U3948 ( .A(n3510), .B(n3511), .Z(n3505) );
  AND U3949 ( .A(n3512), .B(p_input[7605]), .Z(n3511) );
  AND U3950 ( .A(p_input[6605]), .B(p_input[605]), .Z(n3512) );
  AND U3951 ( .A(p_input[9605]), .B(p_input[8605]), .Z(n3510) );
  AND U3952 ( .A(n3513), .B(n3514), .Z(o[604]) );
  AND U3953 ( .A(n3515), .B(n3516), .Z(n3514) );
  AND U3954 ( .A(n3517), .B(p_input[3604]), .Z(n3516) );
  AND U3955 ( .A(p_input[2604]), .B(p_input[1604]), .Z(n3517) );
  AND U3956 ( .A(p_input[5604]), .B(p_input[4604]), .Z(n3515) );
  AND U3957 ( .A(n3518), .B(n3519), .Z(n3513) );
  AND U3958 ( .A(n3520), .B(p_input[7604]), .Z(n3519) );
  AND U3959 ( .A(p_input[6604]), .B(p_input[604]), .Z(n3520) );
  AND U3960 ( .A(p_input[9604]), .B(p_input[8604]), .Z(n3518) );
  AND U3961 ( .A(n3521), .B(n3522), .Z(o[603]) );
  AND U3962 ( .A(n3523), .B(n3524), .Z(n3522) );
  AND U3963 ( .A(n3525), .B(p_input[3603]), .Z(n3524) );
  AND U3964 ( .A(p_input[2603]), .B(p_input[1603]), .Z(n3525) );
  AND U3965 ( .A(p_input[5603]), .B(p_input[4603]), .Z(n3523) );
  AND U3966 ( .A(n3526), .B(n3527), .Z(n3521) );
  AND U3967 ( .A(n3528), .B(p_input[7603]), .Z(n3527) );
  AND U3968 ( .A(p_input[6603]), .B(p_input[603]), .Z(n3528) );
  AND U3969 ( .A(p_input[9603]), .B(p_input[8603]), .Z(n3526) );
  AND U3970 ( .A(n3529), .B(n3530), .Z(o[602]) );
  AND U3971 ( .A(n3531), .B(n3532), .Z(n3530) );
  AND U3972 ( .A(n3533), .B(p_input[3602]), .Z(n3532) );
  AND U3973 ( .A(p_input[2602]), .B(p_input[1602]), .Z(n3533) );
  AND U3974 ( .A(p_input[5602]), .B(p_input[4602]), .Z(n3531) );
  AND U3975 ( .A(n3534), .B(n3535), .Z(n3529) );
  AND U3976 ( .A(n3536), .B(p_input[7602]), .Z(n3535) );
  AND U3977 ( .A(p_input[6602]), .B(p_input[602]), .Z(n3536) );
  AND U3978 ( .A(p_input[9602]), .B(p_input[8602]), .Z(n3534) );
  AND U3979 ( .A(n3537), .B(n3538), .Z(o[601]) );
  AND U3980 ( .A(n3539), .B(n3540), .Z(n3538) );
  AND U3981 ( .A(n3541), .B(p_input[3601]), .Z(n3540) );
  AND U3982 ( .A(p_input[2601]), .B(p_input[1601]), .Z(n3541) );
  AND U3983 ( .A(p_input[5601]), .B(p_input[4601]), .Z(n3539) );
  AND U3984 ( .A(n3542), .B(n3543), .Z(n3537) );
  AND U3985 ( .A(n3544), .B(p_input[7601]), .Z(n3543) );
  AND U3986 ( .A(p_input[6601]), .B(p_input[601]), .Z(n3544) );
  AND U3987 ( .A(p_input[9601]), .B(p_input[8601]), .Z(n3542) );
  AND U3988 ( .A(n3545), .B(n3546), .Z(o[600]) );
  AND U3989 ( .A(n3547), .B(n3548), .Z(n3546) );
  AND U3990 ( .A(n3549), .B(p_input[3600]), .Z(n3548) );
  AND U3991 ( .A(p_input[2600]), .B(p_input[1600]), .Z(n3549) );
  AND U3992 ( .A(p_input[5600]), .B(p_input[4600]), .Z(n3547) );
  AND U3993 ( .A(n3550), .B(n3551), .Z(n3545) );
  AND U3994 ( .A(n3552), .B(p_input[7600]), .Z(n3551) );
  AND U3995 ( .A(p_input[6600]), .B(p_input[600]), .Z(n3552) );
  AND U3996 ( .A(p_input[9600]), .B(p_input[8600]), .Z(n3550) );
  AND U3997 ( .A(n3553), .B(n3554), .Z(o[5]) );
  AND U3998 ( .A(n3555), .B(n3556), .Z(n3554) );
  AND U3999 ( .A(n3557), .B(p_input[3005]), .Z(n3556) );
  AND U4000 ( .A(p_input[2005]), .B(p_input[1005]), .Z(n3557) );
  AND U4001 ( .A(p_input[5005]), .B(p_input[4005]), .Z(n3555) );
  AND U4002 ( .A(n3558), .B(n3559), .Z(n3553) );
  AND U4003 ( .A(n3560), .B(p_input[7005]), .Z(n3559) );
  AND U4004 ( .A(p_input[6005]), .B(p_input[5]), .Z(n3560) );
  AND U4005 ( .A(p_input[9005]), .B(p_input[8005]), .Z(n3558) );
  AND U4006 ( .A(n3561), .B(n3562), .Z(o[59]) );
  AND U4007 ( .A(n3563), .B(n3564), .Z(n3562) );
  AND U4008 ( .A(n3565), .B(p_input[3059]), .Z(n3564) );
  AND U4009 ( .A(p_input[2059]), .B(p_input[1059]), .Z(n3565) );
  AND U4010 ( .A(p_input[5059]), .B(p_input[4059]), .Z(n3563) );
  AND U4011 ( .A(n3566), .B(n3567), .Z(n3561) );
  AND U4012 ( .A(n3568), .B(p_input[7059]), .Z(n3567) );
  AND U4013 ( .A(p_input[6059]), .B(p_input[59]), .Z(n3568) );
  AND U4014 ( .A(p_input[9059]), .B(p_input[8059]), .Z(n3566) );
  AND U4015 ( .A(n3569), .B(n3570), .Z(o[599]) );
  AND U4016 ( .A(n3571), .B(n3572), .Z(n3570) );
  AND U4017 ( .A(n3573), .B(p_input[3599]), .Z(n3572) );
  AND U4018 ( .A(p_input[2599]), .B(p_input[1599]), .Z(n3573) );
  AND U4019 ( .A(p_input[5599]), .B(p_input[4599]), .Z(n3571) );
  AND U4020 ( .A(n3574), .B(n3575), .Z(n3569) );
  AND U4021 ( .A(n3576), .B(p_input[7599]), .Z(n3575) );
  AND U4022 ( .A(p_input[6599]), .B(p_input[599]), .Z(n3576) );
  AND U4023 ( .A(p_input[9599]), .B(p_input[8599]), .Z(n3574) );
  AND U4024 ( .A(n3577), .B(n3578), .Z(o[598]) );
  AND U4025 ( .A(n3579), .B(n3580), .Z(n3578) );
  AND U4026 ( .A(n3581), .B(p_input[3598]), .Z(n3580) );
  AND U4027 ( .A(p_input[2598]), .B(p_input[1598]), .Z(n3581) );
  AND U4028 ( .A(p_input[5598]), .B(p_input[4598]), .Z(n3579) );
  AND U4029 ( .A(n3582), .B(n3583), .Z(n3577) );
  AND U4030 ( .A(n3584), .B(p_input[7598]), .Z(n3583) );
  AND U4031 ( .A(p_input[6598]), .B(p_input[598]), .Z(n3584) );
  AND U4032 ( .A(p_input[9598]), .B(p_input[8598]), .Z(n3582) );
  AND U4033 ( .A(n3585), .B(n3586), .Z(o[597]) );
  AND U4034 ( .A(n3587), .B(n3588), .Z(n3586) );
  AND U4035 ( .A(n3589), .B(p_input[3597]), .Z(n3588) );
  AND U4036 ( .A(p_input[2597]), .B(p_input[1597]), .Z(n3589) );
  AND U4037 ( .A(p_input[5597]), .B(p_input[4597]), .Z(n3587) );
  AND U4038 ( .A(n3590), .B(n3591), .Z(n3585) );
  AND U4039 ( .A(n3592), .B(p_input[7597]), .Z(n3591) );
  AND U4040 ( .A(p_input[6597]), .B(p_input[597]), .Z(n3592) );
  AND U4041 ( .A(p_input[9597]), .B(p_input[8597]), .Z(n3590) );
  AND U4042 ( .A(n3593), .B(n3594), .Z(o[596]) );
  AND U4043 ( .A(n3595), .B(n3596), .Z(n3594) );
  AND U4044 ( .A(n3597), .B(p_input[3596]), .Z(n3596) );
  AND U4045 ( .A(p_input[2596]), .B(p_input[1596]), .Z(n3597) );
  AND U4046 ( .A(p_input[5596]), .B(p_input[4596]), .Z(n3595) );
  AND U4047 ( .A(n3598), .B(n3599), .Z(n3593) );
  AND U4048 ( .A(n3600), .B(p_input[7596]), .Z(n3599) );
  AND U4049 ( .A(p_input[6596]), .B(p_input[596]), .Z(n3600) );
  AND U4050 ( .A(p_input[9596]), .B(p_input[8596]), .Z(n3598) );
  AND U4051 ( .A(n3601), .B(n3602), .Z(o[595]) );
  AND U4052 ( .A(n3603), .B(n3604), .Z(n3602) );
  AND U4053 ( .A(n3605), .B(p_input[3595]), .Z(n3604) );
  AND U4054 ( .A(p_input[2595]), .B(p_input[1595]), .Z(n3605) );
  AND U4055 ( .A(p_input[5595]), .B(p_input[4595]), .Z(n3603) );
  AND U4056 ( .A(n3606), .B(n3607), .Z(n3601) );
  AND U4057 ( .A(n3608), .B(p_input[7595]), .Z(n3607) );
  AND U4058 ( .A(p_input[6595]), .B(p_input[595]), .Z(n3608) );
  AND U4059 ( .A(p_input[9595]), .B(p_input[8595]), .Z(n3606) );
  AND U4060 ( .A(n3609), .B(n3610), .Z(o[594]) );
  AND U4061 ( .A(n3611), .B(n3612), .Z(n3610) );
  AND U4062 ( .A(n3613), .B(p_input[3594]), .Z(n3612) );
  AND U4063 ( .A(p_input[2594]), .B(p_input[1594]), .Z(n3613) );
  AND U4064 ( .A(p_input[5594]), .B(p_input[4594]), .Z(n3611) );
  AND U4065 ( .A(n3614), .B(n3615), .Z(n3609) );
  AND U4066 ( .A(n3616), .B(p_input[7594]), .Z(n3615) );
  AND U4067 ( .A(p_input[6594]), .B(p_input[594]), .Z(n3616) );
  AND U4068 ( .A(p_input[9594]), .B(p_input[8594]), .Z(n3614) );
  AND U4069 ( .A(n3617), .B(n3618), .Z(o[593]) );
  AND U4070 ( .A(n3619), .B(n3620), .Z(n3618) );
  AND U4071 ( .A(n3621), .B(p_input[3593]), .Z(n3620) );
  AND U4072 ( .A(p_input[2593]), .B(p_input[1593]), .Z(n3621) );
  AND U4073 ( .A(p_input[5593]), .B(p_input[4593]), .Z(n3619) );
  AND U4074 ( .A(n3622), .B(n3623), .Z(n3617) );
  AND U4075 ( .A(n3624), .B(p_input[7593]), .Z(n3623) );
  AND U4076 ( .A(p_input[6593]), .B(p_input[593]), .Z(n3624) );
  AND U4077 ( .A(p_input[9593]), .B(p_input[8593]), .Z(n3622) );
  AND U4078 ( .A(n3625), .B(n3626), .Z(o[592]) );
  AND U4079 ( .A(n3627), .B(n3628), .Z(n3626) );
  AND U4080 ( .A(n3629), .B(p_input[3592]), .Z(n3628) );
  AND U4081 ( .A(p_input[2592]), .B(p_input[1592]), .Z(n3629) );
  AND U4082 ( .A(p_input[5592]), .B(p_input[4592]), .Z(n3627) );
  AND U4083 ( .A(n3630), .B(n3631), .Z(n3625) );
  AND U4084 ( .A(n3632), .B(p_input[7592]), .Z(n3631) );
  AND U4085 ( .A(p_input[6592]), .B(p_input[592]), .Z(n3632) );
  AND U4086 ( .A(p_input[9592]), .B(p_input[8592]), .Z(n3630) );
  AND U4087 ( .A(n3633), .B(n3634), .Z(o[591]) );
  AND U4088 ( .A(n3635), .B(n3636), .Z(n3634) );
  AND U4089 ( .A(n3637), .B(p_input[3591]), .Z(n3636) );
  AND U4090 ( .A(p_input[2591]), .B(p_input[1591]), .Z(n3637) );
  AND U4091 ( .A(p_input[5591]), .B(p_input[4591]), .Z(n3635) );
  AND U4092 ( .A(n3638), .B(n3639), .Z(n3633) );
  AND U4093 ( .A(n3640), .B(p_input[7591]), .Z(n3639) );
  AND U4094 ( .A(p_input[6591]), .B(p_input[591]), .Z(n3640) );
  AND U4095 ( .A(p_input[9591]), .B(p_input[8591]), .Z(n3638) );
  AND U4096 ( .A(n3641), .B(n3642), .Z(o[590]) );
  AND U4097 ( .A(n3643), .B(n3644), .Z(n3642) );
  AND U4098 ( .A(n3645), .B(p_input[3590]), .Z(n3644) );
  AND U4099 ( .A(p_input[2590]), .B(p_input[1590]), .Z(n3645) );
  AND U4100 ( .A(p_input[5590]), .B(p_input[4590]), .Z(n3643) );
  AND U4101 ( .A(n3646), .B(n3647), .Z(n3641) );
  AND U4102 ( .A(n3648), .B(p_input[7590]), .Z(n3647) );
  AND U4103 ( .A(p_input[6590]), .B(p_input[590]), .Z(n3648) );
  AND U4104 ( .A(p_input[9590]), .B(p_input[8590]), .Z(n3646) );
  AND U4105 ( .A(n3649), .B(n3650), .Z(o[58]) );
  AND U4106 ( .A(n3651), .B(n3652), .Z(n3650) );
  AND U4107 ( .A(n3653), .B(p_input[3058]), .Z(n3652) );
  AND U4108 ( .A(p_input[2058]), .B(p_input[1058]), .Z(n3653) );
  AND U4109 ( .A(p_input[5058]), .B(p_input[4058]), .Z(n3651) );
  AND U4110 ( .A(n3654), .B(n3655), .Z(n3649) );
  AND U4111 ( .A(n3656), .B(p_input[7058]), .Z(n3655) );
  AND U4112 ( .A(p_input[6058]), .B(p_input[58]), .Z(n3656) );
  AND U4113 ( .A(p_input[9058]), .B(p_input[8058]), .Z(n3654) );
  AND U4114 ( .A(n3657), .B(n3658), .Z(o[589]) );
  AND U4115 ( .A(n3659), .B(n3660), .Z(n3658) );
  AND U4116 ( .A(n3661), .B(p_input[3589]), .Z(n3660) );
  AND U4117 ( .A(p_input[2589]), .B(p_input[1589]), .Z(n3661) );
  AND U4118 ( .A(p_input[5589]), .B(p_input[4589]), .Z(n3659) );
  AND U4119 ( .A(n3662), .B(n3663), .Z(n3657) );
  AND U4120 ( .A(n3664), .B(p_input[7589]), .Z(n3663) );
  AND U4121 ( .A(p_input[6589]), .B(p_input[589]), .Z(n3664) );
  AND U4122 ( .A(p_input[9589]), .B(p_input[8589]), .Z(n3662) );
  AND U4123 ( .A(n3665), .B(n3666), .Z(o[588]) );
  AND U4124 ( .A(n3667), .B(n3668), .Z(n3666) );
  AND U4125 ( .A(n3669), .B(p_input[3588]), .Z(n3668) );
  AND U4126 ( .A(p_input[2588]), .B(p_input[1588]), .Z(n3669) );
  AND U4127 ( .A(p_input[5588]), .B(p_input[4588]), .Z(n3667) );
  AND U4128 ( .A(n3670), .B(n3671), .Z(n3665) );
  AND U4129 ( .A(n3672), .B(p_input[7588]), .Z(n3671) );
  AND U4130 ( .A(p_input[6588]), .B(p_input[588]), .Z(n3672) );
  AND U4131 ( .A(p_input[9588]), .B(p_input[8588]), .Z(n3670) );
  AND U4132 ( .A(n3673), .B(n3674), .Z(o[587]) );
  AND U4133 ( .A(n3675), .B(n3676), .Z(n3674) );
  AND U4134 ( .A(n3677), .B(p_input[3587]), .Z(n3676) );
  AND U4135 ( .A(p_input[2587]), .B(p_input[1587]), .Z(n3677) );
  AND U4136 ( .A(p_input[5587]), .B(p_input[4587]), .Z(n3675) );
  AND U4137 ( .A(n3678), .B(n3679), .Z(n3673) );
  AND U4138 ( .A(n3680), .B(p_input[7587]), .Z(n3679) );
  AND U4139 ( .A(p_input[6587]), .B(p_input[587]), .Z(n3680) );
  AND U4140 ( .A(p_input[9587]), .B(p_input[8587]), .Z(n3678) );
  AND U4141 ( .A(n3681), .B(n3682), .Z(o[586]) );
  AND U4142 ( .A(n3683), .B(n3684), .Z(n3682) );
  AND U4143 ( .A(n3685), .B(p_input[3586]), .Z(n3684) );
  AND U4144 ( .A(p_input[2586]), .B(p_input[1586]), .Z(n3685) );
  AND U4145 ( .A(p_input[5586]), .B(p_input[4586]), .Z(n3683) );
  AND U4146 ( .A(n3686), .B(n3687), .Z(n3681) );
  AND U4147 ( .A(n3688), .B(p_input[7586]), .Z(n3687) );
  AND U4148 ( .A(p_input[6586]), .B(p_input[586]), .Z(n3688) );
  AND U4149 ( .A(p_input[9586]), .B(p_input[8586]), .Z(n3686) );
  AND U4150 ( .A(n3689), .B(n3690), .Z(o[585]) );
  AND U4151 ( .A(n3691), .B(n3692), .Z(n3690) );
  AND U4152 ( .A(n3693), .B(p_input[3585]), .Z(n3692) );
  AND U4153 ( .A(p_input[2585]), .B(p_input[1585]), .Z(n3693) );
  AND U4154 ( .A(p_input[5585]), .B(p_input[4585]), .Z(n3691) );
  AND U4155 ( .A(n3694), .B(n3695), .Z(n3689) );
  AND U4156 ( .A(n3696), .B(p_input[7585]), .Z(n3695) );
  AND U4157 ( .A(p_input[6585]), .B(p_input[585]), .Z(n3696) );
  AND U4158 ( .A(p_input[9585]), .B(p_input[8585]), .Z(n3694) );
  AND U4159 ( .A(n3697), .B(n3698), .Z(o[584]) );
  AND U4160 ( .A(n3699), .B(n3700), .Z(n3698) );
  AND U4161 ( .A(n3701), .B(p_input[3584]), .Z(n3700) );
  AND U4162 ( .A(p_input[2584]), .B(p_input[1584]), .Z(n3701) );
  AND U4163 ( .A(p_input[5584]), .B(p_input[4584]), .Z(n3699) );
  AND U4164 ( .A(n3702), .B(n3703), .Z(n3697) );
  AND U4165 ( .A(n3704), .B(p_input[7584]), .Z(n3703) );
  AND U4166 ( .A(p_input[6584]), .B(p_input[584]), .Z(n3704) );
  AND U4167 ( .A(p_input[9584]), .B(p_input[8584]), .Z(n3702) );
  AND U4168 ( .A(n3705), .B(n3706), .Z(o[583]) );
  AND U4169 ( .A(n3707), .B(n3708), .Z(n3706) );
  AND U4170 ( .A(n3709), .B(p_input[3583]), .Z(n3708) );
  AND U4171 ( .A(p_input[2583]), .B(p_input[1583]), .Z(n3709) );
  AND U4172 ( .A(p_input[5583]), .B(p_input[4583]), .Z(n3707) );
  AND U4173 ( .A(n3710), .B(n3711), .Z(n3705) );
  AND U4174 ( .A(n3712), .B(p_input[7583]), .Z(n3711) );
  AND U4175 ( .A(p_input[6583]), .B(p_input[583]), .Z(n3712) );
  AND U4176 ( .A(p_input[9583]), .B(p_input[8583]), .Z(n3710) );
  AND U4177 ( .A(n3713), .B(n3714), .Z(o[582]) );
  AND U4178 ( .A(n3715), .B(n3716), .Z(n3714) );
  AND U4179 ( .A(n3717), .B(p_input[3582]), .Z(n3716) );
  AND U4180 ( .A(p_input[2582]), .B(p_input[1582]), .Z(n3717) );
  AND U4181 ( .A(p_input[5582]), .B(p_input[4582]), .Z(n3715) );
  AND U4182 ( .A(n3718), .B(n3719), .Z(n3713) );
  AND U4183 ( .A(n3720), .B(p_input[7582]), .Z(n3719) );
  AND U4184 ( .A(p_input[6582]), .B(p_input[582]), .Z(n3720) );
  AND U4185 ( .A(p_input[9582]), .B(p_input[8582]), .Z(n3718) );
  AND U4186 ( .A(n3721), .B(n3722), .Z(o[581]) );
  AND U4187 ( .A(n3723), .B(n3724), .Z(n3722) );
  AND U4188 ( .A(n3725), .B(p_input[3581]), .Z(n3724) );
  AND U4189 ( .A(p_input[2581]), .B(p_input[1581]), .Z(n3725) );
  AND U4190 ( .A(p_input[5581]), .B(p_input[4581]), .Z(n3723) );
  AND U4191 ( .A(n3726), .B(n3727), .Z(n3721) );
  AND U4192 ( .A(n3728), .B(p_input[7581]), .Z(n3727) );
  AND U4193 ( .A(p_input[6581]), .B(p_input[581]), .Z(n3728) );
  AND U4194 ( .A(p_input[9581]), .B(p_input[8581]), .Z(n3726) );
  AND U4195 ( .A(n3729), .B(n3730), .Z(o[580]) );
  AND U4196 ( .A(n3731), .B(n3732), .Z(n3730) );
  AND U4197 ( .A(n3733), .B(p_input[3580]), .Z(n3732) );
  AND U4198 ( .A(p_input[2580]), .B(p_input[1580]), .Z(n3733) );
  AND U4199 ( .A(p_input[5580]), .B(p_input[4580]), .Z(n3731) );
  AND U4200 ( .A(n3734), .B(n3735), .Z(n3729) );
  AND U4201 ( .A(n3736), .B(p_input[7580]), .Z(n3735) );
  AND U4202 ( .A(p_input[6580]), .B(p_input[580]), .Z(n3736) );
  AND U4203 ( .A(p_input[9580]), .B(p_input[8580]), .Z(n3734) );
  AND U4204 ( .A(n3737), .B(n3738), .Z(o[57]) );
  AND U4205 ( .A(n3739), .B(n3740), .Z(n3738) );
  AND U4206 ( .A(n3741), .B(p_input[3057]), .Z(n3740) );
  AND U4207 ( .A(p_input[2057]), .B(p_input[1057]), .Z(n3741) );
  AND U4208 ( .A(p_input[5057]), .B(p_input[4057]), .Z(n3739) );
  AND U4209 ( .A(n3742), .B(n3743), .Z(n3737) );
  AND U4210 ( .A(n3744), .B(p_input[7057]), .Z(n3743) );
  AND U4211 ( .A(p_input[6057]), .B(p_input[57]), .Z(n3744) );
  AND U4212 ( .A(p_input[9057]), .B(p_input[8057]), .Z(n3742) );
  AND U4213 ( .A(n3745), .B(n3746), .Z(o[579]) );
  AND U4214 ( .A(n3747), .B(n3748), .Z(n3746) );
  AND U4215 ( .A(n3749), .B(p_input[3579]), .Z(n3748) );
  AND U4216 ( .A(p_input[2579]), .B(p_input[1579]), .Z(n3749) );
  AND U4217 ( .A(p_input[5579]), .B(p_input[4579]), .Z(n3747) );
  AND U4218 ( .A(n3750), .B(n3751), .Z(n3745) );
  AND U4219 ( .A(n3752), .B(p_input[7579]), .Z(n3751) );
  AND U4220 ( .A(p_input[6579]), .B(p_input[579]), .Z(n3752) );
  AND U4221 ( .A(p_input[9579]), .B(p_input[8579]), .Z(n3750) );
  AND U4222 ( .A(n3753), .B(n3754), .Z(o[578]) );
  AND U4223 ( .A(n3755), .B(n3756), .Z(n3754) );
  AND U4224 ( .A(n3757), .B(p_input[3578]), .Z(n3756) );
  AND U4225 ( .A(p_input[2578]), .B(p_input[1578]), .Z(n3757) );
  AND U4226 ( .A(p_input[5578]), .B(p_input[4578]), .Z(n3755) );
  AND U4227 ( .A(n3758), .B(n3759), .Z(n3753) );
  AND U4228 ( .A(n3760), .B(p_input[7578]), .Z(n3759) );
  AND U4229 ( .A(p_input[6578]), .B(p_input[578]), .Z(n3760) );
  AND U4230 ( .A(p_input[9578]), .B(p_input[8578]), .Z(n3758) );
  AND U4231 ( .A(n3761), .B(n3762), .Z(o[577]) );
  AND U4232 ( .A(n3763), .B(n3764), .Z(n3762) );
  AND U4233 ( .A(n3765), .B(p_input[3577]), .Z(n3764) );
  AND U4234 ( .A(p_input[2577]), .B(p_input[1577]), .Z(n3765) );
  AND U4235 ( .A(p_input[5577]), .B(p_input[4577]), .Z(n3763) );
  AND U4236 ( .A(n3766), .B(n3767), .Z(n3761) );
  AND U4237 ( .A(n3768), .B(p_input[7577]), .Z(n3767) );
  AND U4238 ( .A(p_input[6577]), .B(p_input[577]), .Z(n3768) );
  AND U4239 ( .A(p_input[9577]), .B(p_input[8577]), .Z(n3766) );
  AND U4240 ( .A(n3769), .B(n3770), .Z(o[576]) );
  AND U4241 ( .A(n3771), .B(n3772), .Z(n3770) );
  AND U4242 ( .A(n3773), .B(p_input[3576]), .Z(n3772) );
  AND U4243 ( .A(p_input[2576]), .B(p_input[1576]), .Z(n3773) );
  AND U4244 ( .A(p_input[5576]), .B(p_input[4576]), .Z(n3771) );
  AND U4245 ( .A(n3774), .B(n3775), .Z(n3769) );
  AND U4246 ( .A(n3776), .B(p_input[7576]), .Z(n3775) );
  AND U4247 ( .A(p_input[6576]), .B(p_input[576]), .Z(n3776) );
  AND U4248 ( .A(p_input[9576]), .B(p_input[8576]), .Z(n3774) );
  AND U4249 ( .A(n3777), .B(n3778), .Z(o[575]) );
  AND U4250 ( .A(n3779), .B(n3780), .Z(n3778) );
  AND U4251 ( .A(n3781), .B(p_input[3575]), .Z(n3780) );
  AND U4252 ( .A(p_input[2575]), .B(p_input[1575]), .Z(n3781) );
  AND U4253 ( .A(p_input[5575]), .B(p_input[4575]), .Z(n3779) );
  AND U4254 ( .A(n3782), .B(n3783), .Z(n3777) );
  AND U4255 ( .A(n3784), .B(p_input[7575]), .Z(n3783) );
  AND U4256 ( .A(p_input[6575]), .B(p_input[575]), .Z(n3784) );
  AND U4257 ( .A(p_input[9575]), .B(p_input[8575]), .Z(n3782) );
  AND U4258 ( .A(n3785), .B(n3786), .Z(o[574]) );
  AND U4259 ( .A(n3787), .B(n3788), .Z(n3786) );
  AND U4260 ( .A(n3789), .B(p_input[3574]), .Z(n3788) );
  AND U4261 ( .A(p_input[2574]), .B(p_input[1574]), .Z(n3789) );
  AND U4262 ( .A(p_input[5574]), .B(p_input[4574]), .Z(n3787) );
  AND U4263 ( .A(n3790), .B(n3791), .Z(n3785) );
  AND U4264 ( .A(n3792), .B(p_input[7574]), .Z(n3791) );
  AND U4265 ( .A(p_input[6574]), .B(p_input[574]), .Z(n3792) );
  AND U4266 ( .A(p_input[9574]), .B(p_input[8574]), .Z(n3790) );
  AND U4267 ( .A(n3793), .B(n3794), .Z(o[573]) );
  AND U4268 ( .A(n3795), .B(n3796), .Z(n3794) );
  AND U4269 ( .A(n3797), .B(p_input[3573]), .Z(n3796) );
  AND U4270 ( .A(p_input[2573]), .B(p_input[1573]), .Z(n3797) );
  AND U4271 ( .A(p_input[5573]), .B(p_input[4573]), .Z(n3795) );
  AND U4272 ( .A(n3798), .B(n3799), .Z(n3793) );
  AND U4273 ( .A(n3800), .B(p_input[7573]), .Z(n3799) );
  AND U4274 ( .A(p_input[6573]), .B(p_input[573]), .Z(n3800) );
  AND U4275 ( .A(p_input[9573]), .B(p_input[8573]), .Z(n3798) );
  AND U4276 ( .A(n3801), .B(n3802), .Z(o[572]) );
  AND U4277 ( .A(n3803), .B(n3804), .Z(n3802) );
  AND U4278 ( .A(n3805), .B(p_input[3572]), .Z(n3804) );
  AND U4279 ( .A(p_input[2572]), .B(p_input[1572]), .Z(n3805) );
  AND U4280 ( .A(p_input[5572]), .B(p_input[4572]), .Z(n3803) );
  AND U4281 ( .A(n3806), .B(n3807), .Z(n3801) );
  AND U4282 ( .A(n3808), .B(p_input[7572]), .Z(n3807) );
  AND U4283 ( .A(p_input[6572]), .B(p_input[572]), .Z(n3808) );
  AND U4284 ( .A(p_input[9572]), .B(p_input[8572]), .Z(n3806) );
  AND U4285 ( .A(n3809), .B(n3810), .Z(o[571]) );
  AND U4286 ( .A(n3811), .B(n3812), .Z(n3810) );
  AND U4287 ( .A(n3813), .B(p_input[3571]), .Z(n3812) );
  AND U4288 ( .A(p_input[2571]), .B(p_input[1571]), .Z(n3813) );
  AND U4289 ( .A(p_input[5571]), .B(p_input[4571]), .Z(n3811) );
  AND U4290 ( .A(n3814), .B(n3815), .Z(n3809) );
  AND U4291 ( .A(n3816), .B(p_input[7571]), .Z(n3815) );
  AND U4292 ( .A(p_input[6571]), .B(p_input[571]), .Z(n3816) );
  AND U4293 ( .A(p_input[9571]), .B(p_input[8571]), .Z(n3814) );
  AND U4294 ( .A(n3817), .B(n3818), .Z(o[570]) );
  AND U4295 ( .A(n3819), .B(n3820), .Z(n3818) );
  AND U4296 ( .A(n3821), .B(p_input[3570]), .Z(n3820) );
  AND U4297 ( .A(p_input[2570]), .B(p_input[1570]), .Z(n3821) );
  AND U4298 ( .A(p_input[5570]), .B(p_input[4570]), .Z(n3819) );
  AND U4299 ( .A(n3822), .B(n3823), .Z(n3817) );
  AND U4300 ( .A(n3824), .B(p_input[7570]), .Z(n3823) );
  AND U4301 ( .A(p_input[6570]), .B(p_input[570]), .Z(n3824) );
  AND U4302 ( .A(p_input[9570]), .B(p_input[8570]), .Z(n3822) );
  AND U4303 ( .A(n3825), .B(n3826), .Z(o[56]) );
  AND U4304 ( .A(n3827), .B(n3828), .Z(n3826) );
  AND U4305 ( .A(n3829), .B(p_input[3056]), .Z(n3828) );
  AND U4306 ( .A(p_input[2056]), .B(p_input[1056]), .Z(n3829) );
  AND U4307 ( .A(p_input[5056]), .B(p_input[4056]), .Z(n3827) );
  AND U4308 ( .A(n3830), .B(n3831), .Z(n3825) );
  AND U4309 ( .A(n3832), .B(p_input[7056]), .Z(n3831) );
  AND U4310 ( .A(p_input[6056]), .B(p_input[56]), .Z(n3832) );
  AND U4311 ( .A(p_input[9056]), .B(p_input[8056]), .Z(n3830) );
  AND U4312 ( .A(n3833), .B(n3834), .Z(o[569]) );
  AND U4313 ( .A(n3835), .B(n3836), .Z(n3834) );
  AND U4314 ( .A(n3837), .B(p_input[3569]), .Z(n3836) );
  AND U4315 ( .A(p_input[2569]), .B(p_input[1569]), .Z(n3837) );
  AND U4316 ( .A(p_input[5569]), .B(p_input[4569]), .Z(n3835) );
  AND U4317 ( .A(n3838), .B(n3839), .Z(n3833) );
  AND U4318 ( .A(n3840), .B(p_input[7569]), .Z(n3839) );
  AND U4319 ( .A(p_input[6569]), .B(p_input[569]), .Z(n3840) );
  AND U4320 ( .A(p_input[9569]), .B(p_input[8569]), .Z(n3838) );
  AND U4321 ( .A(n3841), .B(n3842), .Z(o[568]) );
  AND U4322 ( .A(n3843), .B(n3844), .Z(n3842) );
  AND U4323 ( .A(n3845), .B(p_input[3568]), .Z(n3844) );
  AND U4324 ( .A(p_input[2568]), .B(p_input[1568]), .Z(n3845) );
  AND U4325 ( .A(p_input[5568]), .B(p_input[4568]), .Z(n3843) );
  AND U4326 ( .A(n3846), .B(n3847), .Z(n3841) );
  AND U4327 ( .A(n3848), .B(p_input[7568]), .Z(n3847) );
  AND U4328 ( .A(p_input[6568]), .B(p_input[568]), .Z(n3848) );
  AND U4329 ( .A(p_input[9568]), .B(p_input[8568]), .Z(n3846) );
  AND U4330 ( .A(n3849), .B(n3850), .Z(o[567]) );
  AND U4331 ( .A(n3851), .B(n3852), .Z(n3850) );
  AND U4332 ( .A(n3853), .B(p_input[3567]), .Z(n3852) );
  AND U4333 ( .A(p_input[2567]), .B(p_input[1567]), .Z(n3853) );
  AND U4334 ( .A(p_input[5567]), .B(p_input[4567]), .Z(n3851) );
  AND U4335 ( .A(n3854), .B(n3855), .Z(n3849) );
  AND U4336 ( .A(n3856), .B(p_input[7567]), .Z(n3855) );
  AND U4337 ( .A(p_input[6567]), .B(p_input[567]), .Z(n3856) );
  AND U4338 ( .A(p_input[9567]), .B(p_input[8567]), .Z(n3854) );
  AND U4339 ( .A(n3857), .B(n3858), .Z(o[566]) );
  AND U4340 ( .A(n3859), .B(n3860), .Z(n3858) );
  AND U4341 ( .A(n3861), .B(p_input[3566]), .Z(n3860) );
  AND U4342 ( .A(p_input[2566]), .B(p_input[1566]), .Z(n3861) );
  AND U4343 ( .A(p_input[5566]), .B(p_input[4566]), .Z(n3859) );
  AND U4344 ( .A(n3862), .B(n3863), .Z(n3857) );
  AND U4345 ( .A(n3864), .B(p_input[7566]), .Z(n3863) );
  AND U4346 ( .A(p_input[6566]), .B(p_input[566]), .Z(n3864) );
  AND U4347 ( .A(p_input[9566]), .B(p_input[8566]), .Z(n3862) );
  AND U4348 ( .A(n3865), .B(n3866), .Z(o[565]) );
  AND U4349 ( .A(n3867), .B(n3868), .Z(n3866) );
  AND U4350 ( .A(n3869), .B(p_input[3565]), .Z(n3868) );
  AND U4351 ( .A(p_input[2565]), .B(p_input[1565]), .Z(n3869) );
  AND U4352 ( .A(p_input[5565]), .B(p_input[4565]), .Z(n3867) );
  AND U4353 ( .A(n3870), .B(n3871), .Z(n3865) );
  AND U4354 ( .A(n3872), .B(p_input[7565]), .Z(n3871) );
  AND U4355 ( .A(p_input[6565]), .B(p_input[565]), .Z(n3872) );
  AND U4356 ( .A(p_input[9565]), .B(p_input[8565]), .Z(n3870) );
  AND U4357 ( .A(n3873), .B(n3874), .Z(o[564]) );
  AND U4358 ( .A(n3875), .B(n3876), .Z(n3874) );
  AND U4359 ( .A(n3877), .B(p_input[3564]), .Z(n3876) );
  AND U4360 ( .A(p_input[2564]), .B(p_input[1564]), .Z(n3877) );
  AND U4361 ( .A(p_input[5564]), .B(p_input[4564]), .Z(n3875) );
  AND U4362 ( .A(n3878), .B(n3879), .Z(n3873) );
  AND U4363 ( .A(n3880), .B(p_input[7564]), .Z(n3879) );
  AND U4364 ( .A(p_input[6564]), .B(p_input[564]), .Z(n3880) );
  AND U4365 ( .A(p_input[9564]), .B(p_input[8564]), .Z(n3878) );
  AND U4366 ( .A(n3881), .B(n3882), .Z(o[563]) );
  AND U4367 ( .A(n3883), .B(n3884), .Z(n3882) );
  AND U4368 ( .A(n3885), .B(p_input[3563]), .Z(n3884) );
  AND U4369 ( .A(p_input[2563]), .B(p_input[1563]), .Z(n3885) );
  AND U4370 ( .A(p_input[5563]), .B(p_input[4563]), .Z(n3883) );
  AND U4371 ( .A(n3886), .B(n3887), .Z(n3881) );
  AND U4372 ( .A(n3888), .B(p_input[7563]), .Z(n3887) );
  AND U4373 ( .A(p_input[6563]), .B(p_input[563]), .Z(n3888) );
  AND U4374 ( .A(p_input[9563]), .B(p_input[8563]), .Z(n3886) );
  AND U4375 ( .A(n3889), .B(n3890), .Z(o[562]) );
  AND U4376 ( .A(n3891), .B(n3892), .Z(n3890) );
  AND U4377 ( .A(n3893), .B(p_input[3562]), .Z(n3892) );
  AND U4378 ( .A(p_input[2562]), .B(p_input[1562]), .Z(n3893) );
  AND U4379 ( .A(p_input[5562]), .B(p_input[4562]), .Z(n3891) );
  AND U4380 ( .A(n3894), .B(n3895), .Z(n3889) );
  AND U4381 ( .A(n3896), .B(p_input[7562]), .Z(n3895) );
  AND U4382 ( .A(p_input[6562]), .B(p_input[562]), .Z(n3896) );
  AND U4383 ( .A(p_input[9562]), .B(p_input[8562]), .Z(n3894) );
  AND U4384 ( .A(n3897), .B(n3898), .Z(o[561]) );
  AND U4385 ( .A(n3899), .B(n3900), .Z(n3898) );
  AND U4386 ( .A(n3901), .B(p_input[3561]), .Z(n3900) );
  AND U4387 ( .A(p_input[2561]), .B(p_input[1561]), .Z(n3901) );
  AND U4388 ( .A(p_input[5561]), .B(p_input[4561]), .Z(n3899) );
  AND U4389 ( .A(n3902), .B(n3903), .Z(n3897) );
  AND U4390 ( .A(n3904), .B(p_input[7561]), .Z(n3903) );
  AND U4391 ( .A(p_input[6561]), .B(p_input[561]), .Z(n3904) );
  AND U4392 ( .A(p_input[9561]), .B(p_input[8561]), .Z(n3902) );
  AND U4393 ( .A(n3905), .B(n3906), .Z(o[560]) );
  AND U4394 ( .A(n3907), .B(n3908), .Z(n3906) );
  AND U4395 ( .A(n3909), .B(p_input[3560]), .Z(n3908) );
  AND U4396 ( .A(p_input[2560]), .B(p_input[1560]), .Z(n3909) );
  AND U4397 ( .A(p_input[5560]), .B(p_input[4560]), .Z(n3907) );
  AND U4398 ( .A(n3910), .B(n3911), .Z(n3905) );
  AND U4399 ( .A(n3912), .B(p_input[7560]), .Z(n3911) );
  AND U4400 ( .A(p_input[6560]), .B(p_input[560]), .Z(n3912) );
  AND U4401 ( .A(p_input[9560]), .B(p_input[8560]), .Z(n3910) );
  AND U4402 ( .A(n3913), .B(n3914), .Z(o[55]) );
  AND U4403 ( .A(n3915), .B(n3916), .Z(n3914) );
  AND U4404 ( .A(n3917), .B(p_input[3055]), .Z(n3916) );
  AND U4405 ( .A(p_input[2055]), .B(p_input[1055]), .Z(n3917) );
  AND U4406 ( .A(p_input[5055]), .B(p_input[4055]), .Z(n3915) );
  AND U4407 ( .A(n3918), .B(n3919), .Z(n3913) );
  AND U4408 ( .A(n3920), .B(p_input[7055]), .Z(n3919) );
  AND U4409 ( .A(p_input[6055]), .B(p_input[55]), .Z(n3920) );
  AND U4410 ( .A(p_input[9055]), .B(p_input[8055]), .Z(n3918) );
  AND U4411 ( .A(n3921), .B(n3922), .Z(o[559]) );
  AND U4412 ( .A(n3923), .B(n3924), .Z(n3922) );
  AND U4413 ( .A(n3925), .B(p_input[3559]), .Z(n3924) );
  AND U4414 ( .A(p_input[2559]), .B(p_input[1559]), .Z(n3925) );
  AND U4415 ( .A(p_input[5559]), .B(p_input[4559]), .Z(n3923) );
  AND U4416 ( .A(n3926), .B(n3927), .Z(n3921) );
  AND U4417 ( .A(n3928), .B(p_input[7559]), .Z(n3927) );
  AND U4418 ( .A(p_input[6559]), .B(p_input[559]), .Z(n3928) );
  AND U4419 ( .A(p_input[9559]), .B(p_input[8559]), .Z(n3926) );
  AND U4420 ( .A(n3929), .B(n3930), .Z(o[558]) );
  AND U4421 ( .A(n3931), .B(n3932), .Z(n3930) );
  AND U4422 ( .A(n3933), .B(p_input[3558]), .Z(n3932) );
  AND U4423 ( .A(p_input[2558]), .B(p_input[1558]), .Z(n3933) );
  AND U4424 ( .A(p_input[5558]), .B(p_input[4558]), .Z(n3931) );
  AND U4425 ( .A(n3934), .B(n3935), .Z(n3929) );
  AND U4426 ( .A(n3936), .B(p_input[7558]), .Z(n3935) );
  AND U4427 ( .A(p_input[6558]), .B(p_input[558]), .Z(n3936) );
  AND U4428 ( .A(p_input[9558]), .B(p_input[8558]), .Z(n3934) );
  AND U4429 ( .A(n3937), .B(n3938), .Z(o[557]) );
  AND U4430 ( .A(n3939), .B(n3940), .Z(n3938) );
  AND U4431 ( .A(n3941), .B(p_input[3557]), .Z(n3940) );
  AND U4432 ( .A(p_input[2557]), .B(p_input[1557]), .Z(n3941) );
  AND U4433 ( .A(p_input[5557]), .B(p_input[4557]), .Z(n3939) );
  AND U4434 ( .A(n3942), .B(n3943), .Z(n3937) );
  AND U4435 ( .A(n3944), .B(p_input[7557]), .Z(n3943) );
  AND U4436 ( .A(p_input[6557]), .B(p_input[557]), .Z(n3944) );
  AND U4437 ( .A(p_input[9557]), .B(p_input[8557]), .Z(n3942) );
  AND U4438 ( .A(n3945), .B(n3946), .Z(o[556]) );
  AND U4439 ( .A(n3947), .B(n3948), .Z(n3946) );
  AND U4440 ( .A(n3949), .B(p_input[3556]), .Z(n3948) );
  AND U4441 ( .A(p_input[2556]), .B(p_input[1556]), .Z(n3949) );
  AND U4442 ( .A(p_input[5556]), .B(p_input[4556]), .Z(n3947) );
  AND U4443 ( .A(n3950), .B(n3951), .Z(n3945) );
  AND U4444 ( .A(n3952), .B(p_input[7556]), .Z(n3951) );
  AND U4445 ( .A(p_input[6556]), .B(p_input[556]), .Z(n3952) );
  AND U4446 ( .A(p_input[9556]), .B(p_input[8556]), .Z(n3950) );
  AND U4447 ( .A(n3953), .B(n3954), .Z(o[555]) );
  AND U4448 ( .A(n3955), .B(n3956), .Z(n3954) );
  AND U4449 ( .A(n3957), .B(p_input[3555]), .Z(n3956) );
  AND U4450 ( .A(p_input[2555]), .B(p_input[1555]), .Z(n3957) );
  AND U4451 ( .A(p_input[5555]), .B(p_input[4555]), .Z(n3955) );
  AND U4452 ( .A(n3958), .B(n3959), .Z(n3953) );
  AND U4453 ( .A(n3960), .B(p_input[7555]), .Z(n3959) );
  AND U4454 ( .A(p_input[6555]), .B(p_input[555]), .Z(n3960) );
  AND U4455 ( .A(p_input[9555]), .B(p_input[8555]), .Z(n3958) );
  AND U4456 ( .A(n3961), .B(n3962), .Z(o[554]) );
  AND U4457 ( .A(n3963), .B(n3964), .Z(n3962) );
  AND U4458 ( .A(n3965), .B(p_input[3554]), .Z(n3964) );
  AND U4459 ( .A(p_input[2554]), .B(p_input[1554]), .Z(n3965) );
  AND U4460 ( .A(p_input[554]), .B(p_input[4554]), .Z(n3963) );
  AND U4461 ( .A(n3966), .B(n3967), .Z(n3961) );
  AND U4462 ( .A(n3968), .B(p_input[7554]), .Z(n3967) );
  AND U4463 ( .A(p_input[6554]), .B(p_input[5554]), .Z(n3968) );
  AND U4464 ( .A(p_input[9554]), .B(p_input[8554]), .Z(n3966) );
  AND U4465 ( .A(n3969), .B(n3970), .Z(o[553]) );
  AND U4466 ( .A(n3971), .B(n3972), .Z(n3970) );
  AND U4467 ( .A(n3973), .B(p_input[3553]), .Z(n3972) );
  AND U4468 ( .A(p_input[2553]), .B(p_input[1553]), .Z(n3973) );
  AND U4469 ( .A(p_input[553]), .B(p_input[4553]), .Z(n3971) );
  AND U4470 ( .A(n3974), .B(n3975), .Z(n3969) );
  AND U4471 ( .A(n3976), .B(p_input[7553]), .Z(n3975) );
  AND U4472 ( .A(p_input[6553]), .B(p_input[5553]), .Z(n3976) );
  AND U4473 ( .A(p_input[9553]), .B(p_input[8553]), .Z(n3974) );
  AND U4474 ( .A(n3977), .B(n3978), .Z(o[552]) );
  AND U4475 ( .A(n3979), .B(n3980), .Z(n3978) );
  AND U4476 ( .A(n3981), .B(p_input[3552]), .Z(n3980) );
  AND U4477 ( .A(p_input[2552]), .B(p_input[1552]), .Z(n3981) );
  AND U4478 ( .A(p_input[552]), .B(p_input[4552]), .Z(n3979) );
  AND U4479 ( .A(n3982), .B(n3983), .Z(n3977) );
  AND U4480 ( .A(n3984), .B(p_input[7552]), .Z(n3983) );
  AND U4481 ( .A(p_input[6552]), .B(p_input[5552]), .Z(n3984) );
  AND U4482 ( .A(p_input[9552]), .B(p_input[8552]), .Z(n3982) );
  AND U4483 ( .A(n3985), .B(n3986), .Z(o[551]) );
  AND U4484 ( .A(n3987), .B(n3988), .Z(n3986) );
  AND U4485 ( .A(n3989), .B(p_input[3551]), .Z(n3988) );
  AND U4486 ( .A(p_input[2551]), .B(p_input[1551]), .Z(n3989) );
  AND U4487 ( .A(p_input[551]), .B(p_input[4551]), .Z(n3987) );
  AND U4488 ( .A(n3990), .B(n3991), .Z(n3985) );
  AND U4489 ( .A(n3992), .B(p_input[7551]), .Z(n3991) );
  AND U4490 ( .A(p_input[6551]), .B(p_input[5551]), .Z(n3992) );
  AND U4491 ( .A(p_input[9551]), .B(p_input[8551]), .Z(n3990) );
  AND U4492 ( .A(n3993), .B(n3994), .Z(o[550]) );
  AND U4493 ( .A(n3995), .B(n3996), .Z(n3994) );
  AND U4494 ( .A(n3997), .B(p_input[3550]), .Z(n3996) );
  AND U4495 ( .A(p_input[2550]), .B(p_input[1550]), .Z(n3997) );
  AND U4496 ( .A(p_input[550]), .B(p_input[4550]), .Z(n3995) );
  AND U4497 ( .A(n3998), .B(n3999), .Z(n3993) );
  AND U4498 ( .A(n4000), .B(p_input[7550]), .Z(n3999) );
  AND U4499 ( .A(p_input[6550]), .B(p_input[5550]), .Z(n4000) );
  AND U4500 ( .A(p_input[9550]), .B(p_input[8550]), .Z(n3998) );
  AND U4501 ( .A(n4001), .B(n4002), .Z(o[54]) );
  AND U4502 ( .A(n4003), .B(n4004), .Z(n4002) );
  AND U4503 ( .A(n4005), .B(p_input[3054]), .Z(n4004) );
  AND U4504 ( .A(p_input[2054]), .B(p_input[1054]), .Z(n4005) );
  AND U4505 ( .A(p_input[5054]), .B(p_input[4054]), .Z(n4003) );
  AND U4506 ( .A(n4006), .B(n4007), .Z(n4001) );
  AND U4507 ( .A(n4008), .B(p_input[7054]), .Z(n4007) );
  AND U4508 ( .A(p_input[6054]), .B(p_input[54]), .Z(n4008) );
  AND U4509 ( .A(p_input[9054]), .B(p_input[8054]), .Z(n4006) );
  AND U4510 ( .A(n4009), .B(n4010), .Z(o[549]) );
  AND U4511 ( .A(n4011), .B(n4012), .Z(n4010) );
  AND U4512 ( .A(n4013), .B(p_input[3549]), .Z(n4012) );
  AND U4513 ( .A(p_input[2549]), .B(p_input[1549]), .Z(n4013) );
  AND U4514 ( .A(p_input[549]), .B(p_input[4549]), .Z(n4011) );
  AND U4515 ( .A(n4014), .B(n4015), .Z(n4009) );
  AND U4516 ( .A(n4016), .B(p_input[7549]), .Z(n4015) );
  AND U4517 ( .A(p_input[6549]), .B(p_input[5549]), .Z(n4016) );
  AND U4518 ( .A(p_input[9549]), .B(p_input[8549]), .Z(n4014) );
  AND U4519 ( .A(n4017), .B(n4018), .Z(o[548]) );
  AND U4520 ( .A(n4019), .B(n4020), .Z(n4018) );
  AND U4521 ( .A(n4021), .B(p_input[3548]), .Z(n4020) );
  AND U4522 ( .A(p_input[2548]), .B(p_input[1548]), .Z(n4021) );
  AND U4523 ( .A(p_input[548]), .B(p_input[4548]), .Z(n4019) );
  AND U4524 ( .A(n4022), .B(n4023), .Z(n4017) );
  AND U4525 ( .A(n4024), .B(p_input[7548]), .Z(n4023) );
  AND U4526 ( .A(p_input[6548]), .B(p_input[5548]), .Z(n4024) );
  AND U4527 ( .A(p_input[9548]), .B(p_input[8548]), .Z(n4022) );
  AND U4528 ( .A(n4025), .B(n4026), .Z(o[547]) );
  AND U4529 ( .A(n4027), .B(n4028), .Z(n4026) );
  AND U4530 ( .A(n4029), .B(p_input[3547]), .Z(n4028) );
  AND U4531 ( .A(p_input[2547]), .B(p_input[1547]), .Z(n4029) );
  AND U4532 ( .A(p_input[547]), .B(p_input[4547]), .Z(n4027) );
  AND U4533 ( .A(n4030), .B(n4031), .Z(n4025) );
  AND U4534 ( .A(n4032), .B(p_input[7547]), .Z(n4031) );
  AND U4535 ( .A(p_input[6547]), .B(p_input[5547]), .Z(n4032) );
  AND U4536 ( .A(p_input[9547]), .B(p_input[8547]), .Z(n4030) );
  AND U4537 ( .A(n4033), .B(n4034), .Z(o[546]) );
  AND U4538 ( .A(n4035), .B(n4036), .Z(n4034) );
  AND U4539 ( .A(n4037), .B(p_input[3546]), .Z(n4036) );
  AND U4540 ( .A(p_input[2546]), .B(p_input[1546]), .Z(n4037) );
  AND U4541 ( .A(p_input[546]), .B(p_input[4546]), .Z(n4035) );
  AND U4542 ( .A(n4038), .B(n4039), .Z(n4033) );
  AND U4543 ( .A(n4040), .B(p_input[7546]), .Z(n4039) );
  AND U4544 ( .A(p_input[6546]), .B(p_input[5546]), .Z(n4040) );
  AND U4545 ( .A(p_input[9546]), .B(p_input[8546]), .Z(n4038) );
  AND U4546 ( .A(n4041), .B(n4042), .Z(o[545]) );
  AND U4547 ( .A(n4043), .B(n4044), .Z(n4042) );
  AND U4548 ( .A(n4045), .B(p_input[3545]), .Z(n4044) );
  AND U4549 ( .A(p_input[2545]), .B(p_input[1545]), .Z(n4045) );
  AND U4550 ( .A(p_input[545]), .B(p_input[4545]), .Z(n4043) );
  AND U4551 ( .A(n4046), .B(n4047), .Z(n4041) );
  AND U4552 ( .A(n4048), .B(p_input[7545]), .Z(n4047) );
  AND U4553 ( .A(p_input[6545]), .B(p_input[5545]), .Z(n4048) );
  AND U4554 ( .A(p_input[9545]), .B(p_input[8545]), .Z(n4046) );
  AND U4555 ( .A(n4049), .B(n4050), .Z(o[544]) );
  AND U4556 ( .A(n4051), .B(n4052), .Z(n4050) );
  AND U4557 ( .A(n4053), .B(p_input[3544]), .Z(n4052) );
  AND U4558 ( .A(p_input[2544]), .B(p_input[1544]), .Z(n4053) );
  AND U4559 ( .A(p_input[544]), .B(p_input[4544]), .Z(n4051) );
  AND U4560 ( .A(n4054), .B(n4055), .Z(n4049) );
  AND U4561 ( .A(n4056), .B(p_input[7544]), .Z(n4055) );
  AND U4562 ( .A(p_input[6544]), .B(p_input[5544]), .Z(n4056) );
  AND U4563 ( .A(p_input[9544]), .B(p_input[8544]), .Z(n4054) );
  AND U4564 ( .A(n4057), .B(n4058), .Z(o[543]) );
  AND U4565 ( .A(n4059), .B(n4060), .Z(n4058) );
  AND U4566 ( .A(n4061), .B(p_input[3543]), .Z(n4060) );
  AND U4567 ( .A(p_input[2543]), .B(p_input[1543]), .Z(n4061) );
  AND U4568 ( .A(p_input[543]), .B(p_input[4543]), .Z(n4059) );
  AND U4569 ( .A(n4062), .B(n4063), .Z(n4057) );
  AND U4570 ( .A(n4064), .B(p_input[7543]), .Z(n4063) );
  AND U4571 ( .A(p_input[6543]), .B(p_input[5543]), .Z(n4064) );
  AND U4572 ( .A(p_input[9543]), .B(p_input[8543]), .Z(n4062) );
  AND U4573 ( .A(n4065), .B(n4066), .Z(o[542]) );
  AND U4574 ( .A(n4067), .B(n4068), .Z(n4066) );
  AND U4575 ( .A(n4069), .B(p_input[3542]), .Z(n4068) );
  AND U4576 ( .A(p_input[2542]), .B(p_input[1542]), .Z(n4069) );
  AND U4577 ( .A(p_input[542]), .B(p_input[4542]), .Z(n4067) );
  AND U4578 ( .A(n4070), .B(n4071), .Z(n4065) );
  AND U4579 ( .A(n4072), .B(p_input[7542]), .Z(n4071) );
  AND U4580 ( .A(p_input[6542]), .B(p_input[5542]), .Z(n4072) );
  AND U4581 ( .A(p_input[9542]), .B(p_input[8542]), .Z(n4070) );
  AND U4582 ( .A(n4073), .B(n4074), .Z(o[541]) );
  AND U4583 ( .A(n4075), .B(n4076), .Z(n4074) );
  AND U4584 ( .A(n4077), .B(p_input[3541]), .Z(n4076) );
  AND U4585 ( .A(p_input[2541]), .B(p_input[1541]), .Z(n4077) );
  AND U4586 ( .A(p_input[541]), .B(p_input[4541]), .Z(n4075) );
  AND U4587 ( .A(n4078), .B(n4079), .Z(n4073) );
  AND U4588 ( .A(n4080), .B(p_input[7541]), .Z(n4079) );
  AND U4589 ( .A(p_input[6541]), .B(p_input[5541]), .Z(n4080) );
  AND U4590 ( .A(p_input[9541]), .B(p_input[8541]), .Z(n4078) );
  AND U4591 ( .A(n4081), .B(n4082), .Z(o[540]) );
  AND U4592 ( .A(n4083), .B(n4084), .Z(n4082) );
  AND U4593 ( .A(n4085), .B(p_input[3540]), .Z(n4084) );
  AND U4594 ( .A(p_input[2540]), .B(p_input[1540]), .Z(n4085) );
  AND U4595 ( .A(p_input[540]), .B(p_input[4540]), .Z(n4083) );
  AND U4596 ( .A(n4086), .B(n4087), .Z(n4081) );
  AND U4597 ( .A(n4088), .B(p_input[7540]), .Z(n4087) );
  AND U4598 ( .A(p_input[6540]), .B(p_input[5540]), .Z(n4088) );
  AND U4599 ( .A(p_input[9540]), .B(p_input[8540]), .Z(n4086) );
  AND U4600 ( .A(n4089), .B(n4090), .Z(o[53]) );
  AND U4601 ( .A(n4091), .B(n4092), .Z(n4090) );
  AND U4602 ( .A(n4093), .B(p_input[3053]), .Z(n4092) );
  AND U4603 ( .A(p_input[2053]), .B(p_input[1053]), .Z(n4093) );
  AND U4604 ( .A(p_input[5053]), .B(p_input[4053]), .Z(n4091) );
  AND U4605 ( .A(n4094), .B(n4095), .Z(n4089) );
  AND U4606 ( .A(n4096), .B(p_input[7053]), .Z(n4095) );
  AND U4607 ( .A(p_input[6053]), .B(p_input[53]), .Z(n4096) );
  AND U4608 ( .A(p_input[9053]), .B(p_input[8053]), .Z(n4094) );
  AND U4609 ( .A(n4097), .B(n4098), .Z(o[539]) );
  AND U4610 ( .A(n4099), .B(n4100), .Z(n4098) );
  AND U4611 ( .A(n4101), .B(p_input[3539]), .Z(n4100) );
  AND U4612 ( .A(p_input[2539]), .B(p_input[1539]), .Z(n4101) );
  AND U4613 ( .A(p_input[539]), .B(p_input[4539]), .Z(n4099) );
  AND U4614 ( .A(n4102), .B(n4103), .Z(n4097) );
  AND U4615 ( .A(n4104), .B(p_input[7539]), .Z(n4103) );
  AND U4616 ( .A(p_input[6539]), .B(p_input[5539]), .Z(n4104) );
  AND U4617 ( .A(p_input[9539]), .B(p_input[8539]), .Z(n4102) );
  AND U4618 ( .A(n4105), .B(n4106), .Z(o[538]) );
  AND U4619 ( .A(n4107), .B(n4108), .Z(n4106) );
  AND U4620 ( .A(n4109), .B(p_input[3538]), .Z(n4108) );
  AND U4621 ( .A(p_input[2538]), .B(p_input[1538]), .Z(n4109) );
  AND U4622 ( .A(p_input[538]), .B(p_input[4538]), .Z(n4107) );
  AND U4623 ( .A(n4110), .B(n4111), .Z(n4105) );
  AND U4624 ( .A(n4112), .B(p_input[7538]), .Z(n4111) );
  AND U4625 ( .A(p_input[6538]), .B(p_input[5538]), .Z(n4112) );
  AND U4626 ( .A(p_input[9538]), .B(p_input[8538]), .Z(n4110) );
  AND U4627 ( .A(n4113), .B(n4114), .Z(o[537]) );
  AND U4628 ( .A(n4115), .B(n4116), .Z(n4114) );
  AND U4629 ( .A(n4117), .B(p_input[3537]), .Z(n4116) );
  AND U4630 ( .A(p_input[2537]), .B(p_input[1537]), .Z(n4117) );
  AND U4631 ( .A(p_input[537]), .B(p_input[4537]), .Z(n4115) );
  AND U4632 ( .A(n4118), .B(n4119), .Z(n4113) );
  AND U4633 ( .A(n4120), .B(p_input[7537]), .Z(n4119) );
  AND U4634 ( .A(p_input[6537]), .B(p_input[5537]), .Z(n4120) );
  AND U4635 ( .A(p_input[9537]), .B(p_input[8537]), .Z(n4118) );
  AND U4636 ( .A(n4121), .B(n4122), .Z(o[536]) );
  AND U4637 ( .A(n4123), .B(n4124), .Z(n4122) );
  AND U4638 ( .A(n4125), .B(p_input[3536]), .Z(n4124) );
  AND U4639 ( .A(p_input[2536]), .B(p_input[1536]), .Z(n4125) );
  AND U4640 ( .A(p_input[536]), .B(p_input[4536]), .Z(n4123) );
  AND U4641 ( .A(n4126), .B(n4127), .Z(n4121) );
  AND U4642 ( .A(n4128), .B(p_input[7536]), .Z(n4127) );
  AND U4643 ( .A(p_input[6536]), .B(p_input[5536]), .Z(n4128) );
  AND U4644 ( .A(p_input[9536]), .B(p_input[8536]), .Z(n4126) );
  AND U4645 ( .A(n4129), .B(n4130), .Z(o[535]) );
  AND U4646 ( .A(n4131), .B(n4132), .Z(n4130) );
  AND U4647 ( .A(n4133), .B(p_input[3535]), .Z(n4132) );
  AND U4648 ( .A(p_input[2535]), .B(p_input[1535]), .Z(n4133) );
  AND U4649 ( .A(p_input[535]), .B(p_input[4535]), .Z(n4131) );
  AND U4650 ( .A(n4134), .B(n4135), .Z(n4129) );
  AND U4651 ( .A(n4136), .B(p_input[7535]), .Z(n4135) );
  AND U4652 ( .A(p_input[6535]), .B(p_input[5535]), .Z(n4136) );
  AND U4653 ( .A(p_input[9535]), .B(p_input[8535]), .Z(n4134) );
  AND U4654 ( .A(n4137), .B(n4138), .Z(o[534]) );
  AND U4655 ( .A(n4139), .B(n4140), .Z(n4138) );
  AND U4656 ( .A(n4141), .B(p_input[3534]), .Z(n4140) );
  AND U4657 ( .A(p_input[2534]), .B(p_input[1534]), .Z(n4141) );
  AND U4658 ( .A(p_input[534]), .B(p_input[4534]), .Z(n4139) );
  AND U4659 ( .A(n4142), .B(n4143), .Z(n4137) );
  AND U4660 ( .A(n4144), .B(p_input[7534]), .Z(n4143) );
  AND U4661 ( .A(p_input[6534]), .B(p_input[5534]), .Z(n4144) );
  AND U4662 ( .A(p_input[9534]), .B(p_input[8534]), .Z(n4142) );
  AND U4663 ( .A(n4145), .B(n4146), .Z(o[533]) );
  AND U4664 ( .A(n4147), .B(n4148), .Z(n4146) );
  AND U4665 ( .A(n4149), .B(p_input[3533]), .Z(n4148) );
  AND U4666 ( .A(p_input[2533]), .B(p_input[1533]), .Z(n4149) );
  AND U4667 ( .A(p_input[533]), .B(p_input[4533]), .Z(n4147) );
  AND U4668 ( .A(n4150), .B(n4151), .Z(n4145) );
  AND U4669 ( .A(n4152), .B(p_input[7533]), .Z(n4151) );
  AND U4670 ( .A(p_input[6533]), .B(p_input[5533]), .Z(n4152) );
  AND U4671 ( .A(p_input[9533]), .B(p_input[8533]), .Z(n4150) );
  AND U4672 ( .A(n4153), .B(n4154), .Z(o[532]) );
  AND U4673 ( .A(n4155), .B(n4156), .Z(n4154) );
  AND U4674 ( .A(n4157), .B(p_input[3532]), .Z(n4156) );
  AND U4675 ( .A(p_input[2532]), .B(p_input[1532]), .Z(n4157) );
  AND U4676 ( .A(p_input[532]), .B(p_input[4532]), .Z(n4155) );
  AND U4677 ( .A(n4158), .B(n4159), .Z(n4153) );
  AND U4678 ( .A(n4160), .B(p_input[7532]), .Z(n4159) );
  AND U4679 ( .A(p_input[6532]), .B(p_input[5532]), .Z(n4160) );
  AND U4680 ( .A(p_input[9532]), .B(p_input[8532]), .Z(n4158) );
  AND U4681 ( .A(n4161), .B(n4162), .Z(o[531]) );
  AND U4682 ( .A(n4163), .B(n4164), .Z(n4162) );
  AND U4683 ( .A(n4165), .B(p_input[3531]), .Z(n4164) );
  AND U4684 ( .A(p_input[2531]), .B(p_input[1531]), .Z(n4165) );
  AND U4685 ( .A(p_input[531]), .B(p_input[4531]), .Z(n4163) );
  AND U4686 ( .A(n4166), .B(n4167), .Z(n4161) );
  AND U4687 ( .A(n4168), .B(p_input[7531]), .Z(n4167) );
  AND U4688 ( .A(p_input[6531]), .B(p_input[5531]), .Z(n4168) );
  AND U4689 ( .A(p_input[9531]), .B(p_input[8531]), .Z(n4166) );
  AND U4690 ( .A(n4169), .B(n4170), .Z(o[530]) );
  AND U4691 ( .A(n4171), .B(n4172), .Z(n4170) );
  AND U4692 ( .A(n4173), .B(p_input[3530]), .Z(n4172) );
  AND U4693 ( .A(p_input[2530]), .B(p_input[1530]), .Z(n4173) );
  AND U4694 ( .A(p_input[530]), .B(p_input[4530]), .Z(n4171) );
  AND U4695 ( .A(n4174), .B(n4175), .Z(n4169) );
  AND U4696 ( .A(n4176), .B(p_input[7530]), .Z(n4175) );
  AND U4697 ( .A(p_input[6530]), .B(p_input[5530]), .Z(n4176) );
  AND U4698 ( .A(p_input[9530]), .B(p_input[8530]), .Z(n4174) );
  AND U4699 ( .A(n4177), .B(n4178), .Z(o[52]) );
  AND U4700 ( .A(n4179), .B(n4180), .Z(n4178) );
  AND U4701 ( .A(n4181), .B(p_input[3052]), .Z(n4180) );
  AND U4702 ( .A(p_input[2052]), .B(p_input[1052]), .Z(n4181) );
  AND U4703 ( .A(p_input[5052]), .B(p_input[4052]), .Z(n4179) );
  AND U4704 ( .A(n4182), .B(n4183), .Z(n4177) );
  AND U4705 ( .A(n4184), .B(p_input[7052]), .Z(n4183) );
  AND U4706 ( .A(p_input[6052]), .B(p_input[52]), .Z(n4184) );
  AND U4707 ( .A(p_input[9052]), .B(p_input[8052]), .Z(n4182) );
  AND U4708 ( .A(n4185), .B(n4186), .Z(o[529]) );
  AND U4709 ( .A(n4187), .B(n4188), .Z(n4186) );
  AND U4710 ( .A(n4189), .B(p_input[3529]), .Z(n4188) );
  AND U4711 ( .A(p_input[2529]), .B(p_input[1529]), .Z(n4189) );
  AND U4712 ( .A(p_input[529]), .B(p_input[4529]), .Z(n4187) );
  AND U4713 ( .A(n4190), .B(n4191), .Z(n4185) );
  AND U4714 ( .A(n4192), .B(p_input[7529]), .Z(n4191) );
  AND U4715 ( .A(p_input[6529]), .B(p_input[5529]), .Z(n4192) );
  AND U4716 ( .A(p_input[9529]), .B(p_input[8529]), .Z(n4190) );
  AND U4717 ( .A(n4193), .B(n4194), .Z(o[528]) );
  AND U4718 ( .A(n4195), .B(n4196), .Z(n4194) );
  AND U4719 ( .A(n4197), .B(p_input[3528]), .Z(n4196) );
  AND U4720 ( .A(p_input[2528]), .B(p_input[1528]), .Z(n4197) );
  AND U4721 ( .A(p_input[528]), .B(p_input[4528]), .Z(n4195) );
  AND U4722 ( .A(n4198), .B(n4199), .Z(n4193) );
  AND U4723 ( .A(n4200), .B(p_input[7528]), .Z(n4199) );
  AND U4724 ( .A(p_input[6528]), .B(p_input[5528]), .Z(n4200) );
  AND U4725 ( .A(p_input[9528]), .B(p_input[8528]), .Z(n4198) );
  AND U4726 ( .A(n4201), .B(n4202), .Z(o[527]) );
  AND U4727 ( .A(n4203), .B(n4204), .Z(n4202) );
  AND U4728 ( .A(n4205), .B(p_input[3527]), .Z(n4204) );
  AND U4729 ( .A(p_input[2527]), .B(p_input[1527]), .Z(n4205) );
  AND U4730 ( .A(p_input[527]), .B(p_input[4527]), .Z(n4203) );
  AND U4731 ( .A(n4206), .B(n4207), .Z(n4201) );
  AND U4732 ( .A(n4208), .B(p_input[7527]), .Z(n4207) );
  AND U4733 ( .A(p_input[6527]), .B(p_input[5527]), .Z(n4208) );
  AND U4734 ( .A(p_input[9527]), .B(p_input[8527]), .Z(n4206) );
  AND U4735 ( .A(n4209), .B(n4210), .Z(o[526]) );
  AND U4736 ( .A(n4211), .B(n4212), .Z(n4210) );
  AND U4737 ( .A(n4213), .B(p_input[3526]), .Z(n4212) );
  AND U4738 ( .A(p_input[2526]), .B(p_input[1526]), .Z(n4213) );
  AND U4739 ( .A(p_input[526]), .B(p_input[4526]), .Z(n4211) );
  AND U4740 ( .A(n4214), .B(n4215), .Z(n4209) );
  AND U4741 ( .A(n4216), .B(p_input[7526]), .Z(n4215) );
  AND U4742 ( .A(p_input[6526]), .B(p_input[5526]), .Z(n4216) );
  AND U4743 ( .A(p_input[9526]), .B(p_input[8526]), .Z(n4214) );
  AND U4744 ( .A(n4217), .B(n4218), .Z(o[525]) );
  AND U4745 ( .A(n4219), .B(n4220), .Z(n4218) );
  AND U4746 ( .A(n4221), .B(p_input[3525]), .Z(n4220) );
  AND U4747 ( .A(p_input[2525]), .B(p_input[1525]), .Z(n4221) );
  AND U4748 ( .A(p_input[525]), .B(p_input[4525]), .Z(n4219) );
  AND U4749 ( .A(n4222), .B(n4223), .Z(n4217) );
  AND U4750 ( .A(n4224), .B(p_input[7525]), .Z(n4223) );
  AND U4751 ( .A(p_input[6525]), .B(p_input[5525]), .Z(n4224) );
  AND U4752 ( .A(p_input[9525]), .B(p_input[8525]), .Z(n4222) );
  AND U4753 ( .A(n4225), .B(n4226), .Z(o[524]) );
  AND U4754 ( .A(n4227), .B(n4228), .Z(n4226) );
  AND U4755 ( .A(n4229), .B(p_input[3524]), .Z(n4228) );
  AND U4756 ( .A(p_input[2524]), .B(p_input[1524]), .Z(n4229) );
  AND U4757 ( .A(p_input[524]), .B(p_input[4524]), .Z(n4227) );
  AND U4758 ( .A(n4230), .B(n4231), .Z(n4225) );
  AND U4759 ( .A(n4232), .B(p_input[7524]), .Z(n4231) );
  AND U4760 ( .A(p_input[6524]), .B(p_input[5524]), .Z(n4232) );
  AND U4761 ( .A(p_input[9524]), .B(p_input[8524]), .Z(n4230) );
  AND U4762 ( .A(n4233), .B(n4234), .Z(o[523]) );
  AND U4763 ( .A(n4235), .B(n4236), .Z(n4234) );
  AND U4764 ( .A(n4237), .B(p_input[3523]), .Z(n4236) );
  AND U4765 ( .A(p_input[2523]), .B(p_input[1523]), .Z(n4237) );
  AND U4766 ( .A(p_input[523]), .B(p_input[4523]), .Z(n4235) );
  AND U4767 ( .A(n4238), .B(n4239), .Z(n4233) );
  AND U4768 ( .A(n4240), .B(p_input[7523]), .Z(n4239) );
  AND U4769 ( .A(p_input[6523]), .B(p_input[5523]), .Z(n4240) );
  AND U4770 ( .A(p_input[9523]), .B(p_input[8523]), .Z(n4238) );
  AND U4771 ( .A(n4241), .B(n4242), .Z(o[522]) );
  AND U4772 ( .A(n4243), .B(n4244), .Z(n4242) );
  AND U4773 ( .A(n4245), .B(p_input[3522]), .Z(n4244) );
  AND U4774 ( .A(p_input[2522]), .B(p_input[1522]), .Z(n4245) );
  AND U4775 ( .A(p_input[522]), .B(p_input[4522]), .Z(n4243) );
  AND U4776 ( .A(n4246), .B(n4247), .Z(n4241) );
  AND U4777 ( .A(n4248), .B(p_input[7522]), .Z(n4247) );
  AND U4778 ( .A(p_input[6522]), .B(p_input[5522]), .Z(n4248) );
  AND U4779 ( .A(p_input[9522]), .B(p_input[8522]), .Z(n4246) );
  AND U4780 ( .A(n4249), .B(n4250), .Z(o[521]) );
  AND U4781 ( .A(n4251), .B(n4252), .Z(n4250) );
  AND U4782 ( .A(n4253), .B(p_input[3521]), .Z(n4252) );
  AND U4783 ( .A(p_input[2521]), .B(p_input[1521]), .Z(n4253) );
  AND U4784 ( .A(p_input[521]), .B(p_input[4521]), .Z(n4251) );
  AND U4785 ( .A(n4254), .B(n4255), .Z(n4249) );
  AND U4786 ( .A(n4256), .B(p_input[7521]), .Z(n4255) );
  AND U4787 ( .A(p_input[6521]), .B(p_input[5521]), .Z(n4256) );
  AND U4788 ( .A(p_input[9521]), .B(p_input[8521]), .Z(n4254) );
  AND U4789 ( .A(n4257), .B(n4258), .Z(o[520]) );
  AND U4790 ( .A(n4259), .B(n4260), .Z(n4258) );
  AND U4791 ( .A(n4261), .B(p_input[3520]), .Z(n4260) );
  AND U4792 ( .A(p_input[2520]), .B(p_input[1520]), .Z(n4261) );
  AND U4793 ( .A(p_input[520]), .B(p_input[4520]), .Z(n4259) );
  AND U4794 ( .A(n4262), .B(n4263), .Z(n4257) );
  AND U4795 ( .A(n4264), .B(p_input[7520]), .Z(n4263) );
  AND U4796 ( .A(p_input[6520]), .B(p_input[5520]), .Z(n4264) );
  AND U4797 ( .A(p_input[9520]), .B(p_input[8520]), .Z(n4262) );
  AND U4798 ( .A(n4265), .B(n4266), .Z(o[51]) );
  AND U4799 ( .A(n4267), .B(n4268), .Z(n4266) );
  AND U4800 ( .A(n4269), .B(p_input[3051]), .Z(n4268) );
  AND U4801 ( .A(p_input[2051]), .B(p_input[1051]), .Z(n4269) );
  AND U4802 ( .A(p_input[5051]), .B(p_input[4051]), .Z(n4267) );
  AND U4803 ( .A(n4270), .B(n4271), .Z(n4265) );
  AND U4804 ( .A(n4272), .B(p_input[7051]), .Z(n4271) );
  AND U4805 ( .A(p_input[6051]), .B(p_input[51]), .Z(n4272) );
  AND U4806 ( .A(p_input[9051]), .B(p_input[8051]), .Z(n4270) );
  AND U4807 ( .A(n4273), .B(n4274), .Z(o[519]) );
  AND U4808 ( .A(n4275), .B(n4276), .Z(n4274) );
  AND U4809 ( .A(n4277), .B(p_input[3519]), .Z(n4276) );
  AND U4810 ( .A(p_input[2519]), .B(p_input[1519]), .Z(n4277) );
  AND U4811 ( .A(p_input[519]), .B(p_input[4519]), .Z(n4275) );
  AND U4812 ( .A(n4278), .B(n4279), .Z(n4273) );
  AND U4813 ( .A(n4280), .B(p_input[7519]), .Z(n4279) );
  AND U4814 ( .A(p_input[6519]), .B(p_input[5519]), .Z(n4280) );
  AND U4815 ( .A(p_input[9519]), .B(p_input[8519]), .Z(n4278) );
  AND U4816 ( .A(n4281), .B(n4282), .Z(o[518]) );
  AND U4817 ( .A(n4283), .B(n4284), .Z(n4282) );
  AND U4818 ( .A(n4285), .B(p_input[3518]), .Z(n4284) );
  AND U4819 ( .A(p_input[2518]), .B(p_input[1518]), .Z(n4285) );
  AND U4820 ( .A(p_input[518]), .B(p_input[4518]), .Z(n4283) );
  AND U4821 ( .A(n4286), .B(n4287), .Z(n4281) );
  AND U4822 ( .A(n4288), .B(p_input[7518]), .Z(n4287) );
  AND U4823 ( .A(p_input[6518]), .B(p_input[5518]), .Z(n4288) );
  AND U4824 ( .A(p_input[9518]), .B(p_input[8518]), .Z(n4286) );
  AND U4825 ( .A(n4289), .B(n4290), .Z(o[517]) );
  AND U4826 ( .A(n4291), .B(n4292), .Z(n4290) );
  AND U4827 ( .A(n4293), .B(p_input[3517]), .Z(n4292) );
  AND U4828 ( .A(p_input[2517]), .B(p_input[1517]), .Z(n4293) );
  AND U4829 ( .A(p_input[517]), .B(p_input[4517]), .Z(n4291) );
  AND U4830 ( .A(n4294), .B(n4295), .Z(n4289) );
  AND U4831 ( .A(n4296), .B(p_input[7517]), .Z(n4295) );
  AND U4832 ( .A(p_input[6517]), .B(p_input[5517]), .Z(n4296) );
  AND U4833 ( .A(p_input[9517]), .B(p_input[8517]), .Z(n4294) );
  AND U4834 ( .A(n4297), .B(n4298), .Z(o[516]) );
  AND U4835 ( .A(n4299), .B(n4300), .Z(n4298) );
  AND U4836 ( .A(n4301), .B(p_input[3516]), .Z(n4300) );
  AND U4837 ( .A(p_input[2516]), .B(p_input[1516]), .Z(n4301) );
  AND U4838 ( .A(p_input[516]), .B(p_input[4516]), .Z(n4299) );
  AND U4839 ( .A(n4302), .B(n4303), .Z(n4297) );
  AND U4840 ( .A(n4304), .B(p_input[7516]), .Z(n4303) );
  AND U4841 ( .A(p_input[6516]), .B(p_input[5516]), .Z(n4304) );
  AND U4842 ( .A(p_input[9516]), .B(p_input[8516]), .Z(n4302) );
  AND U4843 ( .A(n4305), .B(n4306), .Z(o[515]) );
  AND U4844 ( .A(n4307), .B(n4308), .Z(n4306) );
  AND U4845 ( .A(n4309), .B(p_input[3515]), .Z(n4308) );
  AND U4846 ( .A(p_input[2515]), .B(p_input[1515]), .Z(n4309) );
  AND U4847 ( .A(p_input[515]), .B(p_input[4515]), .Z(n4307) );
  AND U4848 ( .A(n4310), .B(n4311), .Z(n4305) );
  AND U4849 ( .A(n4312), .B(p_input[7515]), .Z(n4311) );
  AND U4850 ( .A(p_input[6515]), .B(p_input[5515]), .Z(n4312) );
  AND U4851 ( .A(p_input[9515]), .B(p_input[8515]), .Z(n4310) );
  AND U4852 ( .A(n4313), .B(n4314), .Z(o[514]) );
  AND U4853 ( .A(n4315), .B(n4316), .Z(n4314) );
  AND U4854 ( .A(n4317), .B(p_input[3514]), .Z(n4316) );
  AND U4855 ( .A(p_input[2514]), .B(p_input[1514]), .Z(n4317) );
  AND U4856 ( .A(p_input[514]), .B(p_input[4514]), .Z(n4315) );
  AND U4857 ( .A(n4318), .B(n4319), .Z(n4313) );
  AND U4858 ( .A(n4320), .B(p_input[7514]), .Z(n4319) );
  AND U4859 ( .A(p_input[6514]), .B(p_input[5514]), .Z(n4320) );
  AND U4860 ( .A(p_input[9514]), .B(p_input[8514]), .Z(n4318) );
  AND U4861 ( .A(n4321), .B(n4322), .Z(o[513]) );
  AND U4862 ( .A(n4323), .B(n4324), .Z(n4322) );
  AND U4863 ( .A(n4325), .B(p_input[3513]), .Z(n4324) );
  AND U4864 ( .A(p_input[2513]), .B(p_input[1513]), .Z(n4325) );
  AND U4865 ( .A(p_input[513]), .B(p_input[4513]), .Z(n4323) );
  AND U4866 ( .A(n4326), .B(n4327), .Z(n4321) );
  AND U4867 ( .A(n4328), .B(p_input[7513]), .Z(n4327) );
  AND U4868 ( .A(p_input[6513]), .B(p_input[5513]), .Z(n4328) );
  AND U4869 ( .A(p_input[9513]), .B(p_input[8513]), .Z(n4326) );
  AND U4870 ( .A(n4329), .B(n4330), .Z(o[512]) );
  AND U4871 ( .A(n4331), .B(n4332), .Z(n4330) );
  AND U4872 ( .A(n4333), .B(p_input[3512]), .Z(n4332) );
  AND U4873 ( .A(p_input[2512]), .B(p_input[1512]), .Z(n4333) );
  AND U4874 ( .A(p_input[512]), .B(p_input[4512]), .Z(n4331) );
  AND U4875 ( .A(n4334), .B(n4335), .Z(n4329) );
  AND U4876 ( .A(n4336), .B(p_input[7512]), .Z(n4335) );
  AND U4877 ( .A(p_input[6512]), .B(p_input[5512]), .Z(n4336) );
  AND U4878 ( .A(p_input[9512]), .B(p_input[8512]), .Z(n4334) );
  AND U4879 ( .A(n4337), .B(n4338), .Z(o[511]) );
  AND U4880 ( .A(n4339), .B(n4340), .Z(n4338) );
  AND U4881 ( .A(n4341), .B(p_input[3511]), .Z(n4340) );
  AND U4882 ( .A(p_input[2511]), .B(p_input[1511]), .Z(n4341) );
  AND U4883 ( .A(p_input[511]), .B(p_input[4511]), .Z(n4339) );
  AND U4884 ( .A(n4342), .B(n4343), .Z(n4337) );
  AND U4885 ( .A(n4344), .B(p_input[7511]), .Z(n4343) );
  AND U4886 ( .A(p_input[6511]), .B(p_input[5511]), .Z(n4344) );
  AND U4887 ( .A(p_input[9511]), .B(p_input[8511]), .Z(n4342) );
  AND U4888 ( .A(n4345), .B(n4346), .Z(o[510]) );
  AND U4889 ( .A(n4347), .B(n4348), .Z(n4346) );
  AND U4890 ( .A(n4349), .B(p_input[3510]), .Z(n4348) );
  AND U4891 ( .A(p_input[2510]), .B(p_input[1510]), .Z(n4349) );
  AND U4892 ( .A(p_input[510]), .B(p_input[4510]), .Z(n4347) );
  AND U4893 ( .A(n4350), .B(n4351), .Z(n4345) );
  AND U4894 ( .A(n4352), .B(p_input[7510]), .Z(n4351) );
  AND U4895 ( .A(p_input[6510]), .B(p_input[5510]), .Z(n4352) );
  AND U4896 ( .A(p_input[9510]), .B(p_input[8510]), .Z(n4350) );
  AND U4897 ( .A(n4353), .B(n4354), .Z(o[50]) );
  AND U4898 ( .A(n4355), .B(n4356), .Z(n4354) );
  AND U4899 ( .A(n4357), .B(p_input[3050]), .Z(n4356) );
  AND U4900 ( .A(p_input[2050]), .B(p_input[1050]), .Z(n4357) );
  AND U4901 ( .A(p_input[5050]), .B(p_input[4050]), .Z(n4355) );
  AND U4902 ( .A(n4358), .B(n4359), .Z(n4353) );
  AND U4903 ( .A(n4360), .B(p_input[7050]), .Z(n4359) );
  AND U4904 ( .A(p_input[6050]), .B(p_input[50]), .Z(n4360) );
  AND U4905 ( .A(p_input[9050]), .B(p_input[8050]), .Z(n4358) );
  AND U4906 ( .A(n4361), .B(n4362), .Z(o[509]) );
  AND U4907 ( .A(n4363), .B(n4364), .Z(n4362) );
  AND U4908 ( .A(n4365), .B(p_input[3509]), .Z(n4364) );
  AND U4909 ( .A(p_input[2509]), .B(p_input[1509]), .Z(n4365) );
  AND U4910 ( .A(p_input[509]), .B(p_input[4509]), .Z(n4363) );
  AND U4911 ( .A(n4366), .B(n4367), .Z(n4361) );
  AND U4912 ( .A(n4368), .B(p_input[7509]), .Z(n4367) );
  AND U4913 ( .A(p_input[6509]), .B(p_input[5509]), .Z(n4368) );
  AND U4914 ( .A(p_input[9509]), .B(p_input[8509]), .Z(n4366) );
  AND U4915 ( .A(n4369), .B(n4370), .Z(o[508]) );
  AND U4916 ( .A(n4371), .B(n4372), .Z(n4370) );
  AND U4917 ( .A(n4373), .B(p_input[3508]), .Z(n4372) );
  AND U4918 ( .A(p_input[2508]), .B(p_input[1508]), .Z(n4373) );
  AND U4919 ( .A(p_input[508]), .B(p_input[4508]), .Z(n4371) );
  AND U4920 ( .A(n4374), .B(n4375), .Z(n4369) );
  AND U4921 ( .A(n4376), .B(p_input[7508]), .Z(n4375) );
  AND U4922 ( .A(p_input[6508]), .B(p_input[5508]), .Z(n4376) );
  AND U4923 ( .A(p_input[9508]), .B(p_input[8508]), .Z(n4374) );
  AND U4924 ( .A(n4377), .B(n4378), .Z(o[507]) );
  AND U4925 ( .A(n4379), .B(n4380), .Z(n4378) );
  AND U4926 ( .A(n4381), .B(p_input[3507]), .Z(n4380) );
  AND U4927 ( .A(p_input[2507]), .B(p_input[1507]), .Z(n4381) );
  AND U4928 ( .A(p_input[507]), .B(p_input[4507]), .Z(n4379) );
  AND U4929 ( .A(n4382), .B(n4383), .Z(n4377) );
  AND U4930 ( .A(n4384), .B(p_input[7507]), .Z(n4383) );
  AND U4931 ( .A(p_input[6507]), .B(p_input[5507]), .Z(n4384) );
  AND U4932 ( .A(p_input[9507]), .B(p_input[8507]), .Z(n4382) );
  AND U4933 ( .A(n4385), .B(n4386), .Z(o[506]) );
  AND U4934 ( .A(n4387), .B(n4388), .Z(n4386) );
  AND U4935 ( .A(n4389), .B(p_input[3506]), .Z(n4388) );
  AND U4936 ( .A(p_input[2506]), .B(p_input[1506]), .Z(n4389) );
  AND U4937 ( .A(p_input[506]), .B(p_input[4506]), .Z(n4387) );
  AND U4938 ( .A(n4390), .B(n4391), .Z(n4385) );
  AND U4939 ( .A(n4392), .B(p_input[7506]), .Z(n4391) );
  AND U4940 ( .A(p_input[6506]), .B(p_input[5506]), .Z(n4392) );
  AND U4941 ( .A(p_input[9506]), .B(p_input[8506]), .Z(n4390) );
  AND U4942 ( .A(n4393), .B(n4394), .Z(o[505]) );
  AND U4943 ( .A(n4395), .B(n4396), .Z(n4394) );
  AND U4944 ( .A(n4397), .B(p_input[3505]), .Z(n4396) );
  AND U4945 ( .A(p_input[2505]), .B(p_input[1505]), .Z(n4397) );
  AND U4946 ( .A(p_input[505]), .B(p_input[4505]), .Z(n4395) );
  AND U4947 ( .A(n4398), .B(n4399), .Z(n4393) );
  AND U4948 ( .A(n4400), .B(p_input[7505]), .Z(n4399) );
  AND U4949 ( .A(p_input[6505]), .B(p_input[5505]), .Z(n4400) );
  AND U4950 ( .A(p_input[9505]), .B(p_input[8505]), .Z(n4398) );
  AND U4951 ( .A(n4401), .B(n4402), .Z(o[504]) );
  AND U4952 ( .A(n4403), .B(n4404), .Z(n4402) );
  AND U4953 ( .A(n4405), .B(p_input[3504]), .Z(n4404) );
  AND U4954 ( .A(p_input[2504]), .B(p_input[1504]), .Z(n4405) );
  AND U4955 ( .A(p_input[504]), .B(p_input[4504]), .Z(n4403) );
  AND U4956 ( .A(n4406), .B(n4407), .Z(n4401) );
  AND U4957 ( .A(n4408), .B(p_input[7504]), .Z(n4407) );
  AND U4958 ( .A(p_input[6504]), .B(p_input[5504]), .Z(n4408) );
  AND U4959 ( .A(p_input[9504]), .B(p_input[8504]), .Z(n4406) );
  AND U4960 ( .A(n4409), .B(n4410), .Z(o[503]) );
  AND U4961 ( .A(n4411), .B(n4412), .Z(n4410) );
  AND U4962 ( .A(n4413), .B(p_input[3503]), .Z(n4412) );
  AND U4963 ( .A(p_input[2503]), .B(p_input[1503]), .Z(n4413) );
  AND U4964 ( .A(p_input[503]), .B(p_input[4503]), .Z(n4411) );
  AND U4965 ( .A(n4414), .B(n4415), .Z(n4409) );
  AND U4966 ( .A(n4416), .B(p_input[7503]), .Z(n4415) );
  AND U4967 ( .A(p_input[6503]), .B(p_input[5503]), .Z(n4416) );
  AND U4968 ( .A(p_input[9503]), .B(p_input[8503]), .Z(n4414) );
  AND U4969 ( .A(n4417), .B(n4418), .Z(o[502]) );
  AND U4970 ( .A(n4419), .B(n4420), .Z(n4418) );
  AND U4971 ( .A(n4421), .B(p_input[3502]), .Z(n4420) );
  AND U4972 ( .A(p_input[2502]), .B(p_input[1502]), .Z(n4421) );
  AND U4973 ( .A(p_input[502]), .B(p_input[4502]), .Z(n4419) );
  AND U4974 ( .A(n4422), .B(n4423), .Z(n4417) );
  AND U4975 ( .A(n4424), .B(p_input[7502]), .Z(n4423) );
  AND U4976 ( .A(p_input[6502]), .B(p_input[5502]), .Z(n4424) );
  AND U4977 ( .A(p_input[9502]), .B(p_input[8502]), .Z(n4422) );
  AND U4978 ( .A(n4425), .B(n4426), .Z(o[501]) );
  AND U4979 ( .A(n4427), .B(n4428), .Z(n4426) );
  AND U4980 ( .A(n4429), .B(p_input[3501]), .Z(n4428) );
  AND U4981 ( .A(p_input[2501]), .B(p_input[1501]), .Z(n4429) );
  AND U4982 ( .A(p_input[501]), .B(p_input[4501]), .Z(n4427) );
  AND U4983 ( .A(n4430), .B(n4431), .Z(n4425) );
  AND U4984 ( .A(n4432), .B(p_input[7501]), .Z(n4431) );
  AND U4985 ( .A(p_input[6501]), .B(p_input[5501]), .Z(n4432) );
  AND U4986 ( .A(p_input[9501]), .B(p_input[8501]), .Z(n4430) );
  AND U4987 ( .A(n4433), .B(n4434), .Z(o[500]) );
  AND U4988 ( .A(n4435), .B(n4436), .Z(n4434) );
  AND U4989 ( .A(n4437), .B(p_input[3500]), .Z(n4436) );
  AND U4990 ( .A(p_input[2500]), .B(p_input[1500]), .Z(n4437) );
  AND U4991 ( .A(p_input[500]), .B(p_input[4500]), .Z(n4435) );
  AND U4992 ( .A(n4438), .B(n4439), .Z(n4433) );
  AND U4993 ( .A(n4440), .B(p_input[7500]), .Z(n4439) );
  AND U4994 ( .A(p_input[6500]), .B(p_input[5500]), .Z(n4440) );
  AND U4995 ( .A(p_input[9500]), .B(p_input[8500]), .Z(n4438) );
  AND U4996 ( .A(n4441), .B(n4442), .Z(o[4]) );
  AND U4997 ( .A(n4443), .B(n4444), .Z(n4442) );
  AND U4998 ( .A(n4445), .B(p_input[3004]), .Z(n4444) );
  AND U4999 ( .A(p_input[2004]), .B(p_input[1004]), .Z(n4445) );
  AND U5000 ( .A(p_input[4]), .B(p_input[4004]), .Z(n4443) );
  AND U5001 ( .A(n4446), .B(n4447), .Z(n4441) );
  AND U5002 ( .A(n4448), .B(p_input[7004]), .Z(n4447) );
  AND U5003 ( .A(p_input[6004]), .B(p_input[5004]), .Z(n4448) );
  AND U5004 ( .A(p_input[9004]), .B(p_input[8004]), .Z(n4446) );
  AND U5005 ( .A(n4449), .B(n4450), .Z(o[49]) );
  AND U5006 ( .A(n4451), .B(n4452), .Z(n4450) );
  AND U5007 ( .A(n4453), .B(p_input[3049]), .Z(n4452) );
  AND U5008 ( .A(p_input[2049]), .B(p_input[1049]), .Z(n4453) );
  AND U5009 ( .A(p_input[49]), .B(p_input[4049]), .Z(n4451) );
  AND U5010 ( .A(n4454), .B(n4455), .Z(n4449) );
  AND U5011 ( .A(n4456), .B(p_input[7049]), .Z(n4455) );
  AND U5012 ( .A(p_input[6049]), .B(p_input[5049]), .Z(n4456) );
  AND U5013 ( .A(p_input[9049]), .B(p_input[8049]), .Z(n4454) );
  AND U5014 ( .A(n4457), .B(n4458), .Z(o[499]) );
  AND U5015 ( .A(n4459), .B(n4460), .Z(n4458) );
  AND U5016 ( .A(n4461), .B(p_input[3499]), .Z(n4460) );
  AND U5017 ( .A(p_input[2499]), .B(p_input[1499]), .Z(n4461) );
  AND U5018 ( .A(p_input[499]), .B(p_input[4499]), .Z(n4459) );
  AND U5019 ( .A(n4462), .B(n4463), .Z(n4457) );
  AND U5020 ( .A(n4464), .B(p_input[7499]), .Z(n4463) );
  AND U5021 ( .A(p_input[6499]), .B(p_input[5499]), .Z(n4464) );
  AND U5022 ( .A(p_input[9499]), .B(p_input[8499]), .Z(n4462) );
  AND U5023 ( .A(n4465), .B(n4466), .Z(o[498]) );
  AND U5024 ( .A(n4467), .B(n4468), .Z(n4466) );
  AND U5025 ( .A(n4469), .B(p_input[3498]), .Z(n4468) );
  AND U5026 ( .A(p_input[2498]), .B(p_input[1498]), .Z(n4469) );
  AND U5027 ( .A(p_input[498]), .B(p_input[4498]), .Z(n4467) );
  AND U5028 ( .A(n4470), .B(n4471), .Z(n4465) );
  AND U5029 ( .A(n4472), .B(p_input[7498]), .Z(n4471) );
  AND U5030 ( .A(p_input[6498]), .B(p_input[5498]), .Z(n4472) );
  AND U5031 ( .A(p_input[9498]), .B(p_input[8498]), .Z(n4470) );
  AND U5032 ( .A(n4473), .B(n4474), .Z(o[497]) );
  AND U5033 ( .A(n4475), .B(n4476), .Z(n4474) );
  AND U5034 ( .A(n4477), .B(p_input[3497]), .Z(n4476) );
  AND U5035 ( .A(p_input[2497]), .B(p_input[1497]), .Z(n4477) );
  AND U5036 ( .A(p_input[497]), .B(p_input[4497]), .Z(n4475) );
  AND U5037 ( .A(n4478), .B(n4479), .Z(n4473) );
  AND U5038 ( .A(n4480), .B(p_input[7497]), .Z(n4479) );
  AND U5039 ( .A(p_input[6497]), .B(p_input[5497]), .Z(n4480) );
  AND U5040 ( .A(p_input[9497]), .B(p_input[8497]), .Z(n4478) );
  AND U5041 ( .A(n4481), .B(n4482), .Z(o[496]) );
  AND U5042 ( .A(n4483), .B(n4484), .Z(n4482) );
  AND U5043 ( .A(n4485), .B(p_input[3496]), .Z(n4484) );
  AND U5044 ( .A(p_input[2496]), .B(p_input[1496]), .Z(n4485) );
  AND U5045 ( .A(p_input[496]), .B(p_input[4496]), .Z(n4483) );
  AND U5046 ( .A(n4486), .B(n4487), .Z(n4481) );
  AND U5047 ( .A(n4488), .B(p_input[7496]), .Z(n4487) );
  AND U5048 ( .A(p_input[6496]), .B(p_input[5496]), .Z(n4488) );
  AND U5049 ( .A(p_input[9496]), .B(p_input[8496]), .Z(n4486) );
  AND U5050 ( .A(n4489), .B(n4490), .Z(o[495]) );
  AND U5051 ( .A(n4491), .B(n4492), .Z(n4490) );
  AND U5052 ( .A(n4493), .B(p_input[3495]), .Z(n4492) );
  AND U5053 ( .A(p_input[2495]), .B(p_input[1495]), .Z(n4493) );
  AND U5054 ( .A(p_input[495]), .B(p_input[4495]), .Z(n4491) );
  AND U5055 ( .A(n4494), .B(n4495), .Z(n4489) );
  AND U5056 ( .A(n4496), .B(p_input[7495]), .Z(n4495) );
  AND U5057 ( .A(p_input[6495]), .B(p_input[5495]), .Z(n4496) );
  AND U5058 ( .A(p_input[9495]), .B(p_input[8495]), .Z(n4494) );
  AND U5059 ( .A(n4497), .B(n4498), .Z(o[494]) );
  AND U5060 ( .A(n4499), .B(n4500), .Z(n4498) );
  AND U5061 ( .A(n4501), .B(p_input[3494]), .Z(n4500) );
  AND U5062 ( .A(p_input[2494]), .B(p_input[1494]), .Z(n4501) );
  AND U5063 ( .A(p_input[494]), .B(p_input[4494]), .Z(n4499) );
  AND U5064 ( .A(n4502), .B(n4503), .Z(n4497) );
  AND U5065 ( .A(n4504), .B(p_input[7494]), .Z(n4503) );
  AND U5066 ( .A(p_input[6494]), .B(p_input[5494]), .Z(n4504) );
  AND U5067 ( .A(p_input[9494]), .B(p_input[8494]), .Z(n4502) );
  AND U5068 ( .A(n4505), .B(n4506), .Z(o[493]) );
  AND U5069 ( .A(n4507), .B(n4508), .Z(n4506) );
  AND U5070 ( .A(n4509), .B(p_input[3493]), .Z(n4508) );
  AND U5071 ( .A(p_input[2493]), .B(p_input[1493]), .Z(n4509) );
  AND U5072 ( .A(p_input[493]), .B(p_input[4493]), .Z(n4507) );
  AND U5073 ( .A(n4510), .B(n4511), .Z(n4505) );
  AND U5074 ( .A(n4512), .B(p_input[7493]), .Z(n4511) );
  AND U5075 ( .A(p_input[6493]), .B(p_input[5493]), .Z(n4512) );
  AND U5076 ( .A(p_input[9493]), .B(p_input[8493]), .Z(n4510) );
  AND U5077 ( .A(n4513), .B(n4514), .Z(o[492]) );
  AND U5078 ( .A(n4515), .B(n4516), .Z(n4514) );
  AND U5079 ( .A(n4517), .B(p_input[3492]), .Z(n4516) );
  AND U5080 ( .A(p_input[2492]), .B(p_input[1492]), .Z(n4517) );
  AND U5081 ( .A(p_input[492]), .B(p_input[4492]), .Z(n4515) );
  AND U5082 ( .A(n4518), .B(n4519), .Z(n4513) );
  AND U5083 ( .A(n4520), .B(p_input[7492]), .Z(n4519) );
  AND U5084 ( .A(p_input[6492]), .B(p_input[5492]), .Z(n4520) );
  AND U5085 ( .A(p_input[9492]), .B(p_input[8492]), .Z(n4518) );
  AND U5086 ( .A(n4521), .B(n4522), .Z(o[491]) );
  AND U5087 ( .A(n4523), .B(n4524), .Z(n4522) );
  AND U5088 ( .A(n4525), .B(p_input[3491]), .Z(n4524) );
  AND U5089 ( .A(p_input[2491]), .B(p_input[1491]), .Z(n4525) );
  AND U5090 ( .A(p_input[491]), .B(p_input[4491]), .Z(n4523) );
  AND U5091 ( .A(n4526), .B(n4527), .Z(n4521) );
  AND U5092 ( .A(n4528), .B(p_input[7491]), .Z(n4527) );
  AND U5093 ( .A(p_input[6491]), .B(p_input[5491]), .Z(n4528) );
  AND U5094 ( .A(p_input[9491]), .B(p_input[8491]), .Z(n4526) );
  AND U5095 ( .A(n4529), .B(n4530), .Z(o[490]) );
  AND U5096 ( .A(n4531), .B(n4532), .Z(n4530) );
  AND U5097 ( .A(n4533), .B(p_input[3490]), .Z(n4532) );
  AND U5098 ( .A(p_input[2490]), .B(p_input[1490]), .Z(n4533) );
  AND U5099 ( .A(p_input[490]), .B(p_input[4490]), .Z(n4531) );
  AND U5100 ( .A(n4534), .B(n4535), .Z(n4529) );
  AND U5101 ( .A(n4536), .B(p_input[7490]), .Z(n4535) );
  AND U5102 ( .A(p_input[6490]), .B(p_input[5490]), .Z(n4536) );
  AND U5103 ( .A(p_input[9490]), .B(p_input[8490]), .Z(n4534) );
  AND U5104 ( .A(n4537), .B(n4538), .Z(o[48]) );
  AND U5105 ( .A(n4539), .B(n4540), .Z(n4538) );
  AND U5106 ( .A(n4541), .B(p_input[3048]), .Z(n4540) );
  AND U5107 ( .A(p_input[2048]), .B(p_input[1048]), .Z(n4541) );
  AND U5108 ( .A(p_input[48]), .B(p_input[4048]), .Z(n4539) );
  AND U5109 ( .A(n4542), .B(n4543), .Z(n4537) );
  AND U5110 ( .A(n4544), .B(p_input[7048]), .Z(n4543) );
  AND U5111 ( .A(p_input[6048]), .B(p_input[5048]), .Z(n4544) );
  AND U5112 ( .A(p_input[9048]), .B(p_input[8048]), .Z(n4542) );
  AND U5113 ( .A(n4545), .B(n4546), .Z(o[489]) );
  AND U5114 ( .A(n4547), .B(n4548), .Z(n4546) );
  AND U5115 ( .A(n4549), .B(p_input[3489]), .Z(n4548) );
  AND U5116 ( .A(p_input[2489]), .B(p_input[1489]), .Z(n4549) );
  AND U5117 ( .A(p_input[489]), .B(p_input[4489]), .Z(n4547) );
  AND U5118 ( .A(n4550), .B(n4551), .Z(n4545) );
  AND U5119 ( .A(n4552), .B(p_input[7489]), .Z(n4551) );
  AND U5120 ( .A(p_input[6489]), .B(p_input[5489]), .Z(n4552) );
  AND U5121 ( .A(p_input[9489]), .B(p_input[8489]), .Z(n4550) );
  AND U5122 ( .A(n4553), .B(n4554), .Z(o[488]) );
  AND U5123 ( .A(n4555), .B(n4556), .Z(n4554) );
  AND U5124 ( .A(n4557), .B(p_input[3488]), .Z(n4556) );
  AND U5125 ( .A(p_input[2488]), .B(p_input[1488]), .Z(n4557) );
  AND U5126 ( .A(p_input[488]), .B(p_input[4488]), .Z(n4555) );
  AND U5127 ( .A(n4558), .B(n4559), .Z(n4553) );
  AND U5128 ( .A(n4560), .B(p_input[7488]), .Z(n4559) );
  AND U5129 ( .A(p_input[6488]), .B(p_input[5488]), .Z(n4560) );
  AND U5130 ( .A(p_input[9488]), .B(p_input[8488]), .Z(n4558) );
  AND U5131 ( .A(n4561), .B(n4562), .Z(o[487]) );
  AND U5132 ( .A(n4563), .B(n4564), .Z(n4562) );
  AND U5133 ( .A(n4565), .B(p_input[3487]), .Z(n4564) );
  AND U5134 ( .A(p_input[2487]), .B(p_input[1487]), .Z(n4565) );
  AND U5135 ( .A(p_input[487]), .B(p_input[4487]), .Z(n4563) );
  AND U5136 ( .A(n4566), .B(n4567), .Z(n4561) );
  AND U5137 ( .A(n4568), .B(p_input[7487]), .Z(n4567) );
  AND U5138 ( .A(p_input[6487]), .B(p_input[5487]), .Z(n4568) );
  AND U5139 ( .A(p_input[9487]), .B(p_input[8487]), .Z(n4566) );
  AND U5140 ( .A(n4569), .B(n4570), .Z(o[486]) );
  AND U5141 ( .A(n4571), .B(n4572), .Z(n4570) );
  AND U5142 ( .A(n4573), .B(p_input[3486]), .Z(n4572) );
  AND U5143 ( .A(p_input[2486]), .B(p_input[1486]), .Z(n4573) );
  AND U5144 ( .A(p_input[486]), .B(p_input[4486]), .Z(n4571) );
  AND U5145 ( .A(n4574), .B(n4575), .Z(n4569) );
  AND U5146 ( .A(n4576), .B(p_input[7486]), .Z(n4575) );
  AND U5147 ( .A(p_input[6486]), .B(p_input[5486]), .Z(n4576) );
  AND U5148 ( .A(p_input[9486]), .B(p_input[8486]), .Z(n4574) );
  AND U5149 ( .A(n4577), .B(n4578), .Z(o[485]) );
  AND U5150 ( .A(n4579), .B(n4580), .Z(n4578) );
  AND U5151 ( .A(n4581), .B(p_input[3485]), .Z(n4580) );
  AND U5152 ( .A(p_input[2485]), .B(p_input[1485]), .Z(n4581) );
  AND U5153 ( .A(p_input[485]), .B(p_input[4485]), .Z(n4579) );
  AND U5154 ( .A(n4582), .B(n4583), .Z(n4577) );
  AND U5155 ( .A(n4584), .B(p_input[7485]), .Z(n4583) );
  AND U5156 ( .A(p_input[6485]), .B(p_input[5485]), .Z(n4584) );
  AND U5157 ( .A(p_input[9485]), .B(p_input[8485]), .Z(n4582) );
  AND U5158 ( .A(n4585), .B(n4586), .Z(o[484]) );
  AND U5159 ( .A(n4587), .B(n4588), .Z(n4586) );
  AND U5160 ( .A(n4589), .B(p_input[3484]), .Z(n4588) );
  AND U5161 ( .A(p_input[2484]), .B(p_input[1484]), .Z(n4589) );
  AND U5162 ( .A(p_input[484]), .B(p_input[4484]), .Z(n4587) );
  AND U5163 ( .A(n4590), .B(n4591), .Z(n4585) );
  AND U5164 ( .A(n4592), .B(p_input[7484]), .Z(n4591) );
  AND U5165 ( .A(p_input[6484]), .B(p_input[5484]), .Z(n4592) );
  AND U5166 ( .A(p_input[9484]), .B(p_input[8484]), .Z(n4590) );
  AND U5167 ( .A(n4593), .B(n4594), .Z(o[483]) );
  AND U5168 ( .A(n4595), .B(n4596), .Z(n4594) );
  AND U5169 ( .A(n4597), .B(p_input[3483]), .Z(n4596) );
  AND U5170 ( .A(p_input[2483]), .B(p_input[1483]), .Z(n4597) );
  AND U5171 ( .A(p_input[483]), .B(p_input[4483]), .Z(n4595) );
  AND U5172 ( .A(n4598), .B(n4599), .Z(n4593) );
  AND U5173 ( .A(n4600), .B(p_input[7483]), .Z(n4599) );
  AND U5174 ( .A(p_input[6483]), .B(p_input[5483]), .Z(n4600) );
  AND U5175 ( .A(p_input[9483]), .B(p_input[8483]), .Z(n4598) );
  AND U5176 ( .A(n4601), .B(n4602), .Z(o[482]) );
  AND U5177 ( .A(n4603), .B(n4604), .Z(n4602) );
  AND U5178 ( .A(n4605), .B(p_input[3482]), .Z(n4604) );
  AND U5179 ( .A(p_input[2482]), .B(p_input[1482]), .Z(n4605) );
  AND U5180 ( .A(p_input[482]), .B(p_input[4482]), .Z(n4603) );
  AND U5181 ( .A(n4606), .B(n4607), .Z(n4601) );
  AND U5182 ( .A(n4608), .B(p_input[7482]), .Z(n4607) );
  AND U5183 ( .A(p_input[6482]), .B(p_input[5482]), .Z(n4608) );
  AND U5184 ( .A(p_input[9482]), .B(p_input[8482]), .Z(n4606) );
  AND U5185 ( .A(n4609), .B(n4610), .Z(o[481]) );
  AND U5186 ( .A(n4611), .B(n4612), .Z(n4610) );
  AND U5187 ( .A(n4613), .B(p_input[3481]), .Z(n4612) );
  AND U5188 ( .A(p_input[2481]), .B(p_input[1481]), .Z(n4613) );
  AND U5189 ( .A(p_input[481]), .B(p_input[4481]), .Z(n4611) );
  AND U5190 ( .A(n4614), .B(n4615), .Z(n4609) );
  AND U5191 ( .A(n4616), .B(p_input[7481]), .Z(n4615) );
  AND U5192 ( .A(p_input[6481]), .B(p_input[5481]), .Z(n4616) );
  AND U5193 ( .A(p_input[9481]), .B(p_input[8481]), .Z(n4614) );
  AND U5194 ( .A(n4617), .B(n4618), .Z(o[480]) );
  AND U5195 ( .A(n4619), .B(n4620), .Z(n4618) );
  AND U5196 ( .A(n4621), .B(p_input[3480]), .Z(n4620) );
  AND U5197 ( .A(p_input[2480]), .B(p_input[1480]), .Z(n4621) );
  AND U5198 ( .A(p_input[480]), .B(p_input[4480]), .Z(n4619) );
  AND U5199 ( .A(n4622), .B(n4623), .Z(n4617) );
  AND U5200 ( .A(n4624), .B(p_input[7480]), .Z(n4623) );
  AND U5201 ( .A(p_input[6480]), .B(p_input[5480]), .Z(n4624) );
  AND U5202 ( .A(p_input[9480]), .B(p_input[8480]), .Z(n4622) );
  AND U5203 ( .A(n4625), .B(n4626), .Z(o[47]) );
  AND U5204 ( .A(n4627), .B(n4628), .Z(n4626) );
  AND U5205 ( .A(n4629), .B(p_input[3047]), .Z(n4628) );
  AND U5206 ( .A(p_input[2047]), .B(p_input[1047]), .Z(n4629) );
  AND U5207 ( .A(p_input[47]), .B(p_input[4047]), .Z(n4627) );
  AND U5208 ( .A(n4630), .B(n4631), .Z(n4625) );
  AND U5209 ( .A(n4632), .B(p_input[7047]), .Z(n4631) );
  AND U5210 ( .A(p_input[6047]), .B(p_input[5047]), .Z(n4632) );
  AND U5211 ( .A(p_input[9047]), .B(p_input[8047]), .Z(n4630) );
  AND U5212 ( .A(n4633), .B(n4634), .Z(o[479]) );
  AND U5213 ( .A(n4635), .B(n4636), .Z(n4634) );
  AND U5214 ( .A(n4637), .B(p_input[3479]), .Z(n4636) );
  AND U5215 ( .A(p_input[2479]), .B(p_input[1479]), .Z(n4637) );
  AND U5216 ( .A(p_input[479]), .B(p_input[4479]), .Z(n4635) );
  AND U5217 ( .A(n4638), .B(n4639), .Z(n4633) );
  AND U5218 ( .A(n4640), .B(p_input[7479]), .Z(n4639) );
  AND U5219 ( .A(p_input[6479]), .B(p_input[5479]), .Z(n4640) );
  AND U5220 ( .A(p_input[9479]), .B(p_input[8479]), .Z(n4638) );
  AND U5221 ( .A(n4641), .B(n4642), .Z(o[478]) );
  AND U5222 ( .A(n4643), .B(n4644), .Z(n4642) );
  AND U5223 ( .A(n4645), .B(p_input[3478]), .Z(n4644) );
  AND U5224 ( .A(p_input[2478]), .B(p_input[1478]), .Z(n4645) );
  AND U5225 ( .A(p_input[478]), .B(p_input[4478]), .Z(n4643) );
  AND U5226 ( .A(n4646), .B(n4647), .Z(n4641) );
  AND U5227 ( .A(n4648), .B(p_input[7478]), .Z(n4647) );
  AND U5228 ( .A(p_input[6478]), .B(p_input[5478]), .Z(n4648) );
  AND U5229 ( .A(p_input[9478]), .B(p_input[8478]), .Z(n4646) );
  AND U5230 ( .A(n4649), .B(n4650), .Z(o[477]) );
  AND U5231 ( .A(n4651), .B(n4652), .Z(n4650) );
  AND U5232 ( .A(n4653), .B(p_input[3477]), .Z(n4652) );
  AND U5233 ( .A(p_input[2477]), .B(p_input[1477]), .Z(n4653) );
  AND U5234 ( .A(p_input[477]), .B(p_input[4477]), .Z(n4651) );
  AND U5235 ( .A(n4654), .B(n4655), .Z(n4649) );
  AND U5236 ( .A(n4656), .B(p_input[7477]), .Z(n4655) );
  AND U5237 ( .A(p_input[6477]), .B(p_input[5477]), .Z(n4656) );
  AND U5238 ( .A(p_input[9477]), .B(p_input[8477]), .Z(n4654) );
  AND U5239 ( .A(n4657), .B(n4658), .Z(o[476]) );
  AND U5240 ( .A(n4659), .B(n4660), .Z(n4658) );
  AND U5241 ( .A(n4661), .B(p_input[3476]), .Z(n4660) );
  AND U5242 ( .A(p_input[2476]), .B(p_input[1476]), .Z(n4661) );
  AND U5243 ( .A(p_input[476]), .B(p_input[4476]), .Z(n4659) );
  AND U5244 ( .A(n4662), .B(n4663), .Z(n4657) );
  AND U5245 ( .A(n4664), .B(p_input[7476]), .Z(n4663) );
  AND U5246 ( .A(p_input[6476]), .B(p_input[5476]), .Z(n4664) );
  AND U5247 ( .A(p_input[9476]), .B(p_input[8476]), .Z(n4662) );
  AND U5248 ( .A(n4665), .B(n4666), .Z(o[475]) );
  AND U5249 ( .A(n4667), .B(n4668), .Z(n4666) );
  AND U5250 ( .A(n4669), .B(p_input[3475]), .Z(n4668) );
  AND U5251 ( .A(p_input[2475]), .B(p_input[1475]), .Z(n4669) );
  AND U5252 ( .A(p_input[475]), .B(p_input[4475]), .Z(n4667) );
  AND U5253 ( .A(n4670), .B(n4671), .Z(n4665) );
  AND U5254 ( .A(n4672), .B(p_input[7475]), .Z(n4671) );
  AND U5255 ( .A(p_input[6475]), .B(p_input[5475]), .Z(n4672) );
  AND U5256 ( .A(p_input[9475]), .B(p_input[8475]), .Z(n4670) );
  AND U5257 ( .A(n4673), .B(n4674), .Z(o[474]) );
  AND U5258 ( .A(n4675), .B(n4676), .Z(n4674) );
  AND U5259 ( .A(n4677), .B(p_input[3474]), .Z(n4676) );
  AND U5260 ( .A(p_input[2474]), .B(p_input[1474]), .Z(n4677) );
  AND U5261 ( .A(p_input[474]), .B(p_input[4474]), .Z(n4675) );
  AND U5262 ( .A(n4678), .B(n4679), .Z(n4673) );
  AND U5263 ( .A(n4680), .B(p_input[7474]), .Z(n4679) );
  AND U5264 ( .A(p_input[6474]), .B(p_input[5474]), .Z(n4680) );
  AND U5265 ( .A(p_input[9474]), .B(p_input[8474]), .Z(n4678) );
  AND U5266 ( .A(n4681), .B(n4682), .Z(o[473]) );
  AND U5267 ( .A(n4683), .B(n4684), .Z(n4682) );
  AND U5268 ( .A(n4685), .B(p_input[3473]), .Z(n4684) );
  AND U5269 ( .A(p_input[2473]), .B(p_input[1473]), .Z(n4685) );
  AND U5270 ( .A(p_input[473]), .B(p_input[4473]), .Z(n4683) );
  AND U5271 ( .A(n4686), .B(n4687), .Z(n4681) );
  AND U5272 ( .A(n4688), .B(p_input[7473]), .Z(n4687) );
  AND U5273 ( .A(p_input[6473]), .B(p_input[5473]), .Z(n4688) );
  AND U5274 ( .A(p_input[9473]), .B(p_input[8473]), .Z(n4686) );
  AND U5275 ( .A(n4689), .B(n4690), .Z(o[472]) );
  AND U5276 ( .A(n4691), .B(n4692), .Z(n4690) );
  AND U5277 ( .A(n4693), .B(p_input[3472]), .Z(n4692) );
  AND U5278 ( .A(p_input[2472]), .B(p_input[1472]), .Z(n4693) );
  AND U5279 ( .A(p_input[472]), .B(p_input[4472]), .Z(n4691) );
  AND U5280 ( .A(n4694), .B(n4695), .Z(n4689) );
  AND U5281 ( .A(n4696), .B(p_input[7472]), .Z(n4695) );
  AND U5282 ( .A(p_input[6472]), .B(p_input[5472]), .Z(n4696) );
  AND U5283 ( .A(p_input[9472]), .B(p_input[8472]), .Z(n4694) );
  AND U5284 ( .A(n4697), .B(n4698), .Z(o[471]) );
  AND U5285 ( .A(n4699), .B(n4700), .Z(n4698) );
  AND U5286 ( .A(n4701), .B(p_input[3471]), .Z(n4700) );
  AND U5287 ( .A(p_input[2471]), .B(p_input[1471]), .Z(n4701) );
  AND U5288 ( .A(p_input[471]), .B(p_input[4471]), .Z(n4699) );
  AND U5289 ( .A(n4702), .B(n4703), .Z(n4697) );
  AND U5290 ( .A(n4704), .B(p_input[7471]), .Z(n4703) );
  AND U5291 ( .A(p_input[6471]), .B(p_input[5471]), .Z(n4704) );
  AND U5292 ( .A(p_input[9471]), .B(p_input[8471]), .Z(n4702) );
  AND U5293 ( .A(n4705), .B(n4706), .Z(o[470]) );
  AND U5294 ( .A(n4707), .B(n4708), .Z(n4706) );
  AND U5295 ( .A(n4709), .B(p_input[3470]), .Z(n4708) );
  AND U5296 ( .A(p_input[2470]), .B(p_input[1470]), .Z(n4709) );
  AND U5297 ( .A(p_input[470]), .B(p_input[4470]), .Z(n4707) );
  AND U5298 ( .A(n4710), .B(n4711), .Z(n4705) );
  AND U5299 ( .A(n4712), .B(p_input[7470]), .Z(n4711) );
  AND U5300 ( .A(p_input[6470]), .B(p_input[5470]), .Z(n4712) );
  AND U5301 ( .A(p_input[9470]), .B(p_input[8470]), .Z(n4710) );
  AND U5302 ( .A(n4713), .B(n4714), .Z(o[46]) );
  AND U5303 ( .A(n4715), .B(n4716), .Z(n4714) );
  AND U5304 ( .A(n4717), .B(p_input[3046]), .Z(n4716) );
  AND U5305 ( .A(p_input[2046]), .B(p_input[1046]), .Z(n4717) );
  AND U5306 ( .A(p_input[46]), .B(p_input[4046]), .Z(n4715) );
  AND U5307 ( .A(n4718), .B(n4719), .Z(n4713) );
  AND U5308 ( .A(n4720), .B(p_input[7046]), .Z(n4719) );
  AND U5309 ( .A(p_input[6046]), .B(p_input[5046]), .Z(n4720) );
  AND U5310 ( .A(p_input[9046]), .B(p_input[8046]), .Z(n4718) );
  AND U5311 ( .A(n4721), .B(n4722), .Z(o[469]) );
  AND U5312 ( .A(n4723), .B(n4724), .Z(n4722) );
  AND U5313 ( .A(n4725), .B(p_input[3469]), .Z(n4724) );
  AND U5314 ( .A(p_input[2469]), .B(p_input[1469]), .Z(n4725) );
  AND U5315 ( .A(p_input[469]), .B(p_input[4469]), .Z(n4723) );
  AND U5316 ( .A(n4726), .B(n4727), .Z(n4721) );
  AND U5317 ( .A(n4728), .B(p_input[7469]), .Z(n4727) );
  AND U5318 ( .A(p_input[6469]), .B(p_input[5469]), .Z(n4728) );
  AND U5319 ( .A(p_input[9469]), .B(p_input[8469]), .Z(n4726) );
  AND U5320 ( .A(n4729), .B(n4730), .Z(o[468]) );
  AND U5321 ( .A(n4731), .B(n4732), .Z(n4730) );
  AND U5322 ( .A(n4733), .B(p_input[3468]), .Z(n4732) );
  AND U5323 ( .A(p_input[2468]), .B(p_input[1468]), .Z(n4733) );
  AND U5324 ( .A(p_input[468]), .B(p_input[4468]), .Z(n4731) );
  AND U5325 ( .A(n4734), .B(n4735), .Z(n4729) );
  AND U5326 ( .A(n4736), .B(p_input[7468]), .Z(n4735) );
  AND U5327 ( .A(p_input[6468]), .B(p_input[5468]), .Z(n4736) );
  AND U5328 ( .A(p_input[9468]), .B(p_input[8468]), .Z(n4734) );
  AND U5329 ( .A(n4737), .B(n4738), .Z(o[467]) );
  AND U5330 ( .A(n4739), .B(n4740), .Z(n4738) );
  AND U5331 ( .A(n4741), .B(p_input[3467]), .Z(n4740) );
  AND U5332 ( .A(p_input[2467]), .B(p_input[1467]), .Z(n4741) );
  AND U5333 ( .A(p_input[467]), .B(p_input[4467]), .Z(n4739) );
  AND U5334 ( .A(n4742), .B(n4743), .Z(n4737) );
  AND U5335 ( .A(n4744), .B(p_input[7467]), .Z(n4743) );
  AND U5336 ( .A(p_input[6467]), .B(p_input[5467]), .Z(n4744) );
  AND U5337 ( .A(p_input[9467]), .B(p_input[8467]), .Z(n4742) );
  AND U5338 ( .A(n4745), .B(n4746), .Z(o[466]) );
  AND U5339 ( .A(n4747), .B(n4748), .Z(n4746) );
  AND U5340 ( .A(n4749), .B(p_input[3466]), .Z(n4748) );
  AND U5341 ( .A(p_input[2466]), .B(p_input[1466]), .Z(n4749) );
  AND U5342 ( .A(p_input[466]), .B(p_input[4466]), .Z(n4747) );
  AND U5343 ( .A(n4750), .B(n4751), .Z(n4745) );
  AND U5344 ( .A(n4752), .B(p_input[7466]), .Z(n4751) );
  AND U5345 ( .A(p_input[6466]), .B(p_input[5466]), .Z(n4752) );
  AND U5346 ( .A(p_input[9466]), .B(p_input[8466]), .Z(n4750) );
  AND U5347 ( .A(n4753), .B(n4754), .Z(o[465]) );
  AND U5348 ( .A(n4755), .B(n4756), .Z(n4754) );
  AND U5349 ( .A(n4757), .B(p_input[3465]), .Z(n4756) );
  AND U5350 ( .A(p_input[2465]), .B(p_input[1465]), .Z(n4757) );
  AND U5351 ( .A(p_input[465]), .B(p_input[4465]), .Z(n4755) );
  AND U5352 ( .A(n4758), .B(n4759), .Z(n4753) );
  AND U5353 ( .A(n4760), .B(p_input[7465]), .Z(n4759) );
  AND U5354 ( .A(p_input[6465]), .B(p_input[5465]), .Z(n4760) );
  AND U5355 ( .A(p_input[9465]), .B(p_input[8465]), .Z(n4758) );
  AND U5356 ( .A(n4761), .B(n4762), .Z(o[464]) );
  AND U5357 ( .A(n4763), .B(n4764), .Z(n4762) );
  AND U5358 ( .A(n4765), .B(p_input[3464]), .Z(n4764) );
  AND U5359 ( .A(p_input[2464]), .B(p_input[1464]), .Z(n4765) );
  AND U5360 ( .A(p_input[464]), .B(p_input[4464]), .Z(n4763) );
  AND U5361 ( .A(n4766), .B(n4767), .Z(n4761) );
  AND U5362 ( .A(n4768), .B(p_input[7464]), .Z(n4767) );
  AND U5363 ( .A(p_input[6464]), .B(p_input[5464]), .Z(n4768) );
  AND U5364 ( .A(p_input[9464]), .B(p_input[8464]), .Z(n4766) );
  AND U5365 ( .A(n4769), .B(n4770), .Z(o[463]) );
  AND U5366 ( .A(n4771), .B(n4772), .Z(n4770) );
  AND U5367 ( .A(n4773), .B(p_input[3463]), .Z(n4772) );
  AND U5368 ( .A(p_input[2463]), .B(p_input[1463]), .Z(n4773) );
  AND U5369 ( .A(p_input[463]), .B(p_input[4463]), .Z(n4771) );
  AND U5370 ( .A(n4774), .B(n4775), .Z(n4769) );
  AND U5371 ( .A(n4776), .B(p_input[7463]), .Z(n4775) );
  AND U5372 ( .A(p_input[6463]), .B(p_input[5463]), .Z(n4776) );
  AND U5373 ( .A(p_input[9463]), .B(p_input[8463]), .Z(n4774) );
  AND U5374 ( .A(n4777), .B(n4778), .Z(o[462]) );
  AND U5375 ( .A(n4779), .B(n4780), .Z(n4778) );
  AND U5376 ( .A(n4781), .B(p_input[3462]), .Z(n4780) );
  AND U5377 ( .A(p_input[2462]), .B(p_input[1462]), .Z(n4781) );
  AND U5378 ( .A(p_input[462]), .B(p_input[4462]), .Z(n4779) );
  AND U5379 ( .A(n4782), .B(n4783), .Z(n4777) );
  AND U5380 ( .A(n4784), .B(p_input[7462]), .Z(n4783) );
  AND U5381 ( .A(p_input[6462]), .B(p_input[5462]), .Z(n4784) );
  AND U5382 ( .A(p_input[9462]), .B(p_input[8462]), .Z(n4782) );
  AND U5383 ( .A(n4785), .B(n4786), .Z(o[461]) );
  AND U5384 ( .A(n4787), .B(n4788), .Z(n4786) );
  AND U5385 ( .A(n4789), .B(p_input[3461]), .Z(n4788) );
  AND U5386 ( .A(p_input[2461]), .B(p_input[1461]), .Z(n4789) );
  AND U5387 ( .A(p_input[461]), .B(p_input[4461]), .Z(n4787) );
  AND U5388 ( .A(n4790), .B(n4791), .Z(n4785) );
  AND U5389 ( .A(n4792), .B(p_input[7461]), .Z(n4791) );
  AND U5390 ( .A(p_input[6461]), .B(p_input[5461]), .Z(n4792) );
  AND U5391 ( .A(p_input[9461]), .B(p_input[8461]), .Z(n4790) );
  AND U5392 ( .A(n4793), .B(n4794), .Z(o[460]) );
  AND U5393 ( .A(n4795), .B(n4796), .Z(n4794) );
  AND U5394 ( .A(n4797), .B(p_input[3460]), .Z(n4796) );
  AND U5395 ( .A(p_input[2460]), .B(p_input[1460]), .Z(n4797) );
  AND U5396 ( .A(p_input[460]), .B(p_input[4460]), .Z(n4795) );
  AND U5397 ( .A(n4798), .B(n4799), .Z(n4793) );
  AND U5398 ( .A(n4800), .B(p_input[7460]), .Z(n4799) );
  AND U5399 ( .A(p_input[6460]), .B(p_input[5460]), .Z(n4800) );
  AND U5400 ( .A(p_input[9460]), .B(p_input[8460]), .Z(n4798) );
  AND U5401 ( .A(n4801), .B(n4802), .Z(o[45]) );
  AND U5402 ( .A(n4803), .B(n4804), .Z(n4802) );
  AND U5403 ( .A(n4805), .B(p_input[3045]), .Z(n4804) );
  AND U5404 ( .A(p_input[2045]), .B(p_input[1045]), .Z(n4805) );
  AND U5405 ( .A(p_input[45]), .B(p_input[4045]), .Z(n4803) );
  AND U5406 ( .A(n4806), .B(n4807), .Z(n4801) );
  AND U5407 ( .A(n4808), .B(p_input[7045]), .Z(n4807) );
  AND U5408 ( .A(p_input[6045]), .B(p_input[5045]), .Z(n4808) );
  AND U5409 ( .A(p_input[9045]), .B(p_input[8045]), .Z(n4806) );
  AND U5410 ( .A(n4809), .B(n4810), .Z(o[459]) );
  AND U5411 ( .A(n4811), .B(n4812), .Z(n4810) );
  AND U5412 ( .A(n4813), .B(p_input[3459]), .Z(n4812) );
  AND U5413 ( .A(p_input[2459]), .B(p_input[1459]), .Z(n4813) );
  AND U5414 ( .A(p_input[459]), .B(p_input[4459]), .Z(n4811) );
  AND U5415 ( .A(n4814), .B(n4815), .Z(n4809) );
  AND U5416 ( .A(n4816), .B(p_input[7459]), .Z(n4815) );
  AND U5417 ( .A(p_input[6459]), .B(p_input[5459]), .Z(n4816) );
  AND U5418 ( .A(p_input[9459]), .B(p_input[8459]), .Z(n4814) );
  AND U5419 ( .A(n4817), .B(n4818), .Z(o[458]) );
  AND U5420 ( .A(n4819), .B(n4820), .Z(n4818) );
  AND U5421 ( .A(n4821), .B(p_input[3458]), .Z(n4820) );
  AND U5422 ( .A(p_input[2458]), .B(p_input[1458]), .Z(n4821) );
  AND U5423 ( .A(p_input[458]), .B(p_input[4458]), .Z(n4819) );
  AND U5424 ( .A(n4822), .B(n4823), .Z(n4817) );
  AND U5425 ( .A(n4824), .B(p_input[7458]), .Z(n4823) );
  AND U5426 ( .A(p_input[6458]), .B(p_input[5458]), .Z(n4824) );
  AND U5427 ( .A(p_input[9458]), .B(p_input[8458]), .Z(n4822) );
  AND U5428 ( .A(n4825), .B(n4826), .Z(o[457]) );
  AND U5429 ( .A(n4827), .B(n4828), .Z(n4826) );
  AND U5430 ( .A(n4829), .B(p_input[3457]), .Z(n4828) );
  AND U5431 ( .A(p_input[2457]), .B(p_input[1457]), .Z(n4829) );
  AND U5432 ( .A(p_input[457]), .B(p_input[4457]), .Z(n4827) );
  AND U5433 ( .A(n4830), .B(n4831), .Z(n4825) );
  AND U5434 ( .A(n4832), .B(p_input[7457]), .Z(n4831) );
  AND U5435 ( .A(p_input[6457]), .B(p_input[5457]), .Z(n4832) );
  AND U5436 ( .A(p_input[9457]), .B(p_input[8457]), .Z(n4830) );
  AND U5437 ( .A(n4833), .B(n4834), .Z(o[456]) );
  AND U5438 ( .A(n4835), .B(n4836), .Z(n4834) );
  AND U5439 ( .A(n4837), .B(p_input[3456]), .Z(n4836) );
  AND U5440 ( .A(p_input[2456]), .B(p_input[1456]), .Z(n4837) );
  AND U5441 ( .A(p_input[456]), .B(p_input[4456]), .Z(n4835) );
  AND U5442 ( .A(n4838), .B(n4839), .Z(n4833) );
  AND U5443 ( .A(n4840), .B(p_input[7456]), .Z(n4839) );
  AND U5444 ( .A(p_input[6456]), .B(p_input[5456]), .Z(n4840) );
  AND U5445 ( .A(p_input[9456]), .B(p_input[8456]), .Z(n4838) );
  AND U5446 ( .A(n4841), .B(n4842), .Z(o[455]) );
  AND U5447 ( .A(n4843), .B(n4844), .Z(n4842) );
  AND U5448 ( .A(n4845), .B(p_input[3455]), .Z(n4844) );
  AND U5449 ( .A(p_input[2455]), .B(p_input[1455]), .Z(n4845) );
  AND U5450 ( .A(p_input[455]), .B(p_input[4455]), .Z(n4843) );
  AND U5451 ( .A(n4846), .B(n4847), .Z(n4841) );
  AND U5452 ( .A(n4848), .B(p_input[7455]), .Z(n4847) );
  AND U5453 ( .A(p_input[6455]), .B(p_input[5455]), .Z(n4848) );
  AND U5454 ( .A(p_input[9455]), .B(p_input[8455]), .Z(n4846) );
  AND U5455 ( .A(n4849), .B(n4850), .Z(o[454]) );
  AND U5456 ( .A(n4851), .B(n4852), .Z(n4850) );
  AND U5457 ( .A(n4853), .B(p_input[3454]), .Z(n4852) );
  AND U5458 ( .A(p_input[2454]), .B(p_input[1454]), .Z(n4853) );
  AND U5459 ( .A(p_input[454]), .B(p_input[4454]), .Z(n4851) );
  AND U5460 ( .A(n4854), .B(n4855), .Z(n4849) );
  AND U5461 ( .A(n4856), .B(p_input[7454]), .Z(n4855) );
  AND U5462 ( .A(p_input[6454]), .B(p_input[5454]), .Z(n4856) );
  AND U5463 ( .A(p_input[9454]), .B(p_input[8454]), .Z(n4854) );
  AND U5464 ( .A(n4857), .B(n4858), .Z(o[453]) );
  AND U5465 ( .A(n4859), .B(n4860), .Z(n4858) );
  AND U5466 ( .A(n4861), .B(p_input[3453]), .Z(n4860) );
  AND U5467 ( .A(p_input[2453]), .B(p_input[1453]), .Z(n4861) );
  AND U5468 ( .A(p_input[453]), .B(p_input[4453]), .Z(n4859) );
  AND U5469 ( .A(n4862), .B(n4863), .Z(n4857) );
  AND U5470 ( .A(n4864), .B(p_input[7453]), .Z(n4863) );
  AND U5471 ( .A(p_input[6453]), .B(p_input[5453]), .Z(n4864) );
  AND U5472 ( .A(p_input[9453]), .B(p_input[8453]), .Z(n4862) );
  AND U5473 ( .A(n4865), .B(n4866), .Z(o[452]) );
  AND U5474 ( .A(n4867), .B(n4868), .Z(n4866) );
  AND U5475 ( .A(n4869), .B(p_input[3452]), .Z(n4868) );
  AND U5476 ( .A(p_input[2452]), .B(p_input[1452]), .Z(n4869) );
  AND U5477 ( .A(p_input[452]), .B(p_input[4452]), .Z(n4867) );
  AND U5478 ( .A(n4870), .B(n4871), .Z(n4865) );
  AND U5479 ( .A(n4872), .B(p_input[7452]), .Z(n4871) );
  AND U5480 ( .A(p_input[6452]), .B(p_input[5452]), .Z(n4872) );
  AND U5481 ( .A(p_input[9452]), .B(p_input[8452]), .Z(n4870) );
  AND U5482 ( .A(n4873), .B(n4874), .Z(o[451]) );
  AND U5483 ( .A(n4875), .B(n4876), .Z(n4874) );
  AND U5484 ( .A(n4877), .B(p_input[3451]), .Z(n4876) );
  AND U5485 ( .A(p_input[2451]), .B(p_input[1451]), .Z(n4877) );
  AND U5486 ( .A(p_input[451]), .B(p_input[4451]), .Z(n4875) );
  AND U5487 ( .A(n4878), .B(n4879), .Z(n4873) );
  AND U5488 ( .A(n4880), .B(p_input[7451]), .Z(n4879) );
  AND U5489 ( .A(p_input[6451]), .B(p_input[5451]), .Z(n4880) );
  AND U5490 ( .A(p_input[9451]), .B(p_input[8451]), .Z(n4878) );
  AND U5491 ( .A(n4881), .B(n4882), .Z(o[450]) );
  AND U5492 ( .A(n4883), .B(n4884), .Z(n4882) );
  AND U5493 ( .A(n4885), .B(p_input[3450]), .Z(n4884) );
  AND U5494 ( .A(p_input[2450]), .B(p_input[1450]), .Z(n4885) );
  AND U5495 ( .A(p_input[450]), .B(p_input[4450]), .Z(n4883) );
  AND U5496 ( .A(n4886), .B(n4887), .Z(n4881) );
  AND U5497 ( .A(n4888), .B(p_input[7450]), .Z(n4887) );
  AND U5498 ( .A(p_input[6450]), .B(p_input[5450]), .Z(n4888) );
  AND U5499 ( .A(p_input[9450]), .B(p_input[8450]), .Z(n4886) );
  AND U5500 ( .A(n4889), .B(n4890), .Z(o[44]) );
  AND U5501 ( .A(n4891), .B(n4892), .Z(n4890) );
  AND U5502 ( .A(n4893), .B(p_input[3044]), .Z(n4892) );
  AND U5503 ( .A(p_input[2044]), .B(p_input[1044]), .Z(n4893) );
  AND U5504 ( .A(p_input[44]), .B(p_input[4044]), .Z(n4891) );
  AND U5505 ( .A(n4894), .B(n4895), .Z(n4889) );
  AND U5506 ( .A(n4896), .B(p_input[7044]), .Z(n4895) );
  AND U5507 ( .A(p_input[6044]), .B(p_input[5044]), .Z(n4896) );
  AND U5508 ( .A(p_input[9044]), .B(p_input[8044]), .Z(n4894) );
  AND U5509 ( .A(n4897), .B(n4898), .Z(o[449]) );
  AND U5510 ( .A(n4899), .B(n4900), .Z(n4898) );
  AND U5511 ( .A(n4901), .B(p_input[3449]), .Z(n4900) );
  AND U5512 ( .A(p_input[2449]), .B(p_input[1449]), .Z(n4901) );
  AND U5513 ( .A(p_input[449]), .B(p_input[4449]), .Z(n4899) );
  AND U5514 ( .A(n4902), .B(n4903), .Z(n4897) );
  AND U5515 ( .A(n4904), .B(p_input[7449]), .Z(n4903) );
  AND U5516 ( .A(p_input[6449]), .B(p_input[5449]), .Z(n4904) );
  AND U5517 ( .A(p_input[9449]), .B(p_input[8449]), .Z(n4902) );
  AND U5518 ( .A(n4905), .B(n4906), .Z(o[448]) );
  AND U5519 ( .A(n4907), .B(n4908), .Z(n4906) );
  AND U5520 ( .A(n4909), .B(p_input[3448]), .Z(n4908) );
  AND U5521 ( .A(p_input[2448]), .B(p_input[1448]), .Z(n4909) );
  AND U5522 ( .A(p_input[448]), .B(p_input[4448]), .Z(n4907) );
  AND U5523 ( .A(n4910), .B(n4911), .Z(n4905) );
  AND U5524 ( .A(n4912), .B(p_input[7448]), .Z(n4911) );
  AND U5525 ( .A(p_input[6448]), .B(p_input[5448]), .Z(n4912) );
  AND U5526 ( .A(p_input[9448]), .B(p_input[8448]), .Z(n4910) );
  AND U5527 ( .A(n4913), .B(n4914), .Z(o[447]) );
  AND U5528 ( .A(n4915), .B(n4916), .Z(n4914) );
  AND U5529 ( .A(n4917), .B(p_input[3447]), .Z(n4916) );
  AND U5530 ( .A(p_input[2447]), .B(p_input[1447]), .Z(n4917) );
  AND U5531 ( .A(p_input[447]), .B(p_input[4447]), .Z(n4915) );
  AND U5532 ( .A(n4918), .B(n4919), .Z(n4913) );
  AND U5533 ( .A(n4920), .B(p_input[7447]), .Z(n4919) );
  AND U5534 ( .A(p_input[6447]), .B(p_input[5447]), .Z(n4920) );
  AND U5535 ( .A(p_input[9447]), .B(p_input[8447]), .Z(n4918) );
  AND U5536 ( .A(n4921), .B(n4922), .Z(o[446]) );
  AND U5537 ( .A(n4923), .B(n4924), .Z(n4922) );
  AND U5538 ( .A(n4925), .B(p_input[3446]), .Z(n4924) );
  AND U5539 ( .A(p_input[2446]), .B(p_input[1446]), .Z(n4925) );
  AND U5540 ( .A(p_input[446]), .B(p_input[4446]), .Z(n4923) );
  AND U5541 ( .A(n4926), .B(n4927), .Z(n4921) );
  AND U5542 ( .A(n4928), .B(p_input[7446]), .Z(n4927) );
  AND U5543 ( .A(p_input[6446]), .B(p_input[5446]), .Z(n4928) );
  AND U5544 ( .A(p_input[9446]), .B(p_input[8446]), .Z(n4926) );
  AND U5545 ( .A(n4929), .B(n4930), .Z(o[445]) );
  AND U5546 ( .A(n4931), .B(n4932), .Z(n4930) );
  AND U5547 ( .A(n4933), .B(p_input[3445]), .Z(n4932) );
  AND U5548 ( .A(p_input[2445]), .B(p_input[1445]), .Z(n4933) );
  AND U5549 ( .A(p_input[445]), .B(p_input[4445]), .Z(n4931) );
  AND U5550 ( .A(n4934), .B(n4935), .Z(n4929) );
  AND U5551 ( .A(n4936), .B(p_input[7445]), .Z(n4935) );
  AND U5552 ( .A(p_input[6445]), .B(p_input[5445]), .Z(n4936) );
  AND U5553 ( .A(p_input[9445]), .B(p_input[8445]), .Z(n4934) );
  AND U5554 ( .A(n4937), .B(n4938), .Z(o[444]) );
  AND U5555 ( .A(n4939), .B(n4940), .Z(n4938) );
  AND U5556 ( .A(n4941), .B(p_input[3444]), .Z(n4940) );
  AND U5557 ( .A(p_input[2444]), .B(p_input[1444]), .Z(n4941) );
  AND U5558 ( .A(p_input[444]), .B(p_input[4444]), .Z(n4939) );
  AND U5559 ( .A(n4942), .B(n4943), .Z(n4937) );
  AND U5560 ( .A(n4944), .B(p_input[7444]), .Z(n4943) );
  AND U5561 ( .A(p_input[6444]), .B(p_input[5444]), .Z(n4944) );
  AND U5562 ( .A(p_input[9444]), .B(p_input[8444]), .Z(n4942) );
  AND U5563 ( .A(n4945), .B(n4946), .Z(o[443]) );
  AND U5564 ( .A(n4947), .B(n4948), .Z(n4946) );
  AND U5565 ( .A(n4949), .B(p_input[3443]), .Z(n4948) );
  AND U5566 ( .A(p_input[2443]), .B(p_input[1443]), .Z(n4949) );
  AND U5567 ( .A(p_input[4443]), .B(p_input[443]), .Z(n4947) );
  AND U5568 ( .A(n4950), .B(n4951), .Z(n4945) );
  AND U5569 ( .A(n4952), .B(p_input[7443]), .Z(n4951) );
  AND U5570 ( .A(p_input[6443]), .B(p_input[5443]), .Z(n4952) );
  AND U5571 ( .A(p_input[9443]), .B(p_input[8443]), .Z(n4950) );
  AND U5572 ( .A(n4953), .B(n4954), .Z(o[442]) );
  AND U5573 ( .A(n4955), .B(n4956), .Z(n4954) );
  AND U5574 ( .A(n4957), .B(p_input[3442]), .Z(n4956) );
  AND U5575 ( .A(p_input[2442]), .B(p_input[1442]), .Z(n4957) );
  AND U5576 ( .A(p_input[4442]), .B(p_input[442]), .Z(n4955) );
  AND U5577 ( .A(n4958), .B(n4959), .Z(n4953) );
  AND U5578 ( .A(n4960), .B(p_input[7442]), .Z(n4959) );
  AND U5579 ( .A(p_input[6442]), .B(p_input[5442]), .Z(n4960) );
  AND U5580 ( .A(p_input[9442]), .B(p_input[8442]), .Z(n4958) );
  AND U5581 ( .A(n4961), .B(n4962), .Z(o[441]) );
  AND U5582 ( .A(n4963), .B(n4964), .Z(n4962) );
  AND U5583 ( .A(n4965), .B(p_input[3441]), .Z(n4964) );
  AND U5584 ( .A(p_input[2441]), .B(p_input[1441]), .Z(n4965) );
  AND U5585 ( .A(p_input[4441]), .B(p_input[441]), .Z(n4963) );
  AND U5586 ( .A(n4966), .B(n4967), .Z(n4961) );
  AND U5587 ( .A(n4968), .B(p_input[7441]), .Z(n4967) );
  AND U5588 ( .A(p_input[6441]), .B(p_input[5441]), .Z(n4968) );
  AND U5589 ( .A(p_input[9441]), .B(p_input[8441]), .Z(n4966) );
  AND U5590 ( .A(n4969), .B(n4970), .Z(o[440]) );
  AND U5591 ( .A(n4971), .B(n4972), .Z(n4970) );
  AND U5592 ( .A(n4973), .B(p_input[3440]), .Z(n4972) );
  AND U5593 ( .A(p_input[2440]), .B(p_input[1440]), .Z(n4973) );
  AND U5594 ( .A(p_input[4440]), .B(p_input[440]), .Z(n4971) );
  AND U5595 ( .A(n4974), .B(n4975), .Z(n4969) );
  AND U5596 ( .A(n4976), .B(p_input[7440]), .Z(n4975) );
  AND U5597 ( .A(p_input[6440]), .B(p_input[5440]), .Z(n4976) );
  AND U5598 ( .A(p_input[9440]), .B(p_input[8440]), .Z(n4974) );
  AND U5599 ( .A(n4977), .B(n4978), .Z(o[43]) );
  AND U5600 ( .A(n4979), .B(n4980), .Z(n4978) );
  AND U5601 ( .A(n4981), .B(p_input[3043]), .Z(n4980) );
  AND U5602 ( .A(p_input[2043]), .B(p_input[1043]), .Z(n4981) );
  AND U5603 ( .A(p_input[43]), .B(p_input[4043]), .Z(n4979) );
  AND U5604 ( .A(n4982), .B(n4983), .Z(n4977) );
  AND U5605 ( .A(n4984), .B(p_input[7043]), .Z(n4983) );
  AND U5606 ( .A(p_input[6043]), .B(p_input[5043]), .Z(n4984) );
  AND U5607 ( .A(p_input[9043]), .B(p_input[8043]), .Z(n4982) );
  AND U5608 ( .A(n4985), .B(n4986), .Z(o[439]) );
  AND U5609 ( .A(n4987), .B(n4988), .Z(n4986) );
  AND U5610 ( .A(n4989), .B(p_input[3439]), .Z(n4988) );
  AND U5611 ( .A(p_input[2439]), .B(p_input[1439]), .Z(n4989) );
  AND U5612 ( .A(p_input[4439]), .B(p_input[439]), .Z(n4987) );
  AND U5613 ( .A(n4990), .B(n4991), .Z(n4985) );
  AND U5614 ( .A(n4992), .B(p_input[7439]), .Z(n4991) );
  AND U5615 ( .A(p_input[6439]), .B(p_input[5439]), .Z(n4992) );
  AND U5616 ( .A(p_input[9439]), .B(p_input[8439]), .Z(n4990) );
  AND U5617 ( .A(n4993), .B(n4994), .Z(o[438]) );
  AND U5618 ( .A(n4995), .B(n4996), .Z(n4994) );
  AND U5619 ( .A(n4997), .B(p_input[3438]), .Z(n4996) );
  AND U5620 ( .A(p_input[2438]), .B(p_input[1438]), .Z(n4997) );
  AND U5621 ( .A(p_input[4438]), .B(p_input[438]), .Z(n4995) );
  AND U5622 ( .A(n4998), .B(n4999), .Z(n4993) );
  AND U5623 ( .A(n5000), .B(p_input[7438]), .Z(n4999) );
  AND U5624 ( .A(p_input[6438]), .B(p_input[5438]), .Z(n5000) );
  AND U5625 ( .A(p_input[9438]), .B(p_input[8438]), .Z(n4998) );
  AND U5626 ( .A(n5001), .B(n5002), .Z(o[437]) );
  AND U5627 ( .A(n5003), .B(n5004), .Z(n5002) );
  AND U5628 ( .A(n5005), .B(p_input[3437]), .Z(n5004) );
  AND U5629 ( .A(p_input[2437]), .B(p_input[1437]), .Z(n5005) );
  AND U5630 ( .A(p_input[4437]), .B(p_input[437]), .Z(n5003) );
  AND U5631 ( .A(n5006), .B(n5007), .Z(n5001) );
  AND U5632 ( .A(n5008), .B(p_input[7437]), .Z(n5007) );
  AND U5633 ( .A(p_input[6437]), .B(p_input[5437]), .Z(n5008) );
  AND U5634 ( .A(p_input[9437]), .B(p_input[8437]), .Z(n5006) );
  AND U5635 ( .A(n5009), .B(n5010), .Z(o[436]) );
  AND U5636 ( .A(n5011), .B(n5012), .Z(n5010) );
  AND U5637 ( .A(n5013), .B(p_input[3436]), .Z(n5012) );
  AND U5638 ( .A(p_input[2436]), .B(p_input[1436]), .Z(n5013) );
  AND U5639 ( .A(p_input[4436]), .B(p_input[436]), .Z(n5011) );
  AND U5640 ( .A(n5014), .B(n5015), .Z(n5009) );
  AND U5641 ( .A(n5016), .B(p_input[7436]), .Z(n5015) );
  AND U5642 ( .A(p_input[6436]), .B(p_input[5436]), .Z(n5016) );
  AND U5643 ( .A(p_input[9436]), .B(p_input[8436]), .Z(n5014) );
  AND U5644 ( .A(n5017), .B(n5018), .Z(o[435]) );
  AND U5645 ( .A(n5019), .B(n5020), .Z(n5018) );
  AND U5646 ( .A(n5021), .B(p_input[3435]), .Z(n5020) );
  AND U5647 ( .A(p_input[2435]), .B(p_input[1435]), .Z(n5021) );
  AND U5648 ( .A(p_input[4435]), .B(p_input[435]), .Z(n5019) );
  AND U5649 ( .A(n5022), .B(n5023), .Z(n5017) );
  AND U5650 ( .A(n5024), .B(p_input[7435]), .Z(n5023) );
  AND U5651 ( .A(p_input[6435]), .B(p_input[5435]), .Z(n5024) );
  AND U5652 ( .A(p_input[9435]), .B(p_input[8435]), .Z(n5022) );
  AND U5653 ( .A(n5025), .B(n5026), .Z(o[434]) );
  AND U5654 ( .A(n5027), .B(n5028), .Z(n5026) );
  AND U5655 ( .A(n5029), .B(p_input[3434]), .Z(n5028) );
  AND U5656 ( .A(p_input[2434]), .B(p_input[1434]), .Z(n5029) );
  AND U5657 ( .A(p_input[4434]), .B(p_input[434]), .Z(n5027) );
  AND U5658 ( .A(n5030), .B(n5031), .Z(n5025) );
  AND U5659 ( .A(n5032), .B(p_input[7434]), .Z(n5031) );
  AND U5660 ( .A(p_input[6434]), .B(p_input[5434]), .Z(n5032) );
  AND U5661 ( .A(p_input[9434]), .B(p_input[8434]), .Z(n5030) );
  AND U5662 ( .A(n5033), .B(n5034), .Z(o[433]) );
  AND U5663 ( .A(n5035), .B(n5036), .Z(n5034) );
  AND U5664 ( .A(n5037), .B(p_input[3433]), .Z(n5036) );
  AND U5665 ( .A(p_input[2433]), .B(p_input[1433]), .Z(n5037) );
  AND U5666 ( .A(p_input[4433]), .B(p_input[433]), .Z(n5035) );
  AND U5667 ( .A(n5038), .B(n5039), .Z(n5033) );
  AND U5668 ( .A(n5040), .B(p_input[7433]), .Z(n5039) );
  AND U5669 ( .A(p_input[6433]), .B(p_input[5433]), .Z(n5040) );
  AND U5670 ( .A(p_input[9433]), .B(p_input[8433]), .Z(n5038) );
  AND U5671 ( .A(n5041), .B(n5042), .Z(o[432]) );
  AND U5672 ( .A(n5043), .B(n5044), .Z(n5042) );
  AND U5673 ( .A(n5045), .B(p_input[3432]), .Z(n5044) );
  AND U5674 ( .A(p_input[2432]), .B(p_input[1432]), .Z(n5045) );
  AND U5675 ( .A(p_input[4432]), .B(p_input[432]), .Z(n5043) );
  AND U5676 ( .A(n5046), .B(n5047), .Z(n5041) );
  AND U5677 ( .A(n5048), .B(p_input[7432]), .Z(n5047) );
  AND U5678 ( .A(p_input[6432]), .B(p_input[5432]), .Z(n5048) );
  AND U5679 ( .A(p_input[9432]), .B(p_input[8432]), .Z(n5046) );
  AND U5680 ( .A(n5049), .B(n5050), .Z(o[431]) );
  AND U5681 ( .A(n5051), .B(n5052), .Z(n5050) );
  AND U5682 ( .A(n5053), .B(p_input[3431]), .Z(n5052) );
  AND U5683 ( .A(p_input[2431]), .B(p_input[1431]), .Z(n5053) );
  AND U5684 ( .A(p_input[4431]), .B(p_input[431]), .Z(n5051) );
  AND U5685 ( .A(n5054), .B(n5055), .Z(n5049) );
  AND U5686 ( .A(n5056), .B(p_input[7431]), .Z(n5055) );
  AND U5687 ( .A(p_input[6431]), .B(p_input[5431]), .Z(n5056) );
  AND U5688 ( .A(p_input[9431]), .B(p_input[8431]), .Z(n5054) );
  AND U5689 ( .A(n5057), .B(n5058), .Z(o[430]) );
  AND U5690 ( .A(n5059), .B(n5060), .Z(n5058) );
  AND U5691 ( .A(n5061), .B(p_input[3430]), .Z(n5060) );
  AND U5692 ( .A(p_input[2430]), .B(p_input[1430]), .Z(n5061) );
  AND U5693 ( .A(p_input[4430]), .B(p_input[430]), .Z(n5059) );
  AND U5694 ( .A(n5062), .B(n5063), .Z(n5057) );
  AND U5695 ( .A(n5064), .B(p_input[7430]), .Z(n5063) );
  AND U5696 ( .A(p_input[6430]), .B(p_input[5430]), .Z(n5064) );
  AND U5697 ( .A(p_input[9430]), .B(p_input[8430]), .Z(n5062) );
  AND U5698 ( .A(n5065), .B(n5066), .Z(o[42]) );
  AND U5699 ( .A(n5067), .B(n5068), .Z(n5066) );
  AND U5700 ( .A(n5069), .B(p_input[3042]), .Z(n5068) );
  AND U5701 ( .A(p_input[2042]), .B(p_input[1042]), .Z(n5069) );
  AND U5702 ( .A(p_input[42]), .B(p_input[4042]), .Z(n5067) );
  AND U5703 ( .A(n5070), .B(n5071), .Z(n5065) );
  AND U5704 ( .A(n5072), .B(p_input[7042]), .Z(n5071) );
  AND U5705 ( .A(p_input[6042]), .B(p_input[5042]), .Z(n5072) );
  AND U5706 ( .A(p_input[9042]), .B(p_input[8042]), .Z(n5070) );
  AND U5707 ( .A(n5073), .B(n5074), .Z(o[429]) );
  AND U5708 ( .A(n5075), .B(n5076), .Z(n5074) );
  AND U5709 ( .A(n5077), .B(p_input[3429]), .Z(n5076) );
  AND U5710 ( .A(p_input[2429]), .B(p_input[1429]), .Z(n5077) );
  AND U5711 ( .A(p_input[4429]), .B(p_input[429]), .Z(n5075) );
  AND U5712 ( .A(n5078), .B(n5079), .Z(n5073) );
  AND U5713 ( .A(n5080), .B(p_input[7429]), .Z(n5079) );
  AND U5714 ( .A(p_input[6429]), .B(p_input[5429]), .Z(n5080) );
  AND U5715 ( .A(p_input[9429]), .B(p_input[8429]), .Z(n5078) );
  AND U5716 ( .A(n5081), .B(n5082), .Z(o[428]) );
  AND U5717 ( .A(n5083), .B(n5084), .Z(n5082) );
  AND U5718 ( .A(n5085), .B(p_input[3428]), .Z(n5084) );
  AND U5719 ( .A(p_input[2428]), .B(p_input[1428]), .Z(n5085) );
  AND U5720 ( .A(p_input[4428]), .B(p_input[428]), .Z(n5083) );
  AND U5721 ( .A(n5086), .B(n5087), .Z(n5081) );
  AND U5722 ( .A(n5088), .B(p_input[7428]), .Z(n5087) );
  AND U5723 ( .A(p_input[6428]), .B(p_input[5428]), .Z(n5088) );
  AND U5724 ( .A(p_input[9428]), .B(p_input[8428]), .Z(n5086) );
  AND U5725 ( .A(n5089), .B(n5090), .Z(o[427]) );
  AND U5726 ( .A(n5091), .B(n5092), .Z(n5090) );
  AND U5727 ( .A(n5093), .B(p_input[3427]), .Z(n5092) );
  AND U5728 ( .A(p_input[2427]), .B(p_input[1427]), .Z(n5093) );
  AND U5729 ( .A(p_input[4427]), .B(p_input[427]), .Z(n5091) );
  AND U5730 ( .A(n5094), .B(n5095), .Z(n5089) );
  AND U5731 ( .A(n5096), .B(p_input[7427]), .Z(n5095) );
  AND U5732 ( .A(p_input[6427]), .B(p_input[5427]), .Z(n5096) );
  AND U5733 ( .A(p_input[9427]), .B(p_input[8427]), .Z(n5094) );
  AND U5734 ( .A(n5097), .B(n5098), .Z(o[426]) );
  AND U5735 ( .A(n5099), .B(n5100), .Z(n5098) );
  AND U5736 ( .A(n5101), .B(p_input[3426]), .Z(n5100) );
  AND U5737 ( .A(p_input[2426]), .B(p_input[1426]), .Z(n5101) );
  AND U5738 ( .A(p_input[4426]), .B(p_input[426]), .Z(n5099) );
  AND U5739 ( .A(n5102), .B(n5103), .Z(n5097) );
  AND U5740 ( .A(n5104), .B(p_input[7426]), .Z(n5103) );
  AND U5741 ( .A(p_input[6426]), .B(p_input[5426]), .Z(n5104) );
  AND U5742 ( .A(p_input[9426]), .B(p_input[8426]), .Z(n5102) );
  AND U5743 ( .A(n5105), .B(n5106), .Z(o[425]) );
  AND U5744 ( .A(n5107), .B(n5108), .Z(n5106) );
  AND U5745 ( .A(n5109), .B(p_input[3425]), .Z(n5108) );
  AND U5746 ( .A(p_input[2425]), .B(p_input[1425]), .Z(n5109) );
  AND U5747 ( .A(p_input[4425]), .B(p_input[425]), .Z(n5107) );
  AND U5748 ( .A(n5110), .B(n5111), .Z(n5105) );
  AND U5749 ( .A(n5112), .B(p_input[7425]), .Z(n5111) );
  AND U5750 ( .A(p_input[6425]), .B(p_input[5425]), .Z(n5112) );
  AND U5751 ( .A(p_input[9425]), .B(p_input[8425]), .Z(n5110) );
  AND U5752 ( .A(n5113), .B(n5114), .Z(o[424]) );
  AND U5753 ( .A(n5115), .B(n5116), .Z(n5114) );
  AND U5754 ( .A(n5117), .B(p_input[3424]), .Z(n5116) );
  AND U5755 ( .A(p_input[2424]), .B(p_input[1424]), .Z(n5117) );
  AND U5756 ( .A(p_input[4424]), .B(p_input[424]), .Z(n5115) );
  AND U5757 ( .A(n5118), .B(n5119), .Z(n5113) );
  AND U5758 ( .A(n5120), .B(p_input[7424]), .Z(n5119) );
  AND U5759 ( .A(p_input[6424]), .B(p_input[5424]), .Z(n5120) );
  AND U5760 ( .A(p_input[9424]), .B(p_input[8424]), .Z(n5118) );
  AND U5761 ( .A(n5121), .B(n5122), .Z(o[423]) );
  AND U5762 ( .A(n5123), .B(n5124), .Z(n5122) );
  AND U5763 ( .A(n5125), .B(p_input[3423]), .Z(n5124) );
  AND U5764 ( .A(p_input[2423]), .B(p_input[1423]), .Z(n5125) );
  AND U5765 ( .A(p_input[4423]), .B(p_input[423]), .Z(n5123) );
  AND U5766 ( .A(n5126), .B(n5127), .Z(n5121) );
  AND U5767 ( .A(n5128), .B(p_input[7423]), .Z(n5127) );
  AND U5768 ( .A(p_input[6423]), .B(p_input[5423]), .Z(n5128) );
  AND U5769 ( .A(p_input[9423]), .B(p_input[8423]), .Z(n5126) );
  AND U5770 ( .A(n5129), .B(n5130), .Z(o[422]) );
  AND U5771 ( .A(n5131), .B(n5132), .Z(n5130) );
  AND U5772 ( .A(n5133), .B(p_input[3422]), .Z(n5132) );
  AND U5773 ( .A(p_input[2422]), .B(p_input[1422]), .Z(n5133) );
  AND U5774 ( .A(p_input[4422]), .B(p_input[422]), .Z(n5131) );
  AND U5775 ( .A(n5134), .B(n5135), .Z(n5129) );
  AND U5776 ( .A(n5136), .B(p_input[7422]), .Z(n5135) );
  AND U5777 ( .A(p_input[6422]), .B(p_input[5422]), .Z(n5136) );
  AND U5778 ( .A(p_input[9422]), .B(p_input[8422]), .Z(n5134) );
  AND U5779 ( .A(n5137), .B(n5138), .Z(o[421]) );
  AND U5780 ( .A(n5139), .B(n5140), .Z(n5138) );
  AND U5781 ( .A(n5141), .B(p_input[3421]), .Z(n5140) );
  AND U5782 ( .A(p_input[2421]), .B(p_input[1421]), .Z(n5141) );
  AND U5783 ( .A(p_input[4421]), .B(p_input[421]), .Z(n5139) );
  AND U5784 ( .A(n5142), .B(n5143), .Z(n5137) );
  AND U5785 ( .A(n5144), .B(p_input[7421]), .Z(n5143) );
  AND U5786 ( .A(p_input[6421]), .B(p_input[5421]), .Z(n5144) );
  AND U5787 ( .A(p_input[9421]), .B(p_input[8421]), .Z(n5142) );
  AND U5788 ( .A(n5145), .B(n5146), .Z(o[420]) );
  AND U5789 ( .A(n5147), .B(n5148), .Z(n5146) );
  AND U5790 ( .A(n5149), .B(p_input[3420]), .Z(n5148) );
  AND U5791 ( .A(p_input[2420]), .B(p_input[1420]), .Z(n5149) );
  AND U5792 ( .A(p_input[4420]), .B(p_input[420]), .Z(n5147) );
  AND U5793 ( .A(n5150), .B(n5151), .Z(n5145) );
  AND U5794 ( .A(n5152), .B(p_input[7420]), .Z(n5151) );
  AND U5795 ( .A(p_input[6420]), .B(p_input[5420]), .Z(n5152) );
  AND U5796 ( .A(p_input[9420]), .B(p_input[8420]), .Z(n5150) );
  AND U5797 ( .A(n5153), .B(n5154), .Z(o[41]) );
  AND U5798 ( .A(n5155), .B(n5156), .Z(n5154) );
  AND U5799 ( .A(n5157), .B(p_input[3041]), .Z(n5156) );
  AND U5800 ( .A(p_input[2041]), .B(p_input[1041]), .Z(n5157) );
  AND U5801 ( .A(p_input[41]), .B(p_input[4041]), .Z(n5155) );
  AND U5802 ( .A(n5158), .B(n5159), .Z(n5153) );
  AND U5803 ( .A(n5160), .B(p_input[7041]), .Z(n5159) );
  AND U5804 ( .A(p_input[6041]), .B(p_input[5041]), .Z(n5160) );
  AND U5805 ( .A(p_input[9041]), .B(p_input[8041]), .Z(n5158) );
  AND U5806 ( .A(n5161), .B(n5162), .Z(o[419]) );
  AND U5807 ( .A(n5163), .B(n5164), .Z(n5162) );
  AND U5808 ( .A(n5165), .B(p_input[3419]), .Z(n5164) );
  AND U5809 ( .A(p_input[2419]), .B(p_input[1419]), .Z(n5165) );
  AND U5810 ( .A(p_input[4419]), .B(p_input[419]), .Z(n5163) );
  AND U5811 ( .A(n5166), .B(n5167), .Z(n5161) );
  AND U5812 ( .A(n5168), .B(p_input[7419]), .Z(n5167) );
  AND U5813 ( .A(p_input[6419]), .B(p_input[5419]), .Z(n5168) );
  AND U5814 ( .A(p_input[9419]), .B(p_input[8419]), .Z(n5166) );
  AND U5815 ( .A(n5169), .B(n5170), .Z(o[418]) );
  AND U5816 ( .A(n5171), .B(n5172), .Z(n5170) );
  AND U5817 ( .A(n5173), .B(p_input[3418]), .Z(n5172) );
  AND U5818 ( .A(p_input[2418]), .B(p_input[1418]), .Z(n5173) );
  AND U5819 ( .A(p_input[4418]), .B(p_input[418]), .Z(n5171) );
  AND U5820 ( .A(n5174), .B(n5175), .Z(n5169) );
  AND U5821 ( .A(n5176), .B(p_input[7418]), .Z(n5175) );
  AND U5822 ( .A(p_input[6418]), .B(p_input[5418]), .Z(n5176) );
  AND U5823 ( .A(p_input[9418]), .B(p_input[8418]), .Z(n5174) );
  AND U5824 ( .A(n5177), .B(n5178), .Z(o[417]) );
  AND U5825 ( .A(n5179), .B(n5180), .Z(n5178) );
  AND U5826 ( .A(n5181), .B(p_input[3417]), .Z(n5180) );
  AND U5827 ( .A(p_input[2417]), .B(p_input[1417]), .Z(n5181) );
  AND U5828 ( .A(p_input[4417]), .B(p_input[417]), .Z(n5179) );
  AND U5829 ( .A(n5182), .B(n5183), .Z(n5177) );
  AND U5830 ( .A(n5184), .B(p_input[7417]), .Z(n5183) );
  AND U5831 ( .A(p_input[6417]), .B(p_input[5417]), .Z(n5184) );
  AND U5832 ( .A(p_input[9417]), .B(p_input[8417]), .Z(n5182) );
  AND U5833 ( .A(n5185), .B(n5186), .Z(o[416]) );
  AND U5834 ( .A(n5187), .B(n5188), .Z(n5186) );
  AND U5835 ( .A(n5189), .B(p_input[3416]), .Z(n5188) );
  AND U5836 ( .A(p_input[2416]), .B(p_input[1416]), .Z(n5189) );
  AND U5837 ( .A(p_input[4416]), .B(p_input[416]), .Z(n5187) );
  AND U5838 ( .A(n5190), .B(n5191), .Z(n5185) );
  AND U5839 ( .A(n5192), .B(p_input[7416]), .Z(n5191) );
  AND U5840 ( .A(p_input[6416]), .B(p_input[5416]), .Z(n5192) );
  AND U5841 ( .A(p_input[9416]), .B(p_input[8416]), .Z(n5190) );
  AND U5842 ( .A(n5193), .B(n5194), .Z(o[415]) );
  AND U5843 ( .A(n5195), .B(n5196), .Z(n5194) );
  AND U5844 ( .A(n5197), .B(p_input[3415]), .Z(n5196) );
  AND U5845 ( .A(p_input[2415]), .B(p_input[1415]), .Z(n5197) );
  AND U5846 ( .A(p_input[4415]), .B(p_input[415]), .Z(n5195) );
  AND U5847 ( .A(n5198), .B(n5199), .Z(n5193) );
  AND U5848 ( .A(n5200), .B(p_input[7415]), .Z(n5199) );
  AND U5849 ( .A(p_input[6415]), .B(p_input[5415]), .Z(n5200) );
  AND U5850 ( .A(p_input[9415]), .B(p_input[8415]), .Z(n5198) );
  AND U5851 ( .A(n5201), .B(n5202), .Z(o[414]) );
  AND U5852 ( .A(n5203), .B(n5204), .Z(n5202) );
  AND U5853 ( .A(n5205), .B(p_input[3414]), .Z(n5204) );
  AND U5854 ( .A(p_input[2414]), .B(p_input[1414]), .Z(n5205) );
  AND U5855 ( .A(p_input[4414]), .B(p_input[414]), .Z(n5203) );
  AND U5856 ( .A(n5206), .B(n5207), .Z(n5201) );
  AND U5857 ( .A(n5208), .B(p_input[7414]), .Z(n5207) );
  AND U5858 ( .A(p_input[6414]), .B(p_input[5414]), .Z(n5208) );
  AND U5859 ( .A(p_input[9414]), .B(p_input[8414]), .Z(n5206) );
  AND U5860 ( .A(n5209), .B(n5210), .Z(o[413]) );
  AND U5861 ( .A(n5211), .B(n5212), .Z(n5210) );
  AND U5862 ( .A(n5213), .B(p_input[3413]), .Z(n5212) );
  AND U5863 ( .A(p_input[2413]), .B(p_input[1413]), .Z(n5213) );
  AND U5864 ( .A(p_input[4413]), .B(p_input[413]), .Z(n5211) );
  AND U5865 ( .A(n5214), .B(n5215), .Z(n5209) );
  AND U5866 ( .A(n5216), .B(p_input[7413]), .Z(n5215) );
  AND U5867 ( .A(p_input[6413]), .B(p_input[5413]), .Z(n5216) );
  AND U5868 ( .A(p_input[9413]), .B(p_input[8413]), .Z(n5214) );
  AND U5869 ( .A(n5217), .B(n5218), .Z(o[412]) );
  AND U5870 ( .A(n5219), .B(n5220), .Z(n5218) );
  AND U5871 ( .A(n5221), .B(p_input[3412]), .Z(n5220) );
  AND U5872 ( .A(p_input[2412]), .B(p_input[1412]), .Z(n5221) );
  AND U5873 ( .A(p_input[4412]), .B(p_input[412]), .Z(n5219) );
  AND U5874 ( .A(n5222), .B(n5223), .Z(n5217) );
  AND U5875 ( .A(n5224), .B(p_input[7412]), .Z(n5223) );
  AND U5876 ( .A(p_input[6412]), .B(p_input[5412]), .Z(n5224) );
  AND U5877 ( .A(p_input[9412]), .B(p_input[8412]), .Z(n5222) );
  AND U5878 ( .A(n5225), .B(n5226), .Z(o[411]) );
  AND U5879 ( .A(n5227), .B(n5228), .Z(n5226) );
  AND U5880 ( .A(n5229), .B(p_input[3411]), .Z(n5228) );
  AND U5881 ( .A(p_input[2411]), .B(p_input[1411]), .Z(n5229) );
  AND U5882 ( .A(p_input[4411]), .B(p_input[411]), .Z(n5227) );
  AND U5883 ( .A(n5230), .B(n5231), .Z(n5225) );
  AND U5884 ( .A(n5232), .B(p_input[7411]), .Z(n5231) );
  AND U5885 ( .A(p_input[6411]), .B(p_input[5411]), .Z(n5232) );
  AND U5886 ( .A(p_input[9411]), .B(p_input[8411]), .Z(n5230) );
  AND U5887 ( .A(n5233), .B(n5234), .Z(o[410]) );
  AND U5888 ( .A(n5235), .B(n5236), .Z(n5234) );
  AND U5889 ( .A(n5237), .B(p_input[3410]), .Z(n5236) );
  AND U5890 ( .A(p_input[2410]), .B(p_input[1410]), .Z(n5237) );
  AND U5891 ( .A(p_input[4410]), .B(p_input[410]), .Z(n5235) );
  AND U5892 ( .A(n5238), .B(n5239), .Z(n5233) );
  AND U5893 ( .A(n5240), .B(p_input[7410]), .Z(n5239) );
  AND U5894 ( .A(p_input[6410]), .B(p_input[5410]), .Z(n5240) );
  AND U5895 ( .A(p_input[9410]), .B(p_input[8410]), .Z(n5238) );
  AND U5896 ( .A(n5241), .B(n5242), .Z(o[40]) );
  AND U5897 ( .A(n5243), .B(n5244), .Z(n5242) );
  AND U5898 ( .A(n5245), .B(p_input[3040]), .Z(n5244) );
  AND U5899 ( .A(p_input[2040]), .B(p_input[1040]), .Z(n5245) );
  AND U5900 ( .A(p_input[40]), .B(p_input[4040]), .Z(n5243) );
  AND U5901 ( .A(n5246), .B(n5247), .Z(n5241) );
  AND U5902 ( .A(n5248), .B(p_input[7040]), .Z(n5247) );
  AND U5903 ( .A(p_input[6040]), .B(p_input[5040]), .Z(n5248) );
  AND U5904 ( .A(p_input[9040]), .B(p_input[8040]), .Z(n5246) );
  AND U5905 ( .A(n5249), .B(n5250), .Z(o[409]) );
  AND U5906 ( .A(n5251), .B(n5252), .Z(n5250) );
  AND U5907 ( .A(n5253), .B(p_input[3409]), .Z(n5252) );
  AND U5908 ( .A(p_input[2409]), .B(p_input[1409]), .Z(n5253) );
  AND U5909 ( .A(p_input[4409]), .B(p_input[409]), .Z(n5251) );
  AND U5910 ( .A(n5254), .B(n5255), .Z(n5249) );
  AND U5911 ( .A(n5256), .B(p_input[7409]), .Z(n5255) );
  AND U5912 ( .A(p_input[6409]), .B(p_input[5409]), .Z(n5256) );
  AND U5913 ( .A(p_input[9409]), .B(p_input[8409]), .Z(n5254) );
  AND U5914 ( .A(n5257), .B(n5258), .Z(o[408]) );
  AND U5915 ( .A(n5259), .B(n5260), .Z(n5258) );
  AND U5916 ( .A(n5261), .B(p_input[3408]), .Z(n5260) );
  AND U5917 ( .A(p_input[2408]), .B(p_input[1408]), .Z(n5261) );
  AND U5918 ( .A(p_input[4408]), .B(p_input[408]), .Z(n5259) );
  AND U5919 ( .A(n5262), .B(n5263), .Z(n5257) );
  AND U5920 ( .A(n5264), .B(p_input[7408]), .Z(n5263) );
  AND U5921 ( .A(p_input[6408]), .B(p_input[5408]), .Z(n5264) );
  AND U5922 ( .A(p_input[9408]), .B(p_input[8408]), .Z(n5262) );
  AND U5923 ( .A(n5265), .B(n5266), .Z(o[407]) );
  AND U5924 ( .A(n5267), .B(n5268), .Z(n5266) );
  AND U5925 ( .A(n5269), .B(p_input[3407]), .Z(n5268) );
  AND U5926 ( .A(p_input[2407]), .B(p_input[1407]), .Z(n5269) );
  AND U5927 ( .A(p_input[4407]), .B(p_input[407]), .Z(n5267) );
  AND U5928 ( .A(n5270), .B(n5271), .Z(n5265) );
  AND U5929 ( .A(n5272), .B(p_input[7407]), .Z(n5271) );
  AND U5930 ( .A(p_input[6407]), .B(p_input[5407]), .Z(n5272) );
  AND U5931 ( .A(p_input[9407]), .B(p_input[8407]), .Z(n5270) );
  AND U5932 ( .A(n5273), .B(n5274), .Z(o[406]) );
  AND U5933 ( .A(n5275), .B(n5276), .Z(n5274) );
  AND U5934 ( .A(n5277), .B(p_input[3406]), .Z(n5276) );
  AND U5935 ( .A(p_input[2406]), .B(p_input[1406]), .Z(n5277) );
  AND U5936 ( .A(p_input[4406]), .B(p_input[406]), .Z(n5275) );
  AND U5937 ( .A(n5278), .B(n5279), .Z(n5273) );
  AND U5938 ( .A(n5280), .B(p_input[7406]), .Z(n5279) );
  AND U5939 ( .A(p_input[6406]), .B(p_input[5406]), .Z(n5280) );
  AND U5940 ( .A(p_input[9406]), .B(p_input[8406]), .Z(n5278) );
  AND U5941 ( .A(n5281), .B(n5282), .Z(o[405]) );
  AND U5942 ( .A(n5283), .B(n5284), .Z(n5282) );
  AND U5943 ( .A(n5285), .B(p_input[3405]), .Z(n5284) );
  AND U5944 ( .A(p_input[2405]), .B(p_input[1405]), .Z(n5285) );
  AND U5945 ( .A(p_input[4405]), .B(p_input[405]), .Z(n5283) );
  AND U5946 ( .A(n5286), .B(n5287), .Z(n5281) );
  AND U5947 ( .A(n5288), .B(p_input[7405]), .Z(n5287) );
  AND U5948 ( .A(p_input[6405]), .B(p_input[5405]), .Z(n5288) );
  AND U5949 ( .A(p_input[9405]), .B(p_input[8405]), .Z(n5286) );
  AND U5950 ( .A(n5289), .B(n5290), .Z(o[404]) );
  AND U5951 ( .A(n5291), .B(n5292), .Z(n5290) );
  AND U5952 ( .A(n5293), .B(p_input[3404]), .Z(n5292) );
  AND U5953 ( .A(p_input[2404]), .B(p_input[1404]), .Z(n5293) );
  AND U5954 ( .A(p_input[4404]), .B(p_input[404]), .Z(n5291) );
  AND U5955 ( .A(n5294), .B(n5295), .Z(n5289) );
  AND U5956 ( .A(n5296), .B(p_input[7404]), .Z(n5295) );
  AND U5957 ( .A(p_input[6404]), .B(p_input[5404]), .Z(n5296) );
  AND U5958 ( .A(p_input[9404]), .B(p_input[8404]), .Z(n5294) );
  AND U5959 ( .A(n5297), .B(n5298), .Z(o[403]) );
  AND U5960 ( .A(n5299), .B(n5300), .Z(n5298) );
  AND U5961 ( .A(n5301), .B(p_input[3403]), .Z(n5300) );
  AND U5962 ( .A(p_input[2403]), .B(p_input[1403]), .Z(n5301) );
  AND U5963 ( .A(p_input[4403]), .B(p_input[403]), .Z(n5299) );
  AND U5964 ( .A(n5302), .B(n5303), .Z(n5297) );
  AND U5965 ( .A(n5304), .B(p_input[7403]), .Z(n5303) );
  AND U5966 ( .A(p_input[6403]), .B(p_input[5403]), .Z(n5304) );
  AND U5967 ( .A(p_input[9403]), .B(p_input[8403]), .Z(n5302) );
  AND U5968 ( .A(n5305), .B(n5306), .Z(o[402]) );
  AND U5969 ( .A(n5307), .B(n5308), .Z(n5306) );
  AND U5970 ( .A(n5309), .B(p_input[3402]), .Z(n5308) );
  AND U5971 ( .A(p_input[2402]), .B(p_input[1402]), .Z(n5309) );
  AND U5972 ( .A(p_input[4402]), .B(p_input[402]), .Z(n5307) );
  AND U5973 ( .A(n5310), .B(n5311), .Z(n5305) );
  AND U5974 ( .A(n5312), .B(p_input[7402]), .Z(n5311) );
  AND U5975 ( .A(p_input[6402]), .B(p_input[5402]), .Z(n5312) );
  AND U5976 ( .A(p_input[9402]), .B(p_input[8402]), .Z(n5310) );
  AND U5977 ( .A(n5313), .B(n5314), .Z(o[401]) );
  AND U5978 ( .A(n5315), .B(n5316), .Z(n5314) );
  AND U5979 ( .A(n5317), .B(p_input[3401]), .Z(n5316) );
  AND U5980 ( .A(p_input[2401]), .B(p_input[1401]), .Z(n5317) );
  AND U5981 ( .A(p_input[4401]), .B(p_input[401]), .Z(n5315) );
  AND U5982 ( .A(n5318), .B(n5319), .Z(n5313) );
  AND U5983 ( .A(n5320), .B(p_input[7401]), .Z(n5319) );
  AND U5984 ( .A(p_input[6401]), .B(p_input[5401]), .Z(n5320) );
  AND U5985 ( .A(p_input[9401]), .B(p_input[8401]), .Z(n5318) );
  AND U5986 ( .A(n5321), .B(n5322), .Z(o[400]) );
  AND U5987 ( .A(n5323), .B(n5324), .Z(n5322) );
  AND U5988 ( .A(n5325), .B(p_input[3400]), .Z(n5324) );
  AND U5989 ( .A(p_input[2400]), .B(p_input[1400]), .Z(n5325) );
  AND U5990 ( .A(p_input[4400]), .B(p_input[400]), .Z(n5323) );
  AND U5991 ( .A(n5326), .B(n5327), .Z(n5321) );
  AND U5992 ( .A(n5328), .B(p_input[7400]), .Z(n5327) );
  AND U5993 ( .A(p_input[6400]), .B(p_input[5400]), .Z(n5328) );
  AND U5994 ( .A(p_input[9400]), .B(p_input[8400]), .Z(n5326) );
  AND U5995 ( .A(n5329), .B(n5330), .Z(o[3]) );
  AND U5996 ( .A(n5331), .B(n5332), .Z(n5330) );
  AND U5997 ( .A(n5333), .B(p_input[3003]), .Z(n5332) );
  AND U5998 ( .A(p_input[2003]), .B(p_input[1003]), .Z(n5333) );
  AND U5999 ( .A(p_input[4003]), .B(p_input[3]), .Z(n5331) );
  AND U6000 ( .A(n5334), .B(n5335), .Z(n5329) );
  AND U6001 ( .A(n5336), .B(p_input[7003]), .Z(n5335) );
  AND U6002 ( .A(p_input[6003]), .B(p_input[5003]), .Z(n5336) );
  AND U6003 ( .A(p_input[9003]), .B(p_input[8003]), .Z(n5334) );
  AND U6004 ( .A(n5337), .B(n5338), .Z(o[39]) );
  AND U6005 ( .A(n5339), .B(n5340), .Z(n5338) );
  AND U6006 ( .A(n5341), .B(p_input[3039]), .Z(n5340) );
  AND U6007 ( .A(p_input[2039]), .B(p_input[1039]), .Z(n5341) );
  AND U6008 ( .A(p_input[4039]), .B(p_input[39]), .Z(n5339) );
  AND U6009 ( .A(n5342), .B(n5343), .Z(n5337) );
  AND U6010 ( .A(n5344), .B(p_input[7039]), .Z(n5343) );
  AND U6011 ( .A(p_input[6039]), .B(p_input[5039]), .Z(n5344) );
  AND U6012 ( .A(p_input[9039]), .B(p_input[8039]), .Z(n5342) );
  AND U6013 ( .A(n5345), .B(n5346), .Z(o[399]) );
  AND U6014 ( .A(n5347), .B(n5348), .Z(n5346) );
  AND U6015 ( .A(n5349), .B(p_input[3399]), .Z(n5348) );
  AND U6016 ( .A(p_input[2399]), .B(p_input[1399]), .Z(n5349) );
  AND U6017 ( .A(p_input[4399]), .B(p_input[399]), .Z(n5347) );
  AND U6018 ( .A(n5350), .B(n5351), .Z(n5345) );
  AND U6019 ( .A(n5352), .B(p_input[7399]), .Z(n5351) );
  AND U6020 ( .A(p_input[6399]), .B(p_input[5399]), .Z(n5352) );
  AND U6021 ( .A(p_input[9399]), .B(p_input[8399]), .Z(n5350) );
  AND U6022 ( .A(n5353), .B(n5354), .Z(o[398]) );
  AND U6023 ( .A(n5355), .B(n5356), .Z(n5354) );
  AND U6024 ( .A(n5357), .B(p_input[3398]), .Z(n5356) );
  AND U6025 ( .A(p_input[2398]), .B(p_input[1398]), .Z(n5357) );
  AND U6026 ( .A(p_input[4398]), .B(p_input[398]), .Z(n5355) );
  AND U6027 ( .A(n5358), .B(n5359), .Z(n5353) );
  AND U6028 ( .A(n5360), .B(p_input[7398]), .Z(n5359) );
  AND U6029 ( .A(p_input[6398]), .B(p_input[5398]), .Z(n5360) );
  AND U6030 ( .A(p_input[9398]), .B(p_input[8398]), .Z(n5358) );
  AND U6031 ( .A(n5361), .B(n5362), .Z(o[397]) );
  AND U6032 ( .A(n5363), .B(n5364), .Z(n5362) );
  AND U6033 ( .A(n5365), .B(p_input[3397]), .Z(n5364) );
  AND U6034 ( .A(p_input[2397]), .B(p_input[1397]), .Z(n5365) );
  AND U6035 ( .A(p_input[4397]), .B(p_input[397]), .Z(n5363) );
  AND U6036 ( .A(n5366), .B(n5367), .Z(n5361) );
  AND U6037 ( .A(n5368), .B(p_input[7397]), .Z(n5367) );
  AND U6038 ( .A(p_input[6397]), .B(p_input[5397]), .Z(n5368) );
  AND U6039 ( .A(p_input[9397]), .B(p_input[8397]), .Z(n5366) );
  AND U6040 ( .A(n5369), .B(n5370), .Z(o[396]) );
  AND U6041 ( .A(n5371), .B(n5372), .Z(n5370) );
  AND U6042 ( .A(n5373), .B(p_input[3396]), .Z(n5372) );
  AND U6043 ( .A(p_input[2396]), .B(p_input[1396]), .Z(n5373) );
  AND U6044 ( .A(p_input[4396]), .B(p_input[396]), .Z(n5371) );
  AND U6045 ( .A(n5374), .B(n5375), .Z(n5369) );
  AND U6046 ( .A(n5376), .B(p_input[7396]), .Z(n5375) );
  AND U6047 ( .A(p_input[6396]), .B(p_input[5396]), .Z(n5376) );
  AND U6048 ( .A(p_input[9396]), .B(p_input[8396]), .Z(n5374) );
  AND U6049 ( .A(n5377), .B(n5378), .Z(o[395]) );
  AND U6050 ( .A(n5379), .B(n5380), .Z(n5378) );
  AND U6051 ( .A(n5381), .B(p_input[3395]), .Z(n5380) );
  AND U6052 ( .A(p_input[2395]), .B(p_input[1395]), .Z(n5381) );
  AND U6053 ( .A(p_input[4395]), .B(p_input[395]), .Z(n5379) );
  AND U6054 ( .A(n5382), .B(n5383), .Z(n5377) );
  AND U6055 ( .A(n5384), .B(p_input[7395]), .Z(n5383) );
  AND U6056 ( .A(p_input[6395]), .B(p_input[5395]), .Z(n5384) );
  AND U6057 ( .A(p_input[9395]), .B(p_input[8395]), .Z(n5382) );
  AND U6058 ( .A(n5385), .B(n5386), .Z(o[394]) );
  AND U6059 ( .A(n5387), .B(n5388), .Z(n5386) );
  AND U6060 ( .A(n5389), .B(p_input[3394]), .Z(n5388) );
  AND U6061 ( .A(p_input[2394]), .B(p_input[1394]), .Z(n5389) );
  AND U6062 ( .A(p_input[4394]), .B(p_input[394]), .Z(n5387) );
  AND U6063 ( .A(n5390), .B(n5391), .Z(n5385) );
  AND U6064 ( .A(n5392), .B(p_input[7394]), .Z(n5391) );
  AND U6065 ( .A(p_input[6394]), .B(p_input[5394]), .Z(n5392) );
  AND U6066 ( .A(p_input[9394]), .B(p_input[8394]), .Z(n5390) );
  AND U6067 ( .A(n5393), .B(n5394), .Z(o[393]) );
  AND U6068 ( .A(n5395), .B(n5396), .Z(n5394) );
  AND U6069 ( .A(n5397), .B(p_input[3393]), .Z(n5396) );
  AND U6070 ( .A(p_input[2393]), .B(p_input[1393]), .Z(n5397) );
  AND U6071 ( .A(p_input[4393]), .B(p_input[393]), .Z(n5395) );
  AND U6072 ( .A(n5398), .B(n5399), .Z(n5393) );
  AND U6073 ( .A(n5400), .B(p_input[7393]), .Z(n5399) );
  AND U6074 ( .A(p_input[6393]), .B(p_input[5393]), .Z(n5400) );
  AND U6075 ( .A(p_input[9393]), .B(p_input[8393]), .Z(n5398) );
  AND U6076 ( .A(n5401), .B(n5402), .Z(o[392]) );
  AND U6077 ( .A(n5403), .B(n5404), .Z(n5402) );
  AND U6078 ( .A(n5405), .B(p_input[3392]), .Z(n5404) );
  AND U6079 ( .A(p_input[2392]), .B(p_input[1392]), .Z(n5405) );
  AND U6080 ( .A(p_input[4392]), .B(p_input[392]), .Z(n5403) );
  AND U6081 ( .A(n5406), .B(n5407), .Z(n5401) );
  AND U6082 ( .A(n5408), .B(p_input[7392]), .Z(n5407) );
  AND U6083 ( .A(p_input[6392]), .B(p_input[5392]), .Z(n5408) );
  AND U6084 ( .A(p_input[9392]), .B(p_input[8392]), .Z(n5406) );
  AND U6085 ( .A(n5409), .B(n5410), .Z(o[391]) );
  AND U6086 ( .A(n5411), .B(n5412), .Z(n5410) );
  AND U6087 ( .A(n5413), .B(p_input[3391]), .Z(n5412) );
  AND U6088 ( .A(p_input[2391]), .B(p_input[1391]), .Z(n5413) );
  AND U6089 ( .A(p_input[4391]), .B(p_input[391]), .Z(n5411) );
  AND U6090 ( .A(n5414), .B(n5415), .Z(n5409) );
  AND U6091 ( .A(n5416), .B(p_input[7391]), .Z(n5415) );
  AND U6092 ( .A(p_input[6391]), .B(p_input[5391]), .Z(n5416) );
  AND U6093 ( .A(p_input[9391]), .B(p_input[8391]), .Z(n5414) );
  AND U6094 ( .A(n5417), .B(n5418), .Z(o[390]) );
  AND U6095 ( .A(n5419), .B(n5420), .Z(n5418) );
  AND U6096 ( .A(n5421), .B(p_input[3390]), .Z(n5420) );
  AND U6097 ( .A(p_input[2390]), .B(p_input[1390]), .Z(n5421) );
  AND U6098 ( .A(p_input[4390]), .B(p_input[390]), .Z(n5419) );
  AND U6099 ( .A(n5422), .B(n5423), .Z(n5417) );
  AND U6100 ( .A(n5424), .B(p_input[7390]), .Z(n5423) );
  AND U6101 ( .A(p_input[6390]), .B(p_input[5390]), .Z(n5424) );
  AND U6102 ( .A(p_input[9390]), .B(p_input[8390]), .Z(n5422) );
  AND U6103 ( .A(n5425), .B(n5426), .Z(o[38]) );
  AND U6104 ( .A(n5427), .B(n5428), .Z(n5426) );
  AND U6105 ( .A(n5429), .B(p_input[3038]), .Z(n5428) );
  AND U6106 ( .A(p_input[2038]), .B(p_input[1038]), .Z(n5429) );
  AND U6107 ( .A(p_input[4038]), .B(p_input[38]), .Z(n5427) );
  AND U6108 ( .A(n5430), .B(n5431), .Z(n5425) );
  AND U6109 ( .A(n5432), .B(p_input[7038]), .Z(n5431) );
  AND U6110 ( .A(p_input[6038]), .B(p_input[5038]), .Z(n5432) );
  AND U6111 ( .A(p_input[9038]), .B(p_input[8038]), .Z(n5430) );
  AND U6112 ( .A(n5433), .B(n5434), .Z(o[389]) );
  AND U6113 ( .A(n5435), .B(n5436), .Z(n5434) );
  AND U6114 ( .A(n5437), .B(p_input[3389]), .Z(n5436) );
  AND U6115 ( .A(p_input[2389]), .B(p_input[1389]), .Z(n5437) );
  AND U6116 ( .A(p_input[4389]), .B(p_input[389]), .Z(n5435) );
  AND U6117 ( .A(n5438), .B(n5439), .Z(n5433) );
  AND U6118 ( .A(n5440), .B(p_input[7389]), .Z(n5439) );
  AND U6119 ( .A(p_input[6389]), .B(p_input[5389]), .Z(n5440) );
  AND U6120 ( .A(p_input[9389]), .B(p_input[8389]), .Z(n5438) );
  AND U6121 ( .A(n5441), .B(n5442), .Z(o[388]) );
  AND U6122 ( .A(n5443), .B(n5444), .Z(n5442) );
  AND U6123 ( .A(n5445), .B(p_input[3388]), .Z(n5444) );
  AND U6124 ( .A(p_input[2388]), .B(p_input[1388]), .Z(n5445) );
  AND U6125 ( .A(p_input[4388]), .B(p_input[388]), .Z(n5443) );
  AND U6126 ( .A(n5446), .B(n5447), .Z(n5441) );
  AND U6127 ( .A(n5448), .B(p_input[7388]), .Z(n5447) );
  AND U6128 ( .A(p_input[6388]), .B(p_input[5388]), .Z(n5448) );
  AND U6129 ( .A(p_input[9388]), .B(p_input[8388]), .Z(n5446) );
  AND U6130 ( .A(n5449), .B(n5450), .Z(o[387]) );
  AND U6131 ( .A(n5451), .B(n5452), .Z(n5450) );
  AND U6132 ( .A(n5453), .B(p_input[3387]), .Z(n5452) );
  AND U6133 ( .A(p_input[2387]), .B(p_input[1387]), .Z(n5453) );
  AND U6134 ( .A(p_input[4387]), .B(p_input[387]), .Z(n5451) );
  AND U6135 ( .A(n5454), .B(n5455), .Z(n5449) );
  AND U6136 ( .A(n5456), .B(p_input[7387]), .Z(n5455) );
  AND U6137 ( .A(p_input[6387]), .B(p_input[5387]), .Z(n5456) );
  AND U6138 ( .A(p_input[9387]), .B(p_input[8387]), .Z(n5454) );
  AND U6139 ( .A(n5457), .B(n5458), .Z(o[386]) );
  AND U6140 ( .A(n5459), .B(n5460), .Z(n5458) );
  AND U6141 ( .A(n5461), .B(p_input[3386]), .Z(n5460) );
  AND U6142 ( .A(p_input[2386]), .B(p_input[1386]), .Z(n5461) );
  AND U6143 ( .A(p_input[4386]), .B(p_input[386]), .Z(n5459) );
  AND U6144 ( .A(n5462), .B(n5463), .Z(n5457) );
  AND U6145 ( .A(n5464), .B(p_input[7386]), .Z(n5463) );
  AND U6146 ( .A(p_input[6386]), .B(p_input[5386]), .Z(n5464) );
  AND U6147 ( .A(p_input[9386]), .B(p_input[8386]), .Z(n5462) );
  AND U6148 ( .A(n5465), .B(n5466), .Z(o[385]) );
  AND U6149 ( .A(n5467), .B(n5468), .Z(n5466) );
  AND U6150 ( .A(n5469), .B(p_input[3385]), .Z(n5468) );
  AND U6151 ( .A(p_input[2385]), .B(p_input[1385]), .Z(n5469) );
  AND U6152 ( .A(p_input[4385]), .B(p_input[385]), .Z(n5467) );
  AND U6153 ( .A(n5470), .B(n5471), .Z(n5465) );
  AND U6154 ( .A(n5472), .B(p_input[7385]), .Z(n5471) );
  AND U6155 ( .A(p_input[6385]), .B(p_input[5385]), .Z(n5472) );
  AND U6156 ( .A(p_input[9385]), .B(p_input[8385]), .Z(n5470) );
  AND U6157 ( .A(n5473), .B(n5474), .Z(o[384]) );
  AND U6158 ( .A(n5475), .B(n5476), .Z(n5474) );
  AND U6159 ( .A(n5477), .B(p_input[3384]), .Z(n5476) );
  AND U6160 ( .A(p_input[2384]), .B(p_input[1384]), .Z(n5477) );
  AND U6161 ( .A(p_input[4384]), .B(p_input[384]), .Z(n5475) );
  AND U6162 ( .A(n5478), .B(n5479), .Z(n5473) );
  AND U6163 ( .A(n5480), .B(p_input[7384]), .Z(n5479) );
  AND U6164 ( .A(p_input[6384]), .B(p_input[5384]), .Z(n5480) );
  AND U6165 ( .A(p_input[9384]), .B(p_input[8384]), .Z(n5478) );
  AND U6166 ( .A(n5481), .B(n5482), .Z(o[383]) );
  AND U6167 ( .A(n5483), .B(n5484), .Z(n5482) );
  AND U6168 ( .A(n5485), .B(p_input[3383]), .Z(n5484) );
  AND U6169 ( .A(p_input[2383]), .B(p_input[1383]), .Z(n5485) );
  AND U6170 ( .A(p_input[4383]), .B(p_input[383]), .Z(n5483) );
  AND U6171 ( .A(n5486), .B(n5487), .Z(n5481) );
  AND U6172 ( .A(n5488), .B(p_input[7383]), .Z(n5487) );
  AND U6173 ( .A(p_input[6383]), .B(p_input[5383]), .Z(n5488) );
  AND U6174 ( .A(p_input[9383]), .B(p_input[8383]), .Z(n5486) );
  AND U6175 ( .A(n5489), .B(n5490), .Z(o[382]) );
  AND U6176 ( .A(n5491), .B(n5492), .Z(n5490) );
  AND U6177 ( .A(n5493), .B(p_input[3382]), .Z(n5492) );
  AND U6178 ( .A(p_input[2382]), .B(p_input[1382]), .Z(n5493) );
  AND U6179 ( .A(p_input[4382]), .B(p_input[382]), .Z(n5491) );
  AND U6180 ( .A(n5494), .B(n5495), .Z(n5489) );
  AND U6181 ( .A(n5496), .B(p_input[7382]), .Z(n5495) );
  AND U6182 ( .A(p_input[6382]), .B(p_input[5382]), .Z(n5496) );
  AND U6183 ( .A(p_input[9382]), .B(p_input[8382]), .Z(n5494) );
  AND U6184 ( .A(n5497), .B(n5498), .Z(o[381]) );
  AND U6185 ( .A(n5499), .B(n5500), .Z(n5498) );
  AND U6186 ( .A(n5501), .B(p_input[3381]), .Z(n5500) );
  AND U6187 ( .A(p_input[2381]), .B(p_input[1381]), .Z(n5501) );
  AND U6188 ( .A(p_input[4381]), .B(p_input[381]), .Z(n5499) );
  AND U6189 ( .A(n5502), .B(n5503), .Z(n5497) );
  AND U6190 ( .A(n5504), .B(p_input[7381]), .Z(n5503) );
  AND U6191 ( .A(p_input[6381]), .B(p_input[5381]), .Z(n5504) );
  AND U6192 ( .A(p_input[9381]), .B(p_input[8381]), .Z(n5502) );
  AND U6193 ( .A(n5505), .B(n5506), .Z(o[380]) );
  AND U6194 ( .A(n5507), .B(n5508), .Z(n5506) );
  AND U6195 ( .A(n5509), .B(p_input[3380]), .Z(n5508) );
  AND U6196 ( .A(p_input[2380]), .B(p_input[1380]), .Z(n5509) );
  AND U6197 ( .A(p_input[4380]), .B(p_input[380]), .Z(n5507) );
  AND U6198 ( .A(n5510), .B(n5511), .Z(n5505) );
  AND U6199 ( .A(n5512), .B(p_input[7380]), .Z(n5511) );
  AND U6200 ( .A(p_input[6380]), .B(p_input[5380]), .Z(n5512) );
  AND U6201 ( .A(p_input[9380]), .B(p_input[8380]), .Z(n5510) );
  AND U6202 ( .A(n5513), .B(n5514), .Z(o[37]) );
  AND U6203 ( .A(n5515), .B(n5516), .Z(n5514) );
  AND U6204 ( .A(n5517), .B(p_input[3037]), .Z(n5516) );
  AND U6205 ( .A(p_input[2037]), .B(p_input[1037]), .Z(n5517) );
  AND U6206 ( .A(p_input[4037]), .B(p_input[37]), .Z(n5515) );
  AND U6207 ( .A(n5518), .B(n5519), .Z(n5513) );
  AND U6208 ( .A(n5520), .B(p_input[7037]), .Z(n5519) );
  AND U6209 ( .A(p_input[6037]), .B(p_input[5037]), .Z(n5520) );
  AND U6210 ( .A(p_input[9037]), .B(p_input[8037]), .Z(n5518) );
  AND U6211 ( .A(n5521), .B(n5522), .Z(o[379]) );
  AND U6212 ( .A(n5523), .B(n5524), .Z(n5522) );
  AND U6213 ( .A(n5525), .B(p_input[3379]), .Z(n5524) );
  AND U6214 ( .A(p_input[2379]), .B(p_input[1379]), .Z(n5525) );
  AND U6215 ( .A(p_input[4379]), .B(p_input[379]), .Z(n5523) );
  AND U6216 ( .A(n5526), .B(n5527), .Z(n5521) );
  AND U6217 ( .A(n5528), .B(p_input[7379]), .Z(n5527) );
  AND U6218 ( .A(p_input[6379]), .B(p_input[5379]), .Z(n5528) );
  AND U6219 ( .A(p_input[9379]), .B(p_input[8379]), .Z(n5526) );
  AND U6220 ( .A(n5529), .B(n5530), .Z(o[378]) );
  AND U6221 ( .A(n5531), .B(n5532), .Z(n5530) );
  AND U6222 ( .A(n5533), .B(p_input[3378]), .Z(n5532) );
  AND U6223 ( .A(p_input[2378]), .B(p_input[1378]), .Z(n5533) );
  AND U6224 ( .A(p_input[4378]), .B(p_input[378]), .Z(n5531) );
  AND U6225 ( .A(n5534), .B(n5535), .Z(n5529) );
  AND U6226 ( .A(n5536), .B(p_input[7378]), .Z(n5535) );
  AND U6227 ( .A(p_input[6378]), .B(p_input[5378]), .Z(n5536) );
  AND U6228 ( .A(p_input[9378]), .B(p_input[8378]), .Z(n5534) );
  AND U6229 ( .A(n5537), .B(n5538), .Z(o[377]) );
  AND U6230 ( .A(n5539), .B(n5540), .Z(n5538) );
  AND U6231 ( .A(n5541), .B(p_input[3377]), .Z(n5540) );
  AND U6232 ( .A(p_input[2377]), .B(p_input[1377]), .Z(n5541) );
  AND U6233 ( .A(p_input[4377]), .B(p_input[377]), .Z(n5539) );
  AND U6234 ( .A(n5542), .B(n5543), .Z(n5537) );
  AND U6235 ( .A(n5544), .B(p_input[7377]), .Z(n5543) );
  AND U6236 ( .A(p_input[6377]), .B(p_input[5377]), .Z(n5544) );
  AND U6237 ( .A(p_input[9377]), .B(p_input[8377]), .Z(n5542) );
  AND U6238 ( .A(n5545), .B(n5546), .Z(o[376]) );
  AND U6239 ( .A(n5547), .B(n5548), .Z(n5546) );
  AND U6240 ( .A(n5549), .B(p_input[3376]), .Z(n5548) );
  AND U6241 ( .A(p_input[2376]), .B(p_input[1376]), .Z(n5549) );
  AND U6242 ( .A(p_input[4376]), .B(p_input[376]), .Z(n5547) );
  AND U6243 ( .A(n5550), .B(n5551), .Z(n5545) );
  AND U6244 ( .A(n5552), .B(p_input[7376]), .Z(n5551) );
  AND U6245 ( .A(p_input[6376]), .B(p_input[5376]), .Z(n5552) );
  AND U6246 ( .A(p_input[9376]), .B(p_input[8376]), .Z(n5550) );
  AND U6247 ( .A(n5553), .B(n5554), .Z(o[375]) );
  AND U6248 ( .A(n5555), .B(n5556), .Z(n5554) );
  AND U6249 ( .A(n5557), .B(p_input[3375]), .Z(n5556) );
  AND U6250 ( .A(p_input[2375]), .B(p_input[1375]), .Z(n5557) );
  AND U6251 ( .A(p_input[4375]), .B(p_input[375]), .Z(n5555) );
  AND U6252 ( .A(n5558), .B(n5559), .Z(n5553) );
  AND U6253 ( .A(n5560), .B(p_input[7375]), .Z(n5559) );
  AND U6254 ( .A(p_input[6375]), .B(p_input[5375]), .Z(n5560) );
  AND U6255 ( .A(p_input[9375]), .B(p_input[8375]), .Z(n5558) );
  AND U6256 ( .A(n5561), .B(n5562), .Z(o[374]) );
  AND U6257 ( .A(n5563), .B(n5564), .Z(n5562) );
  AND U6258 ( .A(n5565), .B(p_input[3374]), .Z(n5564) );
  AND U6259 ( .A(p_input[2374]), .B(p_input[1374]), .Z(n5565) );
  AND U6260 ( .A(p_input[4374]), .B(p_input[374]), .Z(n5563) );
  AND U6261 ( .A(n5566), .B(n5567), .Z(n5561) );
  AND U6262 ( .A(n5568), .B(p_input[7374]), .Z(n5567) );
  AND U6263 ( .A(p_input[6374]), .B(p_input[5374]), .Z(n5568) );
  AND U6264 ( .A(p_input[9374]), .B(p_input[8374]), .Z(n5566) );
  AND U6265 ( .A(n5569), .B(n5570), .Z(o[373]) );
  AND U6266 ( .A(n5571), .B(n5572), .Z(n5570) );
  AND U6267 ( .A(n5573), .B(p_input[3373]), .Z(n5572) );
  AND U6268 ( .A(p_input[2373]), .B(p_input[1373]), .Z(n5573) );
  AND U6269 ( .A(p_input[4373]), .B(p_input[373]), .Z(n5571) );
  AND U6270 ( .A(n5574), .B(n5575), .Z(n5569) );
  AND U6271 ( .A(n5576), .B(p_input[7373]), .Z(n5575) );
  AND U6272 ( .A(p_input[6373]), .B(p_input[5373]), .Z(n5576) );
  AND U6273 ( .A(p_input[9373]), .B(p_input[8373]), .Z(n5574) );
  AND U6274 ( .A(n5577), .B(n5578), .Z(o[372]) );
  AND U6275 ( .A(n5579), .B(n5580), .Z(n5578) );
  AND U6276 ( .A(n5581), .B(p_input[3372]), .Z(n5580) );
  AND U6277 ( .A(p_input[2372]), .B(p_input[1372]), .Z(n5581) );
  AND U6278 ( .A(p_input[4372]), .B(p_input[372]), .Z(n5579) );
  AND U6279 ( .A(n5582), .B(n5583), .Z(n5577) );
  AND U6280 ( .A(n5584), .B(p_input[7372]), .Z(n5583) );
  AND U6281 ( .A(p_input[6372]), .B(p_input[5372]), .Z(n5584) );
  AND U6282 ( .A(p_input[9372]), .B(p_input[8372]), .Z(n5582) );
  AND U6283 ( .A(n5585), .B(n5586), .Z(o[371]) );
  AND U6284 ( .A(n5587), .B(n5588), .Z(n5586) );
  AND U6285 ( .A(n5589), .B(p_input[3371]), .Z(n5588) );
  AND U6286 ( .A(p_input[2371]), .B(p_input[1371]), .Z(n5589) );
  AND U6287 ( .A(p_input[4371]), .B(p_input[371]), .Z(n5587) );
  AND U6288 ( .A(n5590), .B(n5591), .Z(n5585) );
  AND U6289 ( .A(n5592), .B(p_input[7371]), .Z(n5591) );
  AND U6290 ( .A(p_input[6371]), .B(p_input[5371]), .Z(n5592) );
  AND U6291 ( .A(p_input[9371]), .B(p_input[8371]), .Z(n5590) );
  AND U6292 ( .A(n5593), .B(n5594), .Z(o[370]) );
  AND U6293 ( .A(n5595), .B(n5596), .Z(n5594) );
  AND U6294 ( .A(n5597), .B(p_input[3370]), .Z(n5596) );
  AND U6295 ( .A(p_input[2370]), .B(p_input[1370]), .Z(n5597) );
  AND U6296 ( .A(p_input[4370]), .B(p_input[370]), .Z(n5595) );
  AND U6297 ( .A(n5598), .B(n5599), .Z(n5593) );
  AND U6298 ( .A(n5600), .B(p_input[7370]), .Z(n5599) );
  AND U6299 ( .A(p_input[6370]), .B(p_input[5370]), .Z(n5600) );
  AND U6300 ( .A(p_input[9370]), .B(p_input[8370]), .Z(n5598) );
  AND U6301 ( .A(n5601), .B(n5602), .Z(o[36]) );
  AND U6302 ( .A(n5603), .B(n5604), .Z(n5602) );
  AND U6303 ( .A(n5605), .B(p_input[3036]), .Z(n5604) );
  AND U6304 ( .A(p_input[2036]), .B(p_input[1036]), .Z(n5605) );
  AND U6305 ( .A(p_input[4036]), .B(p_input[36]), .Z(n5603) );
  AND U6306 ( .A(n5606), .B(n5607), .Z(n5601) );
  AND U6307 ( .A(n5608), .B(p_input[7036]), .Z(n5607) );
  AND U6308 ( .A(p_input[6036]), .B(p_input[5036]), .Z(n5608) );
  AND U6309 ( .A(p_input[9036]), .B(p_input[8036]), .Z(n5606) );
  AND U6310 ( .A(n5609), .B(n5610), .Z(o[369]) );
  AND U6311 ( .A(n5611), .B(n5612), .Z(n5610) );
  AND U6312 ( .A(n5613), .B(p_input[3369]), .Z(n5612) );
  AND U6313 ( .A(p_input[2369]), .B(p_input[1369]), .Z(n5613) );
  AND U6314 ( .A(p_input[4369]), .B(p_input[369]), .Z(n5611) );
  AND U6315 ( .A(n5614), .B(n5615), .Z(n5609) );
  AND U6316 ( .A(n5616), .B(p_input[7369]), .Z(n5615) );
  AND U6317 ( .A(p_input[6369]), .B(p_input[5369]), .Z(n5616) );
  AND U6318 ( .A(p_input[9369]), .B(p_input[8369]), .Z(n5614) );
  AND U6319 ( .A(n5617), .B(n5618), .Z(o[368]) );
  AND U6320 ( .A(n5619), .B(n5620), .Z(n5618) );
  AND U6321 ( .A(n5621), .B(p_input[3368]), .Z(n5620) );
  AND U6322 ( .A(p_input[2368]), .B(p_input[1368]), .Z(n5621) );
  AND U6323 ( .A(p_input[4368]), .B(p_input[368]), .Z(n5619) );
  AND U6324 ( .A(n5622), .B(n5623), .Z(n5617) );
  AND U6325 ( .A(n5624), .B(p_input[7368]), .Z(n5623) );
  AND U6326 ( .A(p_input[6368]), .B(p_input[5368]), .Z(n5624) );
  AND U6327 ( .A(p_input[9368]), .B(p_input[8368]), .Z(n5622) );
  AND U6328 ( .A(n5625), .B(n5626), .Z(o[367]) );
  AND U6329 ( .A(n5627), .B(n5628), .Z(n5626) );
  AND U6330 ( .A(n5629), .B(p_input[3367]), .Z(n5628) );
  AND U6331 ( .A(p_input[2367]), .B(p_input[1367]), .Z(n5629) );
  AND U6332 ( .A(p_input[4367]), .B(p_input[367]), .Z(n5627) );
  AND U6333 ( .A(n5630), .B(n5631), .Z(n5625) );
  AND U6334 ( .A(n5632), .B(p_input[7367]), .Z(n5631) );
  AND U6335 ( .A(p_input[6367]), .B(p_input[5367]), .Z(n5632) );
  AND U6336 ( .A(p_input[9367]), .B(p_input[8367]), .Z(n5630) );
  AND U6337 ( .A(n5633), .B(n5634), .Z(o[366]) );
  AND U6338 ( .A(n5635), .B(n5636), .Z(n5634) );
  AND U6339 ( .A(n5637), .B(p_input[3366]), .Z(n5636) );
  AND U6340 ( .A(p_input[2366]), .B(p_input[1366]), .Z(n5637) );
  AND U6341 ( .A(p_input[4366]), .B(p_input[366]), .Z(n5635) );
  AND U6342 ( .A(n5638), .B(n5639), .Z(n5633) );
  AND U6343 ( .A(n5640), .B(p_input[7366]), .Z(n5639) );
  AND U6344 ( .A(p_input[6366]), .B(p_input[5366]), .Z(n5640) );
  AND U6345 ( .A(p_input[9366]), .B(p_input[8366]), .Z(n5638) );
  AND U6346 ( .A(n5641), .B(n5642), .Z(o[365]) );
  AND U6347 ( .A(n5643), .B(n5644), .Z(n5642) );
  AND U6348 ( .A(n5645), .B(p_input[3365]), .Z(n5644) );
  AND U6349 ( .A(p_input[2365]), .B(p_input[1365]), .Z(n5645) );
  AND U6350 ( .A(p_input[4365]), .B(p_input[365]), .Z(n5643) );
  AND U6351 ( .A(n5646), .B(n5647), .Z(n5641) );
  AND U6352 ( .A(n5648), .B(p_input[7365]), .Z(n5647) );
  AND U6353 ( .A(p_input[6365]), .B(p_input[5365]), .Z(n5648) );
  AND U6354 ( .A(p_input[9365]), .B(p_input[8365]), .Z(n5646) );
  AND U6355 ( .A(n5649), .B(n5650), .Z(o[364]) );
  AND U6356 ( .A(n5651), .B(n5652), .Z(n5650) );
  AND U6357 ( .A(n5653), .B(p_input[3364]), .Z(n5652) );
  AND U6358 ( .A(p_input[2364]), .B(p_input[1364]), .Z(n5653) );
  AND U6359 ( .A(p_input[4364]), .B(p_input[364]), .Z(n5651) );
  AND U6360 ( .A(n5654), .B(n5655), .Z(n5649) );
  AND U6361 ( .A(n5656), .B(p_input[7364]), .Z(n5655) );
  AND U6362 ( .A(p_input[6364]), .B(p_input[5364]), .Z(n5656) );
  AND U6363 ( .A(p_input[9364]), .B(p_input[8364]), .Z(n5654) );
  AND U6364 ( .A(n5657), .B(n5658), .Z(o[363]) );
  AND U6365 ( .A(n5659), .B(n5660), .Z(n5658) );
  AND U6366 ( .A(n5661), .B(p_input[3363]), .Z(n5660) );
  AND U6367 ( .A(p_input[2363]), .B(p_input[1363]), .Z(n5661) );
  AND U6368 ( .A(p_input[4363]), .B(p_input[363]), .Z(n5659) );
  AND U6369 ( .A(n5662), .B(n5663), .Z(n5657) );
  AND U6370 ( .A(n5664), .B(p_input[7363]), .Z(n5663) );
  AND U6371 ( .A(p_input[6363]), .B(p_input[5363]), .Z(n5664) );
  AND U6372 ( .A(p_input[9363]), .B(p_input[8363]), .Z(n5662) );
  AND U6373 ( .A(n5665), .B(n5666), .Z(o[362]) );
  AND U6374 ( .A(n5667), .B(n5668), .Z(n5666) );
  AND U6375 ( .A(n5669), .B(p_input[3362]), .Z(n5668) );
  AND U6376 ( .A(p_input[2362]), .B(p_input[1362]), .Z(n5669) );
  AND U6377 ( .A(p_input[4362]), .B(p_input[362]), .Z(n5667) );
  AND U6378 ( .A(n5670), .B(n5671), .Z(n5665) );
  AND U6379 ( .A(n5672), .B(p_input[7362]), .Z(n5671) );
  AND U6380 ( .A(p_input[6362]), .B(p_input[5362]), .Z(n5672) );
  AND U6381 ( .A(p_input[9362]), .B(p_input[8362]), .Z(n5670) );
  AND U6382 ( .A(n5673), .B(n5674), .Z(o[361]) );
  AND U6383 ( .A(n5675), .B(n5676), .Z(n5674) );
  AND U6384 ( .A(n5677), .B(p_input[3361]), .Z(n5676) );
  AND U6385 ( .A(p_input[2361]), .B(p_input[1361]), .Z(n5677) );
  AND U6386 ( .A(p_input[4361]), .B(p_input[361]), .Z(n5675) );
  AND U6387 ( .A(n5678), .B(n5679), .Z(n5673) );
  AND U6388 ( .A(n5680), .B(p_input[7361]), .Z(n5679) );
  AND U6389 ( .A(p_input[6361]), .B(p_input[5361]), .Z(n5680) );
  AND U6390 ( .A(p_input[9361]), .B(p_input[8361]), .Z(n5678) );
  AND U6391 ( .A(n5681), .B(n5682), .Z(o[360]) );
  AND U6392 ( .A(n5683), .B(n5684), .Z(n5682) );
  AND U6393 ( .A(n5685), .B(p_input[3360]), .Z(n5684) );
  AND U6394 ( .A(p_input[2360]), .B(p_input[1360]), .Z(n5685) );
  AND U6395 ( .A(p_input[4360]), .B(p_input[360]), .Z(n5683) );
  AND U6396 ( .A(n5686), .B(n5687), .Z(n5681) );
  AND U6397 ( .A(n5688), .B(p_input[7360]), .Z(n5687) );
  AND U6398 ( .A(p_input[6360]), .B(p_input[5360]), .Z(n5688) );
  AND U6399 ( .A(p_input[9360]), .B(p_input[8360]), .Z(n5686) );
  AND U6400 ( .A(n5689), .B(n5690), .Z(o[35]) );
  AND U6401 ( .A(n5691), .B(n5692), .Z(n5690) );
  AND U6402 ( .A(n5693), .B(p_input[3035]), .Z(n5692) );
  AND U6403 ( .A(p_input[2035]), .B(p_input[1035]), .Z(n5693) );
  AND U6404 ( .A(p_input[4035]), .B(p_input[35]), .Z(n5691) );
  AND U6405 ( .A(n5694), .B(n5695), .Z(n5689) );
  AND U6406 ( .A(n5696), .B(p_input[7035]), .Z(n5695) );
  AND U6407 ( .A(p_input[6035]), .B(p_input[5035]), .Z(n5696) );
  AND U6408 ( .A(p_input[9035]), .B(p_input[8035]), .Z(n5694) );
  AND U6409 ( .A(n5697), .B(n5698), .Z(o[359]) );
  AND U6410 ( .A(n5699), .B(n5700), .Z(n5698) );
  AND U6411 ( .A(n5701), .B(p_input[3359]), .Z(n5700) );
  AND U6412 ( .A(p_input[2359]), .B(p_input[1359]), .Z(n5701) );
  AND U6413 ( .A(p_input[4359]), .B(p_input[359]), .Z(n5699) );
  AND U6414 ( .A(n5702), .B(n5703), .Z(n5697) );
  AND U6415 ( .A(n5704), .B(p_input[7359]), .Z(n5703) );
  AND U6416 ( .A(p_input[6359]), .B(p_input[5359]), .Z(n5704) );
  AND U6417 ( .A(p_input[9359]), .B(p_input[8359]), .Z(n5702) );
  AND U6418 ( .A(n5705), .B(n5706), .Z(o[358]) );
  AND U6419 ( .A(n5707), .B(n5708), .Z(n5706) );
  AND U6420 ( .A(n5709), .B(p_input[3358]), .Z(n5708) );
  AND U6421 ( .A(p_input[2358]), .B(p_input[1358]), .Z(n5709) );
  AND U6422 ( .A(p_input[4358]), .B(p_input[358]), .Z(n5707) );
  AND U6423 ( .A(n5710), .B(n5711), .Z(n5705) );
  AND U6424 ( .A(n5712), .B(p_input[7358]), .Z(n5711) );
  AND U6425 ( .A(p_input[6358]), .B(p_input[5358]), .Z(n5712) );
  AND U6426 ( .A(p_input[9358]), .B(p_input[8358]), .Z(n5710) );
  AND U6427 ( .A(n5713), .B(n5714), .Z(o[357]) );
  AND U6428 ( .A(n5715), .B(n5716), .Z(n5714) );
  AND U6429 ( .A(n5717), .B(p_input[3357]), .Z(n5716) );
  AND U6430 ( .A(p_input[2357]), .B(p_input[1357]), .Z(n5717) );
  AND U6431 ( .A(p_input[4357]), .B(p_input[357]), .Z(n5715) );
  AND U6432 ( .A(n5718), .B(n5719), .Z(n5713) );
  AND U6433 ( .A(n5720), .B(p_input[7357]), .Z(n5719) );
  AND U6434 ( .A(p_input[6357]), .B(p_input[5357]), .Z(n5720) );
  AND U6435 ( .A(p_input[9357]), .B(p_input[8357]), .Z(n5718) );
  AND U6436 ( .A(n5721), .B(n5722), .Z(o[356]) );
  AND U6437 ( .A(n5723), .B(n5724), .Z(n5722) );
  AND U6438 ( .A(n5725), .B(p_input[3356]), .Z(n5724) );
  AND U6439 ( .A(p_input[2356]), .B(p_input[1356]), .Z(n5725) );
  AND U6440 ( .A(p_input[4356]), .B(p_input[356]), .Z(n5723) );
  AND U6441 ( .A(n5726), .B(n5727), .Z(n5721) );
  AND U6442 ( .A(n5728), .B(p_input[7356]), .Z(n5727) );
  AND U6443 ( .A(p_input[6356]), .B(p_input[5356]), .Z(n5728) );
  AND U6444 ( .A(p_input[9356]), .B(p_input[8356]), .Z(n5726) );
  AND U6445 ( .A(n5729), .B(n5730), .Z(o[355]) );
  AND U6446 ( .A(n5731), .B(n5732), .Z(n5730) );
  AND U6447 ( .A(n5733), .B(p_input[3355]), .Z(n5732) );
  AND U6448 ( .A(p_input[2355]), .B(p_input[1355]), .Z(n5733) );
  AND U6449 ( .A(p_input[4355]), .B(p_input[355]), .Z(n5731) );
  AND U6450 ( .A(n5734), .B(n5735), .Z(n5729) );
  AND U6451 ( .A(n5736), .B(p_input[7355]), .Z(n5735) );
  AND U6452 ( .A(p_input[6355]), .B(p_input[5355]), .Z(n5736) );
  AND U6453 ( .A(p_input[9355]), .B(p_input[8355]), .Z(n5734) );
  AND U6454 ( .A(n5737), .B(n5738), .Z(o[354]) );
  AND U6455 ( .A(n5739), .B(n5740), .Z(n5738) );
  AND U6456 ( .A(n5741), .B(p_input[3354]), .Z(n5740) );
  AND U6457 ( .A(p_input[2354]), .B(p_input[1354]), .Z(n5741) );
  AND U6458 ( .A(p_input[4354]), .B(p_input[354]), .Z(n5739) );
  AND U6459 ( .A(n5742), .B(n5743), .Z(n5737) );
  AND U6460 ( .A(n5744), .B(p_input[7354]), .Z(n5743) );
  AND U6461 ( .A(p_input[6354]), .B(p_input[5354]), .Z(n5744) );
  AND U6462 ( .A(p_input[9354]), .B(p_input[8354]), .Z(n5742) );
  AND U6463 ( .A(n5745), .B(n5746), .Z(o[353]) );
  AND U6464 ( .A(n5747), .B(n5748), .Z(n5746) );
  AND U6465 ( .A(n5749), .B(p_input[3353]), .Z(n5748) );
  AND U6466 ( .A(p_input[2353]), .B(p_input[1353]), .Z(n5749) );
  AND U6467 ( .A(p_input[4353]), .B(p_input[353]), .Z(n5747) );
  AND U6468 ( .A(n5750), .B(n5751), .Z(n5745) );
  AND U6469 ( .A(n5752), .B(p_input[7353]), .Z(n5751) );
  AND U6470 ( .A(p_input[6353]), .B(p_input[5353]), .Z(n5752) );
  AND U6471 ( .A(p_input[9353]), .B(p_input[8353]), .Z(n5750) );
  AND U6472 ( .A(n5753), .B(n5754), .Z(o[352]) );
  AND U6473 ( .A(n5755), .B(n5756), .Z(n5754) );
  AND U6474 ( .A(n5757), .B(p_input[3352]), .Z(n5756) );
  AND U6475 ( .A(p_input[2352]), .B(p_input[1352]), .Z(n5757) );
  AND U6476 ( .A(p_input[4352]), .B(p_input[352]), .Z(n5755) );
  AND U6477 ( .A(n5758), .B(n5759), .Z(n5753) );
  AND U6478 ( .A(n5760), .B(p_input[7352]), .Z(n5759) );
  AND U6479 ( .A(p_input[6352]), .B(p_input[5352]), .Z(n5760) );
  AND U6480 ( .A(p_input[9352]), .B(p_input[8352]), .Z(n5758) );
  AND U6481 ( .A(n5761), .B(n5762), .Z(o[351]) );
  AND U6482 ( .A(n5763), .B(n5764), .Z(n5762) );
  AND U6483 ( .A(n5765), .B(p_input[3351]), .Z(n5764) );
  AND U6484 ( .A(p_input[2351]), .B(p_input[1351]), .Z(n5765) );
  AND U6485 ( .A(p_input[4351]), .B(p_input[351]), .Z(n5763) );
  AND U6486 ( .A(n5766), .B(n5767), .Z(n5761) );
  AND U6487 ( .A(n5768), .B(p_input[7351]), .Z(n5767) );
  AND U6488 ( .A(p_input[6351]), .B(p_input[5351]), .Z(n5768) );
  AND U6489 ( .A(p_input[9351]), .B(p_input[8351]), .Z(n5766) );
  AND U6490 ( .A(n5769), .B(n5770), .Z(o[350]) );
  AND U6491 ( .A(n5771), .B(n5772), .Z(n5770) );
  AND U6492 ( .A(n5773), .B(p_input[3350]), .Z(n5772) );
  AND U6493 ( .A(p_input[2350]), .B(p_input[1350]), .Z(n5773) );
  AND U6494 ( .A(p_input[4350]), .B(p_input[350]), .Z(n5771) );
  AND U6495 ( .A(n5774), .B(n5775), .Z(n5769) );
  AND U6496 ( .A(n5776), .B(p_input[7350]), .Z(n5775) );
  AND U6497 ( .A(p_input[6350]), .B(p_input[5350]), .Z(n5776) );
  AND U6498 ( .A(p_input[9350]), .B(p_input[8350]), .Z(n5774) );
  AND U6499 ( .A(n5777), .B(n5778), .Z(o[34]) );
  AND U6500 ( .A(n5779), .B(n5780), .Z(n5778) );
  AND U6501 ( .A(n5781), .B(p_input[3034]), .Z(n5780) );
  AND U6502 ( .A(p_input[2034]), .B(p_input[1034]), .Z(n5781) );
  AND U6503 ( .A(p_input[4034]), .B(p_input[34]), .Z(n5779) );
  AND U6504 ( .A(n5782), .B(n5783), .Z(n5777) );
  AND U6505 ( .A(n5784), .B(p_input[7034]), .Z(n5783) );
  AND U6506 ( .A(p_input[6034]), .B(p_input[5034]), .Z(n5784) );
  AND U6507 ( .A(p_input[9034]), .B(p_input[8034]), .Z(n5782) );
  AND U6508 ( .A(n5785), .B(n5786), .Z(o[349]) );
  AND U6509 ( .A(n5787), .B(n5788), .Z(n5786) );
  AND U6510 ( .A(n5789), .B(p_input[3349]), .Z(n5788) );
  AND U6511 ( .A(p_input[2349]), .B(p_input[1349]), .Z(n5789) );
  AND U6512 ( .A(p_input[4349]), .B(p_input[349]), .Z(n5787) );
  AND U6513 ( .A(n5790), .B(n5791), .Z(n5785) );
  AND U6514 ( .A(n5792), .B(p_input[7349]), .Z(n5791) );
  AND U6515 ( .A(p_input[6349]), .B(p_input[5349]), .Z(n5792) );
  AND U6516 ( .A(p_input[9349]), .B(p_input[8349]), .Z(n5790) );
  AND U6517 ( .A(n5793), .B(n5794), .Z(o[348]) );
  AND U6518 ( .A(n5795), .B(n5796), .Z(n5794) );
  AND U6519 ( .A(n5797), .B(p_input[3348]), .Z(n5796) );
  AND U6520 ( .A(p_input[2348]), .B(p_input[1348]), .Z(n5797) );
  AND U6521 ( .A(p_input[4348]), .B(p_input[348]), .Z(n5795) );
  AND U6522 ( .A(n5798), .B(n5799), .Z(n5793) );
  AND U6523 ( .A(n5800), .B(p_input[7348]), .Z(n5799) );
  AND U6524 ( .A(p_input[6348]), .B(p_input[5348]), .Z(n5800) );
  AND U6525 ( .A(p_input[9348]), .B(p_input[8348]), .Z(n5798) );
  AND U6526 ( .A(n5801), .B(n5802), .Z(o[347]) );
  AND U6527 ( .A(n5803), .B(n5804), .Z(n5802) );
  AND U6528 ( .A(n5805), .B(p_input[3347]), .Z(n5804) );
  AND U6529 ( .A(p_input[2347]), .B(p_input[1347]), .Z(n5805) );
  AND U6530 ( .A(p_input[4347]), .B(p_input[347]), .Z(n5803) );
  AND U6531 ( .A(n5806), .B(n5807), .Z(n5801) );
  AND U6532 ( .A(n5808), .B(p_input[7347]), .Z(n5807) );
  AND U6533 ( .A(p_input[6347]), .B(p_input[5347]), .Z(n5808) );
  AND U6534 ( .A(p_input[9347]), .B(p_input[8347]), .Z(n5806) );
  AND U6535 ( .A(n5809), .B(n5810), .Z(o[346]) );
  AND U6536 ( .A(n5811), .B(n5812), .Z(n5810) );
  AND U6537 ( .A(n5813), .B(p_input[3346]), .Z(n5812) );
  AND U6538 ( .A(p_input[2346]), .B(p_input[1346]), .Z(n5813) );
  AND U6539 ( .A(p_input[4346]), .B(p_input[346]), .Z(n5811) );
  AND U6540 ( .A(n5814), .B(n5815), .Z(n5809) );
  AND U6541 ( .A(n5816), .B(p_input[7346]), .Z(n5815) );
  AND U6542 ( .A(p_input[6346]), .B(p_input[5346]), .Z(n5816) );
  AND U6543 ( .A(p_input[9346]), .B(p_input[8346]), .Z(n5814) );
  AND U6544 ( .A(n5817), .B(n5818), .Z(o[345]) );
  AND U6545 ( .A(n5819), .B(n5820), .Z(n5818) );
  AND U6546 ( .A(n5821), .B(p_input[3345]), .Z(n5820) );
  AND U6547 ( .A(p_input[2345]), .B(p_input[1345]), .Z(n5821) );
  AND U6548 ( .A(p_input[4345]), .B(p_input[345]), .Z(n5819) );
  AND U6549 ( .A(n5822), .B(n5823), .Z(n5817) );
  AND U6550 ( .A(n5824), .B(p_input[7345]), .Z(n5823) );
  AND U6551 ( .A(p_input[6345]), .B(p_input[5345]), .Z(n5824) );
  AND U6552 ( .A(p_input[9345]), .B(p_input[8345]), .Z(n5822) );
  AND U6553 ( .A(n5825), .B(n5826), .Z(o[344]) );
  AND U6554 ( .A(n5827), .B(n5828), .Z(n5826) );
  AND U6555 ( .A(n5829), .B(p_input[3344]), .Z(n5828) );
  AND U6556 ( .A(p_input[2344]), .B(p_input[1344]), .Z(n5829) );
  AND U6557 ( .A(p_input[4344]), .B(p_input[344]), .Z(n5827) );
  AND U6558 ( .A(n5830), .B(n5831), .Z(n5825) );
  AND U6559 ( .A(n5832), .B(p_input[7344]), .Z(n5831) );
  AND U6560 ( .A(p_input[6344]), .B(p_input[5344]), .Z(n5832) );
  AND U6561 ( .A(p_input[9344]), .B(p_input[8344]), .Z(n5830) );
  AND U6562 ( .A(n5833), .B(n5834), .Z(o[343]) );
  AND U6563 ( .A(n5835), .B(n5836), .Z(n5834) );
  AND U6564 ( .A(n5837), .B(p_input[3343]), .Z(n5836) );
  AND U6565 ( .A(p_input[2343]), .B(p_input[1343]), .Z(n5837) );
  AND U6566 ( .A(p_input[4343]), .B(p_input[343]), .Z(n5835) );
  AND U6567 ( .A(n5838), .B(n5839), .Z(n5833) );
  AND U6568 ( .A(n5840), .B(p_input[7343]), .Z(n5839) );
  AND U6569 ( .A(p_input[6343]), .B(p_input[5343]), .Z(n5840) );
  AND U6570 ( .A(p_input[9343]), .B(p_input[8343]), .Z(n5838) );
  AND U6571 ( .A(n5841), .B(n5842), .Z(o[342]) );
  AND U6572 ( .A(n5843), .B(n5844), .Z(n5842) );
  AND U6573 ( .A(n5845), .B(p_input[3342]), .Z(n5844) );
  AND U6574 ( .A(p_input[2342]), .B(p_input[1342]), .Z(n5845) );
  AND U6575 ( .A(p_input[4342]), .B(p_input[342]), .Z(n5843) );
  AND U6576 ( .A(n5846), .B(n5847), .Z(n5841) );
  AND U6577 ( .A(n5848), .B(p_input[7342]), .Z(n5847) );
  AND U6578 ( .A(p_input[6342]), .B(p_input[5342]), .Z(n5848) );
  AND U6579 ( .A(p_input[9342]), .B(p_input[8342]), .Z(n5846) );
  AND U6580 ( .A(n5849), .B(n5850), .Z(o[341]) );
  AND U6581 ( .A(n5851), .B(n5852), .Z(n5850) );
  AND U6582 ( .A(n5853), .B(p_input[3341]), .Z(n5852) );
  AND U6583 ( .A(p_input[2341]), .B(p_input[1341]), .Z(n5853) );
  AND U6584 ( .A(p_input[4341]), .B(p_input[341]), .Z(n5851) );
  AND U6585 ( .A(n5854), .B(n5855), .Z(n5849) );
  AND U6586 ( .A(n5856), .B(p_input[7341]), .Z(n5855) );
  AND U6587 ( .A(p_input[6341]), .B(p_input[5341]), .Z(n5856) );
  AND U6588 ( .A(p_input[9341]), .B(p_input[8341]), .Z(n5854) );
  AND U6589 ( .A(n5857), .B(n5858), .Z(o[340]) );
  AND U6590 ( .A(n5859), .B(n5860), .Z(n5858) );
  AND U6591 ( .A(n5861), .B(p_input[3340]), .Z(n5860) );
  AND U6592 ( .A(p_input[2340]), .B(p_input[1340]), .Z(n5861) );
  AND U6593 ( .A(p_input[4340]), .B(p_input[340]), .Z(n5859) );
  AND U6594 ( .A(n5862), .B(n5863), .Z(n5857) );
  AND U6595 ( .A(n5864), .B(p_input[7340]), .Z(n5863) );
  AND U6596 ( .A(p_input[6340]), .B(p_input[5340]), .Z(n5864) );
  AND U6597 ( .A(p_input[9340]), .B(p_input[8340]), .Z(n5862) );
  AND U6598 ( .A(n5865), .B(n5866), .Z(o[33]) );
  AND U6599 ( .A(n5867), .B(n5868), .Z(n5866) );
  AND U6600 ( .A(n5869), .B(p_input[3033]), .Z(n5868) );
  AND U6601 ( .A(p_input[2033]), .B(p_input[1033]), .Z(n5869) );
  AND U6602 ( .A(p_input[4033]), .B(p_input[33]), .Z(n5867) );
  AND U6603 ( .A(n5870), .B(n5871), .Z(n5865) );
  AND U6604 ( .A(n5872), .B(p_input[7033]), .Z(n5871) );
  AND U6605 ( .A(p_input[6033]), .B(p_input[5033]), .Z(n5872) );
  AND U6606 ( .A(p_input[9033]), .B(p_input[8033]), .Z(n5870) );
  AND U6607 ( .A(n5873), .B(n5874), .Z(o[339]) );
  AND U6608 ( .A(n5875), .B(n5876), .Z(n5874) );
  AND U6609 ( .A(n5877), .B(p_input[3339]), .Z(n5876) );
  AND U6610 ( .A(p_input[2339]), .B(p_input[1339]), .Z(n5877) );
  AND U6611 ( .A(p_input[4339]), .B(p_input[339]), .Z(n5875) );
  AND U6612 ( .A(n5878), .B(n5879), .Z(n5873) );
  AND U6613 ( .A(n5880), .B(p_input[7339]), .Z(n5879) );
  AND U6614 ( .A(p_input[6339]), .B(p_input[5339]), .Z(n5880) );
  AND U6615 ( .A(p_input[9339]), .B(p_input[8339]), .Z(n5878) );
  AND U6616 ( .A(n5881), .B(n5882), .Z(o[338]) );
  AND U6617 ( .A(n5883), .B(n5884), .Z(n5882) );
  AND U6618 ( .A(n5885), .B(p_input[3338]), .Z(n5884) );
  AND U6619 ( .A(p_input[2338]), .B(p_input[1338]), .Z(n5885) );
  AND U6620 ( .A(p_input[4338]), .B(p_input[338]), .Z(n5883) );
  AND U6621 ( .A(n5886), .B(n5887), .Z(n5881) );
  AND U6622 ( .A(n5888), .B(p_input[7338]), .Z(n5887) );
  AND U6623 ( .A(p_input[6338]), .B(p_input[5338]), .Z(n5888) );
  AND U6624 ( .A(p_input[9338]), .B(p_input[8338]), .Z(n5886) );
  AND U6625 ( .A(n5889), .B(n5890), .Z(o[337]) );
  AND U6626 ( .A(n5891), .B(n5892), .Z(n5890) );
  AND U6627 ( .A(n5893), .B(p_input[3337]), .Z(n5892) );
  AND U6628 ( .A(p_input[2337]), .B(p_input[1337]), .Z(n5893) );
  AND U6629 ( .A(p_input[4337]), .B(p_input[337]), .Z(n5891) );
  AND U6630 ( .A(n5894), .B(n5895), .Z(n5889) );
  AND U6631 ( .A(n5896), .B(p_input[7337]), .Z(n5895) );
  AND U6632 ( .A(p_input[6337]), .B(p_input[5337]), .Z(n5896) );
  AND U6633 ( .A(p_input[9337]), .B(p_input[8337]), .Z(n5894) );
  AND U6634 ( .A(n5897), .B(n5898), .Z(o[336]) );
  AND U6635 ( .A(n5899), .B(n5900), .Z(n5898) );
  AND U6636 ( .A(n5901), .B(p_input[3336]), .Z(n5900) );
  AND U6637 ( .A(p_input[2336]), .B(p_input[1336]), .Z(n5901) );
  AND U6638 ( .A(p_input[4336]), .B(p_input[336]), .Z(n5899) );
  AND U6639 ( .A(n5902), .B(n5903), .Z(n5897) );
  AND U6640 ( .A(n5904), .B(p_input[7336]), .Z(n5903) );
  AND U6641 ( .A(p_input[6336]), .B(p_input[5336]), .Z(n5904) );
  AND U6642 ( .A(p_input[9336]), .B(p_input[8336]), .Z(n5902) );
  AND U6643 ( .A(n5905), .B(n5906), .Z(o[335]) );
  AND U6644 ( .A(n5907), .B(n5908), .Z(n5906) );
  AND U6645 ( .A(n5909), .B(p_input[3335]), .Z(n5908) );
  AND U6646 ( .A(p_input[2335]), .B(p_input[1335]), .Z(n5909) );
  AND U6647 ( .A(p_input[4335]), .B(p_input[335]), .Z(n5907) );
  AND U6648 ( .A(n5910), .B(n5911), .Z(n5905) );
  AND U6649 ( .A(n5912), .B(p_input[7335]), .Z(n5911) );
  AND U6650 ( .A(p_input[6335]), .B(p_input[5335]), .Z(n5912) );
  AND U6651 ( .A(p_input[9335]), .B(p_input[8335]), .Z(n5910) );
  AND U6652 ( .A(n5913), .B(n5914), .Z(o[334]) );
  AND U6653 ( .A(n5915), .B(n5916), .Z(n5914) );
  AND U6654 ( .A(n5917), .B(p_input[3334]), .Z(n5916) );
  AND U6655 ( .A(p_input[2334]), .B(p_input[1334]), .Z(n5917) );
  AND U6656 ( .A(p_input[4334]), .B(p_input[334]), .Z(n5915) );
  AND U6657 ( .A(n5918), .B(n5919), .Z(n5913) );
  AND U6658 ( .A(n5920), .B(p_input[7334]), .Z(n5919) );
  AND U6659 ( .A(p_input[6334]), .B(p_input[5334]), .Z(n5920) );
  AND U6660 ( .A(p_input[9334]), .B(p_input[8334]), .Z(n5918) );
  AND U6661 ( .A(n5921), .B(n5922), .Z(o[333]) );
  AND U6662 ( .A(n5923), .B(n5924), .Z(n5922) );
  AND U6663 ( .A(n5925), .B(p_input[3333]), .Z(n5924) );
  AND U6664 ( .A(p_input[2333]), .B(p_input[1333]), .Z(n5925) );
  AND U6665 ( .A(p_input[4333]), .B(p_input[333]), .Z(n5923) );
  AND U6666 ( .A(n5926), .B(n5927), .Z(n5921) );
  AND U6667 ( .A(n5928), .B(p_input[7333]), .Z(n5927) );
  AND U6668 ( .A(p_input[6333]), .B(p_input[5333]), .Z(n5928) );
  AND U6669 ( .A(p_input[9333]), .B(p_input[8333]), .Z(n5926) );
  AND U6670 ( .A(n5929), .B(n5930), .Z(o[332]) );
  AND U6671 ( .A(n5931), .B(n5932), .Z(n5930) );
  AND U6672 ( .A(n5933), .B(p_input[332]), .Z(n5932) );
  AND U6673 ( .A(p_input[2332]), .B(p_input[1332]), .Z(n5933) );
  AND U6674 ( .A(p_input[4332]), .B(p_input[3332]), .Z(n5931) );
  AND U6675 ( .A(n5934), .B(n5935), .Z(n5929) );
  AND U6676 ( .A(n5936), .B(p_input[7332]), .Z(n5935) );
  AND U6677 ( .A(p_input[6332]), .B(p_input[5332]), .Z(n5936) );
  AND U6678 ( .A(p_input[9332]), .B(p_input[8332]), .Z(n5934) );
  AND U6679 ( .A(n5937), .B(n5938), .Z(o[331]) );
  AND U6680 ( .A(n5939), .B(n5940), .Z(n5938) );
  AND U6681 ( .A(n5941), .B(p_input[331]), .Z(n5940) );
  AND U6682 ( .A(p_input[2331]), .B(p_input[1331]), .Z(n5941) );
  AND U6683 ( .A(p_input[4331]), .B(p_input[3331]), .Z(n5939) );
  AND U6684 ( .A(n5942), .B(n5943), .Z(n5937) );
  AND U6685 ( .A(n5944), .B(p_input[7331]), .Z(n5943) );
  AND U6686 ( .A(p_input[6331]), .B(p_input[5331]), .Z(n5944) );
  AND U6687 ( .A(p_input[9331]), .B(p_input[8331]), .Z(n5942) );
  AND U6688 ( .A(n5945), .B(n5946), .Z(o[330]) );
  AND U6689 ( .A(n5947), .B(n5948), .Z(n5946) );
  AND U6690 ( .A(n5949), .B(p_input[330]), .Z(n5948) );
  AND U6691 ( .A(p_input[2330]), .B(p_input[1330]), .Z(n5949) );
  AND U6692 ( .A(p_input[4330]), .B(p_input[3330]), .Z(n5947) );
  AND U6693 ( .A(n5950), .B(n5951), .Z(n5945) );
  AND U6694 ( .A(n5952), .B(p_input[7330]), .Z(n5951) );
  AND U6695 ( .A(p_input[6330]), .B(p_input[5330]), .Z(n5952) );
  AND U6696 ( .A(p_input[9330]), .B(p_input[8330]), .Z(n5950) );
  AND U6697 ( .A(n5953), .B(n5954), .Z(o[32]) );
  AND U6698 ( .A(n5955), .B(n5956), .Z(n5954) );
  AND U6699 ( .A(n5957), .B(p_input[3032]), .Z(n5956) );
  AND U6700 ( .A(p_input[2032]), .B(p_input[1032]), .Z(n5957) );
  AND U6701 ( .A(p_input[4032]), .B(p_input[32]), .Z(n5955) );
  AND U6702 ( .A(n5958), .B(n5959), .Z(n5953) );
  AND U6703 ( .A(n5960), .B(p_input[7032]), .Z(n5959) );
  AND U6704 ( .A(p_input[6032]), .B(p_input[5032]), .Z(n5960) );
  AND U6705 ( .A(p_input[9032]), .B(p_input[8032]), .Z(n5958) );
  AND U6706 ( .A(n5961), .B(n5962), .Z(o[329]) );
  AND U6707 ( .A(n5963), .B(n5964), .Z(n5962) );
  AND U6708 ( .A(n5965), .B(p_input[329]), .Z(n5964) );
  AND U6709 ( .A(p_input[2329]), .B(p_input[1329]), .Z(n5965) );
  AND U6710 ( .A(p_input[4329]), .B(p_input[3329]), .Z(n5963) );
  AND U6711 ( .A(n5966), .B(n5967), .Z(n5961) );
  AND U6712 ( .A(n5968), .B(p_input[7329]), .Z(n5967) );
  AND U6713 ( .A(p_input[6329]), .B(p_input[5329]), .Z(n5968) );
  AND U6714 ( .A(p_input[9329]), .B(p_input[8329]), .Z(n5966) );
  AND U6715 ( .A(n5969), .B(n5970), .Z(o[328]) );
  AND U6716 ( .A(n5971), .B(n5972), .Z(n5970) );
  AND U6717 ( .A(n5973), .B(p_input[328]), .Z(n5972) );
  AND U6718 ( .A(p_input[2328]), .B(p_input[1328]), .Z(n5973) );
  AND U6719 ( .A(p_input[4328]), .B(p_input[3328]), .Z(n5971) );
  AND U6720 ( .A(n5974), .B(n5975), .Z(n5969) );
  AND U6721 ( .A(n5976), .B(p_input[7328]), .Z(n5975) );
  AND U6722 ( .A(p_input[6328]), .B(p_input[5328]), .Z(n5976) );
  AND U6723 ( .A(p_input[9328]), .B(p_input[8328]), .Z(n5974) );
  AND U6724 ( .A(n5977), .B(n5978), .Z(o[327]) );
  AND U6725 ( .A(n5979), .B(n5980), .Z(n5978) );
  AND U6726 ( .A(n5981), .B(p_input[327]), .Z(n5980) );
  AND U6727 ( .A(p_input[2327]), .B(p_input[1327]), .Z(n5981) );
  AND U6728 ( .A(p_input[4327]), .B(p_input[3327]), .Z(n5979) );
  AND U6729 ( .A(n5982), .B(n5983), .Z(n5977) );
  AND U6730 ( .A(n5984), .B(p_input[7327]), .Z(n5983) );
  AND U6731 ( .A(p_input[6327]), .B(p_input[5327]), .Z(n5984) );
  AND U6732 ( .A(p_input[9327]), .B(p_input[8327]), .Z(n5982) );
  AND U6733 ( .A(n5985), .B(n5986), .Z(o[326]) );
  AND U6734 ( .A(n5987), .B(n5988), .Z(n5986) );
  AND U6735 ( .A(n5989), .B(p_input[326]), .Z(n5988) );
  AND U6736 ( .A(p_input[2326]), .B(p_input[1326]), .Z(n5989) );
  AND U6737 ( .A(p_input[4326]), .B(p_input[3326]), .Z(n5987) );
  AND U6738 ( .A(n5990), .B(n5991), .Z(n5985) );
  AND U6739 ( .A(n5992), .B(p_input[7326]), .Z(n5991) );
  AND U6740 ( .A(p_input[6326]), .B(p_input[5326]), .Z(n5992) );
  AND U6741 ( .A(p_input[9326]), .B(p_input[8326]), .Z(n5990) );
  AND U6742 ( .A(n5993), .B(n5994), .Z(o[325]) );
  AND U6743 ( .A(n5995), .B(n5996), .Z(n5994) );
  AND U6744 ( .A(n5997), .B(p_input[325]), .Z(n5996) );
  AND U6745 ( .A(p_input[2325]), .B(p_input[1325]), .Z(n5997) );
  AND U6746 ( .A(p_input[4325]), .B(p_input[3325]), .Z(n5995) );
  AND U6747 ( .A(n5998), .B(n5999), .Z(n5993) );
  AND U6748 ( .A(n6000), .B(p_input[7325]), .Z(n5999) );
  AND U6749 ( .A(p_input[6325]), .B(p_input[5325]), .Z(n6000) );
  AND U6750 ( .A(p_input[9325]), .B(p_input[8325]), .Z(n5998) );
  AND U6751 ( .A(n6001), .B(n6002), .Z(o[324]) );
  AND U6752 ( .A(n6003), .B(n6004), .Z(n6002) );
  AND U6753 ( .A(n6005), .B(p_input[324]), .Z(n6004) );
  AND U6754 ( .A(p_input[2324]), .B(p_input[1324]), .Z(n6005) );
  AND U6755 ( .A(p_input[4324]), .B(p_input[3324]), .Z(n6003) );
  AND U6756 ( .A(n6006), .B(n6007), .Z(n6001) );
  AND U6757 ( .A(n6008), .B(p_input[7324]), .Z(n6007) );
  AND U6758 ( .A(p_input[6324]), .B(p_input[5324]), .Z(n6008) );
  AND U6759 ( .A(p_input[9324]), .B(p_input[8324]), .Z(n6006) );
  AND U6760 ( .A(n6009), .B(n6010), .Z(o[323]) );
  AND U6761 ( .A(n6011), .B(n6012), .Z(n6010) );
  AND U6762 ( .A(n6013), .B(p_input[323]), .Z(n6012) );
  AND U6763 ( .A(p_input[2323]), .B(p_input[1323]), .Z(n6013) );
  AND U6764 ( .A(p_input[4323]), .B(p_input[3323]), .Z(n6011) );
  AND U6765 ( .A(n6014), .B(n6015), .Z(n6009) );
  AND U6766 ( .A(n6016), .B(p_input[7323]), .Z(n6015) );
  AND U6767 ( .A(p_input[6323]), .B(p_input[5323]), .Z(n6016) );
  AND U6768 ( .A(p_input[9323]), .B(p_input[8323]), .Z(n6014) );
  AND U6769 ( .A(n6017), .B(n6018), .Z(o[322]) );
  AND U6770 ( .A(n6019), .B(n6020), .Z(n6018) );
  AND U6771 ( .A(n6021), .B(p_input[322]), .Z(n6020) );
  AND U6772 ( .A(p_input[2322]), .B(p_input[1322]), .Z(n6021) );
  AND U6773 ( .A(p_input[4322]), .B(p_input[3322]), .Z(n6019) );
  AND U6774 ( .A(n6022), .B(n6023), .Z(n6017) );
  AND U6775 ( .A(n6024), .B(p_input[7322]), .Z(n6023) );
  AND U6776 ( .A(p_input[6322]), .B(p_input[5322]), .Z(n6024) );
  AND U6777 ( .A(p_input[9322]), .B(p_input[8322]), .Z(n6022) );
  AND U6778 ( .A(n6025), .B(n6026), .Z(o[321]) );
  AND U6779 ( .A(n6027), .B(n6028), .Z(n6026) );
  AND U6780 ( .A(n6029), .B(p_input[321]), .Z(n6028) );
  AND U6781 ( .A(p_input[2321]), .B(p_input[1321]), .Z(n6029) );
  AND U6782 ( .A(p_input[4321]), .B(p_input[3321]), .Z(n6027) );
  AND U6783 ( .A(n6030), .B(n6031), .Z(n6025) );
  AND U6784 ( .A(n6032), .B(p_input[7321]), .Z(n6031) );
  AND U6785 ( .A(p_input[6321]), .B(p_input[5321]), .Z(n6032) );
  AND U6786 ( .A(p_input[9321]), .B(p_input[8321]), .Z(n6030) );
  AND U6787 ( .A(n6033), .B(n6034), .Z(o[320]) );
  AND U6788 ( .A(n6035), .B(n6036), .Z(n6034) );
  AND U6789 ( .A(n6037), .B(p_input[320]), .Z(n6036) );
  AND U6790 ( .A(p_input[2320]), .B(p_input[1320]), .Z(n6037) );
  AND U6791 ( .A(p_input[4320]), .B(p_input[3320]), .Z(n6035) );
  AND U6792 ( .A(n6038), .B(n6039), .Z(n6033) );
  AND U6793 ( .A(n6040), .B(p_input[7320]), .Z(n6039) );
  AND U6794 ( .A(p_input[6320]), .B(p_input[5320]), .Z(n6040) );
  AND U6795 ( .A(p_input[9320]), .B(p_input[8320]), .Z(n6038) );
  AND U6796 ( .A(n6041), .B(n6042), .Z(o[31]) );
  AND U6797 ( .A(n6043), .B(n6044), .Z(n6042) );
  AND U6798 ( .A(n6045), .B(p_input[3031]), .Z(n6044) );
  AND U6799 ( .A(p_input[2031]), .B(p_input[1031]), .Z(n6045) );
  AND U6800 ( .A(p_input[4031]), .B(p_input[31]), .Z(n6043) );
  AND U6801 ( .A(n6046), .B(n6047), .Z(n6041) );
  AND U6802 ( .A(n6048), .B(p_input[7031]), .Z(n6047) );
  AND U6803 ( .A(p_input[6031]), .B(p_input[5031]), .Z(n6048) );
  AND U6804 ( .A(p_input[9031]), .B(p_input[8031]), .Z(n6046) );
  AND U6805 ( .A(n6049), .B(n6050), .Z(o[319]) );
  AND U6806 ( .A(n6051), .B(n6052), .Z(n6050) );
  AND U6807 ( .A(n6053), .B(p_input[319]), .Z(n6052) );
  AND U6808 ( .A(p_input[2319]), .B(p_input[1319]), .Z(n6053) );
  AND U6809 ( .A(p_input[4319]), .B(p_input[3319]), .Z(n6051) );
  AND U6810 ( .A(n6054), .B(n6055), .Z(n6049) );
  AND U6811 ( .A(n6056), .B(p_input[7319]), .Z(n6055) );
  AND U6812 ( .A(p_input[6319]), .B(p_input[5319]), .Z(n6056) );
  AND U6813 ( .A(p_input[9319]), .B(p_input[8319]), .Z(n6054) );
  AND U6814 ( .A(n6057), .B(n6058), .Z(o[318]) );
  AND U6815 ( .A(n6059), .B(n6060), .Z(n6058) );
  AND U6816 ( .A(n6061), .B(p_input[318]), .Z(n6060) );
  AND U6817 ( .A(p_input[2318]), .B(p_input[1318]), .Z(n6061) );
  AND U6818 ( .A(p_input[4318]), .B(p_input[3318]), .Z(n6059) );
  AND U6819 ( .A(n6062), .B(n6063), .Z(n6057) );
  AND U6820 ( .A(n6064), .B(p_input[7318]), .Z(n6063) );
  AND U6821 ( .A(p_input[6318]), .B(p_input[5318]), .Z(n6064) );
  AND U6822 ( .A(p_input[9318]), .B(p_input[8318]), .Z(n6062) );
  AND U6823 ( .A(n6065), .B(n6066), .Z(o[317]) );
  AND U6824 ( .A(n6067), .B(n6068), .Z(n6066) );
  AND U6825 ( .A(n6069), .B(p_input[317]), .Z(n6068) );
  AND U6826 ( .A(p_input[2317]), .B(p_input[1317]), .Z(n6069) );
  AND U6827 ( .A(p_input[4317]), .B(p_input[3317]), .Z(n6067) );
  AND U6828 ( .A(n6070), .B(n6071), .Z(n6065) );
  AND U6829 ( .A(n6072), .B(p_input[7317]), .Z(n6071) );
  AND U6830 ( .A(p_input[6317]), .B(p_input[5317]), .Z(n6072) );
  AND U6831 ( .A(p_input[9317]), .B(p_input[8317]), .Z(n6070) );
  AND U6832 ( .A(n6073), .B(n6074), .Z(o[316]) );
  AND U6833 ( .A(n6075), .B(n6076), .Z(n6074) );
  AND U6834 ( .A(n6077), .B(p_input[316]), .Z(n6076) );
  AND U6835 ( .A(p_input[2316]), .B(p_input[1316]), .Z(n6077) );
  AND U6836 ( .A(p_input[4316]), .B(p_input[3316]), .Z(n6075) );
  AND U6837 ( .A(n6078), .B(n6079), .Z(n6073) );
  AND U6838 ( .A(n6080), .B(p_input[7316]), .Z(n6079) );
  AND U6839 ( .A(p_input[6316]), .B(p_input[5316]), .Z(n6080) );
  AND U6840 ( .A(p_input[9316]), .B(p_input[8316]), .Z(n6078) );
  AND U6841 ( .A(n6081), .B(n6082), .Z(o[315]) );
  AND U6842 ( .A(n6083), .B(n6084), .Z(n6082) );
  AND U6843 ( .A(n6085), .B(p_input[315]), .Z(n6084) );
  AND U6844 ( .A(p_input[2315]), .B(p_input[1315]), .Z(n6085) );
  AND U6845 ( .A(p_input[4315]), .B(p_input[3315]), .Z(n6083) );
  AND U6846 ( .A(n6086), .B(n6087), .Z(n6081) );
  AND U6847 ( .A(n6088), .B(p_input[7315]), .Z(n6087) );
  AND U6848 ( .A(p_input[6315]), .B(p_input[5315]), .Z(n6088) );
  AND U6849 ( .A(p_input[9315]), .B(p_input[8315]), .Z(n6086) );
  AND U6850 ( .A(n6089), .B(n6090), .Z(o[314]) );
  AND U6851 ( .A(n6091), .B(n6092), .Z(n6090) );
  AND U6852 ( .A(n6093), .B(p_input[314]), .Z(n6092) );
  AND U6853 ( .A(p_input[2314]), .B(p_input[1314]), .Z(n6093) );
  AND U6854 ( .A(p_input[4314]), .B(p_input[3314]), .Z(n6091) );
  AND U6855 ( .A(n6094), .B(n6095), .Z(n6089) );
  AND U6856 ( .A(n6096), .B(p_input[7314]), .Z(n6095) );
  AND U6857 ( .A(p_input[6314]), .B(p_input[5314]), .Z(n6096) );
  AND U6858 ( .A(p_input[9314]), .B(p_input[8314]), .Z(n6094) );
  AND U6859 ( .A(n6097), .B(n6098), .Z(o[313]) );
  AND U6860 ( .A(n6099), .B(n6100), .Z(n6098) );
  AND U6861 ( .A(n6101), .B(p_input[313]), .Z(n6100) );
  AND U6862 ( .A(p_input[2313]), .B(p_input[1313]), .Z(n6101) );
  AND U6863 ( .A(p_input[4313]), .B(p_input[3313]), .Z(n6099) );
  AND U6864 ( .A(n6102), .B(n6103), .Z(n6097) );
  AND U6865 ( .A(n6104), .B(p_input[7313]), .Z(n6103) );
  AND U6866 ( .A(p_input[6313]), .B(p_input[5313]), .Z(n6104) );
  AND U6867 ( .A(p_input[9313]), .B(p_input[8313]), .Z(n6102) );
  AND U6868 ( .A(n6105), .B(n6106), .Z(o[312]) );
  AND U6869 ( .A(n6107), .B(n6108), .Z(n6106) );
  AND U6870 ( .A(n6109), .B(p_input[312]), .Z(n6108) );
  AND U6871 ( .A(p_input[2312]), .B(p_input[1312]), .Z(n6109) );
  AND U6872 ( .A(p_input[4312]), .B(p_input[3312]), .Z(n6107) );
  AND U6873 ( .A(n6110), .B(n6111), .Z(n6105) );
  AND U6874 ( .A(n6112), .B(p_input[7312]), .Z(n6111) );
  AND U6875 ( .A(p_input[6312]), .B(p_input[5312]), .Z(n6112) );
  AND U6876 ( .A(p_input[9312]), .B(p_input[8312]), .Z(n6110) );
  AND U6877 ( .A(n6113), .B(n6114), .Z(o[311]) );
  AND U6878 ( .A(n6115), .B(n6116), .Z(n6114) );
  AND U6879 ( .A(n6117), .B(p_input[311]), .Z(n6116) );
  AND U6880 ( .A(p_input[2311]), .B(p_input[1311]), .Z(n6117) );
  AND U6881 ( .A(p_input[4311]), .B(p_input[3311]), .Z(n6115) );
  AND U6882 ( .A(n6118), .B(n6119), .Z(n6113) );
  AND U6883 ( .A(n6120), .B(p_input[7311]), .Z(n6119) );
  AND U6884 ( .A(p_input[6311]), .B(p_input[5311]), .Z(n6120) );
  AND U6885 ( .A(p_input[9311]), .B(p_input[8311]), .Z(n6118) );
  AND U6886 ( .A(n6121), .B(n6122), .Z(o[310]) );
  AND U6887 ( .A(n6123), .B(n6124), .Z(n6122) );
  AND U6888 ( .A(n6125), .B(p_input[310]), .Z(n6124) );
  AND U6889 ( .A(p_input[2310]), .B(p_input[1310]), .Z(n6125) );
  AND U6890 ( .A(p_input[4310]), .B(p_input[3310]), .Z(n6123) );
  AND U6891 ( .A(n6126), .B(n6127), .Z(n6121) );
  AND U6892 ( .A(n6128), .B(p_input[7310]), .Z(n6127) );
  AND U6893 ( .A(p_input[6310]), .B(p_input[5310]), .Z(n6128) );
  AND U6894 ( .A(p_input[9310]), .B(p_input[8310]), .Z(n6126) );
  AND U6895 ( .A(n6129), .B(n6130), .Z(o[30]) );
  AND U6896 ( .A(n6131), .B(n6132), .Z(n6130) );
  AND U6897 ( .A(n6133), .B(p_input[3030]), .Z(n6132) );
  AND U6898 ( .A(p_input[2030]), .B(p_input[1030]), .Z(n6133) );
  AND U6899 ( .A(p_input[4030]), .B(p_input[30]), .Z(n6131) );
  AND U6900 ( .A(n6134), .B(n6135), .Z(n6129) );
  AND U6901 ( .A(n6136), .B(p_input[7030]), .Z(n6135) );
  AND U6902 ( .A(p_input[6030]), .B(p_input[5030]), .Z(n6136) );
  AND U6903 ( .A(p_input[9030]), .B(p_input[8030]), .Z(n6134) );
  AND U6904 ( .A(n6137), .B(n6138), .Z(o[309]) );
  AND U6905 ( .A(n6139), .B(n6140), .Z(n6138) );
  AND U6906 ( .A(n6141), .B(p_input[309]), .Z(n6140) );
  AND U6907 ( .A(p_input[2309]), .B(p_input[1309]), .Z(n6141) );
  AND U6908 ( .A(p_input[4309]), .B(p_input[3309]), .Z(n6139) );
  AND U6909 ( .A(n6142), .B(n6143), .Z(n6137) );
  AND U6910 ( .A(n6144), .B(p_input[7309]), .Z(n6143) );
  AND U6911 ( .A(p_input[6309]), .B(p_input[5309]), .Z(n6144) );
  AND U6912 ( .A(p_input[9309]), .B(p_input[8309]), .Z(n6142) );
  AND U6913 ( .A(n6145), .B(n6146), .Z(o[308]) );
  AND U6914 ( .A(n6147), .B(n6148), .Z(n6146) );
  AND U6915 ( .A(n6149), .B(p_input[308]), .Z(n6148) );
  AND U6916 ( .A(p_input[2308]), .B(p_input[1308]), .Z(n6149) );
  AND U6917 ( .A(p_input[4308]), .B(p_input[3308]), .Z(n6147) );
  AND U6918 ( .A(n6150), .B(n6151), .Z(n6145) );
  AND U6919 ( .A(n6152), .B(p_input[7308]), .Z(n6151) );
  AND U6920 ( .A(p_input[6308]), .B(p_input[5308]), .Z(n6152) );
  AND U6921 ( .A(p_input[9308]), .B(p_input[8308]), .Z(n6150) );
  AND U6922 ( .A(n6153), .B(n6154), .Z(o[307]) );
  AND U6923 ( .A(n6155), .B(n6156), .Z(n6154) );
  AND U6924 ( .A(n6157), .B(p_input[307]), .Z(n6156) );
  AND U6925 ( .A(p_input[2307]), .B(p_input[1307]), .Z(n6157) );
  AND U6926 ( .A(p_input[4307]), .B(p_input[3307]), .Z(n6155) );
  AND U6927 ( .A(n6158), .B(n6159), .Z(n6153) );
  AND U6928 ( .A(n6160), .B(p_input[7307]), .Z(n6159) );
  AND U6929 ( .A(p_input[6307]), .B(p_input[5307]), .Z(n6160) );
  AND U6930 ( .A(p_input[9307]), .B(p_input[8307]), .Z(n6158) );
  AND U6931 ( .A(n6161), .B(n6162), .Z(o[306]) );
  AND U6932 ( .A(n6163), .B(n6164), .Z(n6162) );
  AND U6933 ( .A(n6165), .B(p_input[306]), .Z(n6164) );
  AND U6934 ( .A(p_input[2306]), .B(p_input[1306]), .Z(n6165) );
  AND U6935 ( .A(p_input[4306]), .B(p_input[3306]), .Z(n6163) );
  AND U6936 ( .A(n6166), .B(n6167), .Z(n6161) );
  AND U6937 ( .A(n6168), .B(p_input[7306]), .Z(n6167) );
  AND U6938 ( .A(p_input[6306]), .B(p_input[5306]), .Z(n6168) );
  AND U6939 ( .A(p_input[9306]), .B(p_input[8306]), .Z(n6166) );
  AND U6940 ( .A(n6169), .B(n6170), .Z(o[305]) );
  AND U6941 ( .A(n6171), .B(n6172), .Z(n6170) );
  AND U6942 ( .A(n6173), .B(p_input[305]), .Z(n6172) );
  AND U6943 ( .A(p_input[2305]), .B(p_input[1305]), .Z(n6173) );
  AND U6944 ( .A(p_input[4305]), .B(p_input[3305]), .Z(n6171) );
  AND U6945 ( .A(n6174), .B(n6175), .Z(n6169) );
  AND U6946 ( .A(n6176), .B(p_input[7305]), .Z(n6175) );
  AND U6947 ( .A(p_input[6305]), .B(p_input[5305]), .Z(n6176) );
  AND U6948 ( .A(p_input[9305]), .B(p_input[8305]), .Z(n6174) );
  AND U6949 ( .A(n6177), .B(n6178), .Z(o[304]) );
  AND U6950 ( .A(n6179), .B(n6180), .Z(n6178) );
  AND U6951 ( .A(n6181), .B(p_input[304]), .Z(n6180) );
  AND U6952 ( .A(p_input[2304]), .B(p_input[1304]), .Z(n6181) );
  AND U6953 ( .A(p_input[4304]), .B(p_input[3304]), .Z(n6179) );
  AND U6954 ( .A(n6182), .B(n6183), .Z(n6177) );
  AND U6955 ( .A(n6184), .B(p_input[7304]), .Z(n6183) );
  AND U6956 ( .A(p_input[6304]), .B(p_input[5304]), .Z(n6184) );
  AND U6957 ( .A(p_input[9304]), .B(p_input[8304]), .Z(n6182) );
  AND U6958 ( .A(n6185), .B(n6186), .Z(o[303]) );
  AND U6959 ( .A(n6187), .B(n6188), .Z(n6186) );
  AND U6960 ( .A(n6189), .B(p_input[303]), .Z(n6188) );
  AND U6961 ( .A(p_input[2303]), .B(p_input[1303]), .Z(n6189) );
  AND U6962 ( .A(p_input[4303]), .B(p_input[3303]), .Z(n6187) );
  AND U6963 ( .A(n6190), .B(n6191), .Z(n6185) );
  AND U6964 ( .A(n6192), .B(p_input[7303]), .Z(n6191) );
  AND U6965 ( .A(p_input[6303]), .B(p_input[5303]), .Z(n6192) );
  AND U6966 ( .A(p_input[9303]), .B(p_input[8303]), .Z(n6190) );
  AND U6967 ( .A(n6193), .B(n6194), .Z(o[302]) );
  AND U6968 ( .A(n6195), .B(n6196), .Z(n6194) );
  AND U6969 ( .A(n6197), .B(p_input[302]), .Z(n6196) );
  AND U6970 ( .A(p_input[2302]), .B(p_input[1302]), .Z(n6197) );
  AND U6971 ( .A(p_input[4302]), .B(p_input[3302]), .Z(n6195) );
  AND U6972 ( .A(n6198), .B(n6199), .Z(n6193) );
  AND U6973 ( .A(n6200), .B(p_input[7302]), .Z(n6199) );
  AND U6974 ( .A(p_input[6302]), .B(p_input[5302]), .Z(n6200) );
  AND U6975 ( .A(p_input[9302]), .B(p_input[8302]), .Z(n6198) );
  AND U6976 ( .A(n6201), .B(n6202), .Z(o[301]) );
  AND U6977 ( .A(n6203), .B(n6204), .Z(n6202) );
  AND U6978 ( .A(n6205), .B(p_input[301]), .Z(n6204) );
  AND U6979 ( .A(p_input[2301]), .B(p_input[1301]), .Z(n6205) );
  AND U6980 ( .A(p_input[4301]), .B(p_input[3301]), .Z(n6203) );
  AND U6981 ( .A(n6206), .B(n6207), .Z(n6201) );
  AND U6982 ( .A(n6208), .B(p_input[7301]), .Z(n6207) );
  AND U6983 ( .A(p_input[6301]), .B(p_input[5301]), .Z(n6208) );
  AND U6984 ( .A(p_input[9301]), .B(p_input[8301]), .Z(n6206) );
  AND U6985 ( .A(n6209), .B(n6210), .Z(o[300]) );
  AND U6986 ( .A(n6211), .B(n6212), .Z(n6210) );
  AND U6987 ( .A(n6213), .B(p_input[300]), .Z(n6212) );
  AND U6988 ( .A(p_input[2300]), .B(p_input[1300]), .Z(n6213) );
  AND U6989 ( .A(p_input[4300]), .B(p_input[3300]), .Z(n6211) );
  AND U6990 ( .A(n6214), .B(n6215), .Z(n6209) );
  AND U6991 ( .A(n6216), .B(p_input[7300]), .Z(n6215) );
  AND U6992 ( .A(p_input[6300]), .B(p_input[5300]), .Z(n6216) );
  AND U6993 ( .A(p_input[9300]), .B(p_input[8300]), .Z(n6214) );
  AND U6994 ( .A(n6217), .B(n6218), .Z(o[2]) );
  AND U6995 ( .A(n6219), .B(n6220), .Z(n6218) );
  AND U6996 ( .A(n6221), .B(p_input[2]), .Z(n6220) );
  AND U6997 ( .A(p_input[2002]), .B(p_input[1002]), .Z(n6221) );
  AND U6998 ( .A(p_input[4002]), .B(p_input[3002]), .Z(n6219) );
  AND U6999 ( .A(n6222), .B(n6223), .Z(n6217) );
  AND U7000 ( .A(n6224), .B(p_input[7002]), .Z(n6223) );
  AND U7001 ( .A(p_input[6002]), .B(p_input[5002]), .Z(n6224) );
  AND U7002 ( .A(p_input[9002]), .B(p_input[8002]), .Z(n6222) );
  AND U7003 ( .A(n6225), .B(n6226), .Z(o[29]) );
  AND U7004 ( .A(n6227), .B(n6228), .Z(n6226) );
  AND U7005 ( .A(n6229), .B(p_input[29]), .Z(n6228) );
  AND U7006 ( .A(p_input[2029]), .B(p_input[1029]), .Z(n6229) );
  AND U7007 ( .A(p_input[4029]), .B(p_input[3029]), .Z(n6227) );
  AND U7008 ( .A(n6230), .B(n6231), .Z(n6225) );
  AND U7009 ( .A(n6232), .B(p_input[7029]), .Z(n6231) );
  AND U7010 ( .A(p_input[6029]), .B(p_input[5029]), .Z(n6232) );
  AND U7011 ( .A(p_input[9029]), .B(p_input[8029]), .Z(n6230) );
  AND U7012 ( .A(n6233), .B(n6234), .Z(o[299]) );
  AND U7013 ( .A(n6235), .B(n6236), .Z(n6234) );
  AND U7014 ( .A(n6237), .B(p_input[299]), .Z(n6236) );
  AND U7015 ( .A(p_input[2299]), .B(p_input[1299]), .Z(n6237) );
  AND U7016 ( .A(p_input[4299]), .B(p_input[3299]), .Z(n6235) );
  AND U7017 ( .A(n6238), .B(n6239), .Z(n6233) );
  AND U7018 ( .A(n6240), .B(p_input[7299]), .Z(n6239) );
  AND U7019 ( .A(p_input[6299]), .B(p_input[5299]), .Z(n6240) );
  AND U7020 ( .A(p_input[9299]), .B(p_input[8299]), .Z(n6238) );
  AND U7021 ( .A(n6241), .B(n6242), .Z(o[298]) );
  AND U7022 ( .A(n6243), .B(n6244), .Z(n6242) );
  AND U7023 ( .A(n6245), .B(p_input[298]), .Z(n6244) );
  AND U7024 ( .A(p_input[2298]), .B(p_input[1298]), .Z(n6245) );
  AND U7025 ( .A(p_input[4298]), .B(p_input[3298]), .Z(n6243) );
  AND U7026 ( .A(n6246), .B(n6247), .Z(n6241) );
  AND U7027 ( .A(n6248), .B(p_input[7298]), .Z(n6247) );
  AND U7028 ( .A(p_input[6298]), .B(p_input[5298]), .Z(n6248) );
  AND U7029 ( .A(p_input[9298]), .B(p_input[8298]), .Z(n6246) );
  AND U7030 ( .A(n6249), .B(n6250), .Z(o[297]) );
  AND U7031 ( .A(n6251), .B(n6252), .Z(n6250) );
  AND U7032 ( .A(n6253), .B(p_input[297]), .Z(n6252) );
  AND U7033 ( .A(p_input[2297]), .B(p_input[1297]), .Z(n6253) );
  AND U7034 ( .A(p_input[4297]), .B(p_input[3297]), .Z(n6251) );
  AND U7035 ( .A(n6254), .B(n6255), .Z(n6249) );
  AND U7036 ( .A(n6256), .B(p_input[7297]), .Z(n6255) );
  AND U7037 ( .A(p_input[6297]), .B(p_input[5297]), .Z(n6256) );
  AND U7038 ( .A(p_input[9297]), .B(p_input[8297]), .Z(n6254) );
  AND U7039 ( .A(n6257), .B(n6258), .Z(o[296]) );
  AND U7040 ( .A(n6259), .B(n6260), .Z(n6258) );
  AND U7041 ( .A(n6261), .B(p_input[296]), .Z(n6260) );
  AND U7042 ( .A(p_input[2296]), .B(p_input[1296]), .Z(n6261) );
  AND U7043 ( .A(p_input[4296]), .B(p_input[3296]), .Z(n6259) );
  AND U7044 ( .A(n6262), .B(n6263), .Z(n6257) );
  AND U7045 ( .A(n6264), .B(p_input[7296]), .Z(n6263) );
  AND U7046 ( .A(p_input[6296]), .B(p_input[5296]), .Z(n6264) );
  AND U7047 ( .A(p_input[9296]), .B(p_input[8296]), .Z(n6262) );
  AND U7048 ( .A(n6265), .B(n6266), .Z(o[295]) );
  AND U7049 ( .A(n6267), .B(n6268), .Z(n6266) );
  AND U7050 ( .A(n6269), .B(p_input[295]), .Z(n6268) );
  AND U7051 ( .A(p_input[2295]), .B(p_input[1295]), .Z(n6269) );
  AND U7052 ( .A(p_input[4295]), .B(p_input[3295]), .Z(n6267) );
  AND U7053 ( .A(n6270), .B(n6271), .Z(n6265) );
  AND U7054 ( .A(n6272), .B(p_input[7295]), .Z(n6271) );
  AND U7055 ( .A(p_input[6295]), .B(p_input[5295]), .Z(n6272) );
  AND U7056 ( .A(p_input[9295]), .B(p_input[8295]), .Z(n6270) );
  AND U7057 ( .A(n6273), .B(n6274), .Z(o[294]) );
  AND U7058 ( .A(n6275), .B(n6276), .Z(n6274) );
  AND U7059 ( .A(n6277), .B(p_input[294]), .Z(n6276) );
  AND U7060 ( .A(p_input[2294]), .B(p_input[1294]), .Z(n6277) );
  AND U7061 ( .A(p_input[4294]), .B(p_input[3294]), .Z(n6275) );
  AND U7062 ( .A(n6278), .B(n6279), .Z(n6273) );
  AND U7063 ( .A(n6280), .B(p_input[7294]), .Z(n6279) );
  AND U7064 ( .A(p_input[6294]), .B(p_input[5294]), .Z(n6280) );
  AND U7065 ( .A(p_input[9294]), .B(p_input[8294]), .Z(n6278) );
  AND U7066 ( .A(n6281), .B(n6282), .Z(o[293]) );
  AND U7067 ( .A(n6283), .B(n6284), .Z(n6282) );
  AND U7068 ( .A(n6285), .B(p_input[293]), .Z(n6284) );
  AND U7069 ( .A(p_input[2293]), .B(p_input[1293]), .Z(n6285) );
  AND U7070 ( .A(p_input[4293]), .B(p_input[3293]), .Z(n6283) );
  AND U7071 ( .A(n6286), .B(n6287), .Z(n6281) );
  AND U7072 ( .A(n6288), .B(p_input[7293]), .Z(n6287) );
  AND U7073 ( .A(p_input[6293]), .B(p_input[5293]), .Z(n6288) );
  AND U7074 ( .A(p_input[9293]), .B(p_input[8293]), .Z(n6286) );
  AND U7075 ( .A(n6289), .B(n6290), .Z(o[292]) );
  AND U7076 ( .A(n6291), .B(n6292), .Z(n6290) );
  AND U7077 ( .A(n6293), .B(p_input[292]), .Z(n6292) );
  AND U7078 ( .A(p_input[2292]), .B(p_input[1292]), .Z(n6293) );
  AND U7079 ( .A(p_input[4292]), .B(p_input[3292]), .Z(n6291) );
  AND U7080 ( .A(n6294), .B(n6295), .Z(n6289) );
  AND U7081 ( .A(n6296), .B(p_input[7292]), .Z(n6295) );
  AND U7082 ( .A(p_input[6292]), .B(p_input[5292]), .Z(n6296) );
  AND U7083 ( .A(p_input[9292]), .B(p_input[8292]), .Z(n6294) );
  AND U7084 ( .A(n6297), .B(n6298), .Z(o[291]) );
  AND U7085 ( .A(n6299), .B(n6300), .Z(n6298) );
  AND U7086 ( .A(n6301), .B(p_input[291]), .Z(n6300) );
  AND U7087 ( .A(p_input[2291]), .B(p_input[1291]), .Z(n6301) );
  AND U7088 ( .A(p_input[4291]), .B(p_input[3291]), .Z(n6299) );
  AND U7089 ( .A(n6302), .B(n6303), .Z(n6297) );
  AND U7090 ( .A(n6304), .B(p_input[7291]), .Z(n6303) );
  AND U7091 ( .A(p_input[6291]), .B(p_input[5291]), .Z(n6304) );
  AND U7092 ( .A(p_input[9291]), .B(p_input[8291]), .Z(n6302) );
  AND U7093 ( .A(n6305), .B(n6306), .Z(o[290]) );
  AND U7094 ( .A(n6307), .B(n6308), .Z(n6306) );
  AND U7095 ( .A(n6309), .B(p_input[290]), .Z(n6308) );
  AND U7096 ( .A(p_input[2290]), .B(p_input[1290]), .Z(n6309) );
  AND U7097 ( .A(p_input[4290]), .B(p_input[3290]), .Z(n6307) );
  AND U7098 ( .A(n6310), .B(n6311), .Z(n6305) );
  AND U7099 ( .A(n6312), .B(p_input[7290]), .Z(n6311) );
  AND U7100 ( .A(p_input[6290]), .B(p_input[5290]), .Z(n6312) );
  AND U7101 ( .A(p_input[9290]), .B(p_input[8290]), .Z(n6310) );
  AND U7102 ( .A(n6313), .B(n6314), .Z(o[28]) );
  AND U7103 ( .A(n6315), .B(n6316), .Z(n6314) );
  AND U7104 ( .A(n6317), .B(p_input[28]), .Z(n6316) );
  AND U7105 ( .A(p_input[2028]), .B(p_input[1028]), .Z(n6317) );
  AND U7106 ( .A(p_input[4028]), .B(p_input[3028]), .Z(n6315) );
  AND U7107 ( .A(n6318), .B(n6319), .Z(n6313) );
  AND U7108 ( .A(n6320), .B(p_input[7028]), .Z(n6319) );
  AND U7109 ( .A(p_input[6028]), .B(p_input[5028]), .Z(n6320) );
  AND U7110 ( .A(p_input[9028]), .B(p_input[8028]), .Z(n6318) );
  AND U7111 ( .A(n6321), .B(n6322), .Z(o[289]) );
  AND U7112 ( .A(n6323), .B(n6324), .Z(n6322) );
  AND U7113 ( .A(n6325), .B(p_input[289]), .Z(n6324) );
  AND U7114 ( .A(p_input[2289]), .B(p_input[1289]), .Z(n6325) );
  AND U7115 ( .A(p_input[4289]), .B(p_input[3289]), .Z(n6323) );
  AND U7116 ( .A(n6326), .B(n6327), .Z(n6321) );
  AND U7117 ( .A(n6328), .B(p_input[7289]), .Z(n6327) );
  AND U7118 ( .A(p_input[6289]), .B(p_input[5289]), .Z(n6328) );
  AND U7119 ( .A(p_input[9289]), .B(p_input[8289]), .Z(n6326) );
  AND U7120 ( .A(n6329), .B(n6330), .Z(o[288]) );
  AND U7121 ( .A(n6331), .B(n6332), .Z(n6330) );
  AND U7122 ( .A(n6333), .B(p_input[288]), .Z(n6332) );
  AND U7123 ( .A(p_input[2288]), .B(p_input[1288]), .Z(n6333) );
  AND U7124 ( .A(p_input[4288]), .B(p_input[3288]), .Z(n6331) );
  AND U7125 ( .A(n6334), .B(n6335), .Z(n6329) );
  AND U7126 ( .A(n6336), .B(p_input[7288]), .Z(n6335) );
  AND U7127 ( .A(p_input[6288]), .B(p_input[5288]), .Z(n6336) );
  AND U7128 ( .A(p_input[9288]), .B(p_input[8288]), .Z(n6334) );
  AND U7129 ( .A(n6337), .B(n6338), .Z(o[287]) );
  AND U7130 ( .A(n6339), .B(n6340), .Z(n6338) );
  AND U7131 ( .A(n6341), .B(p_input[287]), .Z(n6340) );
  AND U7132 ( .A(p_input[2287]), .B(p_input[1287]), .Z(n6341) );
  AND U7133 ( .A(p_input[4287]), .B(p_input[3287]), .Z(n6339) );
  AND U7134 ( .A(n6342), .B(n6343), .Z(n6337) );
  AND U7135 ( .A(n6344), .B(p_input[7287]), .Z(n6343) );
  AND U7136 ( .A(p_input[6287]), .B(p_input[5287]), .Z(n6344) );
  AND U7137 ( .A(p_input[9287]), .B(p_input[8287]), .Z(n6342) );
  AND U7138 ( .A(n6345), .B(n6346), .Z(o[286]) );
  AND U7139 ( .A(n6347), .B(n6348), .Z(n6346) );
  AND U7140 ( .A(n6349), .B(p_input[286]), .Z(n6348) );
  AND U7141 ( .A(p_input[2286]), .B(p_input[1286]), .Z(n6349) );
  AND U7142 ( .A(p_input[4286]), .B(p_input[3286]), .Z(n6347) );
  AND U7143 ( .A(n6350), .B(n6351), .Z(n6345) );
  AND U7144 ( .A(n6352), .B(p_input[7286]), .Z(n6351) );
  AND U7145 ( .A(p_input[6286]), .B(p_input[5286]), .Z(n6352) );
  AND U7146 ( .A(p_input[9286]), .B(p_input[8286]), .Z(n6350) );
  AND U7147 ( .A(n6353), .B(n6354), .Z(o[285]) );
  AND U7148 ( .A(n6355), .B(n6356), .Z(n6354) );
  AND U7149 ( .A(n6357), .B(p_input[285]), .Z(n6356) );
  AND U7150 ( .A(p_input[2285]), .B(p_input[1285]), .Z(n6357) );
  AND U7151 ( .A(p_input[4285]), .B(p_input[3285]), .Z(n6355) );
  AND U7152 ( .A(n6358), .B(n6359), .Z(n6353) );
  AND U7153 ( .A(n6360), .B(p_input[7285]), .Z(n6359) );
  AND U7154 ( .A(p_input[6285]), .B(p_input[5285]), .Z(n6360) );
  AND U7155 ( .A(p_input[9285]), .B(p_input[8285]), .Z(n6358) );
  AND U7156 ( .A(n6361), .B(n6362), .Z(o[284]) );
  AND U7157 ( .A(n6363), .B(n6364), .Z(n6362) );
  AND U7158 ( .A(n6365), .B(p_input[284]), .Z(n6364) );
  AND U7159 ( .A(p_input[2284]), .B(p_input[1284]), .Z(n6365) );
  AND U7160 ( .A(p_input[4284]), .B(p_input[3284]), .Z(n6363) );
  AND U7161 ( .A(n6366), .B(n6367), .Z(n6361) );
  AND U7162 ( .A(n6368), .B(p_input[7284]), .Z(n6367) );
  AND U7163 ( .A(p_input[6284]), .B(p_input[5284]), .Z(n6368) );
  AND U7164 ( .A(p_input[9284]), .B(p_input[8284]), .Z(n6366) );
  AND U7165 ( .A(n6369), .B(n6370), .Z(o[283]) );
  AND U7166 ( .A(n6371), .B(n6372), .Z(n6370) );
  AND U7167 ( .A(n6373), .B(p_input[283]), .Z(n6372) );
  AND U7168 ( .A(p_input[2283]), .B(p_input[1283]), .Z(n6373) );
  AND U7169 ( .A(p_input[4283]), .B(p_input[3283]), .Z(n6371) );
  AND U7170 ( .A(n6374), .B(n6375), .Z(n6369) );
  AND U7171 ( .A(n6376), .B(p_input[7283]), .Z(n6375) );
  AND U7172 ( .A(p_input[6283]), .B(p_input[5283]), .Z(n6376) );
  AND U7173 ( .A(p_input[9283]), .B(p_input[8283]), .Z(n6374) );
  AND U7174 ( .A(n6377), .B(n6378), .Z(o[282]) );
  AND U7175 ( .A(n6379), .B(n6380), .Z(n6378) );
  AND U7176 ( .A(n6381), .B(p_input[282]), .Z(n6380) );
  AND U7177 ( .A(p_input[2282]), .B(p_input[1282]), .Z(n6381) );
  AND U7178 ( .A(p_input[4282]), .B(p_input[3282]), .Z(n6379) );
  AND U7179 ( .A(n6382), .B(n6383), .Z(n6377) );
  AND U7180 ( .A(n6384), .B(p_input[7282]), .Z(n6383) );
  AND U7181 ( .A(p_input[6282]), .B(p_input[5282]), .Z(n6384) );
  AND U7182 ( .A(p_input[9282]), .B(p_input[8282]), .Z(n6382) );
  AND U7183 ( .A(n6385), .B(n6386), .Z(o[281]) );
  AND U7184 ( .A(n6387), .B(n6388), .Z(n6386) );
  AND U7185 ( .A(n6389), .B(p_input[281]), .Z(n6388) );
  AND U7186 ( .A(p_input[2281]), .B(p_input[1281]), .Z(n6389) );
  AND U7187 ( .A(p_input[4281]), .B(p_input[3281]), .Z(n6387) );
  AND U7188 ( .A(n6390), .B(n6391), .Z(n6385) );
  AND U7189 ( .A(n6392), .B(p_input[7281]), .Z(n6391) );
  AND U7190 ( .A(p_input[6281]), .B(p_input[5281]), .Z(n6392) );
  AND U7191 ( .A(p_input[9281]), .B(p_input[8281]), .Z(n6390) );
  AND U7192 ( .A(n6393), .B(n6394), .Z(o[280]) );
  AND U7193 ( .A(n6395), .B(n6396), .Z(n6394) );
  AND U7194 ( .A(n6397), .B(p_input[280]), .Z(n6396) );
  AND U7195 ( .A(p_input[2280]), .B(p_input[1280]), .Z(n6397) );
  AND U7196 ( .A(p_input[4280]), .B(p_input[3280]), .Z(n6395) );
  AND U7197 ( .A(n6398), .B(n6399), .Z(n6393) );
  AND U7198 ( .A(n6400), .B(p_input[7280]), .Z(n6399) );
  AND U7199 ( .A(p_input[6280]), .B(p_input[5280]), .Z(n6400) );
  AND U7200 ( .A(p_input[9280]), .B(p_input[8280]), .Z(n6398) );
  AND U7201 ( .A(n6401), .B(n6402), .Z(o[27]) );
  AND U7202 ( .A(n6403), .B(n6404), .Z(n6402) );
  AND U7203 ( .A(n6405), .B(p_input[27]), .Z(n6404) );
  AND U7204 ( .A(p_input[2027]), .B(p_input[1027]), .Z(n6405) );
  AND U7205 ( .A(p_input[4027]), .B(p_input[3027]), .Z(n6403) );
  AND U7206 ( .A(n6406), .B(n6407), .Z(n6401) );
  AND U7207 ( .A(n6408), .B(p_input[7027]), .Z(n6407) );
  AND U7208 ( .A(p_input[6027]), .B(p_input[5027]), .Z(n6408) );
  AND U7209 ( .A(p_input[9027]), .B(p_input[8027]), .Z(n6406) );
  AND U7210 ( .A(n6409), .B(n6410), .Z(o[279]) );
  AND U7211 ( .A(n6411), .B(n6412), .Z(n6410) );
  AND U7212 ( .A(n6413), .B(p_input[279]), .Z(n6412) );
  AND U7213 ( .A(p_input[2279]), .B(p_input[1279]), .Z(n6413) );
  AND U7214 ( .A(p_input[4279]), .B(p_input[3279]), .Z(n6411) );
  AND U7215 ( .A(n6414), .B(n6415), .Z(n6409) );
  AND U7216 ( .A(n6416), .B(p_input[7279]), .Z(n6415) );
  AND U7217 ( .A(p_input[6279]), .B(p_input[5279]), .Z(n6416) );
  AND U7218 ( .A(p_input[9279]), .B(p_input[8279]), .Z(n6414) );
  AND U7219 ( .A(n6417), .B(n6418), .Z(o[278]) );
  AND U7220 ( .A(n6419), .B(n6420), .Z(n6418) );
  AND U7221 ( .A(n6421), .B(p_input[278]), .Z(n6420) );
  AND U7222 ( .A(p_input[2278]), .B(p_input[1278]), .Z(n6421) );
  AND U7223 ( .A(p_input[4278]), .B(p_input[3278]), .Z(n6419) );
  AND U7224 ( .A(n6422), .B(n6423), .Z(n6417) );
  AND U7225 ( .A(n6424), .B(p_input[7278]), .Z(n6423) );
  AND U7226 ( .A(p_input[6278]), .B(p_input[5278]), .Z(n6424) );
  AND U7227 ( .A(p_input[9278]), .B(p_input[8278]), .Z(n6422) );
  AND U7228 ( .A(n6425), .B(n6426), .Z(o[277]) );
  AND U7229 ( .A(n6427), .B(n6428), .Z(n6426) );
  AND U7230 ( .A(n6429), .B(p_input[277]), .Z(n6428) );
  AND U7231 ( .A(p_input[2277]), .B(p_input[1277]), .Z(n6429) );
  AND U7232 ( .A(p_input[4277]), .B(p_input[3277]), .Z(n6427) );
  AND U7233 ( .A(n6430), .B(n6431), .Z(n6425) );
  AND U7234 ( .A(n6432), .B(p_input[7277]), .Z(n6431) );
  AND U7235 ( .A(p_input[6277]), .B(p_input[5277]), .Z(n6432) );
  AND U7236 ( .A(p_input[9277]), .B(p_input[8277]), .Z(n6430) );
  AND U7237 ( .A(n6433), .B(n6434), .Z(o[276]) );
  AND U7238 ( .A(n6435), .B(n6436), .Z(n6434) );
  AND U7239 ( .A(n6437), .B(p_input[276]), .Z(n6436) );
  AND U7240 ( .A(p_input[2276]), .B(p_input[1276]), .Z(n6437) );
  AND U7241 ( .A(p_input[4276]), .B(p_input[3276]), .Z(n6435) );
  AND U7242 ( .A(n6438), .B(n6439), .Z(n6433) );
  AND U7243 ( .A(n6440), .B(p_input[7276]), .Z(n6439) );
  AND U7244 ( .A(p_input[6276]), .B(p_input[5276]), .Z(n6440) );
  AND U7245 ( .A(p_input[9276]), .B(p_input[8276]), .Z(n6438) );
  AND U7246 ( .A(n6441), .B(n6442), .Z(o[275]) );
  AND U7247 ( .A(n6443), .B(n6444), .Z(n6442) );
  AND U7248 ( .A(n6445), .B(p_input[275]), .Z(n6444) );
  AND U7249 ( .A(p_input[2275]), .B(p_input[1275]), .Z(n6445) );
  AND U7250 ( .A(p_input[4275]), .B(p_input[3275]), .Z(n6443) );
  AND U7251 ( .A(n6446), .B(n6447), .Z(n6441) );
  AND U7252 ( .A(n6448), .B(p_input[7275]), .Z(n6447) );
  AND U7253 ( .A(p_input[6275]), .B(p_input[5275]), .Z(n6448) );
  AND U7254 ( .A(p_input[9275]), .B(p_input[8275]), .Z(n6446) );
  AND U7255 ( .A(n6449), .B(n6450), .Z(o[274]) );
  AND U7256 ( .A(n6451), .B(n6452), .Z(n6450) );
  AND U7257 ( .A(n6453), .B(p_input[274]), .Z(n6452) );
  AND U7258 ( .A(p_input[2274]), .B(p_input[1274]), .Z(n6453) );
  AND U7259 ( .A(p_input[4274]), .B(p_input[3274]), .Z(n6451) );
  AND U7260 ( .A(n6454), .B(n6455), .Z(n6449) );
  AND U7261 ( .A(n6456), .B(p_input[7274]), .Z(n6455) );
  AND U7262 ( .A(p_input[6274]), .B(p_input[5274]), .Z(n6456) );
  AND U7263 ( .A(p_input[9274]), .B(p_input[8274]), .Z(n6454) );
  AND U7264 ( .A(n6457), .B(n6458), .Z(o[273]) );
  AND U7265 ( .A(n6459), .B(n6460), .Z(n6458) );
  AND U7266 ( .A(n6461), .B(p_input[273]), .Z(n6460) );
  AND U7267 ( .A(p_input[2273]), .B(p_input[1273]), .Z(n6461) );
  AND U7268 ( .A(p_input[4273]), .B(p_input[3273]), .Z(n6459) );
  AND U7269 ( .A(n6462), .B(n6463), .Z(n6457) );
  AND U7270 ( .A(n6464), .B(p_input[7273]), .Z(n6463) );
  AND U7271 ( .A(p_input[6273]), .B(p_input[5273]), .Z(n6464) );
  AND U7272 ( .A(p_input[9273]), .B(p_input[8273]), .Z(n6462) );
  AND U7273 ( .A(n6465), .B(n6466), .Z(o[272]) );
  AND U7274 ( .A(n6467), .B(n6468), .Z(n6466) );
  AND U7275 ( .A(n6469), .B(p_input[272]), .Z(n6468) );
  AND U7276 ( .A(p_input[2272]), .B(p_input[1272]), .Z(n6469) );
  AND U7277 ( .A(p_input[4272]), .B(p_input[3272]), .Z(n6467) );
  AND U7278 ( .A(n6470), .B(n6471), .Z(n6465) );
  AND U7279 ( .A(n6472), .B(p_input[7272]), .Z(n6471) );
  AND U7280 ( .A(p_input[6272]), .B(p_input[5272]), .Z(n6472) );
  AND U7281 ( .A(p_input[9272]), .B(p_input[8272]), .Z(n6470) );
  AND U7282 ( .A(n6473), .B(n6474), .Z(o[271]) );
  AND U7283 ( .A(n6475), .B(n6476), .Z(n6474) );
  AND U7284 ( .A(n6477), .B(p_input[271]), .Z(n6476) );
  AND U7285 ( .A(p_input[2271]), .B(p_input[1271]), .Z(n6477) );
  AND U7286 ( .A(p_input[4271]), .B(p_input[3271]), .Z(n6475) );
  AND U7287 ( .A(n6478), .B(n6479), .Z(n6473) );
  AND U7288 ( .A(n6480), .B(p_input[7271]), .Z(n6479) );
  AND U7289 ( .A(p_input[6271]), .B(p_input[5271]), .Z(n6480) );
  AND U7290 ( .A(p_input[9271]), .B(p_input[8271]), .Z(n6478) );
  AND U7291 ( .A(n6481), .B(n6482), .Z(o[270]) );
  AND U7292 ( .A(n6483), .B(n6484), .Z(n6482) );
  AND U7293 ( .A(n6485), .B(p_input[270]), .Z(n6484) );
  AND U7294 ( .A(p_input[2270]), .B(p_input[1270]), .Z(n6485) );
  AND U7295 ( .A(p_input[4270]), .B(p_input[3270]), .Z(n6483) );
  AND U7296 ( .A(n6486), .B(n6487), .Z(n6481) );
  AND U7297 ( .A(n6488), .B(p_input[7270]), .Z(n6487) );
  AND U7298 ( .A(p_input[6270]), .B(p_input[5270]), .Z(n6488) );
  AND U7299 ( .A(p_input[9270]), .B(p_input[8270]), .Z(n6486) );
  AND U7300 ( .A(n6489), .B(n6490), .Z(o[26]) );
  AND U7301 ( .A(n6491), .B(n6492), .Z(n6490) );
  AND U7302 ( .A(n6493), .B(p_input[26]), .Z(n6492) );
  AND U7303 ( .A(p_input[2026]), .B(p_input[1026]), .Z(n6493) );
  AND U7304 ( .A(p_input[4026]), .B(p_input[3026]), .Z(n6491) );
  AND U7305 ( .A(n6494), .B(n6495), .Z(n6489) );
  AND U7306 ( .A(n6496), .B(p_input[7026]), .Z(n6495) );
  AND U7307 ( .A(p_input[6026]), .B(p_input[5026]), .Z(n6496) );
  AND U7308 ( .A(p_input[9026]), .B(p_input[8026]), .Z(n6494) );
  AND U7309 ( .A(n6497), .B(n6498), .Z(o[269]) );
  AND U7310 ( .A(n6499), .B(n6500), .Z(n6498) );
  AND U7311 ( .A(n6501), .B(p_input[269]), .Z(n6500) );
  AND U7312 ( .A(p_input[2269]), .B(p_input[1269]), .Z(n6501) );
  AND U7313 ( .A(p_input[4269]), .B(p_input[3269]), .Z(n6499) );
  AND U7314 ( .A(n6502), .B(n6503), .Z(n6497) );
  AND U7315 ( .A(n6504), .B(p_input[7269]), .Z(n6503) );
  AND U7316 ( .A(p_input[6269]), .B(p_input[5269]), .Z(n6504) );
  AND U7317 ( .A(p_input[9269]), .B(p_input[8269]), .Z(n6502) );
  AND U7318 ( .A(n6505), .B(n6506), .Z(o[268]) );
  AND U7319 ( .A(n6507), .B(n6508), .Z(n6506) );
  AND U7320 ( .A(n6509), .B(p_input[268]), .Z(n6508) );
  AND U7321 ( .A(p_input[2268]), .B(p_input[1268]), .Z(n6509) );
  AND U7322 ( .A(p_input[4268]), .B(p_input[3268]), .Z(n6507) );
  AND U7323 ( .A(n6510), .B(n6511), .Z(n6505) );
  AND U7324 ( .A(n6512), .B(p_input[7268]), .Z(n6511) );
  AND U7325 ( .A(p_input[6268]), .B(p_input[5268]), .Z(n6512) );
  AND U7326 ( .A(p_input[9268]), .B(p_input[8268]), .Z(n6510) );
  AND U7327 ( .A(n6513), .B(n6514), .Z(o[267]) );
  AND U7328 ( .A(n6515), .B(n6516), .Z(n6514) );
  AND U7329 ( .A(n6517), .B(p_input[267]), .Z(n6516) );
  AND U7330 ( .A(p_input[2267]), .B(p_input[1267]), .Z(n6517) );
  AND U7331 ( .A(p_input[4267]), .B(p_input[3267]), .Z(n6515) );
  AND U7332 ( .A(n6518), .B(n6519), .Z(n6513) );
  AND U7333 ( .A(n6520), .B(p_input[7267]), .Z(n6519) );
  AND U7334 ( .A(p_input[6267]), .B(p_input[5267]), .Z(n6520) );
  AND U7335 ( .A(p_input[9267]), .B(p_input[8267]), .Z(n6518) );
  AND U7336 ( .A(n6521), .B(n6522), .Z(o[266]) );
  AND U7337 ( .A(n6523), .B(n6524), .Z(n6522) );
  AND U7338 ( .A(n6525), .B(p_input[266]), .Z(n6524) );
  AND U7339 ( .A(p_input[2266]), .B(p_input[1266]), .Z(n6525) );
  AND U7340 ( .A(p_input[4266]), .B(p_input[3266]), .Z(n6523) );
  AND U7341 ( .A(n6526), .B(n6527), .Z(n6521) );
  AND U7342 ( .A(n6528), .B(p_input[7266]), .Z(n6527) );
  AND U7343 ( .A(p_input[6266]), .B(p_input[5266]), .Z(n6528) );
  AND U7344 ( .A(p_input[9266]), .B(p_input[8266]), .Z(n6526) );
  AND U7345 ( .A(n6529), .B(n6530), .Z(o[265]) );
  AND U7346 ( .A(n6531), .B(n6532), .Z(n6530) );
  AND U7347 ( .A(n6533), .B(p_input[265]), .Z(n6532) );
  AND U7348 ( .A(p_input[2265]), .B(p_input[1265]), .Z(n6533) );
  AND U7349 ( .A(p_input[4265]), .B(p_input[3265]), .Z(n6531) );
  AND U7350 ( .A(n6534), .B(n6535), .Z(n6529) );
  AND U7351 ( .A(n6536), .B(p_input[7265]), .Z(n6535) );
  AND U7352 ( .A(p_input[6265]), .B(p_input[5265]), .Z(n6536) );
  AND U7353 ( .A(p_input[9265]), .B(p_input[8265]), .Z(n6534) );
  AND U7354 ( .A(n6537), .B(n6538), .Z(o[264]) );
  AND U7355 ( .A(n6539), .B(n6540), .Z(n6538) );
  AND U7356 ( .A(n6541), .B(p_input[264]), .Z(n6540) );
  AND U7357 ( .A(p_input[2264]), .B(p_input[1264]), .Z(n6541) );
  AND U7358 ( .A(p_input[4264]), .B(p_input[3264]), .Z(n6539) );
  AND U7359 ( .A(n6542), .B(n6543), .Z(n6537) );
  AND U7360 ( .A(n6544), .B(p_input[7264]), .Z(n6543) );
  AND U7361 ( .A(p_input[6264]), .B(p_input[5264]), .Z(n6544) );
  AND U7362 ( .A(p_input[9264]), .B(p_input[8264]), .Z(n6542) );
  AND U7363 ( .A(n6545), .B(n6546), .Z(o[263]) );
  AND U7364 ( .A(n6547), .B(n6548), .Z(n6546) );
  AND U7365 ( .A(n6549), .B(p_input[263]), .Z(n6548) );
  AND U7366 ( .A(p_input[2263]), .B(p_input[1263]), .Z(n6549) );
  AND U7367 ( .A(p_input[4263]), .B(p_input[3263]), .Z(n6547) );
  AND U7368 ( .A(n6550), .B(n6551), .Z(n6545) );
  AND U7369 ( .A(n6552), .B(p_input[7263]), .Z(n6551) );
  AND U7370 ( .A(p_input[6263]), .B(p_input[5263]), .Z(n6552) );
  AND U7371 ( .A(p_input[9263]), .B(p_input[8263]), .Z(n6550) );
  AND U7372 ( .A(n6553), .B(n6554), .Z(o[262]) );
  AND U7373 ( .A(n6555), .B(n6556), .Z(n6554) );
  AND U7374 ( .A(n6557), .B(p_input[262]), .Z(n6556) );
  AND U7375 ( .A(p_input[2262]), .B(p_input[1262]), .Z(n6557) );
  AND U7376 ( .A(p_input[4262]), .B(p_input[3262]), .Z(n6555) );
  AND U7377 ( .A(n6558), .B(n6559), .Z(n6553) );
  AND U7378 ( .A(n6560), .B(p_input[7262]), .Z(n6559) );
  AND U7379 ( .A(p_input[6262]), .B(p_input[5262]), .Z(n6560) );
  AND U7380 ( .A(p_input[9262]), .B(p_input[8262]), .Z(n6558) );
  AND U7381 ( .A(n6561), .B(n6562), .Z(o[261]) );
  AND U7382 ( .A(n6563), .B(n6564), .Z(n6562) );
  AND U7383 ( .A(n6565), .B(p_input[261]), .Z(n6564) );
  AND U7384 ( .A(p_input[2261]), .B(p_input[1261]), .Z(n6565) );
  AND U7385 ( .A(p_input[4261]), .B(p_input[3261]), .Z(n6563) );
  AND U7386 ( .A(n6566), .B(n6567), .Z(n6561) );
  AND U7387 ( .A(n6568), .B(p_input[7261]), .Z(n6567) );
  AND U7388 ( .A(p_input[6261]), .B(p_input[5261]), .Z(n6568) );
  AND U7389 ( .A(p_input[9261]), .B(p_input[8261]), .Z(n6566) );
  AND U7390 ( .A(n6569), .B(n6570), .Z(o[260]) );
  AND U7391 ( .A(n6571), .B(n6572), .Z(n6570) );
  AND U7392 ( .A(n6573), .B(p_input[260]), .Z(n6572) );
  AND U7393 ( .A(p_input[2260]), .B(p_input[1260]), .Z(n6573) );
  AND U7394 ( .A(p_input[4260]), .B(p_input[3260]), .Z(n6571) );
  AND U7395 ( .A(n6574), .B(n6575), .Z(n6569) );
  AND U7396 ( .A(n6576), .B(p_input[7260]), .Z(n6575) );
  AND U7397 ( .A(p_input[6260]), .B(p_input[5260]), .Z(n6576) );
  AND U7398 ( .A(p_input[9260]), .B(p_input[8260]), .Z(n6574) );
  AND U7399 ( .A(n6577), .B(n6578), .Z(o[25]) );
  AND U7400 ( .A(n6579), .B(n6580), .Z(n6578) );
  AND U7401 ( .A(n6581), .B(p_input[25]), .Z(n6580) );
  AND U7402 ( .A(p_input[2025]), .B(p_input[1025]), .Z(n6581) );
  AND U7403 ( .A(p_input[4025]), .B(p_input[3025]), .Z(n6579) );
  AND U7404 ( .A(n6582), .B(n6583), .Z(n6577) );
  AND U7405 ( .A(n6584), .B(p_input[7025]), .Z(n6583) );
  AND U7406 ( .A(p_input[6025]), .B(p_input[5025]), .Z(n6584) );
  AND U7407 ( .A(p_input[9025]), .B(p_input[8025]), .Z(n6582) );
  AND U7408 ( .A(n6585), .B(n6586), .Z(o[259]) );
  AND U7409 ( .A(n6587), .B(n6588), .Z(n6586) );
  AND U7410 ( .A(n6589), .B(p_input[259]), .Z(n6588) );
  AND U7411 ( .A(p_input[2259]), .B(p_input[1259]), .Z(n6589) );
  AND U7412 ( .A(p_input[4259]), .B(p_input[3259]), .Z(n6587) );
  AND U7413 ( .A(n6590), .B(n6591), .Z(n6585) );
  AND U7414 ( .A(n6592), .B(p_input[7259]), .Z(n6591) );
  AND U7415 ( .A(p_input[6259]), .B(p_input[5259]), .Z(n6592) );
  AND U7416 ( .A(p_input[9259]), .B(p_input[8259]), .Z(n6590) );
  AND U7417 ( .A(n6593), .B(n6594), .Z(o[258]) );
  AND U7418 ( .A(n6595), .B(n6596), .Z(n6594) );
  AND U7419 ( .A(n6597), .B(p_input[258]), .Z(n6596) );
  AND U7420 ( .A(p_input[2258]), .B(p_input[1258]), .Z(n6597) );
  AND U7421 ( .A(p_input[4258]), .B(p_input[3258]), .Z(n6595) );
  AND U7422 ( .A(n6598), .B(n6599), .Z(n6593) );
  AND U7423 ( .A(n6600), .B(p_input[7258]), .Z(n6599) );
  AND U7424 ( .A(p_input[6258]), .B(p_input[5258]), .Z(n6600) );
  AND U7425 ( .A(p_input[9258]), .B(p_input[8258]), .Z(n6598) );
  AND U7426 ( .A(n6601), .B(n6602), .Z(o[257]) );
  AND U7427 ( .A(n6603), .B(n6604), .Z(n6602) );
  AND U7428 ( .A(n6605), .B(p_input[257]), .Z(n6604) );
  AND U7429 ( .A(p_input[2257]), .B(p_input[1257]), .Z(n6605) );
  AND U7430 ( .A(p_input[4257]), .B(p_input[3257]), .Z(n6603) );
  AND U7431 ( .A(n6606), .B(n6607), .Z(n6601) );
  AND U7432 ( .A(n6608), .B(p_input[7257]), .Z(n6607) );
  AND U7433 ( .A(p_input[6257]), .B(p_input[5257]), .Z(n6608) );
  AND U7434 ( .A(p_input[9257]), .B(p_input[8257]), .Z(n6606) );
  AND U7435 ( .A(n6609), .B(n6610), .Z(o[256]) );
  AND U7436 ( .A(n6611), .B(n6612), .Z(n6610) );
  AND U7437 ( .A(n6613), .B(p_input[256]), .Z(n6612) );
  AND U7438 ( .A(p_input[2256]), .B(p_input[1256]), .Z(n6613) );
  AND U7439 ( .A(p_input[4256]), .B(p_input[3256]), .Z(n6611) );
  AND U7440 ( .A(n6614), .B(n6615), .Z(n6609) );
  AND U7441 ( .A(n6616), .B(p_input[7256]), .Z(n6615) );
  AND U7442 ( .A(p_input[6256]), .B(p_input[5256]), .Z(n6616) );
  AND U7443 ( .A(p_input[9256]), .B(p_input[8256]), .Z(n6614) );
  AND U7444 ( .A(n6617), .B(n6618), .Z(o[255]) );
  AND U7445 ( .A(n6619), .B(n6620), .Z(n6618) );
  AND U7446 ( .A(n6621), .B(p_input[255]), .Z(n6620) );
  AND U7447 ( .A(p_input[2255]), .B(p_input[1255]), .Z(n6621) );
  AND U7448 ( .A(p_input[4255]), .B(p_input[3255]), .Z(n6619) );
  AND U7449 ( .A(n6622), .B(n6623), .Z(n6617) );
  AND U7450 ( .A(n6624), .B(p_input[7255]), .Z(n6623) );
  AND U7451 ( .A(p_input[6255]), .B(p_input[5255]), .Z(n6624) );
  AND U7452 ( .A(p_input[9255]), .B(p_input[8255]), .Z(n6622) );
  AND U7453 ( .A(n6625), .B(n6626), .Z(o[254]) );
  AND U7454 ( .A(n6627), .B(n6628), .Z(n6626) );
  AND U7455 ( .A(n6629), .B(p_input[254]), .Z(n6628) );
  AND U7456 ( .A(p_input[2254]), .B(p_input[1254]), .Z(n6629) );
  AND U7457 ( .A(p_input[4254]), .B(p_input[3254]), .Z(n6627) );
  AND U7458 ( .A(n6630), .B(n6631), .Z(n6625) );
  AND U7459 ( .A(n6632), .B(p_input[7254]), .Z(n6631) );
  AND U7460 ( .A(p_input[6254]), .B(p_input[5254]), .Z(n6632) );
  AND U7461 ( .A(p_input[9254]), .B(p_input[8254]), .Z(n6630) );
  AND U7462 ( .A(n6633), .B(n6634), .Z(o[253]) );
  AND U7463 ( .A(n6635), .B(n6636), .Z(n6634) );
  AND U7464 ( .A(n6637), .B(p_input[253]), .Z(n6636) );
  AND U7465 ( .A(p_input[2253]), .B(p_input[1253]), .Z(n6637) );
  AND U7466 ( .A(p_input[4253]), .B(p_input[3253]), .Z(n6635) );
  AND U7467 ( .A(n6638), .B(n6639), .Z(n6633) );
  AND U7468 ( .A(n6640), .B(p_input[7253]), .Z(n6639) );
  AND U7469 ( .A(p_input[6253]), .B(p_input[5253]), .Z(n6640) );
  AND U7470 ( .A(p_input[9253]), .B(p_input[8253]), .Z(n6638) );
  AND U7471 ( .A(n6641), .B(n6642), .Z(o[252]) );
  AND U7472 ( .A(n6643), .B(n6644), .Z(n6642) );
  AND U7473 ( .A(n6645), .B(p_input[252]), .Z(n6644) );
  AND U7474 ( .A(p_input[2252]), .B(p_input[1252]), .Z(n6645) );
  AND U7475 ( .A(p_input[4252]), .B(p_input[3252]), .Z(n6643) );
  AND U7476 ( .A(n6646), .B(n6647), .Z(n6641) );
  AND U7477 ( .A(n6648), .B(p_input[7252]), .Z(n6647) );
  AND U7478 ( .A(p_input[6252]), .B(p_input[5252]), .Z(n6648) );
  AND U7479 ( .A(p_input[9252]), .B(p_input[8252]), .Z(n6646) );
  AND U7480 ( .A(n6649), .B(n6650), .Z(o[251]) );
  AND U7481 ( .A(n6651), .B(n6652), .Z(n6650) );
  AND U7482 ( .A(n6653), .B(p_input[251]), .Z(n6652) );
  AND U7483 ( .A(p_input[2251]), .B(p_input[1251]), .Z(n6653) );
  AND U7484 ( .A(p_input[4251]), .B(p_input[3251]), .Z(n6651) );
  AND U7485 ( .A(n6654), .B(n6655), .Z(n6649) );
  AND U7486 ( .A(n6656), .B(p_input[7251]), .Z(n6655) );
  AND U7487 ( .A(p_input[6251]), .B(p_input[5251]), .Z(n6656) );
  AND U7488 ( .A(p_input[9251]), .B(p_input[8251]), .Z(n6654) );
  AND U7489 ( .A(n6657), .B(n6658), .Z(o[250]) );
  AND U7490 ( .A(n6659), .B(n6660), .Z(n6658) );
  AND U7491 ( .A(n6661), .B(p_input[250]), .Z(n6660) );
  AND U7492 ( .A(p_input[2250]), .B(p_input[1250]), .Z(n6661) );
  AND U7493 ( .A(p_input[4250]), .B(p_input[3250]), .Z(n6659) );
  AND U7494 ( .A(n6662), .B(n6663), .Z(n6657) );
  AND U7495 ( .A(n6664), .B(p_input[7250]), .Z(n6663) );
  AND U7496 ( .A(p_input[6250]), .B(p_input[5250]), .Z(n6664) );
  AND U7497 ( .A(p_input[9250]), .B(p_input[8250]), .Z(n6662) );
  AND U7498 ( .A(n6665), .B(n6666), .Z(o[24]) );
  AND U7499 ( .A(n6667), .B(n6668), .Z(n6666) );
  AND U7500 ( .A(n6669), .B(p_input[24]), .Z(n6668) );
  AND U7501 ( .A(p_input[2024]), .B(p_input[1024]), .Z(n6669) );
  AND U7502 ( .A(p_input[4024]), .B(p_input[3024]), .Z(n6667) );
  AND U7503 ( .A(n6670), .B(n6671), .Z(n6665) );
  AND U7504 ( .A(n6672), .B(p_input[7024]), .Z(n6671) );
  AND U7505 ( .A(p_input[6024]), .B(p_input[5024]), .Z(n6672) );
  AND U7506 ( .A(p_input[9024]), .B(p_input[8024]), .Z(n6670) );
  AND U7507 ( .A(n6673), .B(n6674), .Z(o[249]) );
  AND U7508 ( .A(n6675), .B(n6676), .Z(n6674) );
  AND U7509 ( .A(n6677), .B(p_input[249]), .Z(n6676) );
  AND U7510 ( .A(p_input[2249]), .B(p_input[1249]), .Z(n6677) );
  AND U7511 ( .A(p_input[4249]), .B(p_input[3249]), .Z(n6675) );
  AND U7512 ( .A(n6678), .B(n6679), .Z(n6673) );
  AND U7513 ( .A(n6680), .B(p_input[7249]), .Z(n6679) );
  AND U7514 ( .A(p_input[6249]), .B(p_input[5249]), .Z(n6680) );
  AND U7515 ( .A(p_input[9249]), .B(p_input[8249]), .Z(n6678) );
  AND U7516 ( .A(n6681), .B(n6682), .Z(o[248]) );
  AND U7517 ( .A(n6683), .B(n6684), .Z(n6682) );
  AND U7518 ( .A(n6685), .B(p_input[248]), .Z(n6684) );
  AND U7519 ( .A(p_input[2248]), .B(p_input[1248]), .Z(n6685) );
  AND U7520 ( .A(p_input[4248]), .B(p_input[3248]), .Z(n6683) );
  AND U7521 ( .A(n6686), .B(n6687), .Z(n6681) );
  AND U7522 ( .A(n6688), .B(p_input[7248]), .Z(n6687) );
  AND U7523 ( .A(p_input[6248]), .B(p_input[5248]), .Z(n6688) );
  AND U7524 ( .A(p_input[9248]), .B(p_input[8248]), .Z(n6686) );
  AND U7525 ( .A(n6689), .B(n6690), .Z(o[247]) );
  AND U7526 ( .A(n6691), .B(n6692), .Z(n6690) );
  AND U7527 ( .A(n6693), .B(p_input[247]), .Z(n6692) );
  AND U7528 ( .A(p_input[2247]), .B(p_input[1247]), .Z(n6693) );
  AND U7529 ( .A(p_input[4247]), .B(p_input[3247]), .Z(n6691) );
  AND U7530 ( .A(n6694), .B(n6695), .Z(n6689) );
  AND U7531 ( .A(n6696), .B(p_input[7247]), .Z(n6695) );
  AND U7532 ( .A(p_input[6247]), .B(p_input[5247]), .Z(n6696) );
  AND U7533 ( .A(p_input[9247]), .B(p_input[8247]), .Z(n6694) );
  AND U7534 ( .A(n6697), .B(n6698), .Z(o[246]) );
  AND U7535 ( .A(n6699), .B(n6700), .Z(n6698) );
  AND U7536 ( .A(n6701), .B(p_input[246]), .Z(n6700) );
  AND U7537 ( .A(p_input[2246]), .B(p_input[1246]), .Z(n6701) );
  AND U7538 ( .A(p_input[4246]), .B(p_input[3246]), .Z(n6699) );
  AND U7539 ( .A(n6702), .B(n6703), .Z(n6697) );
  AND U7540 ( .A(n6704), .B(p_input[7246]), .Z(n6703) );
  AND U7541 ( .A(p_input[6246]), .B(p_input[5246]), .Z(n6704) );
  AND U7542 ( .A(p_input[9246]), .B(p_input[8246]), .Z(n6702) );
  AND U7543 ( .A(n6705), .B(n6706), .Z(o[245]) );
  AND U7544 ( .A(n6707), .B(n6708), .Z(n6706) );
  AND U7545 ( .A(n6709), .B(p_input[245]), .Z(n6708) );
  AND U7546 ( .A(p_input[2245]), .B(p_input[1245]), .Z(n6709) );
  AND U7547 ( .A(p_input[4245]), .B(p_input[3245]), .Z(n6707) );
  AND U7548 ( .A(n6710), .B(n6711), .Z(n6705) );
  AND U7549 ( .A(n6712), .B(p_input[7245]), .Z(n6711) );
  AND U7550 ( .A(p_input[6245]), .B(p_input[5245]), .Z(n6712) );
  AND U7551 ( .A(p_input[9245]), .B(p_input[8245]), .Z(n6710) );
  AND U7552 ( .A(n6713), .B(n6714), .Z(o[244]) );
  AND U7553 ( .A(n6715), .B(n6716), .Z(n6714) );
  AND U7554 ( .A(n6717), .B(p_input[244]), .Z(n6716) );
  AND U7555 ( .A(p_input[2244]), .B(p_input[1244]), .Z(n6717) );
  AND U7556 ( .A(p_input[4244]), .B(p_input[3244]), .Z(n6715) );
  AND U7557 ( .A(n6718), .B(n6719), .Z(n6713) );
  AND U7558 ( .A(n6720), .B(p_input[7244]), .Z(n6719) );
  AND U7559 ( .A(p_input[6244]), .B(p_input[5244]), .Z(n6720) );
  AND U7560 ( .A(p_input[9244]), .B(p_input[8244]), .Z(n6718) );
  AND U7561 ( .A(n6721), .B(n6722), .Z(o[243]) );
  AND U7562 ( .A(n6723), .B(n6724), .Z(n6722) );
  AND U7563 ( .A(n6725), .B(p_input[243]), .Z(n6724) );
  AND U7564 ( .A(p_input[2243]), .B(p_input[1243]), .Z(n6725) );
  AND U7565 ( .A(p_input[4243]), .B(p_input[3243]), .Z(n6723) );
  AND U7566 ( .A(n6726), .B(n6727), .Z(n6721) );
  AND U7567 ( .A(n6728), .B(p_input[7243]), .Z(n6727) );
  AND U7568 ( .A(p_input[6243]), .B(p_input[5243]), .Z(n6728) );
  AND U7569 ( .A(p_input[9243]), .B(p_input[8243]), .Z(n6726) );
  AND U7570 ( .A(n6729), .B(n6730), .Z(o[242]) );
  AND U7571 ( .A(n6731), .B(n6732), .Z(n6730) );
  AND U7572 ( .A(n6733), .B(p_input[242]), .Z(n6732) );
  AND U7573 ( .A(p_input[2242]), .B(p_input[1242]), .Z(n6733) );
  AND U7574 ( .A(p_input[4242]), .B(p_input[3242]), .Z(n6731) );
  AND U7575 ( .A(n6734), .B(n6735), .Z(n6729) );
  AND U7576 ( .A(n6736), .B(p_input[7242]), .Z(n6735) );
  AND U7577 ( .A(p_input[6242]), .B(p_input[5242]), .Z(n6736) );
  AND U7578 ( .A(p_input[9242]), .B(p_input[8242]), .Z(n6734) );
  AND U7579 ( .A(n6737), .B(n6738), .Z(o[241]) );
  AND U7580 ( .A(n6739), .B(n6740), .Z(n6738) );
  AND U7581 ( .A(n6741), .B(p_input[241]), .Z(n6740) );
  AND U7582 ( .A(p_input[2241]), .B(p_input[1241]), .Z(n6741) );
  AND U7583 ( .A(p_input[4241]), .B(p_input[3241]), .Z(n6739) );
  AND U7584 ( .A(n6742), .B(n6743), .Z(n6737) );
  AND U7585 ( .A(n6744), .B(p_input[7241]), .Z(n6743) );
  AND U7586 ( .A(p_input[6241]), .B(p_input[5241]), .Z(n6744) );
  AND U7587 ( .A(p_input[9241]), .B(p_input[8241]), .Z(n6742) );
  AND U7588 ( .A(n6745), .B(n6746), .Z(o[240]) );
  AND U7589 ( .A(n6747), .B(n6748), .Z(n6746) );
  AND U7590 ( .A(n6749), .B(p_input[240]), .Z(n6748) );
  AND U7591 ( .A(p_input[2240]), .B(p_input[1240]), .Z(n6749) );
  AND U7592 ( .A(p_input[4240]), .B(p_input[3240]), .Z(n6747) );
  AND U7593 ( .A(n6750), .B(n6751), .Z(n6745) );
  AND U7594 ( .A(n6752), .B(p_input[7240]), .Z(n6751) );
  AND U7595 ( .A(p_input[6240]), .B(p_input[5240]), .Z(n6752) );
  AND U7596 ( .A(p_input[9240]), .B(p_input[8240]), .Z(n6750) );
  AND U7597 ( .A(n6753), .B(n6754), .Z(o[23]) );
  AND U7598 ( .A(n6755), .B(n6756), .Z(n6754) );
  AND U7599 ( .A(n6757), .B(p_input[23]), .Z(n6756) );
  AND U7600 ( .A(p_input[2023]), .B(p_input[1023]), .Z(n6757) );
  AND U7601 ( .A(p_input[4023]), .B(p_input[3023]), .Z(n6755) );
  AND U7602 ( .A(n6758), .B(n6759), .Z(n6753) );
  AND U7603 ( .A(n6760), .B(p_input[7023]), .Z(n6759) );
  AND U7604 ( .A(p_input[6023]), .B(p_input[5023]), .Z(n6760) );
  AND U7605 ( .A(p_input[9023]), .B(p_input[8023]), .Z(n6758) );
  AND U7606 ( .A(n6761), .B(n6762), .Z(o[239]) );
  AND U7607 ( .A(n6763), .B(n6764), .Z(n6762) );
  AND U7608 ( .A(n6765), .B(p_input[239]), .Z(n6764) );
  AND U7609 ( .A(p_input[2239]), .B(p_input[1239]), .Z(n6765) );
  AND U7610 ( .A(p_input[4239]), .B(p_input[3239]), .Z(n6763) );
  AND U7611 ( .A(n6766), .B(n6767), .Z(n6761) );
  AND U7612 ( .A(n6768), .B(p_input[7239]), .Z(n6767) );
  AND U7613 ( .A(p_input[6239]), .B(p_input[5239]), .Z(n6768) );
  AND U7614 ( .A(p_input[9239]), .B(p_input[8239]), .Z(n6766) );
  AND U7615 ( .A(n6769), .B(n6770), .Z(o[238]) );
  AND U7616 ( .A(n6771), .B(n6772), .Z(n6770) );
  AND U7617 ( .A(n6773), .B(p_input[238]), .Z(n6772) );
  AND U7618 ( .A(p_input[2238]), .B(p_input[1238]), .Z(n6773) );
  AND U7619 ( .A(p_input[4238]), .B(p_input[3238]), .Z(n6771) );
  AND U7620 ( .A(n6774), .B(n6775), .Z(n6769) );
  AND U7621 ( .A(n6776), .B(p_input[7238]), .Z(n6775) );
  AND U7622 ( .A(p_input[6238]), .B(p_input[5238]), .Z(n6776) );
  AND U7623 ( .A(p_input[9238]), .B(p_input[8238]), .Z(n6774) );
  AND U7624 ( .A(n6777), .B(n6778), .Z(o[237]) );
  AND U7625 ( .A(n6779), .B(n6780), .Z(n6778) );
  AND U7626 ( .A(n6781), .B(p_input[237]), .Z(n6780) );
  AND U7627 ( .A(p_input[2237]), .B(p_input[1237]), .Z(n6781) );
  AND U7628 ( .A(p_input[4237]), .B(p_input[3237]), .Z(n6779) );
  AND U7629 ( .A(n6782), .B(n6783), .Z(n6777) );
  AND U7630 ( .A(n6784), .B(p_input[7237]), .Z(n6783) );
  AND U7631 ( .A(p_input[6237]), .B(p_input[5237]), .Z(n6784) );
  AND U7632 ( .A(p_input[9237]), .B(p_input[8237]), .Z(n6782) );
  AND U7633 ( .A(n6785), .B(n6786), .Z(o[236]) );
  AND U7634 ( .A(n6787), .B(n6788), .Z(n6786) );
  AND U7635 ( .A(n6789), .B(p_input[236]), .Z(n6788) );
  AND U7636 ( .A(p_input[2236]), .B(p_input[1236]), .Z(n6789) );
  AND U7637 ( .A(p_input[4236]), .B(p_input[3236]), .Z(n6787) );
  AND U7638 ( .A(n6790), .B(n6791), .Z(n6785) );
  AND U7639 ( .A(n6792), .B(p_input[7236]), .Z(n6791) );
  AND U7640 ( .A(p_input[6236]), .B(p_input[5236]), .Z(n6792) );
  AND U7641 ( .A(p_input[9236]), .B(p_input[8236]), .Z(n6790) );
  AND U7642 ( .A(n6793), .B(n6794), .Z(o[235]) );
  AND U7643 ( .A(n6795), .B(n6796), .Z(n6794) );
  AND U7644 ( .A(n6797), .B(p_input[235]), .Z(n6796) );
  AND U7645 ( .A(p_input[2235]), .B(p_input[1235]), .Z(n6797) );
  AND U7646 ( .A(p_input[4235]), .B(p_input[3235]), .Z(n6795) );
  AND U7647 ( .A(n6798), .B(n6799), .Z(n6793) );
  AND U7648 ( .A(n6800), .B(p_input[7235]), .Z(n6799) );
  AND U7649 ( .A(p_input[6235]), .B(p_input[5235]), .Z(n6800) );
  AND U7650 ( .A(p_input[9235]), .B(p_input[8235]), .Z(n6798) );
  AND U7651 ( .A(n6801), .B(n6802), .Z(o[234]) );
  AND U7652 ( .A(n6803), .B(n6804), .Z(n6802) );
  AND U7653 ( .A(n6805), .B(p_input[234]), .Z(n6804) );
  AND U7654 ( .A(p_input[2234]), .B(p_input[1234]), .Z(n6805) );
  AND U7655 ( .A(p_input[4234]), .B(p_input[3234]), .Z(n6803) );
  AND U7656 ( .A(n6806), .B(n6807), .Z(n6801) );
  AND U7657 ( .A(n6808), .B(p_input[7234]), .Z(n6807) );
  AND U7658 ( .A(p_input[6234]), .B(p_input[5234]), .Z(n6808) );
  AND U7659 ( .A(p_input[9234]), .B(p_input[8234]), .Z(n6806) );
  AND U7660 ( .A(n6809), .B(n6810), .Z(o[233]) );
  AND U7661 ( .A(n6811), .B(n6812), .Z(n6810) );
  AND U7662 ( .A(n6813), .B(p_input[233]), .Z(n6812) );
  AND U7663 ( .A(p_input[2233]), .B(p_input[1233]), .Z(n6813) );
  AND U7664 ( .A(p_input[4233]), .B(p_input[3233]), .Z(n6811) );
  AND U7665 ( .A(n6814), .B(n6815), .Z(n6809) );
  AND U7666 ( .A(n6816), .B(p_input[7233]), .Z(n6815) );
  AND U7667 ( .A(p_input[6233]), .B(p_input[5233]), .Z(n6816) );
  AND U7668 ( .A(p_input[9233]), .B(p_input[8233]), .Z(n6814) );
  AND U7669 ( .A(n6817), .B(n6818), .Z(o[232]) );
  AND U7670 ( .A(n6819), .B(n6820), .Z(n6818) );
  AND U7671 ( .A(n6821), .B(p_input[232]), .Z(n6820) );
  AND U7672 ( .A(p_input[2232]), .B(p_input[1232]), .Z(n6821) );
  AND U7673 ( .A(p_input[4232]), .B(p_input[3232]), .Z(n6819) );
  AND U7674 ( .A(n6822), .B(n6823), .Z(n6817) );
  AND U7675 ( .A(n6824), .B(p_input[7232]), .Z(n6823) );
  AND U7676 ( .A(p_input[6232]), .B(p_input[5232]), .Z(n6824) );
  AND U7677 ( .A(p_input[9232]), .B(p_input[8232]), .Z(n6822) );
  AND U7678 ( .A(n6825), .B(n6826), .Z(o[231]) );
  AND U7679 ( .A(n6827), .B(n6828), .Z(n6826) );
  AND U7680 ( .A(n6829), .B(p_input[231]), .Z(n6828) );
  AND U7681 ( .A(p_input[2231]), .B(p_input[1231]), .Z(n6829) );
  AND U7682 ( .A(p_input[4231]), .B(p_input[3231]), .Z(n6827) );
  AND U7683 ( .A(n6830), .B(n6831), .Z(n6825) );
  AND U7684 ( .A(n6832), .B(p_input[7231]), .Z(n6831) );
  AND U7685 ( .A(p_input[6231]), .B(p_input[5231]), .Z(n6832) );
  AND U7686 ( .A(p_input[9231]), .B(p_input[8231]), .Z(n6830) );
  AND U7687 ( .A(n6833), .B(n6834), .Z(o[230]) );
  AND U7688 ( .A(n6835), .B(n6836), .Z(n6834) );
  AND U7689 ( .A(n6837), .B(p_input[230]), .Z(n6836) );
  AND U7690 ( .A(p_input[2230]), .B(p_input[1230]), .Z(n6837) );
  AND U7691 ( .A(p_input[4230]), .B(p_input[3230]), .Z(n6835) );
  AND U7692 ( .A(n6838), .B(n6839), .Z(n6833) );
  AND U7693 ( .A(n6840), .B(p_input[7230]), .Z(n6839) );
  AND U7694 ( .A(p_input[6230]), .B(p_input[5230]), .Z(n6840) );
  AND U7695 ( .A(p_input[9230]), .B(p_input[8230]), .Z(n6838) );
  AND U7696 ( .A(n6841), .B(n6842), .Z(o[22]) );
  AND U7697 ( .A(n6843), .B(n6844), .Z(n6842) );
  AND U7698 ( .A(n6845), .B(p_input[22]), .Z(n6844) );
  AND U7699 ( .A(p_input[2022]), .B(p_input[1022]), .Z(n6845) );
  AND U7700 ( .A(p_input[4022]), .B(p_input[3022]), .Z(n6843) );
  AND U7701 ( .A(n6846), .B(n6847), .Z(n6841) );
  AND U7702 ( .A(n6848), .B(p_input[7022]), .Z(n6847) );
  AND U7703 ( .A(p_input[6022]), .B(p_input[5022]), .Z(n6848) );
  AND U7704 ( .A(p_input[9022]), .B(p_input[8022]), .Z(n6846) );
  AND U7705 ( .A(n6849), .B(n6850), .Z(o[229]) );
  AND U7706 ( .A(n6851), .B(n6852), .Z(n6850) );
  AND U7707 ( .A(n6853), .B(p_input[229]), .Z(n6852) );
  AND U7708 ( .A(p_input[2229]), .B(p_input[1229]), .Z(n6853) );
  AND U7709 ( .A(p_input[4229]), .B(p_input[3229]), .Z(n6851) );
  AND U7710 ( .A(n6854), .B(n6855), .Z(n6849) );
  AND U7711 ( .A(n6856), .B(p_input[7229]), .Z(n6855) );
  AND U7712 ( .A(p_input[6229]), .B(p_input[5229]), .Z(n6856) );
  AND U7713 ( .A(p_input[9229]), .B(p_input[8229]), .Z(n6854) );
  AND U7714 ( .A(n6857), .B(n6858), .Z(o[228]) );
  AND U7715 ( .A(n6859), .B(n6860), .Z(n6858) );
  AND U7716 ( .A(n6861), .B(p_input[228]), .Z(n6860) );
  AND U7717 ( .A(p_input[2228]), .B(p_input[1228]), .Z(n6861) );
  AND U7718 ( .A(p_input[4228]), .B(p_input[3228]), .Z(n6859) );
  AND U7719 ( .A(n6862), .B(n6863), .Z(n6857) );
  AND U7720 ( .A(n6864), .B(p_input[7228]), .Z(n6863) );
  AND U7721 ( .A(p_input[6228]), .B(p_input[5228]), .Z(n6864) );
  AND U7722 ( .A(p_input[9228]), .B(p_input[8228]), .Z(n6862) );
  AND U7723 ( .A(n6865), .B(n6866), .Z(o[227]) );
  AND U7724 ( .A(n6867), .B(n6868), .Z(n6866) );
  AND U7725 ( .A(n6869), .B(p_input[227]), .Z(n6868) );
  AND U7726 ( .A(p_input[2227]), .B(p_input[1227]), .Z(n6869) );
  AND U7727 ( .A(p_input[4227]), .B(p_input[3227]), .Z(n6867) );
  AND U7728 ( .A(n6870), .B(n6871), .Z(n6865) );
  AND U7729 ( .A(n6872), .B(p_input[7227]), .Z(n6871) );
  AND U7730 ( .A(p_input[6227]), .B(p_input[5227]), .Z(n6872) );
  AND U7731 ( .A(p_input[9227]), .B(p_input[8227]), .Z(n6870) );
  AND U7732 ( .A(n6873), .B(n6874), .Z(o[226]) );
  AND U7733 ( .A(n6875), .B(n6876), .Z(n6874) );
  AND U7734 ( .A(n6877), .B(p_input[226]), .Z(n6876) );
  AND U7735 ( .A(p_input[2226]), .B(p_input[1226]), .Z(n6877) );
  AND U7736 ( .A(p_input[4226]), .B(p_input[3226]), .Z(n6875) );
  AND U7737 ( .A(n6878), .B(n6879), .Z(n6873) );
  AND U7738 ( .A(n6880), .B(p_input[7226]), .Z(n6879) );
  AND U7739 ( .A(p_input[6226]), .B(p_input[5226]), .Z(n6880) );
  AND U7740 ( .A(p_input[9226]), .B(p_input[8226]), .Z(n6878) );
  AND U7741 ( .A(n6881), .B(n6882), .Z(o[225]) );
  AND U7742 ( .A(n6883), .B(n6884), .Z(n6882) );
  AND U7743 ( .A(n6885), .B(p_input[225]), .Z(n6884) );
  AND U7744 ( .A(p_input[2225]), .B(p_input[1225]), .Z(n6885) );
  AND U7745 ( .A(p_input[4225]), .B(p_input[3225]), .Z(n6883) );
  AND U7746 ( .A(n6886), .B(n6887), .Z(n6881) );
  AND U7747 ( .A(n6888), .B(p_input[7225]), .Z(n6887) );
  AND U7748 ( .A(p_input[6225]), .B(p_input[5225]), .Z(n6888) );
  AND U7749 ( .A(p_input[9225]), .B(p_input[8225]), .Z(n6886) );
  AND U7750 ( .A(n6889), .B(n6890), .Z(o[224]) );
  AND U7751 ( .A(n6891), .B(n6892), .Z(n6890) );
  AND U7752 ( .A(n6893), .B(p_input[224]), .Z(n6892) );
  AND U7753 ( .A(p_input[2224]), .B(p_input[1224]), .Z(n6893) );
  AND U7754 ( .A(p_input[4224]), .B(p_input[3224]), .Z(n6891) );
  AND U7755 ( .A(n6894), .B(n6895), .Z(n6889) );
  AND U7756 ( .A(n6896), .B(p_input[7224]), .Z(n6895) );
  AND U7757 ( .A(p_input[6224]), .B(p_input[5224]), .Z(n6896) );
  AND U7758 ( .A(p_input[9224]), .B(p_input[8224]), .Z(n6894) );
  AND U7759 ( .A(n6897), .B(n6898), .Z(o[223]) );
  AND U7760 ( .A(n6899), .B(n6900), .Z(n6898) );
  AND U7761 ( .A(n6901), .B(p_input[223]), .Z(n6900) );
  AND U7762 ( .A(p_input[2223]), .B(p_input[1223]), .Z(n6901) );
  AND U7763 ( .A(p_input[4223]), .B(p_input[3223]), .Z(n6899) );
  AND U7764 ( .A(n6902), .B(n6903), .Z(n6897) );
  AND U7765 ( .A(n6904), .B(p_input[7223]), .Z(n6903) );
  AND U7766 ( .A(p_input[6223]), .B(p_input[5223]), .Z(n6904) );
  AND U7767 ( .A(p_input[9223]), .B(p_input[8223]), .Z(n6902) );
  AND U7768 ( .A(n6905), .B(n6906), .Z(o[222]) );
  AND U7769 ( .A(n6907), .B(n6908), .Z(n6906) );
  AND U7770 ( .A(n6909), .B(p_input[222]), .Z(n6908) );
  AND U7771 ( .A(p_input[2222]), .B(p_input[1222]), .Z(n6909) );
  AND U7772 ( .A(p_input[4222]), .B(p_input[3222]), .Z(n6907) );
  AND U7773 ( .A(n6910), .B(n6911), .Z(n6905) );
  AND U7774 ( .A(n6912), .B(p_input[7222]), .Z(n6911) );
  AND U7775 ( .A(p_input[6222]), .B(p_input[5222]), .Z(n6912) );
  AND U7776 ( .A(p_input[9222]), .B(p_input[8222]), .Z(n6910) );
  AND U7777 ( .A(n6913), .B(n6914), .Z(o[221]) );
  AND U7778 ( .A(n6915), .B(n6916), .Z(n6914) );
  AND U7779 ( .A(n6917), .B(p_input[2221]), .Z(n6916) );
  AND U7780 ( .A(p_input[221]), .B(p_input[1221]), .Z(n6917) );
  AND U7781 ( .A(p_input[4221]), .B(p_input[3221]), .Z(n6915) );
  AND U7782 ( .A(n6918), .B(n6919), .Z(n6913) );
  AND U7783 ( .A(n6920), .B(p_input[7221]), .Z(n6919) );
  AND U7784 ( .A(p_input[6221]), .B(p_input[5221]), .Z(n6920) );
  AND U7785 ( .A(p_input[9221]), .B(p_input[8221]), .Z(n6918) );
  AND U7786 ( .A(n6921), .B(n6922), .Z(o[220]) );
  AND U7787 ( .A(n6923), .B(n6924), .Z(n6922) );
  AND U7788 ( .A(n6925), .B(p_input[2220]), .Z(n6924) );
  AND U7789 ( .A(p_input[220]), .B(p_input[1220]), .Z(n6925) );
  AND U7790 ( .A(p_input[4220]), .B(p_input[3220]), .Z(n6923) );
  AND U7791 ( .A(n6926), .B(n6927), .Z(n6921) );
  AND U7792 ( .A(n6928), .B(p_input[7220]), .Z(n6927) );
  AND U7793 ( .A(p_input[6220]), .B(p_input[5220]), .Z(n6928) );
  AND U7794 ( .A(p_input[9220]), .B(p_input[8220]), .Z(n6926) );
  AND U7795 ( .A(n6929), .B(n6930), .Z(o[21]) );
  AND U7796 ( .A(n6931), .B(n6932), .Z(n6930) );
  AND U7797 ( .A(n6933), .B(p_input[21]), .Z(n6932) );
  AND U7798 ( .A(p_input[2021]), .B(p_input[1021]), .Z(n6933) );
  AND U7799 ( .A(p_input[4021]), .B(p_input[3021]), .Z(n6931) );
  AND U7800 ( .A(n6934), .B(n6935), .Z(n6929) );
  AND U7801 ( .A(n6936), .B(p_input[7021]), .Z(n6935) );
  AND U7802 ( .A(p_input[6021]), .B(p_input[5021]), .Z(n6936) );
  AND U7803 ( .A(p_input[9021]), .B(p_input[8021]), .Z(n6934) );
  AND U7804 ( .A(n6937), .B(n6938), .Z(o[219]) );
  AND U7805 ( .A(n6939), .B(n6940), .Z(n6938) );
  AND U7806 ( .A(n6941), .B(p_input[2219]), .Z(n6940) );
  AND U7807 ( .A(p_input[219]), .B(p_input[1219]), .Z(n6941) );
  AND U7808 ( .A(p_input[4219]), .B(p_input[3219]), .Z(n6939) );
  AND U7809 ( .A(n6942), .B(n6943), .Z(n6937) );
  AND U7810 ( .A(n6944), .B(p_input[7219]), .Z(n6943) );
  AND U7811 ( .A(p_input[6219]), .B(p_input[5219]), .Z(n6944) );
  AND U7812 ( .A(p_input[9219]), .B(p_input[8219]), .Z(n6942) );
  AND U7813 ( .A(n6945), .B(n6946), .Z(o[218]) );
  AND U7814 ( .A(n6947), .B(n6948), .Z(n6946) );
  AND U7815 ( .A(n6949), .B(p_input[2218]), .Z(n6948) );
  AND U7816 ( .A(p_input[218]), .B(p_input[1218]), .Z(n6949) );
  AND U7817 ( .A(p_input[4218]), .B(p_input[3218]), .Z(n6947) );
  AND U7818 ( .A(n6950), .B(n6951), .Z(n6945) );
  AND U7819 ( .A(n6952), .B(p_input[7218]), .Z(n6951) );
  AND U7820 ( .A(p_input[6218]), .B(p_input[5218]), .Z(n6952) );
  AND U7821 ( .A(p_input[9218]), .B(p_input[8218]), .Z(n6950) );
  AND U7822 ( .A(n6953), .B(n6954), .Z(o[217]) );
  AND U7823 ( .A(n6955), .B(n6956), .Z(n6954) );
  AND U7824 ( .A(n6957), .B(p_input[2217]), .Z(n6956) );
  AND U7825 ( .A(p_input[217]), .B(p_input[1217]), .Z(n6957) );
  AND U7826 ( .A(p_input[4217]), .B(p_input[3217]), .Z(n6955) );
  AND U7827 ( .A(n6958), .B(n6959), .Z(n6953) );
  AND U7828 ( .A(n6960), .B(p_input[7217]), .Z(n6959) );
  AND U7829 ( .A(p_input[6217]), .B(p_input[5217]), .Z(n6960) );
  AND U7830 ( .A(p_input[9217]), .B(p_input[8217]), .Z(n6958) );
  AND U7831 ( .A(n6961), .B(n6962), .Z(o[216]) );
  AND U7832 ( .A(n6963), .B(n6964), .Z(n6962) );
  AND U7833 ( .A(n6965), .B(p_input[2216]), .Z(n6964) );
  AND U7834 ( .A(p_input[216]), .B(p_input[1216]), .Z(n6965) );
  AND U7835 ( .A(p_input[4216]), .B(p_input[3216]), .Z(n6963) );
  AND U7836 ( .A(n6966), .B(n6967), .Z(n6961) );
  AND U7837 ( .A(n6968), .B(p_input[7216]), .Z(n6967) );
  AND U7838 ( .A(p_input[6216]), .B(p_input[5216]), .Z(n6968) );
  AND U7839 ( .A(p_input[9216]), .B(p_input[8216]), .Z(n6966) );
  AND U7840 ( .A(n6969), .B(n6970), .Z(o[215]) );
  AND U7841 ( .A(n6971), .B(n6972), .Z(n6970) );
  AND U7842 ( .A(n6973), .B(p_input[2215]), .Z(n6972) );
  AND U7843 ( .A(p_input[215]), .B(p_input[1215]), .Z(n6973) );
  AND U7844 ( .A(p_input[4215]), .B(p_input[3215]), .Z(n6971) );
  AND U7845 ( .A(n6974), .B(n6975), .Z(n6969) );
  AND U7846 ( .A(n6976), .B(p_input[7215]), .Z(n6975) );
  AND U7847 ( .A(p_input[6215]), .B(p_input[5215]), .Z(n6976) );
  AND U7848 ( .A(p_input[9215]), .B(p_input[8215]), .Z(n6974) );
  AND U7849 ( .A(n6977), .B(n6978), .Z(o[214]) );
  AND U7850 ( .A(n6979), .B(n6980), .Z(n6978) );
  AND U7851 ( .A(n6981), .B(p_input[2214]), .Z(n6980) );
  AND U7852 ( .A(p_input[214]), .B(p_input[1214]), .Z(n6981) );
  AND U7853 ( .A(p_input[4214]), .B(p_input[3214]), .Z(n6979) );
  AND U7854 ( .A(n6982), .B(n6983), .Z(n6977) );
  AND U7855 ( .A(n6984), .B(p_input[7214]), .Z(n6983) );
  AND U7856 ( .A(p_input[6214]), .B(p_input[5214]), .Z(n6984) );
  AND U7857 ( .A(p_input[9214]), .B(p_input[8214]), .Z(n6982) );
  AND U7858 ( .A(n6985), .B(n6986), .Z(o[213]) );
  AND U7859 ( .A(n6987), .B(n6988), .Z(n6986) );
  AND U7860 ( .A(n6989), .B(p_input[2213]), .Z(n6988) );
  AND U7861 ( .A(p_input[213]), .B(p_input[1213]), .Z(n6989) );
  AND U7862 ( .A(p_input[4213]), .B(p_input[3213]), .Z(n6987) );
  AND U7863 ( .A(n6990), .B(n6991), .Z(n6985) );
  AND U7864 ( .A(n6992), .B(p_input[7213]), .Z(n6991) );
  AND U7865 ( .A(p_input[6213]), .B(p_input[5213]), .Z(n6992) );
  AND U7866 ( .A(p_input[9213]), .B(p_input[8213]), .Z(n6990) );
  AND U7867 ( .A(n6993), .B(n6994), .Z(o[212]) );
  AND U7868 ( .A(n6995), .B(n6996), .Z(n6994) );
  AND U7869 ( .A(n6997), .B(p_input[2212]), .Z(n6996) );
  AND U7870 ( .A(p_input[212]), .B(p_input[1212]), .Z(n6997) );
  AND U7871 ( .A(p_input[4212]), .B(p_input[3212]), .Z(n6995) );
  AND U7872 ( .A(n6998), .B(n6999), .Z(n6993) );
  AND U7873 ( .A(n7000), .B(p_input[7212]), .Z(n6999) );
  AND U7874 ( .A(p_input[6212]), .B(p_input[5212]), .Z(n7000) );
  AND U7875 ( .A(p_input[9212]), .B(p_input[8212]), .Z(n6998) );
  AND U7876 ( .A(n7001), .B(n7002), .Z(o[211]) );
  AND U7877 ( .A(n7003), .B(n7004), .Z(n7002) );
  AND U7878 ( .A(n7005), .B(p_input[2211]), .Z(n7004) );
  AND U7879 ( .A(p_input[211]), .B(p_input[1211]), .Z(n7005) );
  AND U7880 ( .A(p_input[4211]), .B(p_input[3211]), .Z(n7003) );
  AND U7881 ( .A(n7006), .B(n7007), .Z(n7001) );
  AND U7882 ( .A(n7008), .B(p_input[7211]), .Z(n7007) );
  AND U7883 ( .A(p_input[6211]), .B(p_input[5211]), .Z(n7008) );
  AND U7884 ( .A(p_input[9211]), .B(p_input[8211]), .Z(n7006) );
  AND U7885 ( .A(n7009), .B(n7010), .Z(o[210]) );
  AND U7886 ( .A(n7011), .B(n7012), .Z(n7010) );
  AND U7887 ( .A(n7013), .B(p_input[2210]), .Z(n7012) );
  AND U7888 ( .A(p_input[210]), .B(p_input[1210]), .Z(n7013) );
  AND U7889 ( .A(p_input[4210]), .B(p_input[3210]), .Z(n7011) );
  AND U7890 ( .A(n7014), .B(n7015), .Z(n7009) );
  AND U7891 ( .A(n7016), .B(p_input[7210]), .Z(n7015) );
  AND U7892 ( .A(p_input[6210]), .B(p_input[5210]), .Z(n7016) );
  AND U7893 ( .A(p_input[9210]), .B(p_input[8210]), .Z(n7014) );
  AND U7894 ( .A(n7017), .B(n7018), .Z(o[20]) );
  AND U7895 ( .A(n7019), .B(n7020), .Z(n7018) );
  AND U7896 ( .A(n7021), .B(p_input[20]), .Z(n7020) );
  AND U7897 ( .A(p_input[2020]), .B(p_input[1020]), .Z(n7021) );
  AND U7898 ( .A(p_input[4020]), .B(p_input[3020]), .Z(n7019) );
  AND U7899 ( .A(n7022), .B(n7023), .Z(n7017) );
  AND U7900 ( .A(n7024), .B(p_input[7020]), .Z(n7023) );
  AND U7901 ( .A(p_input[6020]), .B(p_input[5020]), .Z(n7024) );
  AND U7902 ( .A(p_input[9020]), .B(p_input[8020]), .Z(n7022) );
  AND U7903 ( .A(n7025), .B(n7026), .Z(o[209]) );
  AND U7904 ( .A(n7027), .B(n7028), .Z(n7026) );
  AND U7905 ( .A(n7029), .B(p_input[2209]), .Z(n7028) );
  AND U7906 ( .A(p_input[209]), .B(p_input[1209]), .Z(n7029) );
  AND U7907 ( .A(p_input[4209]), .B(p_input[3209]), .Z(n7027) );
  AND U7908 ( .A(n7030), .B(n7031), .Z(n7025) );
  AND U7909 ( .A(n7032), .B(p_input[7209]), .Z(n7031) );
  AND U7910 ( .A(p_input[6209]), .B(p_input[5209]), .Z(n7032) );
  AND U7911 ( .A(p_input[9209]), .B(p_input[8209]), .Z(n7030) );
  AND U7912 ( .A(n7033), .B(n7034), .Z(o[208]) );
  AND U7913 ( .A(n7035), .B(n7036), .Z(n7034) );
  AND U7914 ( .A(n7037), .B(p_input[2208]), .Z(n7036) );
  AND U7915 ( .A(p_input[208]), .B(p_input[1208]), .Z(n7037) );
  AND U7916 ( .A(p_input[4208]), .B(p_input[3208]), .Z(n7035) );
  AND U7917 ( .A(n7038), .B(n7039), .Z(n7033) );
  AND U7918 ( .A(n7040), .B(p_input[7208]), .Z(n7039) );
  AND U7919 ( .A(p_input[6208]), .B(p_input[5208]), .Z(n7040) );
  AND U7920 ( .A(p_input[9208]), .B(p_input[8208]), .Z(n7038) );
  AND U7921 ( .A(n7041), .B(n7042), .Z(o[207]) );
  AND U7922 ( .A(n7043), .B(n7044), .Z(n7042) );
  AND U7923 ( .A(n7045), .B(p_input[2207]), .Z(n7044) );
  AND U7924 ( .A(p_input[207]), .B(p_input[1207]), .Z(n7045) );
  AND U7925 ( .A(p_input[4207]), .B(p_input[3207]), .Z(n7043) );
  AND U7926 ( .A(n7046), .B(n7047), .Z(n7041) );
  AND U7927 ( .A(n7048), .B(p_input[7207]), .Z(n7047) );
  AND U7928 ( .A(p_input[6207]), .B(p_input[5207]), .Z(n7048) );
  AND U7929 ( .A(p_input[9207]), .B(p_input[8207]), .Z(n7046) );
  AND U7930 ( .A(n7049), .B(n7050), .Z(o[206]) );
  AND U7931 ( .A(n7051), .B(n7052), .Z(n7050) );
  AND U7932 ( .A(n7053), .B(p_input[2206]), .Z(n7052) );
  AND U7933 ( .A(p_input[206]), .B(p_input[1206]), .Z(n7053) );
  AND U7934 ( .A(p_input[4206]), .B(p_input[3206]), .Z(n7051) );
  AND U7935 ( .A(n7054), .B(n7055), .Z(n7049) );
  AND U7936 ( .A(n7056), .B(p_input[7206]), .Z(n7055) );
  AND U7937 ( .A(p_input[6206]), .B(p_input[5206]), .Z(n7056) );
  AND U7938 ( .A(p_input[9206]), .B(p_input[8206]), .Z(n7054) );
  AND U7939 ( .A(n7057), .B(n7058), .Z(o[205]) );
  AND U7940 ( .A(n7059), .B(n7060), .Z(n7058) );
  AND U7941 ( .A(n7061), .B(p_input[2205]), .Z(n7060) );
  AND U7942 ( .A(p_input[205]), .B(p_input[1205]), .Z(n7061) );
  AND U7943 ( .A(p_input[4205]), .B(p_input[3205]), .Z(n7059) );
  AND U7944 ( .A(n7062), .B(n7063), .Z(n7057) );
  AND U7945 ( .A(n7064), .B(p_input[7205]), .Z(n7063) );
  AND U7946 ( .A(p_input[6205]), .B(p_input[5205]), .Z(n7064) );
  AND U7947 ( .A(p_input[9205]), .B(p_input[8205]), .Z(n7062) );
  AND U7948 ( .A(n7065), .B(n7066), .Z(o[204]) );
  AND U7949 ( .A(n7067), .B(n7068), .Z(n7066) );
  AND U7950 ( .A(n7069), .B(p_input[2204]), .Z(n7068) );
  AND U7951 ( .A(p_input[204]), .B(p_input[1204]), .Z(n7069) );
  AND U7952 ( .A(p_input[4204]), .B(p_input[3204]), .Z(n7067) );
  AND U7953 ( .A(n7070), .B(n7071), .Z(n7065) );
  AND U7954 ( .A(n7072), .B(p_input[7204]), .Z(n7071) );
  AND U7955 ( .A(p_input[6204]), .B(p_input[5204]), .Z(n7072) );
  AND U7956 ( .A(p_input[9204]), .B(p_input[8204]), .Z(n7070) );
  AND U7957 ( .A(n7073), .B(n7074), .Z(o[203]) );
  AND U7958 ( .A(n7075), .B(n7076), .Z(n7074) );
  AND U7959 ( .A(n7077), .B(p_input[2203]), .Z(n7076) );
  AND U7960 ( .A(p_input[203]), .B(p_input[1203]), .Z(n7077) );
  AND U7961 ( .A(p_input[4203]), .B(p_input[3203]), .Z(n7075) );
  AND U7962 ( .A(n7078), .B(n7079), .Z(n7073) );
  AND U7963 ( .A(n7080), .B(p_input[7203]), .Z(n7079) );
  AND U7964 ( .A(p_input[6203]), .B(p_input[5203]), .Z(n7080) );
  AND U7965 ( .A(p_input[9203]), .B(p_input[8203]), .Z(n7078) );
  AND U7966 ( .A(n7081), .B(n7082), .Z(o[202]) );
  AND U7967 ( .A(n7083), .B(n7084), .Z(n7082) );
  AND U7968 ( .A(n7085), .B(p_input[2202]), .Z(n7084) );
  AND U7969 ( .A(p_input[202]), .B(p_input[1202]), .Z(n7085) );
  AND U7970 ( .A(p_input[4202]), .B(p_input[3202]), .Z(n7083) );
  AND U7971 ( .A(n7086), .B(n7087), .Z(n7081) );
  AND U7972 ( .A(n7088), .B(p_input[7202]), .Z(n7087) );
  AND U7973 ( .A(p_input[6202]), .B(p_input[5202]), .Z(n7088) );
  AND U7974 ( .A(p_input[9202]), .B(p_input[8202]), .Z(n7086) );
  AND U7975 ( .A(n7089), .B(n7090), .Z(o[201]) );
  AND U7976 ( .A(n7091), .B(n7092), .Z(n7090) );
  AND U7977 ( .A(n7093), .B(p_input[2201]), .Z(n7092) );
  AND U7978 ( .A(p_input[201]), .B(p_input[1201]), .Z(n7093) );
  AND U7979 ( .A(p_input[4201]), .B(p_input[3201]), .Z(n7091) );
  AND U7980 ( .A(n7094), .B(n7095), .Z(n7089) );
  AND U7981 ( .A(n7096), .B(p_input[7201]), .Z(n7095) );
  AND U7982 ( .A(p_input[6201]), .B(p_input[5201]), .Z(n7096) );
  AND U7983 ( .A(p_input[9201]), .B(p_input[8201]), .Z(n7094) );
  AND U7984 ( .A(n7097), .B(n7098), .Z(o[200]) );
  AND U7985 ( .A(n7099), .B(n7100), .Z(n7098) );
  AND U7986 ( .A(n7101), .B(p_input[2200]), .Z(n7100) );
  AND U7987 ( .A(p_input[200]), .B(p_input[1200]), .Z(n7101) );
  AND U7988 ( .A(p_input[4200]), .B(p_input[3200]), .Z(n7099) );
  AND U7989 ( .A(n7102), .B(n7103), .Z(n7097) );
  AND U7990 ( .A(n7104), .B(p_input[7200]), .Z(n7103) );
  AND U7991 ( .A(p_input[6200]), .B(p_input[5200]), .Z(n7104) );
  AND U7992 ( .A(p_input[9200]), .B(p_input[8200]), .Z(n7102) );
  AND U7993 ( .A(n7105), .B(n7106), .Z(o[1]) );
  AND U7994 ( .A(n7107), .B(n7108), .Z(n7106) );
  AND U7995 ( .A(n7109), .B(p_input[2001]), .Z(n7108) );
  AND U7996 ( .A(p_input[1]), .B(p_input[1001]), .Z(n7109) );
  AND U7997 ( .A(p_input[4001]), .B(p_input[3001]), .Z(n7107) );
  AND U7998 ( .A(n7110), .B(n7111), .Z(n7105) );
  AND U7999 ( .A(n7112), .B(p_input[7001]), .Z(n7111) );
  AND U8000 ( .A(p_input[6001]), .B(p_input[5001]), .Z(n7112) );
  AND U8001 ( .A(p_input[9001]), .B(p_input[8001]), .Z(n7110) );
  AND U8002 ( .A(n7113), .B(n7114), .Z(o[19]) );
  AND U8003 ( .A(n7115), .B(n7116), .Z(n7114) );
  AND U8004 ( .A(n7117), .B(p_input[2019]), .Z(n7116) );
  AND U8005 ( .A(p_input[19]), .B(p_input[1019]), .Z(n7117) );
  AND U8006 ( .A(p_input[4019]), .B(p_input[3019]), .Z(n7115) );
  AND U8007 ( .A(n7118), .B(n7119), .Z(n7113) );
  AND U8008 ( .A(n7120), .B(p_input[7019]), .Z(n7119) );
  AND U8009 ( .A(p_input[6019]), .B(p_input[5019]), .Z(n7120) );
  AND U8010 ( .A(p_input[9019]), .B(p_input[8019]), .Z(n7118) );
  AND U8011 ( .A(n7121), .B(n7122), .Z(o[199]) );
  AND U8012 ( .A(n7123), .B(n7124), .Z(n7122) );
  AND U8013 ( .A(n7125), .B(p_input[2199]), .Z(n7124) );
  AND U8014 ( .A(p_input[199]), .B(p_input[1199]), .Z(n7125) );
  AND U8015 ( .A(p_input[4199]), .B(p_input[3199]), .Z(n7123) );
  AND U8016 ( .A(n7126), .B(n7127), .Z(n7121) );
  AND U8017 ( .A(n7128), .B(p_input[7199]), .Z(n7127) );
  AND U8018 ( .A(p_input[6199]), .B(p_input[5199]), .Z(n7128) );
  AND U8019 ( .A(p_input[9199]), .B(p_input[8199]), .Z(n7126) );
  AND U8020 ( .A(n7129), .B(n7130), .Z(o[198]) );
  AND U8021 ( .A(n7131), .B(n7132), .Z(n7130) );
  AND U8022 ( .A(n7133), .B(p_input[2198]), .Z(n7132) );
  AND U8023 ( .A(p_input[198]), .B(p_input[1198]), .Z(n7133) );
  AND U8024 ( .A(p_input[4198]), .B(p_input[3198]), .Z(n7131) );
  AND U8025 ( .A(n7134), .B(n7135), .Z(n7129) );
  AND U8026 ( .A(n7136), .B(p_input[7198]), .Z(n7135) );
  AND U8027 ( .A(p_input[6198]), .B(p_input[5198]), .Z(n7136) );
  AND U8028 ( .A(p_input[9198]), .B(p_input[8198]), .Z(n7134) );
  AND U8029 ( .A(n7137), .B(n7138), .Z(o[197]) );
  AND U8030 ( .A(n7139), .B(n7140), .Z(n7138) );
  AND U8031 ( .A(n7141), .B(p_input[2197]), .Z(n7140) );
  AND U8032 ( .A(p_input[197]), .B(p_input[1197]), .Z(n7141) );
  AND U8033 ( .A(p_input[4197]), .B(p_input[3197]), .Z(n7139) );
  AND U8034 ( .A(n7142), .B(n7143), .Z(n7137) );
  AND U8035 ( .A(n7144), .B(p_input[7197]), .Z(n7143) );
  AND U8036 ( .A(p_input[6197]), .B(p_input[5197]), .Z(n7144) );
  AND U8037 ( .A(p_input[9197]), .B(p_input[8197]), .Z(n7142) );
  AND U8038 ( .A(n7145), .B(n7146), .Z(o[196]) );
  AND U8039 ( .A(n7147), .B(n7148), .Z(n7146) );
  AND U8040 ( .A(n7149), .B(p_input[2196]), .Z(n7148) );
  AND U8041 ( .A(p_input[196]), .B(p_input[1196]), .Z(n7149) );
  AND U8042 ( .A(p_input[4196]), .B(p_input[3196]), .Z(n7147) );
  AND U8043 ( .A(n7150), .B(n7151), .Z(n7145) );
  AND U8044 ( .A(n7152), .B(p_input[7196]), .Z(n7151) );
  AND U8045 ( .A(p_input[6196]), .B(p_input[5196]), .Z(n7152) );
  AND U8046 ( .A(p_input[9196]), .B(p_input[8196]), .Z(n7150) );
  AND U8047 ( .A(n7153), .B(n7154), .Z(o[195]) );
  AND U8048 ( .A(n7155), .B(n7156), .Z(n7154) );
  AND U8049 ( .A(n7157), .B(p_input[2195]), .Z(n7156) );
  AND U8050 ( .A(p_input[195]), .B(p_input[1195]), .Z(n7157) );
  AND U8051 ( .A(p_input[4195]), .B(p_input[3195]), .Z(n7155) );
  AND U8052 ( .A(n7158), .B(n7159), .Z(n7153) );
  AND U8053 ( .A(n7160), .B(p_input[7195]), .Z(n7159) );
  AND U8054 ( .A(p_input[6195]), .B(p_input[5195]), .Z(n7160) );
  AND U8055 ( .A(p_input[9195]), .B(p_input[8195]), .Z(n7158) );
  AND U8056 ( .A(n7161), .B(n7162), .Z(o[194]) );
  AND U8057 ( .A(n7163), .B(n7164), .Z(n7162) );
  AND U8058 ( .A(n7165), .B(p_input[2194]), .Z(n7164) );
  AND U8059 ( .A(p_input[194]), .B(p_input[1194]), .Z(n7165) );
  AND U8060 ( .A(p_input[4194]), .B(p_input[3194]), .Z(n7163) );
  AND U8061 ( .A(n7166), .B(n7167), .Z(n7161) );
  AND U8062 ( .A(n7168), .B(p_input[7194]), .Z(n7167) );
  AND U8063 ( .A(p_input[6194]), .B(p_input[5194]), .Z(n7168) );
  AND U8064 ( .A(p_input[9194]), .B(p_input[8194]), .Z(n7166) );
  AND U8065 ( .A(n7169), .B(n7170), .Z(o[193]) );
  AND U8066 ( .A(n7171), .B(n7172), .Z(n7170) );
  AND U8067 ( .A(n7173), .B(p_input[2193]), .Z(n7172) );
  AND U8068 ( .A(p_input[193]), .B(p_input[1193]), .Z(n7173) );
  AND U8069 ( .A(p_input[4193]), .B(p_input[3193]), .Z(n7171) );
  AND U8070 ( .A(n7174), .B(n7175), .Z(n7169) );
  AND U8071 ( .A(n7176), .B(p_input[7193]), .Z(n7175) );
  AND U8072 ( .A(p_input[6193]), .B(p_input[5193]), .Z(n7176) );
  AND U8073 ( .A(p_input[9193]), .B(p_input[8193]), .Z(n7174) );
  AND U8074 ( .A(n7177), .B(n7178), .Z(o[192]) );
  AND U8075 ( .A(n7179), .B(n7180), .Z(n7178) );
  AND U8076 ( .A(n7181), .B(p_input[2192]), .Z(n7180) );
  AND U8077 ( .A(p_input[192]), .B(p_input[1192]), .Z(n7181) );
  AND U8078 ( .A(p_input[4192]), .B(p_input[3192]), .Z(n7179) );
  AND U8079 ( .A(n7182), .B(n7183), .Z(n7177) );
  AND U8080 ( .A(n7184), .B(p_input[7192]), .Z(n7183) );
  AND U8081 ( .A(p_input[6192]), .B(p_input[5192]), .Z(n7184) );
  AND U8082 ( .A(p_input[9192]), .B(p_input[8192]), .Z(n7182) );
  AND U8083 ( .A(n7185), .B(n7186), .Z(o[191]) );
  AND U8084 ( .A(n7187), .B(n7188), .Z(n7186) );
  AND U8085 ( .A(n7189), .B(p_input[2191]), .Z(n7188) );
  AND U8086 ( .A(p_input[191]), .B(p_input[1191]), .Z(n7189) );
  AND U8087 ( .A(p_input[4191]), .B(p_input[3191]), .Z(n7187) );
  AND U8088 ( .A(n7190), .B(n7191), .Z(n7185) );
  AND U8089 ( .A(n7192), .B(p_input[7191]), .Z(n7191) );
  AND U8090 ( .A(p_input[6191]), .B(p_input[5191]), .Z(n7192) );
  AND U8091 ( .A(p_input[9191]), .B(p_input[8191]), .Z(n7190) );
  AND U8092 ( .A(n7193), .B(n7194), .Z(o[190]) );
  AND U8093 ( .A(n7195), .B(n7196), .Z(n7194) );
  AND U8094 ( .A(n7197), .B(p_input[2190]), .Z(n7196) );
  AND U8095 ( .A(p_input[190]), .B(p_input[1190]), .Z(n7197) );
  AND U8096 ( .A(p_input[4190]), .B(p_input[3190]), .Z(n7195) );
  AND U8097 ( .A(n7198), .B(n7199), .Z(n7193) );
  AND U8098 ( .A(n7200), .B(p_input[7190]), .Z(n7199) );
  AND U8099 ( .A(p_input[6190]), .B(p_input[5190]), .Z(n7200) );
  AND U8100 ( .A(p_input[9190]), .B(p_input[8190]), .Z(n7198) );
  AND U8101 ( .A(n7201), .B(n7202), .Z(o[18]) );
  AND U8102 ( .A(n7203), .B(n7204), .Z(n7202) );
  AND U8103 ( .A(n7205), .B(p_input[2018]), .Z(n7204) );
  AND U8104 ( .A(p_input[18]), .B(p_input[1018]), .Z(n7205) );
  AND U8105 ( .A(p_input[4018]), .B(p_input[3018]), .Z(n7203) );
  AND U8106 ( .A(n7206), .B(n7207), .Z(n7201) );
  AND U8107 ( .A(n7208), .B(p_input[7018]), .Z(n7207) );
  AND U8108 ( .A(p_input[6018]), .B(p_input[5018]), .Z(n7208) );
  AND U8109 ( .A(p_input[9018]), .B(p_input[8018]), .Z(n7206) );
  AND U8110 ( .A(n7209), .B(n7210), .Z(o[189]) );
  AND U8111 ( .A(n7211), .B(n7212), .Z(n7210) );
  AND U8112 ( .A(n7213), .B(p_input[2189]), .Z(n7212) );
  AND U8113 ( .A(p_input[189]), .B(p_input[1189]), .Z(n7213) );
  AND U8114 ( .A(p_input[4189]), .B(p_input[3189]), .Z(n7211) );
  AND U8115 ( .A(n7214), .B(n7215), .Z(n7209) );
  AND U8116 ( .A(n7216), .B(p_input[7189]), .Z(n7215) );
  AND U8117 ( .A(p_input[6189]), .B(p_input[5189]), .Z(n7216) );
  AND U8118 ( .A(p_input[9189]), .B(p_input[8189]), .Z(n7214) );
  AND U8119 ( .A(n7217), .B(n7218), .Z(o[188]) );
  AND U8120 ( .A(n7219), .B(n7220), .Z(n7218) );
  AND U8121 ( .A(n7221), .B(p_input[2188]), .Z(n7220) );
  AND U8122 ( .A(p_input[188]), .B(p_input[1188]), .Z(n7221) );
  AND U8123 ( .A(p_input[4188]), .B(p_input[3188]), .Z(n7219) );
  AND U8124 ( .A(n7222), .B(n7223), .Z(n7217) );
  AND U8125 ( .A(n7224), .B(p_input[7188]), .Z(n7223) );
  AND U8126 ( .A(p_input[6188]), .B(p_input[5188]), .Z(n7224) );
  AND U8127 ( .A(p_input[9188]), .B(p_input[8188]), .Z(n7222) );
  AND U8128 ( .A(n7225), .B(n7226), .Z(o[187]) );
  AND U8129 ( .A(n7227), .B(n7228), .Z(n7226) );
  AND U8130 ( .A(n7229), .B(p_input[2187]), .Z(n7228) );
  AND U8131 ( .A(p_input[187]), .B(p_input[1187]), .Z(n7229) );
  AND U8132 ( .A(p_input[4187]), .B(p_input[3187]), .Z(n7227) );
  AND U8133 ( .A(n7230), .B(n7231), .Z(n7225) );
  AND U8134 ( .A(n7232), .B(p_input[7187]), .Z(n7231) );
  AND U8135 ( .A(p_input[6187]), .B(p_input[5187]), .Z(n7232) );
  AND U8136 ( .A(p_input[9187]), .B(p_input[8187]), .Z(n7230) );
  AND U8137 ( .A(n7233), .B(n7234), .Z(o[186]) );
  AND U8138 ( .A(n7235), .B(n7236), .Z(n7234) );
  AND U8139 ( .A(n7237), .B(p_input[2186]), .Z(n7236) );
  AND U8140 ( .A(p_input[186]), .B(p_input[1186]), .Z(n7237) );
  AND U8141 ( .A(p_input[4186]), .B(p_input[3186]), .Z(n7235) );
  AND U8142 ( .A(n7238), .B(n7239), .Z(n7233) );
  AND U8143 ( .A(n7240), .B(p_input[7186]), .Z(n7239) );
  AND U8144 ( .A(p_input[6186]), .B(p_input[5186]), .Z(n7240) );
  AND U8145 ( .A(p_input[9186]), .B(p_input[8186]), .Z(n7238) );
  AND U8146 ( .A(n7241), .B(n7242), .Z(o[185]) );
  AND U8147 ( .A(n7243), .B(n7244), .Z(n7242) );
  AND U8148 ( .A(n7245), .B(p_input[2185]), .Z(n7244) );
  AND U8149 ( .A(p_input[185]), .B(p_input[1185]), .Z(n7245) );
  AND U8150 ( .A(p_input[4185]), .B(p_input[3185]), .Z(n7243) );
  AND U8151 ( .A(n7246), .B(n7247), .Z(n7241) );
  AND U8152 ( .A(n7248), .B(p_input[7185]), .Z(n7247) );
  AND U8153 ( .A(p_input[6185]), .B(p_input[5185]), .Z(n7248) );
  AND U8154 ( .A(p_input[9185]), .B(p_input[8185]), .Z(n7246) );
  AND U8155 ( .A(n7249), .B(n7250), .Z(o[184]) );
  AND U8156 ( .A(n7251), .B(n7252), .Z(n7250) );
  AND U8157 ( .A(n7253), .B(p_input[2184]), .Z(n7252) );
  AND U8158 ( .A(p_input[184]), .B(p_input[1184]), .Z(n7253) );
  AND U8159 ( .A(p_input[4184]), .B(p_input[3184]), .Z(n7251) );
  AND U8160 ( .A(n7254), .B(n7255), .Z(n7249) );
  AND U8161 ( .A(n7256), .B(p_input[7184]), .Z(n7255) );
  AND U8162 ( .A(p_input[6184]), .B(p_input[5184]), .Z(n7256) );
  AND U8163 ( .A(p_input[9184]), .B(p_input[8184]), .Z(n7254) );
  AND U8164 ( .A(n7257), .B(n7258), .Z(o[183]) );
  AND U8165 ( .A(n7259), .B(n7260), .Z(n7258) );
  AND U8166 ( .A(n7261), .B(p_input[2183]), .Z(n7260) );
  AND U8167 ( .A(p_input[183]), .B(p_input[1183]), .Z(n7261) );
  AND U8168 ( .A(p_input[4183]), .B(p_input[3183]), .Z(n7259) );
  AND U8169 ( .A(n7262), .B(n7263), .Z(n7257) );
  AND U8170 ( .A(n7264), .B(p_input[7183]), .Z(n7263) );
  AND U8171 ( .A(p_input[6183]), .B(p_input[5183]), .Z(n7264) );
  AND U8172 ( .A(p_input[9183]), .B(p_input[8183]), .Z(n7262) );
  AND U8173 ( .A(n7265), .B(n7266), .Z(o[182]) );
  AND U8174 ( .A(n7267), .B(n7268), .Z(n7266) );
  AND U8175 ( .A(n7269), .B(p_input[2182]), .Z(n7268) );
  AND U8176 ( .A(p_input[182]), .B(p_input[1182]), .Z(n7269) );
  AND U8177 ( .A(p_input[4182]), .B(p_input[3182]), .Z(n7267) );
  AND U8178 ( .A(n7270), .B(n7271), .Z(n7265) );
  AND U8179 ( .A(n7272), .B(p_input[7182]), .Z(n7271) );
  AND U8180 ( .A(p_input[6182]), .B(p_input[5182]), .Z(n7272) );
  AND U8181 ( .A(p_input[9182]), .B(p_input[8182]), .Z(n7270) );
  AND U8182 ( .A(n7273), .B(n7274), .Z(o[181]) );
  AND U8183 ( .A(n7275), .B(n7276), .Z(n7274) );
  AND U8184 ( .A(n7277), .B(p_input[2181]), .Z(n7276) );
  AND U8185 ( .A(p_input[181]), .B(p_input[1181]), .Z(n7277) );
  AND U8186 ( .A(p_input[4181]), .B(p_input[3181]), .Z(n7275) );
  AND U8187 ( .A(n7278), .B(n7279), .Z(n7273) );
  AND U8188 ( .A(n7280), .B(p_input[7181]), .Z(n7279) );
  AND U8189 ( .A(p_input[6181]), .B(p_input[5181]), .Z(n7280) );
  AND U8190 ( .A(p_input[9181]), .B(p_input[8181]), .Z(n7278) );
  AND U8191 ( .A(n7281), .B(n7282), .Z(o[180]) );
  AND U8192 ( .A(n7283), .B(n7284), .Z(n7282) );
  AND U8193 ( .A(n7285), .B(p_input[2180]), .Z(n7284) );
  AND U8194 ( .A(p_input[180]), .B(p_input[1180]), .Z(n7285) );
  AND U8195 ( .A(p_input[4180]), .B(p_input[3180]), .Z(n7283) );
  AND U8196 ( .A(n7286), .B(n7287), .Z(n7281) );
  AND U8197 ( .A(n7288), .B(p_input[7180]), .Z(n7287) );
  AND U8198 ( .A(p_input[6180]), .B(p_input[5180]), .Z(n7288) );
  AND U8199 ( .A(p_input[9180]), .B(p_input[8180]), .Z(n7286) );
  AND U8200 ( .A(n7289), .B(n7290), .Z(o[17]) );
  AND U8201 ( .A(n7291), .B(n7292), .Z(n7290) );
  AND U8202 ( .A(n7293), .B(p_input[2017]), .Z(n7292) );
  AND U8203 ( .A(p_input[17]), .B(p_input[1017]), .Z(n7293) );
  AND U8204 ( .A(p_input[4017]), .B(p_input[3017]), .Z(n7291) );
  AND U8205 ( .A(n7294), .B(n7295), .Z(n7289) );
  AND U8206 ( .A(n7296), .B(p_input[7017]), .Z(n7295) );
  AND U8207 ( .A(p_input[6017]), .B(p_input[5017]), .Z(n7296) );
  AND U8208 ( .A(p_input[9017]), .B(p_input[8017]), .Z(n7294) );
  AND U8209 ( .A(n7297), .B(n7298), .Z(o[179]) );
  AND U8210 ( .A(n7299), .B(n7300), .Z(n7298) );
  AND U8211 ( .A(n7301), .B(p_input[2179]), .Z(n7300) );
  AND U8212 ( .A(p_input[179]), .B(p_input[1179]), .Z(n7301) );
  AND U8213 ( .A(p_input[4179]), .B(p_input[3179]), .Z(n7299) );
  AND U8214 ( .A(n7302), .B(n7303), .Z(n7297) );
  AND U8215 ( .A(n7304), .B(p_input[7179]), .Z(n7303) );
  AND U8216 ( .A(p_input[6179]), .B(p_input[5179]), .Z(n7304) );
  AND U8217 ( .A(p_input[9179]), .B(p_input[8179]), .Z(n7302) );
  AND U8218 ( .A(n7305), .B(n7306), .Z(o[178]) );
  AND U8219 ( .A(n7307), .B(n7308), .Z(n7306) );
  AND U8220 ( .A(n7309), .B(p_input[2178]), .Z(n7308) );
  AND U8221 ( .A(p_input[178]), .B(p_input[1178]), .Z(n7309) );
  AND U8222 ( .A(p_input[4178]), .B(p_input[3178]), .Z(n7307) );
  AND U8223 ( .A(n7310), .B(n7311), .Z(n7305) );
  AND U8224 ( .A(n7312), .B(p_input[7178]), .Z(n7311) );
  AND U8225 ( .A(p_input[6178]), .B(p_input[5178]), .Z(n7312) );
  AND U8226 ( .A(p_input[9178]), .B(p_input[8178]), .Z(n7310) );
  AND U8227 ( .A(n7313), .B(n7314), .Z(o[177]) );
  AND U8228 ( .A(n7315), .B(n7316), .Z(n7314) );
  AND U8229 ( .A(n7317), .B(p_input[2177]), .Z(n7316) );
  AND U8230 ( .A(p_input[177]), .B(p_input[1177]), .Z(n7317) );
  AND U8231 ( .A(p_input[4177]), .B(p_input[3177]), .Z(n7315) );
  AND U8232 ( .A(n7318), .B(n7319), .Z(n7313) );
  AND U8233 ( .A(n7320), .B(p_input[7177]), .Z(n7319) );
  AND U8234 ( .A(p_input[6177]), .B(p_input[5177]), .Z(n7320) );
  AND U8235 ( .A(p_input[9177]), .B(p_input[8177]), .Z(n7318) );
  AND U8236 ( .A(n7321), .B(n7322), .Z(o[176]) );
  AND U8237 ( .A(n7323), .B(n7324), .Z(n7322) );
  AND U8238 ( .A(n7325), .B(p_input[2176]), .Z(n7324) );
  AND U8239 ( .A(p_input[176]), .B(p_input[1176]), .Z(n7325) );
  AND U8240 ( .A(p_input[4176]), .B(p_input[3176]), .Z(n7323) );
  AND U8241 ( .A(n7326), .B(n7327), .Z(n7321) );
  AND U8242 ( .A(n7328), .B(p_input[7176]), .Z(n7327) );
  AND U8243 ( .A(p_input[6176]), .B(p_input[5176]), .Z(n7328) );
  AND U8244 ( .A(p_input[9176]), .B(p_input[8176]), .Z(n7326) );
  AND U8245 ( .A(n7329), .B(n7330), .Z(o[175]) );
  AND U8246 ( .A(n7331), .B(n7332), .Z(n7330) );
  AND U8247 ( .A(n7333), .B(p_input[2175]), .Z(n7332) );
  AND U8248 ( .A(p_input[175]), .B(p_input[1175]), .Z(n7333) );
  AND U8249 ( .A(p_input[4175]), .B(p_input[3175]), .Z(n7331) );
  AND U8250 ( .A(n7334), .B(n7335), .Z(n7329) );
  AND U8251 ( .A(n7336), .B(p_input[7175]), .Z(n7335) );
  AND U8252 ( .A(p_input[6175]), .B(p_input[5175]), .Z(n7336) );
  AND U8253 ( .A(p_input[9175]), .B(p_input[8175]), .Z(n7334) );
  AND U8254 ( .A(n7337), .B(n7338), .Z(o[174]) );
  AND U8255 ( .A(n7339), .B(n7340), .Z(n7338) );
  AND U8256 ( .A(n7341), .B(p_input[2174]), .Z(n7340) );
  AND U8257 ( .A(p_input[174]), .B(p_input[1174]), .Z(n7341) );
  AND U8258 ( .A(p_input[4174]), .B(p_input[3174]), .Z(n7339) );
  AND U8259 ( .A(n7342), .B(n7343), .Z(n7337) );
  AND U8260 ( .A(n7344), .B(p_input[7174]), .Z(n7343) );
  AND U8261 ( .A(p_input[6174]), .B(p_input[5174]), .Z(n7344) );
  AND U8262 ( .A(p_input[9174]), .B(p_input[8174]), .Z(n7342) );
  AND U8263 ( .A(n7345), .B(n7346), .Z(o[173]) );
  AND U8264 ( .A(n7347), .B(n7348), .Z(n7346) );
  AND U8265 ( .A(n7349), .B(p_input[2173]), .Z(n7348) );
  AND U8266 ( .A(p_input[173]), .B(p_input[1173]), .Z(n7349) );
  AND U8267 ( .A(p_input[4173]), .B(p_input[3173]), .Z(n7347) );
  AND U8268 ( .A(n7350), .B(n7351), .Z(n7345) );
  AND U8269 ( .A(n7352), .B(p_input[7173]), .Z(n7351) );
  AND U8270 ( .A(p_input[6173]), .B(p_input[5173]), .Z(n7352) );
  AND U8271 ( .A(p_input[9173]), .B(p_input[8173]), .Z(n7350) );
  AND U8272 ( .A(n7353), .B(n7354), .Z(o[172]) );
  AND U8273 ( .A(n7355), .B(n7356), .Z(n7354) );
  AND U8274 ( .A(n7357), .B(p_input[2172]), .Z(n7356) );
  AND U8275 ( .A(p_input[172]), .B(p_input[1172]), .Z(n7357) );
  AND U8276 ( .A(p_input[4172]), .B(p_input[3172]), .Z(n7355) );
  AND U8277 ( .A(n7358), .B(n7359), .Z(n7353) );
  AND U8278 ( .A(n7360), .B(p_input[7172]), .Z(n7359) );
  AND U8279 ( .A(p_input[6172]), .B(p_input[5172]), .Z(n7360) );
  AND U8280 ( .A(p_input[9172]), .B(p_input[8172]), .Z(n7358) );
  AND U8281 ( .A(n7361), .B(n7362), .Z(o[171]) );
  AND U8282 ( .A(n7363), .B(n7364), .Z(n7362) );
  AND U8283 ( .A(n7365), .B(p_input[2171]), .Z(n7364) );
  AND U8284 ( .A(p_input[171]), .B(p_input[1171]), .Z(n7365) );
  AND U8285 ( .A(p_input[4171]), .B(p_input[3171]), .Z(n7363) );
  AND U8286 ( .A(n7366), .B(n7367), .Z(n7361) );
  AND U8287 ( .A(n7368), .B(p_input[7171]), .Z(n7367) );
  AND U8288 ( .A(p_input[6171]), .B(p_input[5171]), .Z(n7368) );
  AND U8289 ( .A(p_input[9171]), .B(p_input[8171]), .Z(n7366) );
  AND U8290 ( .A(n7369), .B(n7370), .Z(o[170]) );
  AND U8291 ( .A(n7371), .B(n7372), .Z(n7370) );
  AND U8292 ( .A(n7373), .B(p_input[2170]), .Z(n7372) );
  AND U8293 ( .A(p_input[170]), .B(p_input[1170]), .Z(n7373) );
  AND U8294 ( .A(p_input[4170]), .B(p_input[3170]), .Z(n7371) );
  AND U8295 ( .A(n7374), .B(n7375), .Z(n7369) );
  AND U8296 ( .A(n7376), .B(p_input[7170]), .Z(n7375) );
  AND U8297 ( .A(p_input[6170]), .B(p_input[5170]), .Z(n7376) );
  AND U8298 ( .A(p_input[9170]), .B(p_input[8170]), .Z(n7374) );
  AND U8299 ( .A(n7377), .B(n7378), .Z(o[16]) );
  AND U8300 ( .A(n7379), .B(n7380), .Z(n7378) );
  AND U8301 ( .A(n7381), .B(p_input[2016]), .Z(n7380) );
  AND U8302 ( .A(p_input[16]), .B(p_input[1016]), .Z(n7381) );
  AND U8303 ( .A(p_input[4016]), .B(p_input[3016]), .Z(n7379) );
  AND U8304 ( .A(n7382), .B(n7383), .Z(n7377) );
  AND U8305 ( .A(n7384), .B(p_input[7016]), .Z(n7383) );
  AND U8306 ( .A(p_input[6016]), .B(p_input[5016]), .Z(n7384) );
  AND U8307 ( .A(p_input[9016]), .B(p_input[8016]), .Z(n7382) );
  AND U8308 ( .A(n7385), .B(n7386), .Z(o[169]) );
  AND U8309 ( .A(n7387), .B(n7388), .Z(n7386) );
  AND U8310 ( .A(n7389), .B(p_input[2169]), .Z(n7388) );
  AND U8311 ( .A(p_input[169]), .B(p_input[1169]), .Z(n7389) );
  AND U8312 ( .A(p_input[4169]), .B(p_input[3169]), .Z(n7387) );
  AND U8313 ( .A(n7390), .B(n7391), .Z(n7385) );
  AND U8314 ( .A(n7392), .B(p_input[7169]), .Z(n7391) );
  AND U8315 ( .A(p_input[6169]), .B(p_input[5169]), .Z(n7392) );
  AND U8316 ( .A(p_input[9169]), .B(p_input[8169]), .Z(n7390) );
  AND U8317 ( .A(n7393), .B(n7394), .Z(o[168]) );
  AND U8318 ( .A(n7395), .B(n7396), .Z(n7394) );
  AND U8319 ( .A(n7397), .B(p_input[2168]), .Z(n7396) );
  AND U8320 ( .A(p_input[168]), .B(p_input[1168]), .Z(n7397) );
  AND U8321 ( .A(p_input[4168]), .B(p_input[3168]), .Z(n7395) );
  AND U8322 ( .A(n7398), .B(n7399), .Z(n7393) );
  AND U8323 ( .A(n7400), .B(p_input[7168]), .Z(n7399) );
  AND U8324 ( .A(p_input[6168]), .B(p_input[5168]), .Z(n7400) );
  AND U8325 ( .A(p_input[9168]), .B(p_input[8168]), .Z(n7398) );
  AND U8326 ( .A(n7401), .B(n7402), .Z(o[167]) );
  AND U8327 ( .A(n7403), .B(n7404), .Z(n7402) );
  AND U8328 ( .A(n7405), .B(p_input[2167]), .Z(n7404) );
  AND U8329 ( .A(p_input[167]), .B(p_input[1167]), .Z(n7405) );
  AND U8330 ( .A(p_input[4167]), .B(p_input[3167]), .Z(n7403) );
  AND U8331 ( .A(n7406), .B(n7407), .Z(n7401) );
  AND U8332 ( .A(n7408), .B(p_input[7167]), .Z(n7407) );
  AND U8333 ( .A(p_input[6167]), .B(p_input[5167]), .Z(n7408) );
  AND U8334 ( .A(p_input[9167]), .B(p_input[8167]), .Z(n7406) );
  AND U8335 ( .A(n7409), .B(n7410), .Z(o[166]) );
  AND U8336 ( .A(n7411), .B(n7412), .Z(n7410) );
  AND U8337 ( .A(n7413), .B(p_input[2166]), .Z(n7412) );
  AND U8338 ( .A(p_input[166]), .B(p_input[1166]), .Z(n7413) );
  AND U8339 ( .A(p_input[4166]), .B(p_input[3166]), .Z(n7411) );
  AND U8340 ( .A(n7414), .B(n7415), .Z(n7409) );
  AND U8341 ( .A(n7416), .B(p_input[7166]), .Z(n7415) );
  AND U8342 ( .A(p_input[6166]), .B(p_input[5166]), .Z(n7416) );
  AND U8343 ( .A(p_input[9166]), .B(p_input[8166]), .Z(n7414) );
  AND U8344 ( .A(n7417), .B(n7418), .Z(o[165]) );
  AND U8345 ( .A(n7419), .B(n7420), .Z(n7418) );
  AND U8346 ( .A(n7421), .B(p_input[2165]), .Z(n7420) );
  AND U8347 ( .A(p_input[165]), .B(p_input[1165]), .Z(n7421) );
  AND U8348 ( .A(p_input[4165]), .B(p_input[3165]), .Z(n7419) );
  AND U8349 ( .A(n7422), .B(n7423), .Z(n7417) );
  AND U8350 ( .A(n7424), .B(p_input[7165]), .Z(n7423) );
  AND U8351 ( .A(p_input[6165]), .B(p_input[5165]), .Z(n7424) );
  AND U8352 ( .A(p_input[9165]), .B(p_input[8165]), .Z(n7422) );
  AND U8353 ( .A(n7425), .B(n7426), .Z(o[164]) );
  AND U8354 ( .A(n7427), .B(n7428), .Z(n7426) );
  AND U8355 ( .A(n7429), .B(p_input[2164]), .Z(n7428) );
  AND U8356 ( .A(p_input[164]), .B(p_input[1164]), .Z(n7429) );
  AND U8357 ( .A(p_input[4164]), .B(p_input[3164]), .Z(n7427) );
  AND U8358 ( .A(n7430), .B(n7431), .Z(n7425) );
  AND U8359 ( .A(n7432), .B(p_input[7164]), .Z(n7431) );
  AND U8360 ( .A(p_input[6164]), .B(p_input[5164]), .Z(n7432) );
  AND U8361 ( .A(p_input[9164]), .B(p_input[8164]), .Z(n7430) );
  AND U8362 ( .A(n7433), .B(n7434), .Z(o[163]) );
  AND U8363 ( .A(n7435), .B(n7436), .Z(n7434) );
  AND U8364 ( .A(n7437), .B(p_input[2163]), .Z(n7436) );
  AND U8365 ( .A(p_input[163]), .B(p_input[1163]), .Z(n7437) );
  AND U8366 ( .A(p_input[4163]), .B(p_input[3163]), .Z(n7435) );
  AND U8367 ( .A(n7438), .B(n7439), .Z(n7433) );
  AND U8368 ( .A(n7440), .B(p_input[7163]), .Z(n7439) );
  AND U8369 ( .A(p_input[6163]), .B(p_input[5163]), .Z(n7440) );
  AND U8370 ( .A(p_input[9163]), .B(p_input[8163]), .Z(n7438) );
  AND U8371 ( .A(n7441), .B(n7442), .Z(o[162]) );
  AND U8372 ( .A(n7443), .B(n7444), .Z(n7442) );
  AND U8373 ( .A(n7445), .B(p_input[2162]), .Z(n7444) );
  AND U8374 ( .A(p_input[162]), .B(p_input[1162]), .Z(n7445) );
  AND U8375 ( .A(p_input[4162]), .B(p_input[3162]), .Z(n7443) );
  AND U8376 ( .A(n7446), .B(n7447), .Z(n7441) );
  AND U8377 ( .A(n7448), .B(p_input[7162]), .Z(n7447) );
  AND U8378 ( .A(p_input[6162]), .B(p_input[5162]), .Z(n7448) );
  AND U8379 ( .A(p_input[9162]), .B(p_input[8162]), .Z(n7446) );
  AND U8380 ( .A(n7449), .B(n7450), .Z(o[161]) );
  AND U8381 ( .A(n7451), .B(n7452), .Z(n7450) );
  AND U8382 ( .A(n7453), .B(p_input[2161]), .Z(n7452) );
  AND U8383 ( .A(p_input[161]), .B(p_input[1161]), .Z(n7453) );
  AND U8384 ( .A(p_input[4161]), .B(p_input[3161]), .Z(n7451) );
  AND U8385 ( .A(n7454), .B(n7455), .Z(n7449) );
  AND U8386 ( .A(n7456), .B(p_input[7161]), .Z(n7455) );
  AND U8387 ( .A(p_input[6161]), .B(p_input[5161]), .Z(n7456) );
  AND U8388 ( .A(p_input[9161]), .B(p_input[8161]), .Z(n7454) );
  AND U8389 ( .A(n7457), .B(n7458), .Z(o[160]) );
  AND U8390 ( .A(n7459), .B(n7460), .Z(n7458) );
  AND U8391 ( .A(n7461), .B(p_input[2160]), .Z(n7460) );
  AND U8392 ( .A(p_input[160]), .B(p_input[1160]), .Z(n7461) );
  AND U8393 ( .A(p_input[4160]), .B(p_input[3160]), .Z(n7459) );
  AND U8394 ( .A(n7462), .B(n7463), .Z(n7457) );
  AND U8395 ( .A(n7464), .B(p_input[7160]), .Z(n7463) );
  AND U8396 ( .A(p_input[6160]), .B(p_input[5160]), .Z(n7464) );
  AND U8397 ( .A(p_input[9160]), .B(p_input[8160]), .Z(n7462) );
  AND U8398 ( .A(n7465), .B(n7466), .Z(o[15]) );
  AND U8399 ( .A(n7467), .B(n7468), .Z(n7466) );
  AND U8400 ( .A(n7469), .B(p_input[2015]), .Z(n7468) );
  AND U8401 ( .A(p_input[15]), .B(p_input[1015]), .Z(n7469) );
  AND U8402 ( .A(p_input[4015]), .B(p_input[3015]), .Z(n7467) );
  AND U8403 ( .A(n7470), .B(n7471), .Z(n7465) );
  AND U8404 ( .A(n7472), .B(p_input[7015]), .Z(n7471) );
  AND U8405 ( .A(p_input[6015]), .B(p_input[5015]), .Z(n7472) );
  AND U8406 ( .A(p_input[9015]), .B(p_input[8015]), .Z(n7470) );
  AND U8407 ( .A(n7473), .B(n7474), .Z(o[159]) );
  AND U8408 ( .A(n7475), .B(n7476), .Z(n7474) );
  AND U8409 ( .A(n7477), .B(p_input[2159]), .Z(n7476) );
  AND U8410 ( .A(p_input[159]), .B(p_input[1159]), .Z(n7477) );
  AND U8411 ( .A(p_input[4159]), .B(p_input[3159]), .Z(n7475) );
  AND U8412 ( .A(n7478), .B(n7479), .Z(n7473) );
  AND U8413 ( .A(n7480), .B(p_input[7159]), .Z(n7479) );
  AND U8414 ( .A(p_input[6159]), .B(p_input[5159]), .Z(n7480) );
  AND U8415 ( .A(p_input[9159]), .B(p_input[8159]), .Z(n7478) );
  AND U8416 ( .A(n7481), .B(n7482), .Z(o[158]) );
  AND U8417 ( .A(n7483), .B(n7484), .Z(n7482) );
  AND U8418 ( .A(n7485), .B(p_input[2158]), .Z(n7484) );
  AND U8419 ( .A(p_input[158]), .B(p_input[1158]), .Z(n7485) );
  AND U8420 ( .A(p_input[4158]), .B(p_input[3158]), .Z(n7483) );
  AND U8421 ( .A(n7486), .B(n7487), .Z(n7481) );
  AND U8422 ( .A(n7488), .B(p_input[7158]), .Z(n7487) );
  AND U8423 ( .A(p_input[6158]), .B(p_input[5158]), .Z(n7488) );
  AND U8424 ( .A(p_input[9158]), .B(p_input[8158]), .Z(n7486) );
  AND U8425 ( .A(n7489), .B(n7490), .Z(o[157]) );
  AND U8426 ( .A(n7491), .B(n7492), .Z(n7490) );
  AND U8427 ( .A(n7493), .B(p_input[2157]), .Z(n7492) );
  AND U8428 ( .A(p_input[157]), .B(p_input[1157]), .Z(n7493) );
  AND U8429 ( .A(p_input[4157]), .B(p_input[3157]), .Z(n7491) );
  AND U8430 ( .A(n7494), .B(n7495), .Z(n7489) );
  AND U8431 ( .A(n7496), .B(p_input[7157]), .Z(n7495) );
  AND U8432 ( .A(p_input[6157]), .B(p_input[5157]), .Z(n7496) );
  AND U8433 ( .A(p_input[9157]), .B(p_input[8157]), .Z(n7494) );
  AND U8434 ( .A(n7497), .B(n7498), .Z(o[156]) );
  AND U8435 ( .A(n7499), .B(n7500), .Z(n7498) );
  AND U8436 ( .A(n7501), .B(p_input[2156]), .Z(n7500) );
  AND U8437 ( .A(p_input[156]), .B(p_input[1156]), .Z(n7501) );
  AND U8438 ( .A(p_input[4156]), .B(p_input[3156]), .Z(n7499) );
  AND U8439 ( .A(n7502), .B(n7503), .Z(n7497) );
  AND U8440 ( .A(n7504), .B(p_input[7156]), .Z(n7503) );
  AND U8441 ( .A(p_input[6156]), .B(p_input[5156]), .Z(n7504) );
  AND U8442 ( .A(p_input[9156]), .B(p_input[8156]), .Z(n7502) );
  AND U8443 ( .A(n7505), .B(n7506), .Z(o[155]) );
  AND U8444 ( .A(n7507), .B(n7508), .Z(n7506) );
  AND U8445 ( .A(n7509), .B(p_input[2155]), .Z(n7508) );
  AND U8446 ( .A(p_input[155]), .B(p_input[1155]), .Z(n7509) );
  AND U8447 ( .A(p_input[4155]), .B(p_input[3155]), .Z(n7507) );
  AND U8448 ( .A(n7510), .B(n7511), .Z(n7505) );
  AND U8449 ( .A(n7512), .B(p_input[7155]), .Z(n7511) );
  AND U8450 ( .A(p_input[6155]), .B(p_input[5155]), .Z(n7512) );
  AND U8451 ( .A(p_input[9155]), .B(p_input[8155]), .Z(n7510) );
  AND U8452 ( .A(n7513), .B(n7514), .Z(o[154]) );
  AND U8453 ( .A(n7515), .B(n7516), .Z(n7514) );
  AND U8454 ( .A(n7517), .B(p_input[2154]), .Z(n7516) );
  AND U8455 ( .A(p_input[154]), .B(p_input[1154]), .Z(n7517) );
  AND U8456 ( .A(p_input[4154]), .B(p_input[3154]), .Z(n7515) );
  AND U8457 ( .A(n7518), .B(n7519), .Z(n7513) );
  AND U8458 ( .A(n7520), .B(p_input[7154]), .Z(n7519) );
  AND U8459 ( .A(p_input[6154]), .B(p_input[5154]), .Z(n7520) );
  AND U8460 ( .A(p_input[9154]), .B(p_input[8154]), .Z(n7518) );
  AND U8461 ( .A(n7521), .B(n7522), .Z(o[153]) );
  AND U8462 ( .A(n7523), .B(n7524), .Z(n7522) );
  AND U8463 ( .A(n7525), .B(p_input[2153]), .Z(n7524) );
  AND U8464 ( .A(p_input[153]), .B(p_input[1153]), .Z(n7525) );
  AND U8465 ( .A(p_input[4153]), .B(p_input[3153]), .Z(n7523) );
  AND U8466 ( .A(n7526), .B(n7527), .Z(n7521) );
  AND U8467 ( .A(n7528), .B(p_input[7153]), .Z(n7527) );
  AND U8468 ( .A(p_input[6153]), .B(p_input[5153]), .Z(n7528) );
  AND U8469 ( .A(p_input[9153]), .B(p_input[8153]), .Z(n7526) );
  AND U8470 ( .A(n7529), .B(n7530), .Z(o[152]) );
  AND U8471 ( .A(n7531), .B(n7532), .Z(n7530) );
  AND U8472 ( .A(n7533), .B(p_input[2152]), .Z(n7532) );
  AND U8473 ( .A(p_input[152]), .B(p_input[1152]), .Z(n7533) );
  AND U8474 ( .A(p_input[4152]), .B(p_input[3152]), .Z(n7531) );
  AND U8475 ( .A(n7534), .B(n7535), .Z(n7529) );
  AND U8476 ( .A(n7536), .B(p_input[7152]), .Z(n7535) );
  AND U8477 ( .A(p_input[6152]), .B(p_input[5152]), .Z(n7536) );
  AND U8478 ( .A(p_input[9152]), .B(p_input[8152]), .Z(n7534) );
  AND U8479 ( .A(n7537), .B(n7538), .Z(o[151]) );
  AND U8480 ( .A(n7539), .B(n7540), .Z(n7538) );
  AND U8481 ( .A(n7541), .B(p_input[2151]), .Z(n7540) );
  AND U8482 ( .A(p_input[151]), .B(p_input[1151]), .Z(n7541) );
  AND U8483 ( .A(p_input[4151]), .B(p_input[3151]), .Z(n7539) );
  AND U8484 ( .A(n7542), .B(n7543), .Z(n7537) );
  AND U8485 ( .A(n7544), .B(p_input[7151]), .Z(n7543) );
  AND U8486 ( .A(p_input[6151]), .B(p_input[5151]), .Z(n7544) );
  AND U8487 ( .A(p_input[9151]), .B(p_input[8151]), .Z(n7542) );
  AND U8488 ( .A(n7545), .B(n7546), .Z(o[150]) );
  AND U8489 ( .A(n7547), .B(n7548), .Z(n7546) );
  AND U8490 ( .A(n7549), .B(p_input[2150]), .Z(n7548) );
  AND U8491 ( .A(p_input[150]), .B(p_input[1150]), .Z(n7549) );
  AND U8492 ( .A(p_input[4150]), .B(p_input[3150]), .Z(n7547) );
  AND U8493 ( .A(n7550), .B(n7551), .Z(n7545) );
  AND U8494 ( .A(n7552), .B(p_input[7150]), .Z(n7551) );
  AND U8495 ( .A(p_input[6150]), .B(p_input[5150]), .Z(n7552) );
  AND U8496 ( .A(p_input[9150]), .B(p_input[8150]), .Z(n7550) );
  AND U8497 ( .A(n7553), .B(n7554), .Z(o[14]) );
  AND U8498 ( .A(n7555), .B(n7556), .Z(n7554) );
  AND U8499 ( .A(n7557), .B(p_input[2014]), .Z(n7556) );
  AND U8500 ( .A(p_input[14]), .B(p_input[1014]), .Z(n7557) );
  AND U8501 ( .A(p_input[4014]), .B(p_input[3014]), .Z(n7555) );
  AND U8502 ( .A(n7558), .B(n7559), .Z(n7553) );
  AND U8503 ( .A(n7560), .B(p_input[7014]), .Z(n7559) );
  AND U8504 ( .A(p_input[6014]), .B(p_input[5014]), .Z(n7560) );
  AND U8505 ( .A(p_input[9014]), .B(p_input[8014]), .Z(n7558) );
  AND U8506 ( .A(n7561), .B(n7562), .Z(o[149]) );
  AND U8507 ( .A(n7563), .B(n7564), .Z(n7562) );
  AND U8508 ( .A(n7565), .B(p_input[2149]), .Z(n7564) );
  AND U8509 ( .A(p_input[149]), .B(p_input[1149]), .Z(n7565) );
  AND U8510 ( .A(p_input[4149]), .B(p_input[3149]), .Z(n7563) );
  AND U8511 ( .A(n7566), .B(n7567), .Z(n7561) );
  AND U8512 ( .A(n7568), .B(p_input[7149]), .Z(n7567) );
  AND U8513 ( .A(p_input[6149]), .B(p_input[5149]), .Z(n7568) );
  AND U8514 ( .A(p_input[9149]), .B(p_input[8149]), .Z(n7566) );
  AND U8515 ( .A(n7569), .B(n7570), .Z(o[148]) );
  AND U8516 ( .A(n7571), .B(n7572), .Z(n7570) );
  AND U8517 ( .A(n7573), .B(p_input[2148]), .Z(n7572) );
  AND U8518 ( .A(p_input[148]), .B(p_input[1148]), .Z(n7573) );
  AND U8519 ( .A(p_input[4148]), .B(p_input[3148]), .Z(n7571) );
  AND U8520 ( .A(n7574), .B(n7575), .Z(n7569) );
  AND U8521 ( .A(n7576), .B(p_input[7148]), .Z(n7575) );
  AND U8522 ( .A(p_input[6148]), .B(p_input[5148]), .Z(n7576) );
  AND U8523 ( .A(p_input[9148]), .B(p_input[8148]), .Z(n7574) );
  AND U8524 ( .A(n7577), .B(n7578), .Z(o[147]) );
  AND U8525 ( .A(n7579), .B(n7580), .Z(n7578) );
  AND U8526 ( .A(n7581), .B(p_input[2147]), .Z(n7580) );
  AND U8527 ( .A(p_input[147]), .B(p_input[1147]), .Z(n7581) );
  AND U8528 ( .A(p_input[4147]), .B(p_input[3147]), .Z(n7579) );
  AND U8529 ( .A(n7582), .B(n7583), .Z(n7577) );
  AND U8530 ( .A(n7584), .B(p_input[7147]), .Z(n7583) );
  AND U8531 ( .A(p_input[6147]), .B(p_input[5147]), .Z(n7584) );
  AND U8532 ( .A(p_input[9147]), .B(p_input[8147]), .Z(n7582) );
  AND U8533 ( .A(n7585), .B(n7586), .Z(o[146]) );
  AND U8534 ( .A(n7587), .B(n7588), .Z(n7586) );
  AND U8535 ( .A(n7589), .B(p_input[2146]), .Z(n7588) );
  AND U8536 ( .A(p_input[146]), .B(p_input[1146]), .Z(n7589) );
  AND U8537 ( .A(p_input[4146]), .B(p_input[3146]), .Z(n7587) );
  AND U8538 ( .A(n7590), .B(n7591), .Z(n7585) );
  AND U8539 ( .A(n7592), .B(p_input[7146]), .Z(n7591) );
  AND U8540 ( .A(p_input[6146]), .B(p_input[5146]), .Z(n7592) );
  AND U8541 ( .A(p_input[9146]), .B(p_input[8146]), .Z(n7590) );
  AND U8542 ( .A(n7593), .B(n7594), .Z(o[145]) );
  AND U8543 ( .A(n7595), .B(n7596), .Z(n7594) );
  AND U8544 ( .A(n7597), .B(p_input[2145]), .Z(n7596) );
  AND U8545 ( .A(p_input[145]), .B(p_input[1145]), .Z(n7597) );
  AND U8546 ( .A(p_input[4145]), .B(p_input[3145]), .Z(n7595) );
  AND U8547 ( .A(n7598), .B(n7599), .Z(n7593) );
  AND U8548 ( .A(n7600), .B(p_input[7145]), .Z(n7599) );
  AND U8549 ( .A(p_input[6145]), .B(p_input[5145]), .Z(n7600) );
  AND U8550 ( .A(p_input[9145]), .B(p_input[8145]), .Z(n7598) );
  AND U8551 ( .A(n7601), .B(n7602), .Z(o[144]) );
  AND U8552 ( .A(n7603), .B(n7604), .Z(n7602) );
  AND U8553 ( .A(n7605), .B(p_input[2144]), .Z(n7604) );
  AND U8554 ( .A(p_input[144]), .B(p_input[1144]), .Z(n7605) );
  AND U8555 ( .A(p_input[4144]), .B(p_input[3144]), .Z(n7603) );
  AND U8556 ( .A(n7606), .B(n7607), .Z(n7601) );
  AND U8557 ( .A(n7608), .B(p_input[7144]), .Z(n7607) );
  AND U8558 ( .A(p_input[6144]), .B(p_input[5144]), .Z(n7608) );
  AND U8559 ( .A(p_input[9144]), .B(p_input[8144]), .Z(n7606) );
  AND U8560 ( .A(n7609), .B(n7610), .Z(o[143]) );
  AND U8561 ( .A(n7611), .B(n7612), .Z(n7610) );
  AND U8562 ( .A(n7613), .B(p_input[2143]), .Z(n7612) );
  AND U8563 ( .A(p_input[143]), .B(p_input[1143]), .Z(n7613) );
  AND U8564 ( .A(p_input[4143]), .B(p_input[3143]), .Z(n7611) );
  AND U8565 ( .A(n7614), .B(n7615), .Z(n7609) );
  AND U8566 ( .A(n7616), .B(p_input[7143]), .Z(n7615) );
  AND U8567 ( .A(p_input[6143]), .B(p_input[5143]), .Z(n7616) );
  AND U8568 ( .A(p_input[9143]), .B(p_input[8143]), .Z(n7614) );
  AND U8569 ( .A(n7617), .B(n7618), .Z(o[142]) );
  AND U8570 ( .A(n7619), .B(n7620), .Z(n7618) );
  AND U8571 ( .A(n7621), .B(p_input[2142]), .Z(n7620) );
  AND U8572 ( .A(p_input[142]), .B(p_input[1142]), .Z(n7621) );
  AND U8573 ( .A(p_input[4142]), .B(p_input[3142]), .Z(n7619) );
  AND U8574 ( .A(n7622), .B(n7623), .Z(n7617) );
  AND U8575 ( .A(n7624), .B(p_input[7142]), .Z(n7623) );
  AND U8576 ( .A(p_input[6142]), .B(p_input[5142]), .Z(n7624) );
  AND U8577 ( .A(p_input[9142]), .B(p_input[8142]), .Z(n7622) );
  AND U8578 ( .A(n7625), .B(n7626), .Z(o[141]) );
  AND U8579 ( .A(n7627), .B(n7628), .Z(n7626) );
  AND U8580 ( .A(n7629), .B(p_input[2141]), .Z(n7628) );
  AND U8581 ( .A(p_input[141]), .B(p_input[1141]), .Z(n7629) );
  AND U8582 ( .A(p_input[4141]), .B(p_input[3141]), .Z(n7627) );
  AND U8583 ( .A(n7630), .B(n7631), .Z(n7625) );
  AND U8584 ( .A(n7632), .B(p_input[7141]), .Z(n7631) );
  AND U8585 ( .A(p_input[6141]), .B(p_input[5141]), .Z(n7632) );
  AND U8586 ( .A(p_input[9141]), .B(p_input[8141]), .Z(n7630) );
  AND U8587 ( .A(n7633), .B(n7634), .Z(o[140]) );
  AND U8588 ( .A(n7635), .B(n7636), .Z(n7634) );
  AND U8589 ( .A(n7637), .B(p_input[2140]), .Z(n7636) );
  AND U8590 ( .A(p_input[140]), .B(p_input[1140]), .Z(n7637) );
  AND U8591 ( .A(p_input[4140]), .B(p_input[3140]), .Z(n7635) );
  AND U8592 ( .A(n7638), .B(n7639), .Z(n7633) );
  AND U8593 ( .A(n7640), .B(p_input[7140]), .Z(n7639) );
  AND U8594 ( .A(p_input[6140]), .B(p_input[5140]), .Z(n7640) );
  AND U8595 ( .A(p_input[9140]), .B(p_input[8140]), .Z(n7638) );
  AND U8596 ( .A(n7641), .B(n7642), .Z(o[13]) );
  AND U8597 ( .A(n7643), .B(n7644), .Z(n7642) );
  AND U8598 ( .A(n7645), .B(p_input[2013]), .Z(n7644) );
  AND U8599 ( .A(p_input[13]), .B(p_input[1013]), .Z(n7645) );
  AND U8600 ( .A(p_input[4013]), .B(p_input[3013]), .Z(n7643) );
  AND U8601 ( .A(n7646), .B(n7647), .Z(n7641) );
  AND U8602 ( .A(n7648), .B(p_input[7013]), .Z(n7647) );
  AND U8603 ( .A(p_input[6013]), .B(p_input[5013]), .Z(n7648) );
  AND U8604 ( .A(p_input[9013]), .B(p_input[8013]), .Z(n7646) );
  AND U8605 ( .A(n7649), .B(n7650), .Z(o[139]) );
  AND U8606 ( .A(n7651), .B(n7652), .Z(n7650) );
  AND U8607 ( .A(n7653), .B(p_input[2139]), .Z(n7652) );
  AND U8608 ( .A(p_input[139]), .B(p_input[1139]), .Z(n7653) );
  AND U8609 ( .A(p_input[4139]), .B(p_input[3139]), .Z(n7651) );
  AND U8610 ( .A(n7654), .B(n7655), .Z(n7649) );
  AND U8611 ( .A(n7656), .B(p_input[7139]), .Z(n7655) );
  AND U8612 ( .A(p_input[6139]), .B(p_input[5139]), .Z(n7656) );
  AND U8613 ( .A(p_input[9139]), .B(p_input[8139]), .Z(n7654) );
  AND U8614 ( .A(n7657), .B(n7658), .Z(o[138]) );
  AND U8615 ( .A(n7659), .B(n7660), .Z(n7658) );
  AND U8616 ( .A(n7661), .B(p_input[2138]), .Z(n7660) );
  AND U8617 ( .A(p_input[138]), .B(p_input[1138]), .Z(n7661) );
  AND U8618 ( .A(p_input[4138]), .B(p_input[3138]), .Z(n7659) );
  AND U8619 ( .A(n7662), .B(n7663), .Z(n7657) );
  AND U8620 ( .A(n7664), .B(p_input[7138]), .Z(n7663) );
  AND U8621 ( .A(p_input[6138]), .B(p_input[5138]), .Z(n7664) );
  AND U8622 ( .A(p_input[9138]), .B(p_input[8138]), .Z(n7662) );
  AND U8623 ( .A(n7665), .B(n7666), .Z(o[137]) );
  AND U8624 ( .A(n7667), .B(n7668), .Z(n7666) );
  AND U8625 ( .A(n7669), .B(p_input[2137]), .Z(n7668) );
  AND U8626 ( .A(p_input[137]), .B(p_input[1137]), .Z(n7669) );
  AND U8627 ( .A(p_input[4137]), .B(p_input[3137]), .Z(n7667) );
  AND U8628 ( .A(n7670), .B(n7671), .Z(n7665) );
  AND U8629 ( .A(n7672), .B(p_input[7137]), .Z(n7671) );
  AND U8630 ( .A(p_input[6137]), .B(p_input[5137]), .Z(n7672) );
  AND U8631 ( .A(p_input[9137]), .B(p_input[8137]), .Z(n7670) );
  AND U8632 ( .A(n7673), .B(n7674), .Z(o[136]) );
  AND U8633 ( .A(n7675), .B(n7676), .Z(n7674) );
  AND U8634 ( .A(n7677), .B(p_input[2136]), .Z(n7676) );
  AND U8635 ( .A(p_input[136]), .B(p_input[1136]), .Z(n7677) );
  AND U8636 ( .A(p_input[4136]), .B(p_input[3136]), .Z(n7675) );
  AND U8637 ( .A(n7678), .B(n7679), .Z(n7673) );
  AND U8638 ( .A(n7680), .B(p_input[7136]), .Z(n7679) );
  AND U8639 ( .A(p_input[6136]), .B(p_input[5136]), .Z(n7680) );
  AND U8640 ( .A(p_input[9136]), .B(p_input[8136]), .Z(n7678) );
  AND U8641 ( .A(n7681), .B(n7682), .Z(o[135]) );
  AND U8642 ( .A(n7683), .B(n7684), .Z(n7682) );
  AND U8643 ( .A(n7685), .B(p_input[2135]), .Z(n7684) );
  AND U8644 ( .A(p_input[135]), .B(p_input[1135]), .Z(n7685) );
  AND U8645 ( .A(p_input[4135]), .B(p_input[3135]), .Z(n7683) );
  AND U8646 ( .A(n7686), .B(n7687), .Z(n7681) );
  AND U8647 ( .A(n7688), .B(p_input[7135]), .Z(n7687) );
  AND U8648 ( .A(p_input[6135]), .B(p_input[5135]), .Z(n7688) );
  AND U8649 ( .A(p_input[9135]), .B(p_input[8135]), .Z(n7686) );
  AND U8650 ( .A(n7689), .B(n7690), .Z(o[134]) );
  AND U8651 ( .A(n7691), .B(n7692), .Z(n7690) );
  AND U8652 ( .A(n7693), .B(p_input[2134]), .Z(n7692) );
  AND U8653 ( .A(p_input[134]), .B(p_input[1134]), .Z(n7693) );
  AND U8654 ( .A(p_input[4134]), .B(p_input[3134]), .Z(n7691) );
  AND U8655 ( .A(n7694), .B(n7695), .Z(n7689) );
  AND U8656 ( .A(n7696), .B(p_input[7134]), .Z(n7695) );
  AND U8657 ( .A(p_input[6134]), .B(p_input[5134]), .Z(n7696) );
  AND U8658 ( .A(p_input[9134]), .B(p_input[8134]), .Z(n7694) );
  AND U8659 ( .A(n7697), .B(n7698), .Z(o[133]) );
  AND U8660 ( .A(n7699), .B(n7700), .Z(n7698) );
  AND U8661 ( .A(n7701), .B(p_input[2133]), .Z(n7700) );
  AND U8662 ( .A(p_input[133]), .B(p_input[1133]), .Z(n7701) );
  AND U8663 ( .A(p_input[4133]), .B(p_input[3133]), .Z(n7699) );
  AND U8664 ( .A(n7702), .B(n7703), .Z(n7697) );
  AND U8665 ( .A(n7704), .B(p_input[7133]), .Z(n7703) );
  AND U8666 ( .A(p_input[6133]), .B(p_input[5133]), .Z(n7704) );
  AND U8667 ( .A(p_input[9133]), .B(p_input[8133]), .Z(n7702) );
  AND U8668 ( .A(n7705), .B(n7706), .Z(o[132]) );
  AND U8669 ( .A(n7707), .B(n7708), .Z(n7706) );
  AND U8670 ( .A(n7709), .B(p_input[2132]), .Z(n7708) );
  AND U8671 ( .A(p_input[132]), .B(p_input[1132]), .Z(n7709) );
  AND U8672 ( .A(p_input[4132]), .B(p_input[3132]), .Z(n7707) );
  AND U8673 ( .A(n7710), .B(n7711), .Z(n7705) );
  AND U8674 ( .A(n7712), .B(p_input[7132]), .Z(n7711) );
  AND U8675 ( .A(p_input[6132]), .B(p_input[5132]), .Z(n7712) );
  AND U8676 ( .A(p_input[9132]), .B(p_input[8132]), .Z(n7710) );
  AND U8677 ( .A(n7713), .B(n7714), .Z(o[131]) );
  AND U8678 ( .A(n7715), .B(n7716), .Z(n7714) );
  AND U8679 ( .A(n7717), .B(p_input[2131]), .Z(n7716) );
  AND U8680 ( .A(p_input[131]), .B(p_input[1131]), .Z(n7717) );
  AND U8681 ( .A(p_input[4131]), .B(p_input[3131]), .Z(n7715) );
  AND U8682 ( .A(n7718), .B(n7719), .Z(n7713) );
  AND U8683 ( .A(n7720), .B(p_input[7131]), .Z(n7719) );
  AND U8684 ( .A(p_input[6131]), .B(p_input[5131]), .Z(n7720) );
  AND U8685 ( .A(p_input[9131]), .B(p_input[8131]), .Z(n7718) );
  AND U8686 ( .A(n7721), .B(n7722), .Z(o[130]) );
  AND U8687 ( .A(n7723), .B(n7724), .Z(n7722) );
  AND U8688 ( .A(n7725), .B(p_input[2130]), .Z(n7724) );
  AND U8689 ( .A(p_input[130]), .B(p_input[1130]), .Z(n7725) );
  AND U8690 ( .A(p_input[4130]), .B(p_input[3130]), .Z(n7723) );
  AND U8691 ( .A(n7726), .B(n7727), .Z(n7721) );
  AND U8692 ( .A(n7728), .B(p_input[7130]), .Z(n7727) );
  AND U8693 ( .A(p_input[6130]), .B(p_input[5130]), .Z(n7728) );
  AND U8694 ( .A(p_input[9130]), .B(p_input[8130]), .Z(n7726) );
  AND U8695 ( .A(n7729), .B(n7730), .Z(o[12]) );
  AND U8696 ( .A(n7731), .B(n7732), .Z(n7730) );
  AND U8697 ( .A(n7733), .B(p_input[2012]), .Z(n7732) );
  AND U8698 ( .A(p_input[12]), .B(p_input[1012]), .Z(n7733) );
  AND U8699 ( .A(p_input[4012]), .B(p_input[3012]), .Z(n7731) );
  AND U8700 ( .A(n7734), .B(n7735), .Z(n7729) );
  AND U8701 ( .A(n7736), .B(p_input[7012]), .Z(n7735) );
  AND U8702 ( .A(p_input[6012]), .B(p_input[5012]), .Z(n7736) );
  AND U8703 ( .A(p_input[9012]), .B(p_input[8012]), .Z(n7734) );
  AND U8704 ( .A(n7737), .B(n7738), .Z(o[129]) );
  AND U8705 ( .A(n7739), .B(n7740), .Z(n7738) );
  AND U8706 ( .A(n7741), .B(p_input[2129]), .Z(n7740) );
  AND U8707 ( .A(p_input[129]), .B(p_input[1129]), .Z(n7741) );
  AND U8708 ( .A(p_input[4129]), .B(p_input[3129]), .Z(n7739) );
  AND U8709 ( .A(n7742), .B(n7743), .Z(n7737) );
  AND U8710 ( .A(n7744), .B(p_input[7129]), .Z(n7743) );
  AND U8711 ( .A(p_input[6129]), .B(p_input[5129]), .Z(n7744) );
  AND U8712 ( .A(p_input[9129]), .B(p_input[8129]), .Z(n7742) );
  AND U8713 ( .A(n7745), .B(n7746), .Z(o[128]) );
  AND U8714 ( .A(n7747), .B(n7748), .Z(n7746) );
  AND U8715 ( .A(n7749), .B(p_input[2128]), .Z(n7748) );
  AND U8716 ( .A(p_input[128]), .B(p_input[1128]), .Z(n7749) );
  AND U8717 ( .A(p_input[4128]), .B(p_input[3128]), .Z(n7747) );
  AND U8718 ( .A(n7750), .B(n7751), .Z(n7745) );
  AND U8719 ( .A(n7752), .B(p_input[7128]), .Z(n7751) );
  AND U8720 ( .A(p_input[6128]), .B(p_input[5128]), .Z(n7752) );
  AND U8721 ( .A(p_input[9128]), .B(p_input[8128]), .Z(n7750) );
  AND U8722 ( .A(n7753), .B(n7754), .Z(o[127]) );
  AND U8723 ( .A(n7755), .B(n7756), .Z(n7754) );
  AND U8724 ( .A(n7757), .B(p_input[2127]), .Z(n7756) );
  AND U8725 ( .A(p_input[127]), .B(p_input[1127]), .Z(n7757) );
  AND U8726 ( .A(p_input[4127]), .B(p_input[3127]), .Z(n7755) );
  AND U8727 ( .A(n7758), .B(n7759), .Z(n7753) );
  AND U8728 ( .A(n7760), .B(p_input[7127]), .Z(n7759) );
  AND U8729 ( .A(p_input[6127]), .B(p_input[5127]), .Z(n7760) );
  AND U8730 ( .A(p_input[9127]), .B(p_input[8127]), .Z(n7758) );
  AND U8731 ( .A(n7761), .B(n7762), .Z(o[126]) );
  AND U8732 ( .A(n7763), .B(n7764), .Z(n7762) );
  AND U8733 ( .A(n7765), .B(p_input[2126]), .Z(n7764) );
  AND U8734 ( .A(p_input[126]), .B(p_input[1126]), .Z(n7765) );
  AND U8735 ( .A(p_input[4126]), .B(p_input[3126]), .Z(n7763) );
  AND U8736 ( .A(n7766), .B(n7767), .Z(n7761) );
  AND U8737 ( .A(n7768), .B(p_input[7126]), .Z(n7767) );
  AND U8738 ( .A(p_input[6126]), .B(p_input[5126]), .Z(n7768) );
  AND U8739 ( .A(p_input[9126]), .B(p_input[8126]), .Z(n7766) );
  AND U8740 ( .A(n7769), .B(n7770), .Z(o[125]) );
  AND U8741 ( .A(n7771), .B(n7772), .Z(n7770) );
  AND U8742 ( .A(n7773), .B(p_input[2125]), .Z(n7772) );
  AND U8743 ( .A(p_input[125]), .B(p_input[1125]), .Z(n7773) );
  AND U8744 ( .A(p_input[4125]), .B(p_input[3125]), .Z(n7771) );
  AND U8745 ( .A(n7774), .B(n7775), .Z(n7769) );
  AND U8746 ( .A(n7776), .B(p_input[7125]), .Z(n7775) );
  AND U8747 ( .A(p_input[6125]), .B(p_input[5125]), .Z(n7776) );
  AND U8748 ( .A(p_input[9125]), .B(p_input[8125]), .Z(n7774) );
  AND U8749 ( .A(n7777), .B(n7778), .Z(o[124]) );
  AND U8750 ( .A(n7779), .B(n7780), .Z(n7778) );
  AND U8751 ( .A(n7781), .B(p_input[2124]), .Z(n7780) );
  AND U8752 ( .A(p_input[124]), .B(p_input[1124]), .Z(n7781) );
  AND U8753 ( .A(p_input[4124]), .B(p_input[3124]), .Z(n7779) );
  AND U8754 ( .A(n7782), .B(n7783), .Z(n7777) );
  AND U8755 ( .A(n7784), .B(p_input[7124]), .Z(n7783) );
  AND U8756 ( .A(p_input[6124]), .B(p_input[5124]), .Z(n7784) );
  AND U8757 ( .A(p_input[9124]), .B(p_input[8124]), .Z(n7782) );
  AND U8758 ( .A(n7785), .B(n7786), .Z(o[123]) );
  AND U8759 ( .A(n7787), .B(n7788), .Z(n7786) );
  AND U8760 ( .A(n7789), .B(p_input[2123]), .Z(n7788) );
  AND U8761 ( .A(p_input[123]), .B(p_input[1123]), .Z(n7789) );
  AND U8762 ( .A(p_input[4123]), .B(p_input[3123]), .Z(n7787) );
  AND U8763 ( .A(n7790), .B(n7791), .Z(n7785) );
  AND U8764 ( .A(n7792), .B(p_input[7123]), .Z(n7791) );
  AND U8765 ( .A(p_input[6123]), .B(p_input[5123]), .Z(n7792) );
  AND U8766 ( .A(p_input[9123]), .B(p_input[8123]), .Z(n7790) );
  AND U8767 ( .A(n7793), .B(n7794), .Z(o[122]) );
  AND U8768 ( .A(n7795), .B(n7796), .Z(n7794) );
  AND U8769 ( .A(n7797), .B(p_input[2122]), .Z(n7796) );
  AND U8770 ( .A(p_input[122]), .B(p_input[1122]), .Z(n7797) );
  AND U8771 ( .A(p_input[4122]), .B(p_input[3122]), .Z(n7795) );
  AND U8772 ( .A(n7798), .B(n7799), .Z(n7793) );
  AND U8773 ( .A(n7800), .B(p_input[7122]), .Z(n7799) );
  AND U8774 ( .A(p_input[6122]), .B(p_input[5122]), .Z(n7800) );
  AND U8775 ( .A(p_input[9122]), .B(p_input[8122]), .Z(n7798) );
  AND U8776 ( .A(n7801), .B(n7802), .Z(o[121]) );
  AND U8777 ( .A(n7803), .B(n7804), .Z(n7802) );
  AND U8778 ( .A(n7805), .B(p_input[2121]), .Z(n7804) );
  AND U8779 ( .A(p_input[121]), .B(p_input[1121]), .Z(n7805) );
  AND U8780 ( .A(p_input[4121]), .B(p_input[3121]), .Z(n7803) );
  AND U8781 ( .A(n7806), .B(n7807), .Z(n7801) );
  AND U8782 ( .A(n7808), .B(p_input[7121]), .Z(n7807) );
  AND U8783 ( .A(p_input[6121]), .B(p_input[5121]), .Z(n7808) );
  AND U8784 ( .A(p_input[9121]), .B(p_input[8121]), .Z(n7806) );
  AND U8785 ( .A(n7809), .B(n7810), .Z(o[120]) );
  AND U8786 ( .A(n7811), .B(n7812), .Z(n7810) );
  AND U8787 ( .A(n7813), .B(p_input[2120]), .Z(n7812) );
  AND U8788 ( .A(p_input[120]), .B(p_input[1120]), .Z(n7813) );
  AND U8789 ( .A(p_input[4120]), .B(p_input[3120]), .Z(n7811) );
  AND U8790 ( .A(n7814), .B(n7815), .Z(n7809) );
  AND U8791 ( .A(n7816), .B(p_input[7120]), .Z(n7815) );
  AND U8792 ( .A(p_input[6120]), .B(p_input[5120]), .Z(n7816) );
  AND U8793 ( .A(p_input[9120]), .B(p_input[8120]), .Z(n7814) );
  AND U8794 ( .A(n7817), .B(n7818), .Z(o[11]) );
  AND U8795 ( .A(n7819), .B(n7820), .Z(n7818) );
  AND U8796 ( .A(n7821), .B(p_input[2011]), .Z(n7820) );
  AND U8797 ( .A(p_input[11]), .B(p_input[1011]), .Z(n7821) );
  AND U8798 ( .A(p_input[4011]), .B(p_input[3011]), .Z(n7819) );
  AND U8799 ( .A(n7822), .B(n7823), .Z(n7817) );
  AND U8800 ( .A(n7824), .B(p_input[7011]), .Z(n7823) );
  AND U8801 ( .A(p_input[6011]), .B(p_input[5011]), .Z(n7824) );
  AND U8802 ( .A(p_input[9011]), .B(p_input[8011]), .Z(n7822) );
  AND U8803 ( .A(n7825), .B(n7826), .Z(o[119]) );
  AND U8804 ( .A(n7827), .B(n7828), .Z(n7826) );
  AND U8805 ( .A(n7829), .B(p_input[2119]), .Z(n7828) );
  AND U8806 ( .A(p_input[119]), .B(p_input[1119]), .Z(n7829) );
  AND U8807 ( .A(p_input[4119]), .B(p_input[3119]), .Z(n7827) );
  AND U8808 ( .A(n7830), .B(n7831), .Z(n7825) );
  AND U8809 ( .A(n7832), .B(p_input[7119]), .Z(n7831) );
  AND U8810 ( .A(p_input[6119]), .B(p_input[5119]), .Z(n7832) );
  AND U8811 ( .A(p_input[9119]), .B(p_input[8119]), .Z(n7830) );
  AND U8812 ( .A(n7833), .B(n7834), .Z(o[118]) );
  AND U8813 ( .A(n7835), .B(n7836), .Z(n7834) );
  AND U8814 ( .A(n7837), .B(p_input[2118]), .Z(n7836) );
  AND U8815 ( .A(p_input[118]), .B(p_input[1118]), .Z(n7837) );
  AND U8816 ( .A(p_input[4118]), .B(p_input[3118]), .Z(n7835) );
  AND U8817 ( .A(n7838), .B(n7839), .Z(n7833) );
  AND U8818 ( .A(n7840), .B(p_input[7118]), .Z(n7839) );
  AND U8819 ( .A(p_input[6118]), .B(p_input[5118]), .Z(n7840) );
  AND U8820 ( .A(p_input[9118]), .B(p_input[8118]), .Z(n7838) );
  AND U8821 ( .A(n7841), .B(n7842), .Z(o[117]) );
  AND U8822 ( .A(n7843), .B(n7844), .Z(n7842) );
  AND U8823 ( .A(n7845), .B(p_input[2117]), .Z(n7844) );
  AND U8824 ( .A(p_input[117]), .B(p_input[1117]), .Z(n7845) );
  AND U8825 ( .A(p_input[4117]), .B(p_input[3117]), .Z(n7843) );
  AND U8826 ( .A(n7846), .B(n7847), .Z(n7841) );
  AND U8827 ( .A(n7848), .B(p_input[7117]), .Z(n7847) );
  AND U8828 ( .A(p_input[6117]), .B(p_input[5117]), .Z(n7848) );
  AND U8829 ( .A(p_input[9117]), .B(p_input[8117]), .Z(n7846) );
  AND U8830 ( .A(n7849), .B(n7850), .Z(o[116]) );
  AND U8831 ( .A(n7851), .B(n7852), .Z(n7850) );
  AND U8832 ( .A(n7853), .B(p_input[2116]), .Z(n7852) );
  AND U8833 ( .A(p_input[116]), .B(p_input[1116]), .Z(n7853) );
  AND U8834 ( .A(p_input[4116]), .B(p_input[3116]), .Z(n7851) );
  AND U8835 ( .A(n7854), .B(n7855), .Z(n7849) );
  AND U8836 ( .A(n7856), .B(p_input[7116]), .Z(n7855) );
  AND U8837 ( .A(p_input[6116]), .B(p_input[5116]), .Z(n7856) );
  AND U8838 ( .A(p_input[9116]), .B(p_input[8116]), .Z(n7854) );
  AND U8839 ( .A(n7857), .B(n7858), .Z(o[115]) );
  AND U8840 ( .A(n7859), .B(n7860), .Z(n7858) );
  AND U8841 ( .A(n7861), .B(p_input[2115]), .Z(n7860) );
  AND U8842 ( .A(p_input[115]), .B(p_input[1115]), .Z(n7861) );
  AND U8843 ( .A(p_input[4115]), .B(p_input[3115]), .Z(n7859) );
  AND U8844 ( .A(n7862), .B(n7863), .Z(n7857) );
  AND U8845 ( .A(n7864), .B(p_input[7115]), .Z(n7863) );
  AND U8846 ( .A(p_input[6115]), .B(p_input[5115]), .Z(n7864) );
  AND U8847 ( .A(p_input[9115]), .B(p_input[8115]), .Z(n7862) );
  AND U8848 ( .A(n7865), .B(n7866), .Z(o[114]) );
  AND U8849 ( .A(n7867), .B(n7868), .Z(n7866) );
  AND U8850 ( .A(n7869), .B(p_input[2114]), .Z(n7868) );
  AND U8851 ( .A(p_input[114]), .B(p_input[1114]), .Z(n7869) );
  AND U8852 ( .A(p_input[4114]), .B(p_input[3114]), .Z(n7867) );
  AND U8853 ( .A(n7870), .B(n7871), .Z(n7865) );
  AND U8854 ( .A(n7872), .B(p_input[7114]), .Z(n7871) );
  AND U8855 ( .A(p_input[6114]), .B(p_input[5114]), .Z(n7872) );
  AND U8856 ( .A(p_input[9114]), .B(p_input[8114]), .Z(n7870) );
  AND U8857 ( .A(n7873), .B(n7874), .Z(o[113]) );
  AND U8858 ( .A(n7875), .B(n7876), .Z(n7874) );
  AND U8859 ( .A(n7877), .B(p_input[2113]), .Z(n7876) );
  AND U8860 ( .A(p_input[113]), .B(p_input[1113]), .Z(n7877) );
  AND U8861 ( .A(p_input[4113]), .B(p_input[3113]), .Z(n7875) );
  AND U8862 ( .A(n7878), .B(n7879), .Z(n7873) );
  AND U8863 ( .A(n7880), .B(p_input[7113]), .Z(n7879) );
  AND U8864 ( .A(p_input[6113]), .B(p_input[5113]), .Z(n7880) );
  AND U8865 ( .A(p_input[9113]), .B(p_input[8113]), .Z(n7878) );
  AND U8866 ( .A(n7881), .B(n7882), .Z(o[112]) );
  AND U8867 ( .A(n7883), .B(n7884), .Z(n7882) );
  AND U8868 ( .A(n7885), .B(p_input[2112]), .Z(n7884) );
  AND U8869 ( .A(p_input[112]), .B(p_input[1112]), .Z(n7885) );
  AND U8870 ( .A(p_input[4112]), .B(p_input[3112]), .Z(n7883) );
  AND U8871 ( .A(n7886), .B(n7887), .Z(n7881) );
  AND U8872 ( .A(n7888), .B(p_input[7112]), .Z(n7887) );
  AND U8873 ( .A(p_input[6112]), .B(p_input[5112]), .Z(n7888) );
  AND U8874 ( .A(p_input[9112]), .B(p_input[8112]), .Z(n7886) );
  AND U8875 ( .A(n7889), .B(n7890), .Z(o[111]) );
  AND U8876 ( .A(n7891), .B(n7892), .Z(n7890) );
  AND U8877 ( .A(n7893), .B(p_input[2111]), .Z(n7892) );
  AND U8878 ( .A(p_input[111]), .B(p_input[1111]), .Z(n7893) );
  AND U8879 ( .A(p_input[4111]), .B(p_input[3111]), .Z(n7891) );
  AND U8880 ( .A(n7894), .B(n7895), .Z(n7889) );
  AND U8881 ( .A(n7896), .B(p_input[7111]), .Z(n7895) );
  AND U8882 ( .A(p_input[6111]), .B(p_input[5111]), .Z(n7896) );
  AND U8883 ( .A(p_input[9111]), .B(p_input[8111]), .Z(n7894) );
  AND U8884 ( .A(n7897), .B(n7898), .Z(o[110]) );
  AND U8885 ( .A(n7899), .B(n7900), .Z(n7898) );
  AND U8886 ( .A(n7901), .B(p_input[2110]), .Z(n7900) );
  AND U8887 ( .A(p_input[1110]), .B(p_input[110]), .Z(n7901) );
  AND U8888 ( .A(p_input[4110]), .B(p_input[3110]), .Z(n7899) );
  AND U8889 ( .A(n7902), .B(n7903), .Z(n7897) );
  AND U8890 ( .A(n7904), .B(p_input[7110]), .Z(n7903) );
  AND U8891 ( .A(p_input[6110]), .B(p_input[5110]), .Z(n7904) );
  AND U8892 ( .A(p_input[9110]), .B(p_input[8110]), .Z(n7902) );
  AND U8893 ( .A(n7905), .B(n7906), .Z(o[10]) );
  AND U8894 ( .A(n7907), .B(n7908), .Z(n7906) );
  AND U8895 ( .A(n7909), .B(p_input[2010]), .Z(n7908) );
  AND U8896 ( .A(p_input[10]), .B(p_input[1010]), .Z(n7909) );
  AND U8897 ( .A(p_input[4010]), .B(p_input[3010]), .Z(n7907) );
  AND U8898 ( .A(n7910), .B(n7911), .Z(n7905) );
  AND U8899 ( .A(n7912), .B(p_input[7010]), .Z(n7911) );
  AND U8900 ( .A(p_input[6010]), .B(p_input[5010]), .Z(n7912) );
  AND U8901 ( .A(p_input[9010]), .B(p_input[8010]), .Z(n7910) );
  AND U8902 ( .A(n7913), .B(n7914), .Z(o[109]) );
  AND U8903 ( .A(n7915), .B(n7916), .Z(n7914) );
  AND U8904 ( .A(n7917), .B(p_input[2109]), .Z(n7916) );
  AND U8905 ( .A(p_input[1109]), .B(p_input[109]), .Z(n7917) );
  AND U8906 ( .A(p_input[4109]), .B(p_input[3109]), .Z(n7915) );
  AND U8907 ( .A(n7918), .B(n7919), .Z(n7913) );
  AND U8908 ( .A(n7920), .B(p_input[7109]), .Z(n7919) );
  AND U8909 ( .A(p_input[6109]), .B(p_input[5109]), .Z(n7920) );
  AND U8910 ( .A(p_input[9109]), .B(p_input[8109]), .Z(n7918) );
  AND U8911 ( .A(n7921), .B(n7922), .Z(o[108]) );
  AND U8912 ( .A(n7923), .B(n7924), .Z(n7922) );
  AND U8913 ( .A(n7925), .B(p_input[2108]), .Z(n7924) );
  AND U8914 ( .A(p_input[1108]), .B(p_input[108]), .Z(n7925) );
  AND U8915 ( .A(p_input[4108]), .B(p_input[3108]), .Z(n7923) );
  AND U8916 ( .A(n7926), .B(n7927), .Z(n7921) );
  AND U8917 ( .A(n7928), .B(p_input[7108]), .Z(n7927) );
  AND U8918 ( .A(p_input[6108]), .B(p_input[5108]), .Z(n7928) );
  AND U8919 ( .A(p_input[9108]), .B(p_input[8108]), .Z(n7926) );
  AND U8920 ( .A(n7929), .B(n7930), .Z(o[107]) );
  AND U8921 ( .A(n7931), .B(n7932), .Z(n7930) );
  AND U8922 ( .A(n7933), .B(p_input[2107]), .Z(n7932) );
  AND U8923 ( .A(p_input[1107]), .B(p_input[107]), .Z(n7933) );
  AND U8924 ( .A(p_input[4107]), .B(p_input[3107]), .Z(n7931) );
  AND U8925 ( .A(n7934), .B(n7935), .Z(n7929) );
  AND U8926 ( .A(n7936), .B(p_input[7107]), .Z(n7935) );
  AND U8927 ( .A(p_input[6107]), .B(p_input[5107]), .Z(n7936) );
  AND U8928 ( .A(p_input[9107]), .B(p_input[8107]), .Z(n7934) );
  AND U8929 ( .A(n7937), .B(n7938), .Z(o[106]) );
  AND U8930 ( .A(n7939), .B(n7940), .Z(n7938) );
  AND U8931 ( .A(n7941), .B(p_input[2106]), .Z(n7940) );
  AND U8932 ( .A(p_input[1106]), .B(p_input[106]), .Z(n7941) );
  AND U8933 ( .A(p_input[4106]), .B(p_input[3106]), .Z(n7939) );
  AND U8934 ( .A(n7942), .B(n7943), .Z(n7937) );
  AND U8935 ( .A(n7944), .B(p_input[7106]), .Z(n7943) );
  AND U8936 ( .A(p_input[6106]), .B(p_input[5106]), .Z(n7944) );
  AND U8937 ( .A(p_input[9106]), .B(p_input[8106]), .Z(n7942) );
  AND U8938 ( .A(n7945), .B(n7946), .Z(o[105]) );
  AND U8939 ( .A(n7947), .B(n7948), .Z(n7946) );
  AND U8940 ( .A(n7949), .B(p_input[2105]), .Z(n7948) );
  AND U8941 ( .A(p_input[1105]), .B(p_input[105]), .Z(n7949) );
  AND U8942 ( .A(p_input[4105]), .B(p_input[3105]), .Z(n7947) );
  AND U8943 ( .A(n7950), .B(n7951), .Z(n7945) );
  AND U8944 ( .A(n7952), .B(p_input[7105]), .Z(n7951) );
  AND U8945 ( .A(p_input[6105]), .B(p_input[5105]), .Z(n7952) );
  AND U8946 ( .A(p_input[9105]), .B(p_input[8105]), .Z(n7950) );
  AND U8947 ( .A(n7953), .B(n7954), .Z(o[104]) );
  AND U8948 ( .A(n7955), .B(n7956), .Z(n7954) );
  AND U8949 ( .A(n7957), .B(p_input[2104]), .Z(n7956) );
  AND U8950 ( .A(p_input[1104]), .B(p_input[104]), .Z(n7957) );
  AND U8951 ( .A(p_input[4104]), .B(p_input[3104]), .Z(n7955) );
  AND U8952 ( .A(n7958), .B(n7959), .Z(n7953) );
  AND U8953 ( .A(n7960), .B(p_input[7104]), .Z(n7959) );
  AND U8954 ( .A(p_input[6104]), .B(p_input[5104]), .Z(n7960) );
  AND U8955 ( .A(p_input[9104]), .B(p_input[8104]), .Z(n7958) );
  AND U8956 ( .A(n7961), .B(n7962), .Z(o[103]) );
  AND U8957 ( .A(n7963), .B(n7964), .Z(n7962) );
  AND U8958 ( .A(n7965), .B(p_input[2103]), .Z(n7964) );
  AND U8959 ( .A(p_input[1103]), .B(p_input[103]), .Z(n7965) );
  AND U8960 ( .A(p_input[4103]), .B(p_input[3103]), .Z(n7963) );
  AND U8961 ( .A(n7966), .B(n7967), .Z(n7961) );
  AND U8962 ( .A(n7968), .B(p_input[7103]), .Z(n7967) );
  AND U8963 ( .A(p_input[6103]), .B(p_input[5103]), .Z(n7968) );
  AND U8964 ( .A(p_input[9103]), .B(p_input[8103]), .Z(n7966) );
  AND U8965 ( .A(n7969), .B(n7970), .Z(o[102]) );
  AND U8966 ( .A(n7971), .B(n7972), .Z(n7970) );
  AND U8967 ( .A(n7973), .B(p_input[2102]), .Z(n7972) );
  AND U8968 ( .A(p_input[1102]), .B(p_input[102]), .Z(n7973) );
  AND U8969 ( .A(p_input[4102]), .B(p_input[3102]), .Z(n7971) );
  AND U8970 ( .A(n7974), .B(n7975), .Z(n7969) );
  AND U8971 ( .A(n7976), .B(p_input[7102]), .Z(n7975) );
  AND U8972 ( .A(p_input[6102]), .B(p_input[5102]), .Z(n7976) );
  AND U8973 ( .A(p_input[9102]), .B(p_input[8102]), .Z(n7974) );
  AND U8974 ( .A(n7977), .B(n7978), .Z(o[101]) );
  AND U8975 ( .A(n7979), .B(n7980), .Z(n7978) );
  AND U8976 ( .A(n7981), .B(p_input[2101]), .Z(n7980) );
  AND U8977 ( .A(p_input[1101]), .B(p_input[101]), .Z(n7981) );
  AND U8978 ( .A(p_input[4101]), .B(p_input[3101]), .Z(n7979) );
  AND U8979 ( .A(n7982), .B(n7983), .Z(n7977) );
  AND U8980 ( .A(n7984), .B(p_input[7101]), .Z(n7983) );
  AND U8981 ( .A(p_input[6101]), .B(p_input[5101]), .Z(n7984) );
  AND U8982 ( .A(p_input[9101]), .B(p_input[8101]), .Z(n7982) );
  AND U8983 ( .A(n7985), .B(n7986), .Z(o[100]) );
  AND U8984 ( .A(n7987), .B(n7988), .Z(n7986) );
  AND U8985 ( .A(n7989), .B(p_input[2100]), .Z(n7988) );
  AND U8986 ( .A(p_input[1100]), .B(p_input[100]), .Z(n7989) );
  AND U8987 ( .A(p_input[4100]), .B(p_input[3100]), .Z(n7987) );
  AND U8988 ( .A(n7990), .B(n7991), .Z(n7985) );
  AND U8989 ( .A(n7992), .B(p_input[7100]), .Z(n7991) );
  AND U8990 ( .A(p_input[6100]), .B(p_input[5100]), .Z(n7992) );
  AND U8991 ( .A(p_input[9100]), .B(p_input[8100]), .Z(n7990) );
  AND U8992 ( .A(n7993), .B(n7994), .Z(o[0]) );
  AND U8993 ( .A(n7995), .B(n7996), .Z(n7994) );
  AND U8994 ( .A(n7997), .B(p_input[2000]), .Z(n7996) );
  AND U8995 ( .A(p_input[1000]), .B(p_input[0]), .Z(n7997) );
  AND U8996 ( .A(p_input[4000]), .B(p_input[3000]), .Z(n7995) );
  AND U8997 ( .A(n7998), .B(n7999), .Z(n7993) );
  AND U8998 ( .A(n8000), .B(p_input[7000]), .Z(n7999) );
  AND U8999 ( .A(p_input[6000]), .B(p_input[5000]), .Z(n8000) );
  AND U9000 ( .A(p_input[9000]), .B(p_input[8000]), .Z(n7998) );
endmodule

