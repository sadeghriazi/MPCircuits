
module auction_BMR_N5_W16 ( p_input, o );
  input [511:0] p_input;
  output [20:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537;

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(o[4]), .B(n3), .Z(n1) );
  XOR U3 ( .A(n2), .B(n4), .Z(n3) );
  XOR U4 ( .A(n5), .B(n6), .Z(o[8]) );
  AND U5 ( .A(o[4]), .B(n7), .Z(n5) );
  XOR U6 ( .A(n8), .B(n9), .Z(n7) );
  XOR U7 ( .A(n10), .B(n11), .Z(o[7]) );
  AND U8 ( .A(o[4]), .B(n12), .Z(n10) );
  XOR U9 ( .A(n13), .B(n14), .Z(n12) );
  XOR U10 ( .A(n15), .B(n16), .Z(o[6]) );
  AND U11 ( .A(o[4]), .B(n17), .Z(n15) );
  XOR U12 ( .A(n18), .B(n19), .Z(n17) );
  XNOR U13 ( .A(n20), .B(n21), .Z(o[5]) );
  AND U14 ( .A(o[4]), .B(n22), .Z(n20) );
  XNOR U15 ( .A(n23), .B(n21), .Z(n22) );
  XNOR U16 ( .A(n24), .B(n25), .Z(o[20]) );
  AND U17 ( .A(o[4]), .B(n26), .Z(n24) );
  XOR U18 ( .A(n27), .B(n25), .Z(n26) );
  XOR U19 ( .A(n28), .B(n29), .Z(o[19]) );
  AND U20 ( .A(o[4]), .B(n30), .Z(n28) );
  XOR U21 ( .A(n31), .B(n32), .Z(n30) );
  XOR U22 ( .A(n33), .B(n34), .Z(o[18]) );
  AND U23 ( .A(o[4]), .B(n35), .Z(n33) );
  XOR U24 ( .A(n36), .B(n37), .Z(n35) );
  XOR U25 ( .A(n38), .B(n39), .Z(o[17]) );
  AND U26 ( .A(o[4]), .B(n40), .Z(n38) );
  XOR U27 ( .A(n41), .B(n42), .Z(n40) );
  XOR U28 ( .A(n43), .B(n44), .Z(o[16]) );
  AND U29 ( .A(o[4]), .B(n45), .Z(n43) );
  XOR U30 ( .A(n46), .B(n47), .Z(n45) );
  XOR U31 ( .A(n48), .B(n49), .Z(o[15]) );
  AND U32 ( .A(o[4]), .B(n50), .Z(n48) );
  XOR U33 ( .A(n51), .B(n52), .Z(n50) );
  XOR U34 ( .A(n53), .B(n54), .Z(o[14]) );
  AND U35 ( .A(o[4]), .B(n55), .Z(n53) );
  XOR U36 ( .A(n56), .B(n57), .Z(n55) );
  XOR U37 ( .A(n58), .B(n59), .Z(o[13]) );
  AND U38 ( .A(o[4]), .B(n60), .Z(n58) );
  XOR U39 ( .A(n61), .B(n62), .Z(n60) );
  XOR U40 ( .A(n63), .B(n64), .Z(o[12]) );
  AND U41 ( .A(o[4]), .B(n65), .Z(n63) );
  XOR U42 ( .A(n66), .B(n67), .Z(n65) );
  XOR U43 ( .A(n68), .B(n69), .Z(o[11]) );
  AND U44 ( .A(o[4]), .B(n70), .Z(n68) );
  XOR U45 ( .A(n71), .B(n72), .Z(n70) );
  XOR U46 ( .A(n73), .B(n74), .Z(o[10]) );
  AND U47 ( .A(o[4]), .B(n75), .Z(n73) );
  XOR U48 ( .A(n76), .B(n77), .Z(n75) );
  XOR U49 ( .A(n78), .B(n79), .Z(o[0]) );
  AND U50 ( .A(o[1]), .B(n80), .Z(n79) );
  XNOR U51 ( .A(n81), .B(n82), .Z(n80) );
  XNOR U52 ( .A(n83), .B(n78), .Z(n82) );
  AND U53 ( .A(o[2]), .B(n84), .Z(n83) );
  XNOR U54 ( .A(n85), .B(n86), .Z(n84) );
  XNOR U55 ( .A(n87), .B(n81), .Z(n86) );
  AND U56 ( .A(o[3]), .B(n88), .Z(n87) );
  XNOR U57 ( .A(n85), .B(n89), .Z(n88) );
  XNOR U58 ( .A(n90), .B(n91), .Z(n89) );
  AND U59 ( .A(o[4]), .B(n92), .Z(n90) );
  XOR U60 ( .A(n91), .B(n93), .Z(n92) );
  XOR U61 ( .A(n94), .B(n95), .Z(n85) );
  AND U62 ( .A(o[4]), .B(n96), .Z(n95) );
  XOR U63 ( .A(n94), .B(n97), .Z(n96) );
  XOR U64 ( .A(n98), .B(n99), .Z(n81) );
  AND U65 ( .A(o[3]), .B(n100), .Z(n99) );
  XNOR U66 ( .A(n98), .B(n101), .Z(n100) );
  XNOR U67 ( .A(n102), .B(n103), .Z(n101) );
  AND U68 ( .A(o[4]), .B(n104), .Z(n102) );
  XOR U69 ( .A(n103), .B(n105), .Z(n104) );
  XOR U70 ( .A(n106), .B(n107), .Z(n98) );
  AND U71 ( .A(o[4]), .B(n108), .Z(n107) );
  XOR U72 ( .A(n106), .B(n109), .Z(n108) );
  XOR U73 ( .A(n110), .B(n111), .Z(o[1]) );
  AND U74 ( .A(o[2]), .B(n112), .Z(n111) );
  XNOR U75 ( .A(n113), .B(n114), .Z(n112) );
  XNOR U76 ( .A(n115), .B(n110), .Z(n114) );
  AND U77 ( .A(o[3]), .B(n116), .Z(n115) );
  XNOR U78 ( .A(n113), .B(n117), .Z(n116) );
  XNOR U79 ( .A(n118), .B(n119), .Z(n117) );
  AND U80 ( .A(o[4]), .B(n120), .Z(n118) );
  XOR U81 ( .A(n119), .B(n121), .Z(n120) );
  XOR U82 ( .A(n122), .B(n123), .Z(n113) );
  AND U83 ( .A(o[4]), .B(n124), .Z(n123) );
  XOR U84 ( .A(n122), .B(n125), .Z(n124) );
  XOR U85 ( .A(n126), .B(n127), .Z(n110) );
  AND U86 ( .A(o[3]), .B(n128), .Z(n127) );
  XNOR U87 ( .A(n126), .B(n129), .Z(n128) );
  XNOR U88 ( .A(n130), .B(n131), .Z(n129) );
  AND U89 ( .A(o[4]), .B(n132), .Z(n130) );
  XOR U90 ( .A(n131), .B(n133), .Z(n132) );
  XOR U91 ( .A(n134), .B(n135), .Z(n126) );
  AND U92 ( .A(o[4]), .B(n136), .Z(n135) );
  XOR U93 ( .A(n134), .B(n137), .Z(n136) );
  XOR U94 ( .A(n138), .B(n139), .Z(n78) );
  AND U95 ( .A(o[2]), .B(n140), .Z(n139) );
  XNOR U96 ( .A(n141), .B(n142), .Z(n140) );
  XNOR U97 ( .A(n143), .B(n138), .Z(n142) );
  AND U98 ( .A(o[3]), .B(n144), .Z(n143) );
  XNOR U99 ( .A(n141), .B(n145), .Z(n144) );
  XNOR U100 ( .A(n146), .B(n147), .Z(n145) );
  AND U101 ( .A(o[4]), .B(n148), .Z(n146) );
  XOR U102 ( .A(n147), .B(n149), .Z(n148) );
  XOR U103 ( .A(n150), .B(n151), .Z(n141) );
  AND U104 ( .A(o[4]), .B(n152), .Z(n151) );
  XOR U105 ( .A(n150), .B(n153), .Z(n152) );
  XOR U106 ( .A(n154), .B(n155), .Z(o[2]) );
  AND U107 ( .A(o[3]), .B(n156), .Z(n155) );
  XNOR U108 ( .A(n154), .B(n157), .Z(n156) );
  XNOR U109 ( .A(n158), .B(n159), .Z(n157) );
  AND U110 ( .A(o[4]), .B(n160), .Z(n158) );
  XOR U111 ( .A(n159), .B(n161), .Z(n160) );
  XOR U112 ( .A(n162), .B(n163), .Z(n154) );
  AND U113 ( .A(o[4]), .B(n164), .Z(n163) );
  XOR U114 ( .A(n162), .B(n165), .Z(n164) );
  XOR U115 ( .A(n166), .B(n167), .Z(n138) );
  AND U116 ( .A(o[3]), .B(n168), .Z(n167) );
  XNOR U117 ( .A(n166), .B(n169), .Z(n168) );
  XNOR U118 ( .A(n170), .B(n171), .Z(n169) );
  AND U119 ( .A(o[4]), .B(n172), .Z(n170) );
  XOR U120 ( .A(n171), .B(n173), .Z(n172) );
  XOR U121 ( .A(n174), .B(n175), .Z(o[3]) );
  AND U122 ( .A(o[4]), .B(n176), .Z(n175) );
  XOR U123 ( .A(n174), .B(n177), .Z(n176) );
  XOR U124 ( .A(n178), .B(n179), .Z(n166) );
  AND U125 ( .A(o[4]), .B(n180), .Z(n179) );
  XOR U126 ( .A(n178), .B(n181), .Z(n180) );
  XOR U127 ( .A(n182), .B(n183), .Z(o[4]) );
  AND U128 ( .A(n184), .B(n185), .Z(n183) );
  XOR U129 ( .A(n182), .B(n27), .Z(n185) );
  XNOR U130 ( .A(n186), .B(n187), .Z(n27) );
  AND U131 ( .A(n188), .B(n177), .Z(n187) );
  AND U132 ( .A(n186), .B(n189), .Z(n188) );
  XNOR U133 ( .A(n25), .B(n182), .Z(n184) );
  XOR U134 ( .A(n190), .B(n191), .Z(n25) );
  AND U135 ( .A(n192), .B(n174), .Z(n191) );
  NOR U136 ( .A(n190), .B(n193), .Z(n192) );
  XOR U137 ( .A(n194), .B(n195), .Z(n182) );
  AND U138 ( .A(n196), .B(n197), .Z(n195) );
  XOR U139 ( .A(n194), .B(n31), .Z(n197) );
  XOR U140 ( .A(n198), .B(n199), .Z(n31) );
  AND U141 ( .A(n177), .B(n200), .Z(n199) );
  XOR U142 ( .A(n201), .B(n198), .Z(n200) );
  XNOR U143 ( .A(n32), .B(n194), .Z(n196) );
  IV U144 ( .A(n29), .Z(n32) );
  XNOR U145 ( .A(n202), .B(n203), .Z(n29) );
  AND U146 ( .A(n174), .B(n204), .Z(n203) );
  XOR U147 ( .A(n205), .B(n202), .Z(n204) );
  XOR U148 ( .A(n206), .B(n207), .Z(n194) );
  AND U149 ( .A(n208), .B(n209), .Z(n207) );
  XOR U150 ( .A(n206), .B(n36), .Z(n209) );
  XOR U151 ( .A(n210), .B(n211), .Z(n36) );
  AND U152 ( .A(n177), .B(n212), .Z(n211) );
  XOR U153 ( .A(n213), .B(n210), .Z(n212) );
  XNOR U154 ( .A(n37), .B(n206), .Z(n208) );
  IV U155 ( .A(n34), .Z(n37) );
  XNOR U156 ( .A(n214), .B(n215), .Z(n34) );
  AND U157 ( .A(n174), .B(n216), .Z(n215) );
  XOR U158 ( .A(n217), .B(n214), .Z(n216) );
  XOR U159 ( .A(n218), .B(n219), .Z(n206) );
  AND U160 ( .A(n220), .B(n221), .Z(n219) );
  XOR U161 ( .A(n218), .B(n41), .Z(n221) );
  XOR U162 ( .A(n222), .B(n223), .Z(n41) );
  AND U163 ( .A(n177), .B(n224), .Z(n223) );
  XOR U164 ( .A(n225), .B(n222), .Z(n224) );
  XNOR U165 ( .A(n42), .B(n218), .Z(n220) );
  IV U166 ( .A(n39), .Z(n42) );
  XNOR U167 ( .A(n226), .B(n227), .Z(n39) );
  AND U168 ( .A(n174), .B(n228), .Z(n227) );
  XOR U169 ( .A(n229), .B(n226), .Z(n228) );
  XOR U170 ( .A(n230), .B(n231), .Z(n218) );
  AND U171 ( .A(n232), .B(n233), .Z(n231) );
  XOR U172 ( .A(n230), .B(n46), .Z(n233) );
  XOR U173 ( .A(n234), .B(n235), .Z(n46) );
  AND U174 ( .A(n177), .B(n236), .Z(n235) );
  XOR U175 ( .A(n237), .B(n234), .Z(n236) );
  XNOR U176 ( .A(n47), .B(n230), .Z(n232) );
  IV U177 ( .A(n44), .Z(n47) );
  XNOR U178 ( .A(n238), .B(n239), .Z(n44) );
  AND U179 ( .A(n174), .B(n240), .Z(n239) );
  XOR U180 ( .A(n241), .B(n238), .Z(n240) );
  XOR U181 ( .A(n242), .B(n243), .Z(n230) );
  AND U182 ( .A(n244), .B(n245), .Z(n243) );
  XOR U183 ( .A(n242), .B(n51), .Z(n245) );
  XOR U184 ( .A(n246), .B(n247), .Z(n51) );
  AND U185 ( .A(n177), .B(n248), .Z(n247) );
  XOR U186 ( .A(n249), .B(n246), .Z(n248) );
  XNOR U187 ( .A(n52), .B(n242), .Z(n244) );
  IV U188 ( .A(n49), .Z(n52) );
  XNOR U189 ( .A(n250), .B(n251), .Z(n49) );
  AND U190 ( .A(n174), .B(n252), .Z(n251) );
  XOR U191 ( .A(n253), .B(n250), .Z(n252) );
  XOR U192 ( .A(n254), .B(n255), .Z(n242) );
  AND U193 ( .A(n256), .B(n257), .Z(n255) );
  XOR U194 ( .A(n254), .B(n56), .Z(n257) );
  XOR U195 ( .A(n258), .B(n259), .Z(n56) );
  AND U196 ( .A(n177), .B(n260), .Z(n259) );
  XOR U197 ( .A(n261), .B(n258), .Z(n260) );
  XNOR U198 ( .A(n57), .B(n254), .Z(n256) );
  IV U199 ( .A(n54), .Z(n57) );
  XNOR U200 ( .A(n262), .B(n263), .Z(n54) );
  AND U201 ( .A(n174), .B(n264), .Z(n263) );
  XOR U202 ( .A(n265), .B(n262), .Z(n264) );
  XOR U203 ( .A(n266), .B(n267), .Z(n254) );
  AND U204 ( .A(n268), .B(n269), .Z(n267) );
  XOR U205 ( .A(n266), .B(n61), .Z(n269) );
  XOR U206 ( .A(n270), .B(n271), .Z(n61) );
  AND U207 ( .A(n177), .B(n272), .Z(n271) );
  XOR U208 ( .A(n273), .B(n270), .Z(n272) );
  XNOR U209 ( .A(n62), .B(n266), .Z(n268) );
  IV U210 ( .A(n59), .Z(n62) );
  XNOR U211 ( .A(n274), .B(n275), .Z(n59) );
  AND U212 ( .A(n174), .B(n276), .Z(n275) );
  XOR U213 ( .A(n277), .B(n274), .Z(n276) );
  XOR U214 ( .A(n278), .B(n279), .Z(n266) );
  AND U215 ( .A(n280), .B(n281), .Z(n279) );
  XOR U216 ( .A(n278), .B(n66), .Z(n281) );
  XOR U217 ( .A(n282), .B(n283), .Z(n66) );
  AND U218 ( .A(n177), .B(n284), .Z(n283) );
  XOR U219 ( .A(n285), .B(n282), .Z(n284) );
  XNOR U220 ( .A(n67), .B(n278), .Z(n280) );
  IV U221 ( .A(n64), .Z(n67) );
  XNOR U222 ( .A(n286), .B(n287), .Z(n64) );
  AND U223 ( .A(n174), .B(n288), .Z(n287) );
  XOR U224 ( .A(n289), .B(n286), .Z(n288) );
  XOR U225 ( .A(n290), .B(n291), .Z(n278) );
  AND U226 ( .A(n292), .B(n293), .Z(n291) );
  XOR U227 ( .A(n290), .B(n71), .Z(n293) );
  XOR U228 ( .A(n294), .B(n295), .Z(n71) );
  AND U229 ( .A(n177), .B(n296), .Z(n295) );
  XOR U230 ( .A(n297), .B(n294), .Z(n296) );
  XNOR U231 ( .A(n72), .B(n290), .Z(n292) );
  IV U232 ( .A(n69), .Z(n72) );
  XNOR U233 ( .A(n298), .B(n299), .Z(n69) );
  AND U234 ( .A(n174), .B(n300), .Z(n299) );
  XOR U235 ( .A(n301), .B(n298), .Z(n300) );
  XOR U236 ( .A(n302), .B(n303), .Z(n290) );
  AND U237 ( .A(n304), .B(n305), .Z(n303) );
  XOR U238 ( .A(n302), .B(n76), .Z(n305) );
  XOR U239 ( .A(n306), .B(n307), .Z(n76) );
  AND U240 ( .A(n177), .B(n308), .Z(n307) );
  XOR U241 ( .A(n309), .B(n306), .Z(n308) );
  XNOR U242 ( .A(n77), .B(n302), .Z(n304) );
  IV U243 ( .A(n74), .Z(n77) );
  XNOR U244 ( .A(n310), .B(n311), .Z(n74) );
  AND U245 ( .A(n174), .B(n312), .Z(n311) );
  XOR U246 ( .A(n313), .B(n310), .Z(n312) );
  XOR U247 ( .A(n314), .B(n315), .Z(n302) );
  AND U248 ( .A(n316), .B(n317), .Z(n315) );
  XOR U249 ( .A(n4), .B(n314), .Z(n317) );
  XOR U250 ( .A(n318), .B(n319), .Z(n4) );
  AND U251 ( .A(n177), .B(n320), .Z(n319) );
  XOR U252 ( .A(n318), .B(n321), .Z(n320) );
  XNOR U253 ( .A(n314), .B(n2), .Z(n316) );
  XOR U254 ( .A(n322), .B(n323), .Z(n2) );
  AND U255 ( .A(n174), .B(n324), .Z(n323) );
  XOR U256 ( .A(n322), .B(n325), .Z(n324) );
  XOR U257 ( .A(n326), .B(n327), .Z(n314) );
  AND U258 ( .A(n328), .B(n329), .Z(n327) );
  XOR U259 ( .A(n326), .B(n8), .Z(n329) );
  XOR U260 ( .A(n330), .B(n331), .Z(n8) );
  AND U261 ( .A(n177), .B(n332), .Z(n331) );
  XOR U262 ( .A(n333), .B(n330), .Z(n332) );
  XNOR U263 ( .A(n9), .B(n326), .Z(n328) );
  IV U264 ( .A(n6), .Z(n9) );
  XNOR U265 ( .A(n334), .B(n335), .Z(n6) );
  AND U266 ( .A(n174), .B(n336), .Z(n335) );
  XOR U267 ( .A(n337), .B(n334), .Z(n336) );
  XOR U268 ( .A(n338), .B(n339), .Z(n326) );
  AND U269 ( .A(n340), .B(n341), .Z(n339) );
  XOR U270 ( .A(n338), .B(n13), .Z(n341) );
  XOR U271 ( .A(n342), .B(n343), .Z(n13) );
  AND U272 ( .A(n177), .B(n344), .Z(n343) );
  XOR U273 ( .A(n345), .B(n342), .Z(n344) );
  XNOR U274 ( .A(n14), .B(n338), .Z(n340) );
  IV U275 ( .A(n11), .Z(n14) );
  XNOR U276 ( .A(n346), .B(n347), .Z(n11) );
  AND U277 ( .A(n174), .B(n348), .Z(n347) );
  XOR U278 ( .A(n349), .B(n346), .Z(n348) );
  XNOR U279 ( .A(n350), .B(n351), .Z(n338) );
  AND U280 ( .A(n352), .B(n353), .Z(n351) );
  XNOR U281 ( .A(n350), .B(n18), .Z(n353) );
  XOR U282 ( .A(n354), .B(n355), .Z(n18) );
  AND U283 ( .A(n177), .B(n356), .Z(n355) );
  XOR U284 ( .A(n357), .B(n354), .Z(n356) );
  XOR U285 ( .A(n19), .B(n350), .Z(n352) );
  IV U286 ( .A(n16), .Z(n19) );
  XNOR U287 ( .A(n358), .B(n359), .Z(n16) );
  AND U288 ( .A(n174), .B(n360), .Z(n359) );
  XOR U289 ( .A(n361), .B(n358), .Z(n360) );
  AND U290 ( .A(n21), .B(n23), .Z(n350) );
  XNOR U291 ( .A(n362), .B(n363), .Z(n23) );
  AND U292 ( .A(n177), .B(n364), .Z(n363) );
  XNOR U293 ( .A(n365), .B(n362), .Z(n364) );
  XOR U294 ( .A(n366), .B(n367), .Z(n177) );
  AND U295 ( .A(n368), .B(n369), .Z(n367) );
  XOR U296 ( .A(n189), .B(n366), .Z(n369) );
  IV U297 ( .A(n370), .Z(n189) );
  AND U298 ( .A(n371), .B(n372), .Z(n370) );
  XOR U299 ( .A(n366), .B(n186), .Z(n368) );
  AND U300 ( .A(n373), .B(n374), .Z(n186) );
  XOR U301 ( .A(n375), .B(n376), .Z(n366) );
  AND U302 ( .A(n377), .B(n378), .Z(n376) );
  XOR U303 ( .A(n375), .B(n201), .Z(n378) );
  XOR U304 ( .A(n379), .B(n380), .Z(n201) );
  AND U305 ( .A(n161), .B(n381), .Z(n380) );
  XOR U306 ( .A(n382), .B(n379), .Z(n381) );
  XNOR U307 ( .A(n198), .B(n375), .Z(n377) );
  XOR U308 ( .A(n383), .B(n384), .Z(n198) );
  AND U309 ( .A(n159), .B(n385), .Z(n384) );
  XOR U310 ( .A(n386), .B(n383), .Z(n385) );
  XOR U311 ( .A(n387), .B(n388), .Z(n375) );
  AND U312 ( .A(n389), .B(n390), .Z(n388) );
  XOR U313 ( .A(n387), .B(n213), .Z(n390) );
  XOR U314 ( .A(n391), .B(n392), .Z(n213) );
  AND U315 ( .A(n161), .B(n393), .Z(n392) );
  XOR U316 ( .A(n394), .B(n391), .Z(n393) );
  XNOR U317 ( .A(n210), .B(n387), .Z(n389) );
  XOR U318 ( .A(n395), .B(n396), .Z(n210) );
  AND U319 ( .A(n159), .B(n397), .Z(n396) );
  XOR U320 ( .A(n398), .B(n395), .Z(n397) );
  XOR U321 ( .A(n399), .B(n400), .Z(n387) );
  AND U322 ( .A(n401), .B(n402), .Z(n400) );
  XOR U323 ( .A(n399), .B(n225), .Z(n402) );
  XOR U324 ( .A(n403), .B(n404), .Z(n225) );
  AND U325 ( .A(n161), .B(n405), .Z(n404) );
  XOR U326 ( .A(n406), .B(n403), .Z(n405) );
  XNOR U327 ( .A(n222), .B(n399), .Z(n401) );
  XOR U328 ( .A(n407), .B(n408), .Z(n222) );
  AND U329 ( .A(n159), .B(n409), .Z(n408) );
  XOR U330 ( .A(n410), .B(n407), .Z(n409) );
  XOR U331 ( .A(n411), .B(n412), .Z(n399) );
  AND U332 ( .A(n413), .B(n414), .Z(n412) );
  XOR U333 ( .A(n411), .B(n237), .Z(n414) );
  XOR U334 ( .A(n415), .B(n416), .Z(n237) );
  AND U335 ( .A(n161), .B(n417), .Z(n416) );
  XOR U336 ( .A(n418), .B(n415), .Z(n417) );
  XNOR U337 ( .A(n234), .B(n411), .Z(n413) );
  XOR U338 ( .A(n419), .B(n420), .Z(n234) );
  AND U339 ( .A(n159), .B(n421), .Z(n420) );
  XOR U340 ( .A(n422), .B(n419), .Z(n421) );
  XOR U341 ( .A(n423), .B(n424), .Z(n411) );
  AND U342 ( .A(n425), .B(n426), .Z(n424) );
  XOR U343 ( .A(n423), .B(n249), .Z(n426) );
  XOR U344 ( .A(n427), .B(n428), .Z(n249) );
  AND U345 ( .A(n161), .B(n429), .Z(n428) );
  XOR U346 ( .A(n430), .B(n427), .Z(n429) );
  XNOR U347 ( .A(n246), .B(n423), .Z(n425) );
  XOR U348 ( .A(n431), .B(n432), .Z(n246) );
  AND U349 ( .A(n159), .B(n433), .Z(n432) );
  XOR U350 ( .A(n434), .B(n431), .Z(n433) );
  XOR U351 ( .A(n435), .B(n436), .Z(n423) );
  AND U352 ( .A(n437), .B(n438), .Z(n436) );
  XOR U353 ( .A(n435), .B(n261), .Z(n438) );
  XOR U354 ( .A(n439), .B(n440), .Z(n261) );
  AND U355 ( .A(n161), .B(n441), .Z(n440) );
  XOR U356 ( .A(n442), .B(n439), .Z(n441) );
  XNOR U357 ( .A(n258), .B(n435), .Z(n437) );
  XOR U358 ( .A(n443), .B(n444), .Z(n258) );
  AND U359 ( .A(n159), .B(n445), .Z(n444) );
  XOR U360 ( .A(n446), .B(n443), .Z(n445) );
  XOR U361 ( .A(n447), .B(n448), .Z(n435) );
  AND U362 ( .A(n449), .B(n450), .Z(n448) );
  XOR U363 ( .A(n447), .B(n273), .Z(n450) );
  XOR U364 ( .A(n451), .B(n452), .Z(n273) );
  AND U365 ( .A(n161), .B(n453), .Z(n452) );
  XOR U366 ( .A(n454), .B(n451), .Z(n453) );
  XNOR U367 ( .A(n270), .B(n447), .Z(n449) );
  XOR U368 ( .A(n455), .B(n456), .Z(n270) );
  AND U369 ( .A(n159), .B(n457), .Z(n456) );
  XOR U370 ( .A(n458), .B(n455), .Z(n457) );
  XOR U371 ( .A(n459), .B(n460), .Z(n447) );
  AND U372 ( .A(n461), .B(n462), .Z(n460) );
  XOR U373 ( .A(n459), .B(n285), .Z(n462) );
  XOR U374 ( .A(n463), .B(n464), .Z(n285) );
  AND U375 ( .A(n161), .B(n465), .Z(n464) );
  XOR U376 ( .A(n466), .B(n463), .Z(n465) );
  XNOR U377 ( .A(n282), .B(n459), .Z(n461) );
  XOR U378 ( .A(n467), .B(n468), .Z(n282) );
  AND U379 ( .A(n159), .B(n469), .Z(n468) );
  XOR U380 ( .A(n470), .B(n467), .Z(n469) );
  XOR U381 ( .A(n471), .B(n472), .Z(n459) );
  AND U382 ( .A(n473), .B(n474), .Z(n472) );
  XOR U383 ( .A(n471), .B(n297), .Z(n474) );
  XOR U384 ( .A(n475), .B(n476), .Z(n297) );
  AND U385 ( .A(n161), .B(n477), .Z(n476) );
  XOR U386 ( .A(n478), .B(n475), .Z(n477) );
  XNOR U387 ( .A(n294), .B(n471), .Z(n473) );
  XOR U388 ( .A(n479), .B(n480), .Z(n294) );
  AND U389 ( .A(n159), .B(n481), .Z(n480) );
  XOR U390 ( .A(n482), .B(n479), .Z(n481) );
  XOR U391 ( .A(n483), .B(n484), .Z(n471) );
  AND U392 ( .A(n485), .B(n486), .Z(n484) );
  XOR U393 ( .A(n483), .B(n309), .Z(n486) );
  XOR U394 ( .A(n487), .B(n488), .Z(n309) );
  AND U395 ( .A(n161), .B(n489), .Z(n488) );
  XOR U396 ( .A(n490), .B(n487), .Z(n489) );
  XNOR U397 ( .A(n306), .B(n483), .Z(n485) );
  XOR U398 ( .A(n491), .B(n492), .Z(n306) );
  AND U399 ( .A(n159), .B(n493), .Z(n492) );
  XOR U400 ( .A(n494), .B(n491), .Z(n493) );
  XOR U401 ( .A(n495), .B(n496), .Z(n483) );
  AND U402 ( .A(n497), .B(n498), .Z(n496) );
  XOR U403 ( .A(n321), .B(n495), .Z(n498) );
  XOR U404 ( .A(n499), .B(n500), .Z(n321) );
  AND U405 ( .A(n161), .B(n501), .Z(n500) );
  XOR U406 ( .A(n499), .B(n502), .Z(n501) );
  XNOR U407 ( .A(n495), .B(n318), .Z(n497) );
  XOR U408 ( .A(n503), .B(n504), .Z(n318) );
  AND U409 ( .A(n159), .B(n505), .Z(n504) );
  XOR U410 ( .A(n503), .B(n506), .Z(n505) );
  XOR U411 ( .A(n507), .B(n508), .Z(n495) );
  AND U412 ( .A(n509), .B(n510), .Z(n508) );
  XOR U413 ( .A(n507), .B(n333), .Z(n510) );
  XOR U414 ( .A(n511), .B(n512), .Z(n333) );
  AND U415 ( .A(n161), .B(n513), .Z(n512) );
  XOR U416 ( .A(n514), .B(n511), .Z(n513) );
  XNOR U417 ( .A(n330), .B(n507), .Z(n509) );
  XOR U418 ( .A(n515), .B(n516), .Z(n330) );
  AND U419 ( .A(n159), .B(n517), .Z(n516) );
  XOR U420 ( .A(n518), .B(n515), .Z(n517) );
  XOR U421 ( .A(n519), .B(n520), .Z(n507) );
  AND U422 ( .A(n521), .B(n522), .Z(n520) );
  XOR U423 ( .A(n519), .B(n345), .Z(n522) );
  XOR U424 ( .A(n523), .B(n524), .Z(n345) );
  AND U425 ( .A(n161), .B(n525), .Z(n524) );
  XOR U426 ( .A(n526), .B(n523), .Z(n525) );
  XNOR U427 ( .A(n342), .B(n519), .Z(n521) );
  XOR U428 ( .A(n527), .B(n528), .Z(n342) );
  AND U429 ( .A(n159), .B(n529), .Z(n528) );
  XOR U430 ( .A(n530), .B(n527), .Z(n529) );
  XOR U431 ( .A(n531), .B(n532), .Z(n519) );
  AND U432 ( .A(n533), .B(n534), .Z(n532) );
  XNOR U433 ( .A(n535), .B(n357), .Z(n534) );
  XOR U434 ( .A(n536), .B(n537), .Z(n357) );
  AND U435 ( .A(n161), .B(n538), .Z(n537) );
  XOR U436 ( .A(n539), .B(n536), .Z(n538) );
  XNOR U437 ( .A(n354), .B(n531), .Z(n533) );
  XOR U438 ( .A(n540), .B(n541), .Z(n354) );
  AND U439 ( .A(n159), .B(n542), .Z(n541) );
  XOR U440 ( .A(n543), .B(n540), .Z(n542) );
  IV U441 ( .A(n535), .Z(n531) );
  AND U442 ( .A(n362), .B(n365), .Z(n535) );
  XNOR U443 ( .A(n544), .B(n545), .Z(n365) );
  AND U444 ( .A(n161), .B(n546), .Z(n545) );
  XNOR U445 ( .A(n547), .B(n544), .Z(n546) );
  XOR U446 ( .A(n548), .B(n549), .Z(n161) );
  AND U447 ( .A(n550), .B(n551), .Z(n549) );
  XNOR U448 ( .A(n371), .B(n548), .Z(n551) );
  AND U449 ( .A(n552), .B(n553), .Z(n371) );
  XOR U450 ( .A(n548), .B(n372), .Z(n550) );
  AND U451 ( .A(n554), .B(n555), .Z(n372) );
  XOR U452 ( .A(n556), .B(n557), .Z(n548) );
  AND U453 ( .A(n558), .B(n559), .Z(n557) );
  XOR U454 ( .A(n556), .B(n382), .Z(n559) );
  XOR U455 ( .A(n560), .B(n561), .Z(n382) );
  AND U456 ( .A(n121), .B(n562), .Z(n561) );
  XOR U457 ( .A(n563), .B(n560), .Z(n562) );
  XNOR U458 ( .A(n379), .B(n556), .Z(n558) );
  XOR U459 ( .A(n564), .B(n565), .Z(n379) );
  AND U460 ( .A(n119), .B(n566), .Z(n565) );
  XOR U461 ( .A(n567), .B(n564), .Z(n566) );
  XOR U462 ( .A(n568), .B(n569), .Z(n556) );
  AND U463 ( .A(n570), .B(n571), .Z(n569) );
  XOR U464 ( .A(n568), .B(n394), .Z(n571) );
  XOR U465 ( .A(n572), .B(n573), .Z(n394) );
  AND U466 ( .A(n121), .B(n574), .Z(n573) );
  XOR U467 ( .A(n575), .B(n572), .Z(n574) );
  XNOR U468 ( .A(n391), .B(n568), .Z(n570) );
  XOR U469 ( .A(n576), .B(n577), .Z(n391) );
  AND U470 ( .A(n119), .B(n578), .Z(n577) );
  XOR U471 ( .A(n579), .B(n576), .Z(n578) );
  XOR U472 ( .A(n580), .B(n581), .Z(n568) );
  AND U473 ( .A(n582), .B(n583), .Z(n581) );
  XOR U474 ( .A(n580), .B(n406), .Z(n583) );
  XOR U475 ( .A(n584), .B(n585), .Z(n406) );
  AND U476 ( .A(n121), .B(n586), .Z(n585) );
  XOR U477 ( .A(n587), .B(n584), .Z(n586) );
  XNOR U478 ( .A(n403), .B(n580), .Z(n582) );
  XOR U479 ( .A(n588), .B(n589), .Z(n403) );
  AND U480 ( .A(n119), .B(n590), .Z(n589) );
  XOR U481 ( .A(n591), .B(n588), .Z(n590) );
  XOR U482 ( .A(n592), .B(n593), .Z(n580) );
  AND U483 ( .A(n594), .B(n595), .Z(n593) );
  XOR U484 ( .A(n592), .B(n418), .Z(n595) );
  XOR U485 ( .A(n596), .B(n597), .Z(n418) );
  AND U486 ( .A(n121), .B(n598), .Z(n597) );
  XOR U487 ( .A(n599), .B(n596), .Z(n598) );
  XNOR U488 ( .A(n415), .B(n592), .Z(n594) );
  XOR U489 ( .A(n600), .B(n601), .Z(n415) );
  AND U490 ( .A(n119), .B(n602), .Z(n601) );
  XOR U491 ( .A(n603), .B(n600), .Z(n602) );
  XOR U492 ( .A(n604), .B(n605), .Z(n592) );
  AND U493 ( .A(n606), .B(n607), .Z(n605) );
  XOR U494 ( .A(n604), .B(n430), .Z(n607) );
  XOR U495 ( .A(n608), .B(n609), .Z(n430) );
  AND U496 ( .A(n121), .B(n610), .Z(n609) );
  XOR U497 ( .A(n611), .B(n608), .Z(n610) );
  XNOR U498 ( .A(n427), .B(n604), .Z(n606) );
  XOR U499 ( .A(n612), .B(n613), .Z(n427) );
  AND U500 ( .A(n119), .B(n614), .Z(n613) );
  XOR U501 ( .A(n615), .B(n612), .Z(n614) );
  XOR U502 ( .A(n616), .B(n617), .Z(n604) );
  AND U503 ( .A(n618), .B(n619), .Z(n617) );
  XOR U504 ( .A(n616), .B(n442), .Z(n619) );
  XOR U505 ( .A(n620), .B(n621), .Z(n442) );
  AND U506 ( .A(n121), .B(n622), .Z(n621) );
  XOR U507 ( .A(n623), .B(n620), .Z(n622) );
  XNOR U508 ( .A(n439), .B(n616), .Z(n618) );
  XOR U509 ( .A(n624), .B(n625), .Z(n439) );
  AND U510 ( .A(n119), .B(n626), .Z(n625) );
  XOR U511 ( .A(n627), .B(n624), .Z(n626) );
  XOR U512 ( .A(n628), .B(n629), .Z(n616) );
  AND U513 ( .A(n630), .B(n631), .Z(n629) );
  XOR U514 ( .A(n628), .B(n454), .Z(n631) );
  XOR U515 ( .A(n632), .B(n633), .Z(n454) );
  AND U516 ( .A(n121), .B(n634), .Z(n633) );
  XOR U517 ( .A(n635), .B(n632), .Z(n634) );
  XNOR U518 ( .A(n451), .B(n628), .Z(n630) );
  XOR U519 ( .A(n636), .B(n637), .Z(n451) );
  AND U520 ( .A(n119), .B(n638), .Z(n637) );
  XOR U521 ( .A(n639), .B(n636), .Z(n638) );
  XOR U522 ( .A(n640), .B(n641), .Z(n628) );
  AND U523 ( .A(n642), .B(n643), .Z(n641) );
  XOR U524 ( .A(n640), .B(n466), .Z(n643) );
  XOR U525 ( .A(n644), .B(n645), .Z(n466) );
  AND U526 ( .A(n121), .B(n646), .Z(n645) );
  XOR U527 ( .A(n647), .B(n644), .Z(n646) );
  XNOR U528 ( .A(n463), .B(n640), .Z(n642) );
  XOR U529 ( .A(n648), .B(n649), .Z(n463) );
  AND U530 ( .A(n119), .B(n650), .Z(n649) );
  XOR U531 ( .A(n651), .B(n648), .Z(n650) );
  XOR U532 ( .A(n652), .B(n653), .Z(n640) );
  AND U533 ( .A(n654), .B(n655), .Z(n653) );
  XOR U534 ( .A(n652), .B(n478), .Z(n655) );
  XOR U535 ( .A(n656), .B(n657), .Z(n478) );
  AND U536 ( .A(n121), .B(n658), .Z(n657) );
  XOR U537 ( .A(n659), .B(n656), .Z(n658) );
  XNOR U538 ( .A(n475), .B(n652), .Z(n654) );
  XOR U539 ( .A(n660), .B(n661), .Z(n475) );
  AND U540 ( .A(n119), .B(n662), .Z(n661) );
  XOR U541 ( .A(n663), .B(n660), .Z(n662) );
  XOR U542 ( .A(n664), .B(n665), .Z(n652) );
  AND U543 ( .A(n666), .B(n667), .Z(n665) );
  XOR U544 ( .A(n664), .B(n490), .Z(n667) );
  XOR U545 ( .A(n668), .B(n669), .Z(n490) );
  AND U546 ( .A(n121), .B(n670), .Z(n669) );
  XOR U547 ( .A(n671), .B(n668), .Z(n670) );
  XNOR U548 ( .A(n487), .B(n664), .Z(n666) );
  XOR U549 ( .A(n672), .B(n673), .Z(n487) );
  AND U550 ( .A(n119), .B(n674), .Z(n673) );
  XOR U551 ( .A(n675), .B(n672), .Z(n674) );
  XOR U552 ( .A(n676), .B(n677), .Z(n664) );
  AND U553 ( .A(n678), .B(n679), .Z(n677) );
  XOR U554 ( .A(n502), .B(n676), .Z(n679) );
  XOR U555 ( .A(n680), .B(n681), .Z(n502) );
  AND U556 ( .A(n121), .B(n682), .Z(n681) );
  XOR U557 ( .A(n680), .B(n683), .Z(n682) );
  XNOR U558 ( .A(n676), .B(n499), .Z(n678) );
  XOR U559 ( .A(n684), .B(n685), .Z(n499) );
  AND U560 ( .A(n119), .B(n686), .Z(n685) );
  XOR U561 ( .A(n684), .B(n687), .Z(n686) );
  XOR U562 ( .A(n688), .B(n689), .Z(n676) );
  AND U563 ( .A(n690), .B(n691), .Z(n689) );
  XOR U564 ( .A(n688), .B(n514), .Z(n691) );
  XOR U565 ( .A(n692), .B(n693), .Z(n514) );
  AND U566 ( .A(n121), .B(n694), .Z(n693) );
  XOR U567 ( .A(n695), .B(n692), .Z(n694) );
  XNOR U568 ( .A(n511), .B(n688), .Z(n690) );
  XOR U569 ( .A(n696), .B(n697), .Z(n511) );
  AND U570 ( .A(n119), .B(n698), .Z(n697) );
  XOR U571 ( .A(n699), .B(n696), .Z(n698) );
  XOR U572 ( .A(n700), .B(n701), .Z(n688) );
  AND U573 ( .A(n702), .B(n703), .Z(n701) );
  XOR U574 ( .A(n700), .B(n526), .Z(n703) );
  XOR U575 ( .A(n704), .B(n705), .Z(n526) );
  AND U576 ( .A(n121), .B(n706), .Z(n705) );
  XOR U577 ( .A(n707), .B(n704), .Z(n706) );
  XNOR U578 ( .A(n523), .B(n700), .Z(n702) );
  XOR U579 ( .A(n708), .B(n709), .Z(n523) );
  AND U580 ( .A(n119), .B(n710), .Z(n709) );
  XOR U581 ( .A(n711), .B(n708), .Z(n710) );
  XOR U582 ( .A(n712), .B(n713), .Z(n700) );
  AND U583 ( .A(n714), .B(n715), .Z(n713) );
  XNOR U584 ( .A(n716), .B(n539), .Z(n715) );
  XOR U585 ( .A(n717), .B(n718), .Z(n539) );
  AND U586 ( .A(n121), .B(n719), .Z(n718) );
  XOR U587 ( .A(n720), .B(n717), .Z(n719) );
  XNOR U588 ( .A(n536), .B(n712), .Z(n714) );
  XOR U589 ( .A(n721), .B(n722), .Z(n536) );
  AND U590 ( .A(n119), .B(n723), .Z(n722) );
  XOR U591 ( .A(n724), .B(n721), .Z(n723) );
  IV U592 ( .A(n716), .Z(n712) );
  AND U593 ( .A(n544), .B(n547), .Z(n716) );
  XNOR U594 ( .A(n725), .B(n726), .Z(n547) );
  AND U595 ( .A(n121), .B(n727), .Z(n726) );
  XNOR U596 ( .A(n728), .B(n725), .Z(n727) );
  XOR U597 ( .A(n729), .B(n730), .Z(n121) );
  AND U598 ( .A(n731), .B(n732), .Z(n730) );
  XNOR U599 ( .A(n552), .B(n729), .Z(n732) );
  AND U600 ( .A(p_input[511]), .B(p_input[495]), .Z(n552) );
  XOR U601 ( .A(n729), .B(n553), .Z(n731) );
  AND U602 ( .A(p_input[479]), .B(p_input[463]), .Z(n553) );
  XOR U603 ( .A(n733), .B(n734), .Z(n729) );
  AND U604 ( .A(n735), .B(n736), .Z(n734) );
  XOR U605 ( .A(n733), .B(n563), .Z(n736) );
  XNOR U606 ( .A(p_input[494]), .B(n737), .Z(n563) );
  AND U607 ( .A(n93), .B(n738), .Z(n737) );
  XOR U608 ( .A(p_input[510]), .B(p_input[494]), .Z(n738) );
  XNOR U609 ( .A(n560), .B(n733), .Z(n735) );
  XOR U610 ( .A(n739), .B(n740), .Z(n560) );
  AND U611 ( .A(n91), .B(n741), .Z(n740) );
  XOR U612 ( .A(p_input[478]), .B(p_input[462]), .Z(n741) );
  XOR U613 ( .A(n742), .B(n743), .Z(n733) );
  AND U614 ( .A(n744), .B(n745), .Z(n743) );
  XOR U615 ( .A(n742), .B(n575), .Z(n745) );
  XNOR U616 ( .A(p_input[493]), .B(n746), .Z(n575) );
  AND U617 ( .A(n93), .B(n747), .Z(n746) );
  XOR U618 ( .A(p_input[509]), .B(p_input[493]), .Z(n747) );
  XNOR U619 ( .A(n572), .B(n742), .Z(n744) );
  XOR U620 ( .A(n748), .B(n749), .Z(n572) );
  AND U621 ( .A(n91), .B(n750), .Z(n749) );
  XOR U622 ( .A(p_input[477]), .B(p_input[461]), .Z(n750) );
  XOR U623 ( .A(n751), .B(n752), .Z(n742) );
  AND U624 ( .A(n753), .B(n754), .Z(n752) );
  XOR U625 ( .A(n751), .B(n587), .Z(n754) );
  XNOR U626 ( .A(p_input[492]), .B(n755), .Z(n587) );
  AND U627 ( .A(n93), .B(n756), .Z(n755) );
  XOR U628 ( .A(p_input[508]), .B(p_input[492]), .Z(n756) );
  XNOR U629 ( .A(n584), .B(n751), .Z(n753) );
  XOR U630 ( .A(n757), .B(n758), .Z(n584) );
  AND U631 ( .A(n91), .B(n759), .Z(n758) );
  XOR U632 ( .A(p_input[476]), .B(p_input[460]), .Z(n759) );
  XOR U633 ( .A(n760), .B(n761), .Z(n751) );
  AND U634 ( .A(n762), .B(n763), .Z(n761) );
  XOR U635 ( .A(n760), .B(n599), .Z(n763) );
  XNOR U636 ( .A(p_input[491]), .B(n764), .Z(n599) );
  AND U637 ( .A(n93), .B(n765), .Z(n764) );
  XOR U638 ( .A(p_input[507]), .B(p_input[491]), .Z(n765) );
  XNOR U639 ( .A(n596), .B(n760), .Z(n762) );
  XOR U640 ( .A(n766), .B(n767), .Z(n596) );
  AND U641 ( .A(n91), .B(n768), .Z(n767) );
  XOR U642 ( .A(p_input[475]), .B(p_input[459]), .Z(n768) );
  XOR U643 ( .A(n769), .B(n770), .Z(n760) );
  AND U644 ( .A(n771), .B(n772), .Z(n770) );
  XOR U645 ( .A(n769), .B(n611), .Z(n772) );
  XNOR U646 ( .A(p_input[490]), .B(n773), .Z(n611) );
  AND U647 ( .A(n93), .B(n774), .Z(n773) );
  XOR U648 ( .A(p_input[506]), .B(p_input[490]), .Z(n774) );
  XNOR U649 ( .A(n608), .B(n769), .Z(n771) );
  XOR U650 ( .A(n775), .B(n776), .Z(n608) );
  AND U651 ( .A(n91), .B(n777), .Z(n776) );
  XOR U652 ( .A(p_input[474]), .B(p_input[458]), .Z(n777) );
  XOR U653 ( .A(n778), .B(n779), .Z(n769) );
  AND U654 ( .A(n780), .B(n781), .Z(n779) );
  XOR U655 ( .A(n778), .B(n623), .Z(n781) );
  XNOR U656 ( .A(p_input[489]), .B(n782), .Z(n623) );
  AND U657 ( .A(n93), .B(n783), .Z(n782) );
  XOR U658 ( .A(p_input[505]), .B(p_input[489]), .Z(n783) );
  XNOR U659 ( .A(n620), .B(n778), .Z(n780) );
  XOR U660 ( .A(n784), .B(n785), .Z(n620) );
  AND U661 ( .A(n91), .B(n786), .Z(n785) );
  XOR U662 ( .A(p_input[473]), .B(p_input[457]), .Z(n786) );
  XOR U663 ( .A(n787), .B(n788), .Z(n778) );
  AND U664 ( .A(n789), .B(n790), .Z(n788) );
  XOR U665 ( .A(n787), .B(n635), .Z(n790) );
  XNOR U666 ( .A(p_input[488]), .B(n791), .Z(n635) );
  AND U667 ( .A(n93), .B(n792), .Z(n791) );
  XOR U668 ( .A(p_input[504]), .B(p_input[488]), .Z(n792) );
  XNOR U669 ( .A(n632), .B(n787), .Z(n789) );
  XOR U670 ( .A(n793), .B(n794), .Z(n632) );
  AND U671 ( .A(n91), .B(n795), .Z(n794) );
  XOR U672 ( .A(p_input[472]), .B(p_input[456]), .Z(n795) );
  XOR U673 ( .A(n796), .B(n797), .Z(n787) );
  AND U674 ( .A(n798), .B(n799), .Z(n797) );
  XOR U675 ( .A(n796), .B(n647), .Z(n799) );
  XNOR U676 ( .A(p_input[487]), .B(n800), .Z(n647) );
  AND U677 ( .A(n93), .B(n801), .Z(n800) );
  XOR U678 ( .A(p_input[503]), .B(p_input[487]), .Z(n801) );
  XNOR U679 ( .A(n644), .B(n796), .Z(n798) );
  XOR U680 ( .A(n802), .B(n803), .Z(n644) );
  AND U681 ( .A(n91), .B(n804), .Z(n803) );
  XOR U682 ( .A(p_input[471]), .B(p_input[455]), .Z(n804) );
  XOR U683 ( .A(n805), .B(n806), .Z(n796) );
  AND U684 ( .A(n807), .B(n808), .Z(n806) );
  XOR U685 ( .A(n805), .B(n659), .Z(n808) );
  XNOR U686 ( .A(p_input[486]), .B(n809), .Z(n659) );
  AND U687 ( .A(n93), .B(n810), .Z(n809) );
  XOR U688 ( .A(p_input[502]), .B(p_input[486]), .Z(n810) );
  XNOR U689 ( .A(n656), .B(n805), .Z(n807) );
  XOR U690 ( .A(n811), .B(n812), .Z(n656) );
  AND U691 ( .A(n91), .B(n813), .Z(n812) );
  XOR U692 ( .A(p_input[470]), .B(p_input[454]), .Z(n813) );
  XOR U693 ( .A(n814), .B(n815), .Z(n805) );
  AND U694 ( .A(n816), .B(n817), .Z(n815) );
  XOR U695 ( .A(n814), .B(n671), .Z(n817) );
  XNOR U696 ( .A(p_input[485]), .B(n818), .Z(n671) );
  AND U697 ( .A(n93), .B(n819), .Z(n818) );
  XOR U698 ( .A(p_input[501]), .B(p_input[485]), .Z(n819) );
  XNOR U699 ( .A(n668), .B(n814), .Z(n816) );
  XOR U700 ( .A(n820), .B(n821), .Z(n668) );
  AND U701 ( .A(n91), .B(n822), .Z(n821) );
  XOR U702 ( .A(p_input[469]), .B(p_input[453]), .Z(n822) );
  XOR U703 ( .A(n823), .B(n824), .Z(n814) );
  AND U704 ( .A(n825), .B(n826), .Z(n824) );
  XOR U705 ( .A(n683), .B(n823), .Z(n826) );
  XNOR U706 ( .A(p_input[484]), .B(n827), .Z(n683) );
  AND U707 ( .A(n93), .B(n828), .Z(n827) );
  XOR U708 ( .A(p_input[500]), .B(p_input[484]), .Z(n828) );
  XNOR U709 ( .A(n823), .B(n680), .Z(n825) );
  XOR U710 ( .A(n829), .B(n830), .Z(n680) );
  AND U711 ( .A(n91), .B(n831), .Z(n830) );
  XOR U712 ( .A(p_input[468]), .B(p_input[452]), .Z(n831) );
  XOR U713 ( .A(n832), .B(n833), .Z(n823) );
  AND U714 ( .A(n834), .B(n835), .Z(n833) );
  XOR U715 ( .A(n832), .B(n695), .Z(n835) );
  XNOR U716 ( .A(p_input[483]), .B(n836), .Z(n695) );
  AND U717 ( .A(n93), .B(n837), .Z(n836) );
  XOR U718 ( .A(p_input[499]), .B(p_input[483]), .Z(n837) );
  XNOR U719 ( .A(n692), .B(n832), .Z(n834) );
  XOR U720 ( .A(n838), .B(n839), .Z(n692) );
  AND U721 ( .A(n91), .B(n840), .Z(n839) );
  XOR U722 ( .A(p_input[467]), .B(p_input[451]), .Z(n840) );
  XOR U723 ( .A(n841), .B(n842), .Z(n832) );
  AND U724 ( .A(n843), .B(n844), .Z(n842) );
  XOR U725 ( .A(n841), .B(n707), .Z(n844) );
  XNOR U726 ( .A(p_input[482]), .B(n845), .Z(n707) );
  AND U727 ( .A(n93), .B(n846), .Z(n845) );
  XOR U728 ( .A(p_input[498]), .B(p_input[482]), .Z(n846) );
  XNOR U729 ( .A(n704), .B(n841), .Z(n843) );
  XOR U730 ( .A(n847), .B(n848), .Z(n704) );
  AND U731 ( .A(n91), .B(n849), .Z(n848) );
  XOR U732 ( .A(p_input[466]), .B(p_input[450]), .Z(n849) );
  XOR U733 ( .A(n850), .B(n851), .Z(n841) );
  AND U734 ( .A(n852), .B(n853), .Z(n851) );
  XNOR U735 ( .A(n854), .B(n720), .Z(n853) );
  XNOR U736 ( .A(p_input[481]), .B(n855), .Z(n720) );
  AND U737 ( .A(n93), .B(n856), .Z(n855) );
  XNOR U738 ( .A(p_input[497]), .B(n857), .Z(n856) );
  IV U739 ( .A(p_input[481]), .Z(n857) );
  XNOR U740 ( .A(n717), .B(n850), .Z(n852) );
  XNOR U741 ( .A(p_input[449]), .B(n858), .Z(n717) );
  AND U742 ( .A(n91), .B(n859), .Z(n858) );
  XOR U743 ( .A(p_input[465]), .B(p_input[449]), .Z(n859) );
  IV U744 ( .A(n854), .Z(n850) );
  AND U745 ( .A(n725), .B(n728), .Z(n854) );
  XOR U746 ( .A(p_input[480]), .B(n860), .Z(n728) );
  AND U747 ( .A(n93), .B(n861), .Z(n860) );
  XOR U748 ( .A(p_input[496]), .B(p_input[480]), .Z(n861) );
  XOR U749 ( .A(n862), .B(n863), .Z(n93) );
  AND U750 ( .A(n864), .B(n865), .Z(n863) );
  XNOR U751 ( .A(p_input[511]), .B(n862), .Z(n865) );
  XOR U752 ( .A(n862), .B(p_input[495]), .Z(n864) );
  XOR U753 ( .A(n866), .B(n867), .Z(n862) );
  AND U754 ( .A(n868), .B(n869), .Z(n867) );
  XNOR U755 ( .A(p_input[510]), .B(n866), .Z(n869) );
  XOR U756 ( .A(n866), .B(p_input[494]), .Z(n868) );
  XOR U757 ( .A(n870), .B(n871), .Z(n866) );
  AND U758 ( .A(n872), .B(n873), .Z(n871) );
  XNOR U759 ( .A(p_input[509]), .B(n870), .Z(n873) );
  XOR U760 ( .A(n870), .B(p_input[493]), .Z(n872) );
  XOR U761 ( .A(n874), .B(n875), .Z(n870) );
  AND U762 ( .A(n876), .B(n877), .Z(n875) );
  XNOR U763 ( .A(p_input[508]), .B(n874), .Z(n877) );
  XOR U764 ( .A(n874), .B(p_input[492]), .Z(n876) );
  XOR U765 ( .A(n878), .B(n879), .Z(n874) );
  AND U766 ( .A(n880), .B(n881), .Z(n879) );
  XNOR U767 ( .A(p_input[507]), .B(n878), .Z(n881) );
  XOR U768 ( .A(n878), .B(p_input[491]), .Z(n880) );
  XOR U769 ( .A(n882), .B(n883), .Z(n878) );
  AND U770 ( .A(n884), .B(n885), .Z(n883) );
  XNOR U771 ( .A(p_input[506]), .B(n882), .Z(n885) );
  XOR U772 ( .A(n882), .B(p_input[490]), .Z(n884) );
  XOR U773 ( .A(n886), .B(n887), .Z(n882) );
  AND U774 ( .A(n888), .B(n889), .Z(n887) );
  XNOR U775 ( .A(p_input[505]), .B(n886), .Z(n889) );
  XOR U776 ( .A(n886), .B(p_input[489]), .Z(n888) );
  XOR U777 ( .A(n890), .B(n891), .Z(n886) );
  AND U778 ( .A(n892), .B(n893), .Z(n891) );
  XNOR U779 ( .A(p_input[504]), .B(n890), .Z(n893) );
  XOR U780 ( .A(n890), .B(p_input[488]), .Z(n892) );
  XOR U781 ( .A(n894), .B(n895), .Z(n890) );
  AND U782 ( .A(n896), .B(n897), .Z(n895) );
  XNOR U783 ( .A(p_input[503]), .B(n894), .Z(n897) );
  XOR U784 ( .A(n894), .B(p_input[487]), .Z(n896) );
  XOR U785 ( .A(n898), .B(n899), .Z(n894) );
  AND U786 ( .A(n900), .B(n901), .Z(n899) );
  XNOR U787 ( .A(p_input[502]), .B(n898), .Z(n901) );
  XOR U788 ( .A(n898), .B(p_input[486]), .Z(n900) );
  XOR U789 ( .A(n902), .B(n903), .Z(n898) );
  AND U790 ( .A(n904), .B(n905), .Z(n903) );
  XNOR U791 ( .A(p_input[501]), .B(n902), .Z(n905) );
  XOR U792 ( .A(n902), .B(p_input[485]), .Z(n904) );
  XOR U793 ( .A(n906), .B(n907), .Z(n902) );
  AND U794 ( .A(n908), .B(n909), .Z(n907) );
  XNOR U795 ( .A(p_input[500]), .B(n906), .Z(n909) );
  XOR U796 ( .A(n906), .B(p_input[484]), .Z(n908) );
  XOR U797 ( .A(n910), .B(n911), .Z(n906) );
  AND U798 ( .A(n912), .B(n913), .Z(n911) );
  XNOR U799 ( .A(p_input[499]), .B(n910), .Z(n913) );
  XOR U800 ( .A(n910), .B(p_input[483]), .Z(n912) );
  XOR U801 ( .A(n914), .B(n915), .Z(n910) );
  AND U802 ( .A(n916), .B(n917), .Z(n915) );
  XNOR U803 ( .A(p_input[498]), .B(n914), .Z(n917) );
  XOR U804 ( .A(n914), .B(p_input[482]), .Z(n916) );
  XNOR U805 ( .A(n918), .B(n919), .Z(n914) );
  AND U806 ( .A(n920), .B(n921), .Z(n919) );
  XOR U807 ( .A(p_input[497]), .B(n918), .Z(n921) );
  XNOR U808 ( .A(p_input[481]), .B(n918), .Z(n920) );
  AND U809 ( .A(p_input[496]), .B(n922), .Z(n918) );
  IV U810 ( .A(p_input[480]), .Z(n922) );
  XNOR U811 ( .A(p_input[448]), .B(n923), .Z(n725) );
  AND U812 ( .A(n91), .B(n924), .Z(n923) );
  XOR U813 ( .A(p_input[464]), .B(p_input[448]), .Z(n924) );
  XOR U814 ( .A(n925), .B(n926), .Z(n91) );
  AND U815 ( .A(n927), .B(n928), .Z(n926) );
  XNOR U816 ( .A(p_input[479]), .B(n925), .Z(n928) );
  XOR U817 ( .A(n925), .B(p_input[463]), .Z(n927) );
  XOR U818 ( .A(n929), .B(n930), .Z(n925) );
  AND U819 ( .A(n931), .B(n932), .Z(n930) );
  XNOR U820 ( .A(p_input[478]), .B(n929), .Z(n932) );
  XNOR U821 ( .A(n929), .B(n739), .Z(n931) );
  IV U822 ( .A(p_input[462]), .Z(n739) );
  XOR U823 ( .A(n933), .B(n934), .Z(n929) );
  AND U824 ( .A(n935), .B(n936), .Z(n934) );
  XNOR U825 ( .A(p_input[477]), .B(n933), .Z(n936) );
  XNOR U826 ( .A(n933), .B(n748), .Z(n935) );
  IV U827 ( .A(p_input[461]), .Z(n748) );
  XOR U828 ( .A(n937), .B(n938), .Z(n933) );
  AND U829 ( .A(n939), .B(n940), .Z(n938) );
  XNOR U830 ( .A(p_input[476]), .B(n937), .Z(n940) );
  XNOR U831 ( .A(n937), .B(n757), .Z(n939) );
  IV U832 ( .A(p_input[460]), .Z(n757) );
  XOR U833 ( .A(n941), .B(n942), .Z(n937) );
  AND U834 ( .A(n943), .B(n944), .Z(n942) );
  XNOR U835 ( .A(p_input[475]), .B(n941), .Z(n944) );
  XNOR U836 ( .A(n941), .B(n766), .Z(n943) );
  IV U837 ( .A(p_input[459]), .Z(n766) );
  XOR U838 ( .A(n945), .B(n946), .Z(n941) );
  AND U839 ( .A(n947), .B(n948), .Z(n946) );
  XNOR U840 ( .A(p_input[474]), .B(n945), .Z(n948) );
  XNOR U841 ( .A(n945), .B(n775), .Z(n947) );
  IV U842 ( .A(p_input[458]), .Z(n775) );
  XOR U843 ( .A(n949), .B(n950), .Z(n945) );
  AND U844 ( .A(n951), .B(n952), .Z(n950) );
  XNOR U845 ( .A(p_input[473]), .B(n949), .Z(n952) );
  XNOR U846 ( .A(n949), .B(n784), .Z(n951) );
  IV U847 ( .A(p_input[457]), .Z(n784) );
  XOR U848 ( .A(n953), .B(n954), .Z(n949) );
  AND U849 ( .A(n955), .B(n956), .Z(n954) );
  XNOR U850 ( .A(p_input[472]), .B(n953), .Z(n956) );
  XNOR U851 ( .A(n953), .B(n793), .Z(n955) );
  IV U852 ( .A(p_input[456]), .Z(n793) );
  XOR U853 ( .A(n957), .B(n958), .Z(n953) );
  AND U854 ( .A(n959), .B(n960), .Z(n958) );
  XNOR U855 ( .A(p_input[471]), .B(n957), .Z(n960) );
  XNOR U856 ( .A(n957), .B(n802), .Z(n959) );
  IV U857 ( .A(p_input[455]), .Z(n802) );
  XOR U858 ( .A(n961), .B(n962), .Z(n957) );
  AND U859 ( .A(n963), .B(n964), .Z(n962) );
  XNOR U860 ( .A(p_input[470]), .B(n961), .Z(n964) );
  XNOR U861 ( .A(n961), .B(n811), .Z(n963) );
  IV U862 ( .A(p_input[454]), .Z(n811) );
  XOR U863 ( .A(n965), .B(n966), .Z(n961) );
  AND U864 ( .A(n967), .B(n968), .Z(n966) );
  XNOR U865 ( .A(p_input[469]), .B(n965), .Z(n968) );
  XNOR U866 ( .A(n965), .B(n820), .Z(n967) );
  IV U867 ( .A(p_input[453]), .Z(n820) );
  XOR U868 ( .A(n969), .B(n970), .Z(n965) );
  AND U869 ( .A(n971), .B(n972), .Z(n970) );
  XNOR U870 ( .A(p_input[468]), .B(n969), .Z(n972) );
  XNOR U871 ( .A(n969), .B(n829), .Z(n971) );
  IV U872 ( .A(p_input[452]), .Z(n829) );
  XOR U873 ( .A(n973), .B(n974), .Z(n969) );
  AND U874 ( .A(n975), .B(n976), .Z(n974) );
  XNOR U875 ( .A(p_input[467]), .B(n973), .Z(n976) );
  XNOR U876 ( .A(n973), .B(n838), .Z(n975) );
  IV U877 ( .A(p_input[451]), .Z(n838) );
  XOR U878 ( .A(n977), .B(n978), .Z(n973) );
  AND U879 ( .A(n979), .B(n980), .Z(n978) );
  XNOR U880 ( .A(p_input[466]), .B(n977), .Z(n980) );
  XNOR U881 ( .A(n977), .B(n847), .Z(n979) );
  IV U882 ( .A(p_input[450]), .Z(n847) );
  XNOR U883 ( .A(n981), .B(n982), .Z(n977) );
  AND U884 ( .A(n983), .B(n984), .Z(n982) );
  XOR U885 ( .A(p_input[465]), .B(n981), .Z(n984) );
  XNOR U886 ( .A(p_input[449]), .B(n981), .Z(n983) );
  AND U887 ( .A(p_input[464]), .B(n985), .Z(n981) );
  IV U888 ( .A(p_input[448]), .Z(n985) );
  XOR U889 ( .A(n986), .B(n987), .Z(n544) );
  AND U890 ( .A(n119), .B(n988), .Z(n987) );
  XNOR U891 ( .A(n989), .B(n986), .Z(n988) );
  XOR U892 ( .A(n990), .B(n991), .Z(n119) );
  AND U893 ( .A(n992), .B(n993), .Z(n991) );
  XNOR U894 ( .A(n554), .B(n990), .Z(n993) );
  AND U895 ( .A(p_input[447]), .B(p_input[431]), .Z(n554) );
  XOR U896 ( .A(n990), .B(n555), .Z(n992) );
  AND U897 ( .A(p_input[415]), .B(p_input[399]), .Z(n555) );
  XOR U898 ( .A(n994), .B(n995), .Z(n990) );
  AND U899 ( .A(n996), .B(n997), .Z(n995) );
  XOR U900 ( .A(n994), .B(n567), .Z(n997) );
  XNOR U901 ( .A(p_input[430]), .B(n998), .Z(n567) );
  AND U902 ( .A(n97), .B(n999), .Z(n998) );
  XOR U903 ( .A(p_input[446]), .B(p_input[430]), .Z(n999) );
  XNOR U904 ( .A(n564), .B(n994), .Z(n996) );
  XOR U905 ( .A(n1000), .B(n1001), .Z(n564) );
  AND U906 ( .A(n94), .B(n1002), .Z(n1001) );
  XOR U907 ( .A(p_input[414]), .B(p_input[398]), .Z(n1002) );
  XOR U908 ( .A(n1003), .B(n1004), .Z(n994) );
  AND U909 ( .A(n1005), .B(n1006), .Z(n1004) );
  XOR U910 ( .A(n1003), .B(n579), .Z(n1006) );
  XNOR U911 ( .A(p_input[429]), .B(n1007), .Z(n579) );
  AND U912 ( .A(n97), .B(n1008), .Z(n1007) );
  XOR U913 ( .A(p_input[445]), .B(p_input[429]), .Z(n1008) );
  XNOR U914 ( .A(n576), .B(n1003), .Z(n1005) );
  XOR U915 ( .A(n1009), .B(n1010), .Z(n576) );
  AND U916 ( .A(n94), .B(n1011), .Z(n1010) );
  XOR U917 ( .A(p_input[413]), .B(p_input[397]), .Z(n1011) );
  XOR U918 ( .A(n1012), .B(n1013), .Z(n1003) );
  AND U919 ( .A(n1014), .B(n1015), .Z(n1013) );
  XOR U920 ( .A(n1012), .B(n591), .Z(n1015) );
  XNOR U921 ( .A(p_input[428]), .B(n1016), .Z(n591) );
  AND U922 ( .A(n97), .B(n1017), .Z(n1016) );
  XOR U923 ( .A(p_input[444]), .B(p_input[428]), .Z(n1017) );
  XNOR U924 ( .A(n588), .B(n1012), .Z(n1014) );
  XOR U925 ( .A(n1018), .B(n1019), .Z(n588) );
  AND U926 ( .A(n94), .B(n1020), .Z(n1019) );
  XOR U927 ( .A(p_input[412]), .B(p_input[396]), .Z(n1020) );
  XOR U928 ( .A(n1021), .B(n1022), .Z(n1012) );
  AND U929 ( .A(n1023), .B(n1024), .Z(n1022) );
  XOR U930 ( .A(n1021), .B(n603), .Z(n1024) );
  XNOR U931 ( .A(p_input[427]), .B(n1025), .Z(n603) );
  AND U932 ( .A(n97), .B(n1026), .Z(n1025) );
  XOR U933 ( .A(p_input[443]), .B(p_input[427]), .Z(n1026) );
  XNOR U934 ( .A(n600), .B(n1021), .Z(n1023) );
  XOR U935 ( .A(n1027), .B(n1028), .Z(n600) );
  AND U936 ( .A(n94), .B(n1029), .Z(n1028) );
  XOR U937 ( .A(p_input[411]), .B(p_input[395]), .Z(n1029) );
  XOR U938 ( .A(n1030), .B(n1031), .Z(n1021) );
  AND U939 ( .A(n1032), .B(n1033), .Z(n1031) );
  XOR U940 ( .A(n1030), .B(n615), .Z(n1033) );
  XNOR U941 ( .A(p_input[426]), .B(n1034), .Z(n615) );
  AND U942 ( .A(n97), .B(n1035), .Z(n1034) );
  XOR U943 ( .A(p_input[442]), .B(p_input[426]), .Z(n1035) );
  XNOR U944 ( .A(n612), .B(n1030), .Z(n1032) );
  XOR U945 ( .A(n1036), .B(n1037), .Z(n612) );
  AND U946 ( .A(n94), .B(n1038), .Z(n1037) );
  XOR U947 ( .A(p_input[410]), .B(p_input[394]), .Z(n1038) );
  XOR U948 ( .A(n1039), .B(n1040), .Z(n1030) );
  AND U949 ( .A(n1041), .B(n1042), .Z(n1040) );
  XOR U950 ( .A(n1039), .B(n627), .Z(n1042) );
  XNOR U951 ( .A(p_input[425]), .B(n1043), .Z(n627) );
  AND U952 ( .A(n97), .B(n1044), .Z(n1043) );
  XOR U953 ( .A(p_input[441]), .B(p_input[425]), .Z(n1044) );
  XNOR U954 ( .A(n624), .B(n1039), .Z(n1041) );
  XOR U955 ( .A(n1045), .B(n1046), .Z(n624) );
  AND U956 ( .A(n94), .B(n1047), .Z(n1046) );
  XOR U957 ( .A(p_input[409]), .B(p_input[393]), .Z(n1047) );
  XOR U958 ( .A(n1048), .B(n1049), .Z(n1039) );
  AND U959 ( .A(n1050), .B(n1051), .Z(n1049) );
  XOR U960 ( .A(n1048), .B(n639), .Z(n1051) );
  XNOR U961 ( .A(p_input[424]), .B(n1052), .Z(n639) );
  AND U962 ( .A(n97), .B(n1053), .Z(n1052) );
  XOR U963 ( .A(p_input[440]), .B(p_input[424]), .Z(n1053) );
  XNOR U964 ( .A(n636), .B(n1048), .Z(n1050) );
  XOR U965 ( .A(n1054), .B(n1055), .Z(n636) );
  AND U966 ( .A(n94), .B(n1056), .Z(n1055) );
  XOR U967 ( .A(p_input[408]), .B(p_input[392]), .Z(n1056) );
  XOR U968 ( .A(n1057), .B(n1058), .Z(n1048) );
  AND U969 ( .A(n1059), .B(n1060), .Z(n1058) );
  XOR U970 ( .A(n1057), .B(n651), .Z(n1060) );
  XNOR U971 ( .A(p_input[423]), .B(n1061), .Z(n651) );
  AND U972 ( .A(n97), .B(n1062), .Z(n1061) );
  XOR U973 ( .A(p_input[439]), .B(p_input[423]), .Z(n1062) );
  XNOR U974 ( .A(n648), .B(n1057), .Z(n1059) );
  XOR U975 ( .A(n1063), .B(n1064), .Z(n648) );
  AND U976 ( .A(n94), .B(n1065), .Z(n1064) );
  XOR U977 ( .A(p_input[407]), .B(p_input[391]), .Z(n1065) );
  XOR U978 ( .A(n1066), .B(n1067), .Z(n1057) );
  AND U979 ( .A(n1068), .B(n1069), .Z(n1067) );
  XOR U980 ( .A(n1066), .B(n663), .Z(n1069) );
  XNOR U981 ( .A(p_input[422]), .B(n1070), .Z(n663) );
  AND U982 ( .A(n97), .B(n1071), .Z(n1070) );
  XOR U983 ( .A(p_input[438]), .B(p_input[422]), .Z(n1071) );
  XNOR U984 ( .A(n660), .B(n1066), .Z(n1068) );
  XOR U985 ( .A(n1072), .B(n1073), .Z(n660) );
  AND U986 ( .A(n94), .B(n1074), .Z(n1073) );
  XOR U987 ( .A(p_input[406]), .B(p_input[390]), .Z(n1074) );
  XOR U988 ( .A(n1075), .B(n1076), .Z(n1066) );
  AND U989 ( .A(n1077), .B(n1078), .Z(n1076) );
  XOR U990 ( .A(n1075), .B(n675), .Z(n1078) );
  XNOR U991 ( .A(p_input[421]), .B(n1079), .Z(n675) );
  AND U992 ( .A(n97), .B(n1080), .Z(n1079) );
  XOR U993 ( .A(p_input[437]), .B(p_input[421]), .Z(n1080) );
  XNOR U994 ( .A(n672), .B(n1075), .Z(n1077) );
  XOR U995 ( .A(n1081), .B(n1082), .Z(n672) );
  AND U996 ( .A(n94), .B(n1083), .Z(n1082) );
  XOR U997 ( .A(p_input[405]), .B(p_input[389]), .Z(n1083) );
  XOR U998 ( .A(n1084), .B(n1085), .Z(n1075) );
  AND U999 ( .A(n1086), .B(n1087), .Z(n1085) );
  XOR U1000 ( .A(n687), .B(n1084), .Z(n1087) );
  XNOR U1001 ( .A(p_input[420]), .B(n1088), .Z(n687) );
  AND U1002 ( .A(n97), .B(n1089), .Z(n1088) );
  XOR U1003 ( .A(p_input[436]), .B(p_input[420]), .Z(n1089) );
  XNOR U1004 ( .A(n1084), .B(n684), .Z(n1086) );
  XOR U1005 ( .A(n1090), .B(n1091), .Z(n684) );
  AND U1006 ( .A(n94), .B(n1092), .Z(n1091) );
  XOR U1007 ( .A(p_input[404]), .B(p_input[388]), .Z(n1092) );
  XOR U1008 ( .A(n1093), .B(n1094), .Z(n1084) );
  AND U1009 ( .A(n1095), .B(n1096), .Z(n1094) );
  XOR U1010 ( .A(n1093), .B(n699), .Z(n1096) );
  XNOR U1011 ( .A(p_input[419]), .B(n1097), .Z(n699) );
  AND U1012 ( .A(n97), .B(n1098), .Z(n1097) );
  XOR U1013 ( .A(p_input[435]), .B(p_input[419]), .Z(n1098) );
  XNOR U1014 ( .A(n696), .B(n1093), .Z(n1095) );
  XOR U1015 ( .A(n1099), .B(n1100), .Z(n696) );
  AND U1016 ( .A(n94), .B(n1101), .Z(n1100) );
  XOR U1017 ( .A(p_input[403]), .B(p_input[387]), .Z(n1101) );
  XOR U1018 ( .A(n1102), .B(n1103), .Z(n1093) );
  AND U1019 ( .A(n1104), .B(n1105), .Z(n1103) );
  XOR U1020 ( .A(n1102), .B(n711), .Z(n1105) );
  XNOR U1021 ( .A(p_input[418]), .B(n1106), .Z(n711) );
  AND U1022 ( .A(n97), .B(n1107), .Z(n1106) );
  XOR U1023 ( .A(p_input[434]), .B(p_input[418]), .Z(n1107) );
  XNOR U1024 ( .A(n708), .B(n1102), .Z(n1104) );
  XOR U1025 ( .A(n1108), .B(n1109), .Z(n708) );
  AND U1026 ( .A(n94), .B(n1110), .Z(n1109) );
  XOR U1027 ( .A(p_input[402]), .B(p_input[386]), .Z(n1110) );
  XOR U1028 ( .A(n1111), .B(n1112), .Z(n1102) );
  AND U1029 ( .A(n1113), .B(n1114), .Z(n1112) );
  XNOR U1030 ( .A(n1115), .B(n724), .Z(n1114) );
  XNOR U1031 ( .A(p_input[417]), .B(n1116), .Z(n724) );
  AND U1032 ( .A(n97), .B(n1117), .Z(n1116) );
  XNOR U1033 ( .A(p_input[433]), .B(n1118), .Z(n1117) );
  IV U1034 ( .A(p_input[417]), .Z(n1118) );
  XNOR U1035 ( .A(n721), .B(n1111), .Z(n1113) );
  XNOR U1036 ( .A(p_input[385]), .B(n1119), .Z(n721) );
  AND U1037 ( .A(n94), .B(n1120), .Z(n1119) );
  XOR U1038 ( .A(p_input[401]), .B(p_input[385]), .Z(n1120) );
  IV U1039 ( .A(n1115), .Z(n1111) );
  AND U1040 ( .A(n986), .B(n989), .Z(n1115) );
  XOR U1041 ( .A(p_input[416]), .B(n1121), .Z(n989) );
  AND U1042 ( .A(n97), .B(n1122), .Z(n1121) );
  XOR U1043 ( .A(p_input[432]), .B(p_input[416]), .Z(n1122) );
  XOR U1044 ( .A(n1123), .B(n1124), .Z(n97) );
  AND U1045 ( .A(n1125), .B(n1126), .Z(n1124) );
  XNOR U1046 ( .A(p_input[447]), .B(n1123), .Z(n1126) );
  XOR U1047 ( .A(n1123), .B(p_input[431]), .Z(n1125) );
  XOR U1048 ( .A(n1127), .B(n1128), .Z(n1123) );
  AND U1049 ( .A(n1129), .B(n1130), .Z(n1128) );
  XNOR U1050 ( .A(p_input[446]), .B(n1127), .Z(n1130) );
  XOR U1051 ( .A(n1127), .B(p_input[430]), .Z(n1129) );
  XOR U1052 ( .A(n1131), .B(n1132), .Z(n1127) );
  AND U1053 ( .A(n1133), .B(n1134), .Z(n1132) );
  XNOR U1054 ( .A(p_input[445]), .B(n1131), .Z(n1134) );
  XOR U1055 ( .A(n1131), .B(p_input[429]), .Z(n1133) );
  XOR U1056 ( .A(n1135), .B(n1136), .Z(n1131) );
  AND U1057 ( .A(n1137), .B(n1138), .Z(n1136) );
  XNOR U1058 ( .A(p_input[444]), .B(n1135), .Z(n1138) );
  XOR U1059 ( .A(n1135), .B(p_input[428]), .Z(n1137) );
  XOR U1060 ( .A(n1139), .B(n1140), .Z(n1135) );
  AND U1061 ( .A(n1141), .B(n1142), .Z(n1140) );
  XNOR U1062 ( .A(p_input[443]), .B(n1139), .Z(n1142) );
  XOR U1063 ( .A(n1139), .B(p_input[427]), .Z(n1141) );
  XOR U1064 ( .A(n1143), .B(n1144), .Z(n1139) );
  AND U1065 ( .A(n1145), .B(n1146), .Z(n1144) );
  XNOR U1066 ( .A(p_input[442]), .B(n1143), .Z(n1146) );
  XOR U1067 ( .A(n1143), .B(p_input[426]), .Z(n1145) );
  XOR U1068 ( .A(n1147), .B(n1148), .Z(n1143) );
  AND U1069 ( .A(n1149), .B(n1150), .Z(n1148) );
  XNOR U1070 ( .A(p_input[441]), .B(n1147), .Z(n1150) );
  XOR U1071 ( .A(n1147), .B(p_input[425]), .Z(n1149) );
  XOR U1072 ( .A(n1151), .B(n1152), .Z(n1147) );
  AND U1073 ( .A(n1153), .B(n1154), .Z(n1152) );
  XNOR U1074 ( .A(p_input[440]), .B(n1151), .Z(n1154) );
  XOR U1075 ( .A(n1151), .B(p_input[424]), .Z(n1153) );
  XOR U1076 ( .A(n1155), .B(n1156), .Z(n1151) );
  AND U1077 ( .A(n1157), .B(n1158), .Z(n1156) );
  XNOR U1078 ( .A(p_input[439]), .B(n1155), .Z(n1158) );
  XOR U1079 ( .A(n1155), .B(p_input[423]), .Z(n1157) );
  XOR U1080 ( .A(n1159), .B(n1160), .Z(n1155) );
  AND U1081 ( .A(n1161), .B(n1162), .Z(n1160) );
  XNOR U1082 ( .A(p_input[438]), .B(n1159), .Z(n1162) );
  XOR U1083 ( .A(n1159), .B(p_input[422]), .Z(n1161) );
  XOR U1084 ( .A(n1163), .B(n1164), .Z(n1159) );
  AND U1085 ( .A(n1165), .B(n1166), .Z(n1164) );
  XNOR U1086 ( .A(p_input[437]), .B(n1163), .Z(n1166) );
  XOR U1087 ( .A(n1163), .B(p_input[421]), .Z(n1165) );
  XOR U1088 ( .A(n1167), .B(n1168), .Z(n1163) );
  AND U1089 ( .A(n1169), .B(n1170), .Z(n1168) );
  XNOR U1090 ( .A(p_input[436]), .B(n1167), .Z(n1170) );
  XOR U1091 ( .A(n1167), .B(p_input[420]), .Z(n1169) );
  XOR U1092 ( .A(n1171), .B(n1172), .Z(n1167) );
  AND U1093 ( .A(n1173), .B(n1174), .Z(n1172) );
  XNOR U1094 ( .A(p_input[435]), .B(n1171), .Z(n1174) );
  XOR U1095 ( .A(n1171), .B(p_input[419]), .Z(n1173) );
  XOR U1096 ( .A(n1175), .B(n1176), .Z(n1171) );
  AND U1097 ( .A(n1177), .B(n1178), .Z(n1176) );
  XNOR U1098 ( .A(p_input[434]), .B(n1175), .Z(n1178) );
  XOR U1099 ( .A(n1175), .B(p_input[418]), .Z(n1177) );
  XNOR U1100 ( .A(n1179), .B(n1180), .Z(n1175) );
  AND U1101 ( .A(n1181), .B(n1182), .Z(n1180) );
  XOR U1102 ( .A(p_input[433]), .B(n1179), .Z(n1182) );
  XNOR U1103 ( .A(p_input[417]), .B(n1179), .Z(n1181) );
  AND U1104 ( .A(p_input[432]), .B(n1183), .Z(n1179) );
  IV U1105 ( .A(p_input[416]), .Z(n1183) );
  XNOR U1106 ( .A(p_input[384]), .B(n1184), .Z(n986) );
  AND U1107 ( .A(n94), .B(n1185), .Z(n1184) );
  XOR U1108 ( .A(p_input[400]), .B(p_input[384]), .Z(n1185) );
  XOR U1109 ( .A(n1186), .B(n1187), .Z(n94) );
  AND U1110 ( .A(n1188), .B(n1189), .Z(n1187) );
  XNOR U1111 ( .A(p_input[415]), .B(n1186), .Z(n1189) );
  XOR U1112 ( .A(n1186), .B(p_input[399]), .Z(n1188) );
  XOR U1113 ( .A(n1190), .B(n1191), .Z(n1186) );
  AND U1114 ( .A(n1192), .B(n1193), .Z(n1191) );
  XNOR U1115 ( .A(p_input[414]), .B(n1190), .Z(n1193) );
  XNOR U1116 ( .A(n1190), .B(n1000), .Z(n1192) );
  IV U1117 ( .A(p_input[398]), .Z(n1000) );
  XOR U1118 ( .A(n1194), .B(n1195), .Z(n1190) );
  AND U1119 ( .A(n1196), .B(n1197), .Z(n1195) );
  XNOR U1120 ( .A(p_input[413]), .B(n1194), .Z(n1197) );
  XNOR U1121 ( .A(n1194), .B(n1009), .Z(n1196) );
  IV U1122 ( .A(p_input[397]), .Z(n1009) );
  XOR U1123 ( .A(n1198), .B(n1199), .Z(n1194) );
  AND U1124 ( .A(n1200), .B(n1201), .Z(n1199) );
  XNOR U1125 ( .A(p_input[412]), .B(n1198), .Z(n1201) );
  XNOR U1126 ( .A(n1198), .B(n1018), .Z(n1200) );
  IV U1127 ( .A(p_input[396]), .Z(n1018) );
  XOR U1128 ( .A(n1202), .B(n1203), .Z(n1198) );
  AND U1129 ( .A(n1204), .B(n1205), .Z(n1203) );
  XNOR U1130 ( .A(p_input[411]), .B(n1202), .Z(n1205) );
  XNOR U1131 ( .A(n1202), .B(n1027), .Z(n1204) );
  IV U1132 ( .A(p_input[395]), .Z(n1027) );
  XOR U1133 ( .A(n1206), .B(n1207), .Z(n1202) );
  AND U1134 ( .A(n1208), .B(n1209), .Z(n1207) );
  XNOR U1135 ( .A(p_input[410]), .B(n1206), .Z(n1209) );
  XNOR U1136 ( .A(n1206), .B(n1036), .Z(n1208) );
  IV U1137 ( .A(p_input[394]), .Z(n1036) );
  XOR U1138 ( .A(n1210), .B(n1211), .Z(n1206) );
  AND U1139 ( .A(n1212), .B(n1213), .Z(n1211) );
  XNOR U1140 ( .A(p_input[409]), .B(n1210), .Z(n1213) );
  XNOR U1141 ( .A(n1210), .B(n1045), .Z(n1212) );
  IV U1142 ( .A(p_input[393]), .Z(n1045) );
  XOR U1143 ( .A(n1214), .B(n1215), .Z(n1210) );
  AND U1144 ( .A(n1216), .B(n1217), .Z(n1215) );
  XNOR U1145 ( .A(p_input[408]), .B(n1214), .Z(n1217) );
  XNOR U1146 ( .A(n1214), .B(n1054), .Z(n1216) );
  IV U1147 ( .A(p_input[392]), .Z(n1054) );
  XOR U1148 ( .A(n1218), .B(n1219), .Z(n1214) );
  AND U1149 ( .A(n1220), .B(n1221), .Z(n1219) );
  XNOR U1150 ( .A(p_input[407]), .B(n1218), .Z(n1221) );
  XNOR U1151 ( .A(n1218), .B(n1063), .Z(n1220) );
  IV U1152 ( .A(p_input[391]), .Z(n1063) );
  XOR U1153 ( .A(n1222), .B(n1223), .Z(n1218) );
  AND U1154 ( .A(n1224), .B(n1225), .Z(n1223) );
  XNOR U1155 ( .A(p_input[406]), .B(n1222), .Z(n1225) );
  XNOR U1156 ( .A(n1222), .B(n1072), .Z(n1224) );
  IV U1157 ( .A(p_input[390]), .Z(n1072) );
  XOR U1158 ( .A(n1226), .B(n1227), .Z(n1222) );
  AND U1159 ( .A(n1228), .B(n1229), .Z(n1227) );
  XNOR U1160 ( .A(p_input[405]), .B(n1226), .Z(n1229) );
  XNOR U1161 ( .A(n1226), .B(n1081), .Z(n1228) );
  IV U1162 ( .A(p_input[389]), .Z(n1081) );
  XOR U1163 ( .A(n1230), .B(n1231), .Z(n1226) );
  AND U1164 ( .A(n1232), .B(n1233), .Z(n1231) );
  XNOR U1165 ( .A(p_input[404]), .B(n1230), .Z(n1233) );
  XNOR U1166 ( .A(n1230), .B(n1090), .Z(n1232) );
  IV U1167 ( .A(p_input[388]), .Z(n1090) );
  XOR U1168 ( .A(n1234), .B(n1235), .Z(n1230) );
  AND U1169 ( .A(n1236), .B(n1237), .Z(n1235) );
  XNOR U1170 ( .A(p_input[403]), .B(n1234), .Z(n1237) );
  XNOR U1171 ( .A(n1234), .B(n1099), .Z(n1236) );
  IV U1172 ( .A(p_input[387]), .Z(n1099) );
  XOR U1173 ( .A(n1238), .B(n1239), .Z(n1234) );
  AND U1174 ( .A(n1240), .B(n1241), .Z(n1239) );
  XNOR U1175 ( .A(p_input[402]), .B(n1238), .Z(n1241) );
  XNOR U1176 ( .A(n1238), .B(n1108), .Z(n1240) );
  IV U1177 ( .A(p_input[386]), .Z(n1108) );
  XNOR U1178 ( .A(n1242), .B(n1243), .Z(n1238) );
  AND U1179 ( .A(n1244), .B(n1245), .Z(n1243) );
  XOR U1180 ( .A(p_input[401]), .B(n1242), .Z(n1245) );
  XNOR U1181 ( .A(p_input[385]), .B(n1242), .Z(n1244) );
  AND U1182 ( .A(p_input[400]), .B(n1246), .Z(n1242) );
  IV U1183 ( .A(p_input[384]), .Z(n1246) );
  XOR U1184 ( .A(n1247), .B(n1248), .Z(n362) );
  AND U1185 ( .A(n159), .B(n1249), .Z(n1248) );
  XNOR U1186 ( .A(n1250), .B(n1247), .Z(n1249) );
  XOR U1187 ( .A(n1251), .B(n1252), .Z(n159) );
  AND U1188 ( .A(n1253), .B(n1254), .Z(n1252) );
  XNOR U1189 ( .A(n374), .B(n1251), .Z(n1254) );
  AND U1190 ( .A(n1255), .B(n1256), .Z(n374) );
  XOR U1191 ( .A(n1251), .B(n373), .Z(n1253) );
  AND U1192 ( .A(n1257), .B(n1258), .Z(n373) );
  XOR U1193 ( .A(n1259), .B(n1260), .Z(n1251) );
  AND U1194 ( .A(n1261), .B(n1262), .Z(n1260) );
  XOR U1195 ( .A(n1259), .B(n386), .Z(n1262) );
  XOR U1196 ( .A(n1263), .B(n1264), .Z(n386) );
  AND U1197 ( .A(n125), .B(n1265), .Z(n1264) );
  XOR U1198 ( .A(n1266), .B(n1263), .Z(n1265) );
  XNOR U1199 ( .A(n383), .B(n1259), .Z(n1261) );
  XOR U1200 ( .A(n1267), .B(n1268), .Z(n383) );
  AND U1201 ( .A(n122), .B(n1269), .Z(n1268) );
  XOR U1202 ( .A(n1270), .B(n1267), .Z(n1269) );
  XOR U1203 ( .A(n1271), .B(n1272), .Z(n1259) );
  AND U1204 ( .A(n1273), .B(n1274), .Z(n1272) );
  XOR U1205 ( .A(n1271), .B(n398), .Z(n1274) );
  XOR U1206 ( .A(n1275), .B(n1276), .Z(n398) );
  AND U1207 ( .A(n125), .B(n1277), .Z(n1276) );
  XOR U1208 ( .A(n1278), .B(n1275), .Z(n1277) );
  XNOR U1209 ( .A(n395), .B(n1271), .Z(n1273) );
  XOR U1210 ( .A(n1279), .B(n1280), .Z(n395) );
  AND U1211 ( .A(n122), .B(n1281), .Z(n1280) );
  XOR U1212 ( .A(n1282), .B(n1279), .Z(n1281) );
  XOR U1213 ( .A(n1283), .B(n1284), .Z(n1271) );
  AND U1214 ( .A(n1285), .B(n1286), .Z(n1284) );
  XOR U1215 ( .A(n1283), .B(n410), .Z(n1286) );
  XOR U1216 ( .A(n1287), .B(n1288), .Z(n410) );
  AND U1217 ( .A(n125), .B(n1289), .Z(n1288) );
  XOR U1218 ( .A(n1290), .B(n1287), .Z(n1289) );
  XNOR U1219 ( .A(n407), .B(n1283), .Z(n1285) );
  XOR U1220 ( .A(n1291), .B(n1292), .Z(n407) );
  AND U1221 ( .A(n122), .B(n1293), .Z(n1292) );
  XOR U1222 ( .A(n1294), .B(n1291), .Z(n1293) );
  XOR U1223 ( .A(n1295), .B(n1296), .Z(n1283) );
  AND U1224 ( .A(n1297), .B(n1298), .Z(n1296) );
  XOR U1225 ( .A(n1295), .B(n422), .Z(n1298) );
  XOR U1226 ( .A(n1299), .B(n1300), .Z(n422) );
  AND U1227 ( .A(n125), .B(n1301), .Z(n1300) );
  XOR U1228 ( .A(n1302), .B(n1299), .Z(n1301) );
  XNOR U1229 ( .A(n419), .B(n1295), .Z(n1297) );
  XOR U1230 ( .A(n1303), .B(n1304), .Z(n419) );
  AND U1231 ( .A(n122), .B(n1305), .Z(n1304) );
  XOR U1232 ( .A(n1306), .B(n1303), .Z(n1305) );
  XOR U1233 ( .A(n1307), .B(n1308), .Z(n1295) );
  AND U1234 ( .A(n1309), .B(n1310), .Z(n1308) );
  XOR U1235 ( .A(n1307), .B(n434), .Z(n1310) );
  XOR U1236 ( .A(n1311), .B(n1312), .Z(n434) );
  AND U1237 ( .A(n125), .B(n1313), .Z(n1312) );
  XOR U1238 ( .A(n1314), .B(n1311), .Z(n1313) );
  XNOR U1239 ( .A(n431), .B(n1307), .Z(n1309) );
  XOR U1240 ( .A(n1315), .B(n1316), .Z(n431) );
  AND U1241 ( .A(n122), .B(n1317), .Z(n1316) );
  XOR U1242 ( .A(n1318), .B(n1315), .Z(n1317) );
  XOR U1243 ( .A(n1319), .B(n1320), .Z(n1307) );
  AND U1244 ( .A(n1321), .B(n1322), .Z(n1320) );
  XOR U1245 ( .A(n1319), .B(n446), .Z(n1322) );
  XOR U1246 ( .A(n1323), .B(n1324), .Z(n446) );
  AND U1247 ( .A(n125), .B(n1325), .Z(n1324) );
  XOR U1248 ( .A(n1326), .B(n1323), .Z(n1325) );
  XNOR U1249 ( .A(n443), .B(n1319), .Z(n1321) );
  XOR U1250 ( .A(n1327), .B(n1328), .Z(n443) );
  AND U1251 ( .A(n122), .B(n1329), .Z(n1328) );
  XOR U1252 ( .A(n1330), .B(n1327), .Z(n1329) );
  XOR U1253 ( .A(n1331), .B(n1332), .Z(n1319) );
  AND U1254 ( .A(n1333), .B(n1334), .Z(n1332) );
  XOR U1255 ( .A(n1331), .B(n458), .Z(n1334) );
  XOR U1256 ( .A(n1335), .B(n1336), .Z(n458) );
  AND U1257 ( .A(n125), .B(n1337), .Z(n1336) );
  XOR U1258 ( .A(n1338), .B(n1335), .Z(n1337) );
  XNOR U1259 ( .A(n455), .B(n1331), .Z(n1333) );
  XOR U1260 ( .A(n1339), .B(n1340), .Z(n455) );
  AND U1261 ( .A(n122), .B(n1341), .Z(n1340) );
  XOR U1262 ( .A(n1342), .B(n1339), .Z(n1341) );
  XOR U1263 ( .A(n1343), .B(n1344), .Z(n1331) );
  AND U1264 ( .A(n1345), .B(n1346), .Z(n1344) );
  XOR U1265 ( .A(n1343), .B(n470), .Z(n1346) );
  XOR U1266 ( .A(n1347), .B(n1348), .Z(n470) );
  AND U1267 ( .A(n125), .B(n1349), .Z(n1348) );
  XOR U1268 ( .A(n1350), .B(n1347), .Z(n1349) );
  XNOR U1269 ( .A(n467), .B(n1343), .Z(n1345) );
  XOR U1270 ( .A(n1351), .B(n1352), .Z(n467) );
  AND U1271 ( .A(n122), .B(n1353), .Z(n1352) );
  XOR U1272 ( .A(n1354), .B(n1351), .Z(n1353) );
  XOR U1273 ( .A(n1355), .B(n1356), .Z(n1343) );
  AND U1274 ( .A(n1357), .B(n1358), .Z(n1356) );
  XOR U1275 ( .A(n1355), .B(n482), .Z(n1358) );
  XOR U1276 ( .A(n1359), .B(n1360), .Z(n482) );
  AND U1277 ( .A(n125), .B(n1361), .Z(n1360) );
  XOR U1278 ( .A(n1362), .B(n1359), .Z(n1361) );
  XNOR U1279 ( .A(n479), .B(n1355), .Z(n1357) );
  XOR U1280 ( .A(n1363), .B(n1364), .Z(n479) );
  AND U1281 ( .A(n122), .B(n1365), .Z(n1364) );
  XOR U1282 ( .A(n1366), .B(n1363), .Z(n1365) );
  XOR U1283 ( .A(n1367), .B(n1368), .Z(n1355) );
  AND U1284 ( .A(n1369), .B(n1370), .Z(n1368) );
  XOR U1285 ( .A(n1367), .B(n494), .Z(n1370) );
  XOR U1286 ( .A(n1371), .B(n1372), .Z(n494) );
  AND U1287 ( .A(n125), .B(n1373), .Z(n1372) );
  XOR U1288 ( .A(n1374), .B(n1371), .Z(n1373) );
  XNOR U1289 ( .A(n491), .B(n1367), .Z(n1369) );
  XOR U1290 ( .A(n1375), .B(n1376), .Z(n491) );
  AND U1291 ( .A(n122), .B(n1377), .Z(n1376) );
  XOR U1292 ( .A(n1378), .B(n1375), .Z(n1377) );
  XOR U1293 ( .A(n1379), .B(n1380), .Z(n1367) );
  AND U1294 ( .A(n1381), .B(n1382), .Z(n1380) );
  XOR U1295 ( .A(n506), .B(n1379), .Z(n1382) );
  XOR U1296 ( .A(n1383), .B(n1384), .Z(n506) );
  AND U1297 ( .A(n125), .B(n1385), .Z(n1384) );
  XOR U1298 ( .A(n1383), .B(n1386), .Z(n1385) );
  XNOR U1299 ( .A(n1379), .B(n503), .Z(n1381) );
  XOR U1300 ( .A(n1387), .B(n1388), .Z(n503) );
  AND U1301 ( .A(n122), .B(n1389), .Z(n1388) );
  XOR U1302 ( .A(n1387), .B(n1390), .Z(n1389) );
  XOR U1303 ( .A(n1391), .B(n1392), .Z(n1379) );
  AND U1304 ( .A(n1393), .B(n1394), .Z(n1392) );
  XOR U1305 ( .A(n1391), .B(n518), .Z(n1394) );
  XOR U1306 ( .A(n1395), .B(n1396), .Z(n518) );
  AND U1307 ( .A(n125), .B(n1397), .Z(n1396) );
  XOR U1308 ( .A(n1398), .B(n1395), .Z(n1397) );
  XNOR U1309 ( .A(n515), .B(n1391), .Z(n1393) );
  XOR U1310 ( .A(n1399), .B(n1400), .Z(n515) );
  AND U1311 ( .A(n122), .B(n1401), .Z(n1400) );
  XOR U1312 ( .A(n1402), .B(n1399), .Z(n1401) );
  XOR U1313 ( .A(n1403), .B(n1404), .Z(n1391) );
  AND U1314 ( .A(n1405), .B(n1406), .Z(n1404) );
  XOR U1315 ( .A(n1403), .B(n530), .Z(n1406) );
  XOR U1316 ( .A(n1407), .B(n1408), .Z(n530) );
  AND U1317 ( .A(n125), .B(n1409), .Z(n1408) );
  XOR U1318 ( .A(n1410), .B(n1407), .Z(n1409) );
  XNOR U1319 ( .A(n527), .B(n1403), .Z(n1405) );
  XOR U1320 ( .A(n1411), .B(n1412), .Z(n527) );
  AND U1321 ( .A(n122), .B(n1413), .Z(n1412) );
  XOR U1322 ( .A(n1414), .B(n1411), .Z(n1413) );
  XOR U1323 ( .A(n1415), .B(n1416), .Z(n1403) );
  AND U1324 ( .A(n1417), .B(n1418), .Z(n1416) );
  XNOR U1325 ( .A(n1419), .B(n543), .Z(n1418) );
  XOR U1326 ( .A(n1420), .B(n1421), .Z(n543) );
  AND U1327 ( .A(n125), .B(n1422), .Z(n1421) );
  XOR U1328 ( .A(n1423), .B(n1420), .Z(n1422) );
  XNOR U1329 ( .A(n540), .B(n1415), .Z(n1417) );
  XOR U1330 ( .A(n1424), .B(n1425), .Z(n540) );
  AND U1331 ( .A(n122), .B(n1426), .Z(n1425) );
  XOR U1332 ( .A(n1427), .B(n1424), .Z(n1426) );
  IV U1333 ( .A(n1419), .Z(n1415) );
  AND U1334 ( .A(n1247), .B(n1250), .Z(n1419) );
  XNOR U1335 ( .A(n1428), .B(n1429), .Z(n1250) );
  AND U1336 ( .A(n125), .B(n1430), .Z(n1429) );
  XNOR U1337 ( .A(n1431), .B(n1428), .Z(n1430) );
  XOR U1338 ( .A(n1432), .B(n1433), .Z(n125) );
  AND U1339 ( .A(n1434), .B(n1435), .Z(n1433) );
  XNOR U1340 ( .A(n1255), .B(n1432), .Z(n1435) );
  AND U1341 ( .A(p_input[383]), .B(p_input[367]), .Z(n1255) );
  XOR U1342 ( .A(n1432), .B(n1256), .Z(n1434) );
  AND U1343 ( .A(p_input[351]), .B(p_input[335]), .Z(n1256) );
  XOR U1344 ( .A(n1436), .B(n1437), .Z(n1432) );
  AND U1345 ( .A(n1438), .B(n1439), .Z(n1437) );
  XOR U1346 ( .A(n1436), .B(n1266), .Z(n1439) );
  XNOR U1347 ( .A(p_input[366]), .B(n1440), .Z(n1266) );
  AND U1348 ( .A(n105), .B(n1441), .Z(n1440) );
  XOR U1349 ( .A(p_input[382]), .B(p_input[366]), .Z(n1441) );
  XNOR U1350 ( .A(n1263), .B(n1436), .Z(n1438) );
  XOR U1351 ( .A(n1442), .B(n1443), .Z(n1263) );
  AND U1352 ( .A(n103), .B(n1444), .Z(n1443) );
  XOR U1353 ( .A(p_input[350]), .B(p_input[334]), .Z(n1444) );
  XOR U1354 ( .A(n1445), .B(n1446), .Z(n1436) );
  AND U1355 ( .A(n1447), .B(n1448), .Z(n1446) );
  XOR U1356 ( .A(n1445), .B(n1278), .Z(n1448) );
  XNOR U1357 ( .A(p_input[365]), .B(n1449), .Z(n1278) );
  AND U1358 ( .A(n105), .B(n1450), .Z(n1449) );
  XOR U1359 ( .A(p_input[381]), .B(p_input[365]), .Z(n1450) );
  XNOR U1360 ( .A(n1275), .B(n1445), .Z(n1447) );
  XOR U1361 ( .A(n1451), .B(n1452), .Z(n1275) );
  AND U1362 ( .A(n103), .B(n1453), .Z(n1452) );
  XOR U1363 ( .A(p_input[349]), .B(p_input[333]), .Z(n1453) );
  XOR U1364 ( .A(n1454), .B(n1455), .Z(n1445) );
  AND U1365 ( .A(n1456), .B(n1457), .Z(n1455) );
  XOR U1366 ( .A(n1454), .B(n1290), .Z(n1457) );
  XNOR U1367 ( .A(p_input[364]), .B(n1458), .Z(n1290) );
  AND U1368 ( .A(n105), .B(n1459), .Z(n1458) );
  XOR U1369 ( .A(p_input[380]), .B(p_input[364]), .Z(n1459) );
  XNOR U1370 ( .A(n1287), .B(n1454), .Z(n1456) );
  XOR U1371 ( .A(n1460), .B(n1461), .Z(n1287) );
  AND U1372 ( .A(n103), .B(n1462), .Z(n1461) );
  XOR U1373 ( .A(p_input[348]), .B(p_input[332]), .Z(n1462) );
  XOR U1374 ( .A(n1463), .B(n1464), .Z(n1454) );
  AND U1375 ( .A(n1465), .B(n1466), .Z(n1464) );
  XOR U1376 ( .A(n1463), .B(n1302), .Z(n1466) );
  XNOR U1377 ( .A(p_input[363]), .B(n1467), .Z(n1302) );
  AND U1378 ( .A(n105), .B(n1468), .Z(n1467) );
  XOR U1379 ( .A(p_input[379]), .B(p_input[363]), .Z(n1468) );
  XNOR U1380 ( .A(n1299), .B(n1463), .Z(n1465) );
  XOR U1381 ( .A(n1469), .B(n1470), .Z(n1299) );
  AND U1382 ( .A(n103), .B(n1471), .Z(n1470) );
  XOR U1383 ( .A(p_input[347]), .B(p_input[331]), .Z(n1471) );
  XOR U1384 ( .A(n1472), .B(n1473), .Z(n1463) );
  AND U1385 ( .A(n1474), .B(n1475), .Z(n1473) );
  XOR U1386 ( .A(n1472), .B(n1314), .Z(n1475) );
  XNOR U1387 ( .A(p_input[362]), .B(n1476), .Z(n1314) );
  AND U1388 ( .A(n105), .B(n1477), .Z(n1476) );
  XOR U1389 ( .A(p_input[378]), .B(p_input[362]), .Z(n1477) );
  XNOR U1390 ( .A(n1311), .B(n1472), .Z(n1474) );
  XOR U1391 ( .A(n1478), .B(n1479), .Z(n1311) );
  AND U1392 ( .A(n103), .B(n1480), .Z(n1479) );
  XOR U1393 ( .A(p_input[346]), .B(p_input[330]), .Z(n1480) );
  XOR U1394 ( .A(n1481), .B(n1482), .Z(n1472) );
  AND U1395 ( .A(n1483), .B(n1484), .Z(n1482) );
  XOR U1396 ( .A(n1481), .B(n1326), .Z(n1484) );
  XNOR U1397 ( .A(p_input[361]), .B(n1485), .Z(n1326) );
  AND U1398 ( .A(n105), .B(n1486), .Z(n1485) );
  XOR U1399 ( .A(p_input[377]), .B(p_input[361]), .Z(n1486) );
  XNOR U1400 ( .A(n1323), .B(n1481), .Z(n1483) );
  XOR U1401 ( .A(n1487), .B(n1488), .Z(n1323) );
  AND U1402 ( .A(n103), .B(n1489), .Z(n1488) );
  XOR U1403 ( .A(p_input[345]), .B(p_input[329]), .Z(n1489) );
  XOR U1404 ( .A(n1490), .B(n1491), .Z(n1481) );
  AND U1405 ( .A(n1492), .B(n1493), .Z(n1491) );
  XOR U1406 ( .A(n1490), .B(n1338), .Z(n1493) );
  XNOR U1407 ( .A(p_input[360]), .B(n1494), .Z(n1338) );
  AND U1408 ( .A(n105), .B(n1495), .Z(n1494) );
  XOR U1409 ( .A(p_input[376]), .B(p_input[360]), .Z(n1495) );
  XNOR U1410 ( .A(n1335), .B(n1490), .Z(n1492) );
  XOR U1411 ( .A(n1496), .B(n1497), .Z(n1335) );
  AND U1412 ( .A(n103), .B(n1498), .Z(n1497) );
  XOR U1413 ( .A(p_input[344]), .B(p_input[328]), .Z(n1498) );
  XOR U1414 ( .A(n1499), .B(n1500), .Z(n1490) );
  AND U1415 ( .A(n1501), .B(n1502), .Z(n1500) );
  XOR U1416 ( .A(n1499), .B(n1350), .Z(n1502) );
  XNOR U1417 ( .A(p_input[359]), .B(n1503), .Z(n1350) );
  AND U1418 ( .A(n105), .B(n1504), .Z(n1503) );
  XOR U1419 ( .A(p_input[375]), .B(p_input[359]), .Z(n1504) );
  XNOR U1420 ( .A(n1347), .B(n1499), .Z(n1501) );
  XOR U1421 ( .A(n1505), .B(n1506), .Z(n1347) );
  AND U1422 ( .A(n103), .B(n1507), .Z(n1506) );
  XOR U1423 ( .A(p_input[343]), .B(p_input[327]), .Z(n1507) );
  XOR U1424 ( .A(n1508), .B(n1509), .Z(n1499) );
  AND U1425 ( .A(n1510), .B(n1511), .Z(n1509) );
  XOR U1426 ( .A(n1508), .B(n1362), .Z(n1511) );
  XNOR U1427 ( .A(p_input[358]), .B(n1512), .Z(n1362) );
  AND U1428 ( .A(n105), .B(n1513), .Z(n1512) );
  XOR U1429 ( .A(p_input[374]), .B(p_input[358]), .Z(n1513) );
  XNOR U1430 ( .A(n1359), .B(n1508), .Z(n1510) );
  XOR U1431 ( .A(n1514), .B(n1515), .Z(n1359) );
  AND U1432 ( .A(n103), .B(n1516), .Z(n1515) );
  XOR U1433 ( .A(p_input[342]), .B(p_input[326]), .Z(n1516) );
  XOR U1434 ( .A(n1517), .B(n1518), .Z(n1508) );
  AND U1435 ( .A(n1519), .B(n1520), .Z(n1518) );
  XOR U1436 ( .A(n1517), .B(n1374), .Z(n1520) );
  XNOR U1437 ( .A(p_input[357]), .B(n1521), .Z(n1374) );
  AND U1438 ( .A(n105), .B(n1522), .Z(n1521) );
  XOR U1439 ( .A(p_input[373]), .B(p_input[357]), .Z(n1522) );
  XNOR U1440 ( .A(n1371), .B(n1517), .Z(n1519) );
  XOR U1441 ( .A(n1523), .B(n1524), .Z(n1371) );
  AND U1442 ( .A(n103), .B(n1525), .Z(n1524) );
  XOR U1443 ( .A(p_input[341]), .B(p_input[325]), .Z(n1525) );
  XOR U1444 ( .A(n1526), .B(n1527), .Z(n1517) );
  AND U1445 ( .A(n1528), .B(n1529), .Z(n1527) );
  XOR U1446 ( .A(n1386), .B(n1526), .Z(n1529) );
  XNOR U1447 ( .A(p_input[356]), .B(n1530), .Z(n1386) );
  AND U1448 ( .A(n105), .B(n1531), .Z(n1530) );
  XOR U1449 ( .A(p_input[372]), .B(p_input[356]), .Z(n1531) );
  XNOR U1450 ( .A(n1526), .B(n1383), .Z(n1528) );
  XOR U1451 ( .A(n1532), .B(n1533), .Z(n1383) );
  AND U1452 ( .A(n103), .B(n1534), .Z(n1533) );
  XOR U1453 ( .A(p_input[340]), .B(p_input[324]), .Z(n1534) );
  XOR U1454 ( .A(n1535), .B(n1536), .Z(n1526) );
  AND U1455 ( .A(n1537), .B(n1538), .Z(n1536) );
  XOR U1456 ( .A(n1535), .B(n1398), .Z(n1538) );
  XNOR U1457 ( .A(p_input[355]), .B(n1539), .Z(n1398) );
  AND U1458 ( .A(n105), .B(n1540), .Z(n1539) );
  XOR U1459 ( .A(p_input[371]), .B(p_input[355]), .Z(n1540) );
  XNOR U1460 ( .A(n1395), .B(n1535), .Z(n1537) );
  XOR U1461 ( .A(n1541), .B(n1542), .Z(n1395) );
  AND U1462 ( .A(n103), .B(n1543), .Z(n1542) );
  XOR U1463 ( .A(p_input[339]), .B(p_input[323]), .Z(n1543) );
  XOR U1464 ( .A(n1544), .B(n1545), .Z(n1535) );
  AND U1465 ( .A(n1546), .B(n1547), .Z(n1545) );
  XOR U1466 ( .A(n1544), .B(n1410), .Z(n1547) );
  XNOR U1467 ( .A(p_input[354]), .B(n1548), .Z(n1410) );
  AND U1468 ( .A(n105), .B(n1549), .Z(n1548) );
  XOR U1469 ( .A(p_input[370]), .B(p_input[354]), .Z(n1549) );
  XNOR U1470 ( .A(n1407), .B(n1544), .Z(n1546) );
  XOR U1471 ( .A(n1550), .B(n1551), .Z(n1407) );
  AND U1472 ( .A(n103), .B(n1552), .Z(n1551) );
  XOR U1473 ( .A(p_input[338]), .B(p_input[322]), .Z(n1552) );
  XOR U1474 ( .A(n1553), .B(n1554), .Z(n1544) );
  AND U1475 ( .A(n1555), .B(n1556), .Z(n1554) );
  XNOR U1476 ( .A(n1557), .B(n1423), .Z(n1556) );
  XNOR U1477 ( .A(p_input[353]), .B(n1558), .Z(n1423) );
  AND U1478 ( .A(n105), .B(n1559), .Z(n1558) );
  XNOR U1479 ( .A(p_input[369]), .B(n1560), .Z(n1559) );
  IV U1480 ( .A(p_input[353]), .Z(n1560) );
  XNOR U1481 ( .A(n1420), .B(n1553), .Z(n1555) );
  XNOR U1482 ( .A(p_input[321]), .B(n1561), .Z(n1420) );
  AND U1483 ( .A(n103), .B(n1562), .Z(n1561) );
  XOR U1484 ( .A(p_input[337]), .B(p_input[321]), .Z(n1562) );
  IV U1485 ( .A(n1557), .Z(n1553) );
  AND U1486 ( .A(n1428), .B(n1431), .Z(n1557) );
  XOR U1487 ( .A(p_input[352]), .B(n1563), .Z(n1431) );
  AND U1488 ( .A(n105), .B(n1564), .Z(n1563) );
  XOR U1489 ( .A(p_input[368]), .B(p_input[352]), .Z(n1564) );
  XOR U1490 ( .A(n1565), .B(n1566), .Z(n105) );
  AND U1491 ( .A(n1567), .B(n1568), .Z(n1566) );
  XNOR U1492 ( .A(p_input[383]), .B(n1565), .Z(n1568) );
  XOR U1493 ( .A(n1565), .B(p_input[367]), .Z(n1567) );
  XOR U1494 ( .A(n1569), .B(n1570), .Z(n1565) );
  AND U1495 ( .A(n1571), .B(n1572), .Z(n1570) );
  XNOR U1496 ( .A(p_input[382]), .B(n1569), .Z(n1572) );
  XOR U1497 ( .A(n1569), .B(p_input[366]), .Z(n1571) );
  XOR U1498 ( .A(n1573), .B(n1574), .Z(n1569) );
  AND U1499 ( .A(n1575), .B(n1576), .Z(n1574) );
  XNOR U1500 ( .A(p_input[381]), .B(n1573), .Z(n1576) );
  XOR U1501 ( .A(n1573), .B(p_input[365]), .Z(n1575) );
  XOR U1502 ( .A(n1577), .B(n1578), .Z(n1573) );
  AND U1503 ( .A(n1579), .B(n1580), .Z(n1578) );
  XNOR U1504 ( .A(p_input[380]), .B(n1577), .Z(n1580) );
  XOR U1505 ( .A(n1577), .B(p_input[364]), .Z(n1579) );
  XOR U1506 ( .A(n1581), .B(n1582), .Z(n1577) );
  AND U1507 ( .A(n1583), .B(n1584), .Z(n1582) );
  XNOR U1508 ( .A(p_input[379]), .B(n1581), .Z(n1584) );
  XOR U1509 ( .A(n1581), .B(p_input[363]), .Z(n1583) );
  XOR U1510 ( .A(n1585), .B(n1586), .Z(n1581) );
  AND U1511 ( .A(n1587), .B(n1588), .Z(n1586) );
  XNOR U1512 ( .A(p_input[378]), .B(n1585), .Z(n1588) );
  XOR U1513 ( .A(n1585), .B(p_input[362]), .Z(n1587) );
  XOR U1514 ( .A(n1589), .B(n1590), .Z(n1585) );
  AND U1515 ( .A(n1591), .B(n1592), .Z(n1590) );
  XNOR U1516 ( .A(p_input[377]), .B(n1589), .Z(n1592) );
  XOR U1517 ( .A(n1589), .B(p_input[361]), .Z(n1591) );
  XOR U1518 ( .A(n1593), .B(n1594), .Z(n1589) );
  AND U1519 ( .A(n1595), .B(n1596), .Z(n1594) );
  XNOR U1520 ( .A(p_input[376]), .B(n1593), .Z(n1596) );
  XOR U1521 ( .A(n1593), .B(p_input[360]), .Z(n1595) );
  XOR U1522 ( .A(n1597), .B(n1598), .Z(n1593) );
  AND U1523 ( .A(n1599), .B(n1600), .Z(n1598) );
  XNOR U1524 ( .A(p_input[375]), .B(n1597), .Z(n1600) );
  XOR U1525 ( .A(n1597), .B(p_input[359]), .Z(n1599) );
  XOR U1526 ( .A(n1601), .B(n1602), .Z(n1597) );
  AND U1527 ( .A(n1603), .B(n1604), .Z(n1602) );
  XNOR U1528 ( .A(p_input[374]), .B(n1601), .Z(n1604) );
  XOR U1529 ( .A(n1601), .B(p_input[358]), .Z(n1603) );
  XOR U1530 ( .A(n1605), .B(n1606), .Z(n1601) );
  AND U1531 ( .A(n1607), .B(n1608), .Z(n1606) );
  XNOR U1532 ( .A(p_input[373]), .B(n1605), .Z(n1608) );
  XOR U1533 ( .A(n1605), .B(p_input[357]), .Z(n1607) );
  XOR U1534 ( .A(n1609), .B(n1610), .Z(n1605) );
  AND U1535 ( .A(n1611), .B(n1612), .Z(n1610) );
  XNOR U1536 ( .A(p_input[372]), .B(n1609), .Z(n1612) );
  XOR U1537 ( .A(n1609), .B(p_input[356]), .Z(n1611) );
  XOR U1538 ( .A(n1613), .B(n1614), .Z(n1609) );
  AND U1539 ( .A(n1615), .B(n1616), .Z(n1614) );
  XNOR U1540 ( .A(p_input[371]), .B(n1613), .Z(n1616) );
  XOR U1541 ( .A(n1613), .B(p_input[355]), .Z(n1615) );
  XOR U1542 ( .A(n1617), .B(n1618), .Z(n1613) );
  AND U1543 ( .A(n1619), .B(n1620), .Z(n1618) );
  XNOR U1544 ( .A(p_input[370]), .B(n1617), .Z(n1620) );
  XOR U1545 ( .A(n1617), .B(p_input[354]), .Z(n1619) );
  XNOR U1546 ( .A(n1621), .B(n1622), .Z(n1617) );
  AND U1547 ( .A(n1623), .B(n1624), .Z(n1622) );
  XOR U1548 ( .A(p_input[369]), .B(n1621), .Z(n1624) );
  XNOR U1549 ( .A(p_input[353]), .B(n1621), .Z(n1623) );
  AND U1550 ( .A(p_input[368]), .B(n1625), .Z(n1621) );
  IV U1551 ( .A(p_input[352]), .Z(n1625) );
  XNOR U1552 ( .A(p_input[320]), .B(n1626), .Z(n1428) );
  AND U1553 ( .A(n103), .B(n1627), .Z(n1626) );
  XOR U1554 ( .A(p_input[336]), .B(p_input[320]), .Z(n1627) );
  XOR U1555 ( .A(n1628), .B(n1629), .Z(n103) );
  AND U1556 ( .A(n1630), .B(n1631), .Z(n1629) );
  XNOR U1557 ( .A(p_input[351]), .B(n1628), .Z(n1631) );
  XOR U1558 ( .A(n1628), .B(p_input[335]), .Z(n1630) );
  XOR U1559 ( .A(n1632), .B(n1633), .Z(n1628) );
  AND U1560 ( .A(n1634), .B(n1635), .Z(n1633) );
  XNOR U1561 ( .A(p_input[350]), .B(n1632), .Z(n1635) );
  XNOR U1562 ( .A(n1632), .B(n1442), .Z(n1634) );
  IV U1563 ( .A(p_input[334]), .Z(n1442) );
  XOR U1564 ( .A(n1636), .B(n1637), .Z(n1632) );
  AND U1565 ( .A(n1638), .B(n1639), .Z(n1637) );
  XNOR U1566 ( .A(p_input[349]), .B(n1636), .Z(n1639) );
  XNOR U1567 ( .A(n1636), .B(n1451), .Z(n1638) );
  IV U1568 ( .A(p_input[333]), .Z(n1451) );
  XOR U1569 ( .A(n1640), .B(n1641), .Z(n1636) );
  AND U1570 ( .A(n1642), .B(n1643), .Z(n1641) );
  XNOR U1571 ( .A(p_input[348]), .B(n1640), .Z(n1643) );
  XNOR U1572 ( .A(n1640), .B(n1460), .Z(n1642) );
  IV U1573 ( .A(p_input[332]), .Z(n1460) );
  XOR U1574 ( .A(n1644), .B(n1645), .Z(n1640) );
  AND U1575 ( .A(n1646), .B(n1647), .Z(n1645) );
  XNOR U1576 ( .A(p_input[347]), .B(n1644), .Z(n1647) );
  XNOR U1577 ( .A(n1644), .B(n1469), .Z(n1646) );
  IV U1578 ( .A(p_input[331]), .Z(n1469) );
  XOR U1579 ( .A(n1648), .B(n1649), .Z(n1644) );
  AND U1580 ( .A(n1650), .B(n1651), .Z(n1649) );
  XNOR U1581 ( .A(p_input[346]), .B(n1648), .Z(n1651) );
  XNOR U1582 ( .A(n1648), .B(n1478), .Z(n1650) );
  IV U1583 ( .A(p_input[330]), .Z(n1478) );
  XOR U1584 ( .A(n1652), .B(n1653), .Z(n1648) );
  AND U1585 ( .A(n1654), .B(n1655), .Z(n1653) );
  XNOR U1586 ( .A(p_input[345]), .B(n1652), .Z(n1655) );
  XNOR U1587 ( .A(n1652), .B(n1487), .Z(n1654) );
  IV U1588 ( .A(p_input[329]), .Z(n1487) );
  XOR U1589 ( .A(n1656), .B(n1657), .Z(n1652) );
  AND U1590 ( .A(n1658), .B(n1659), .Z(n1657) );
  XNOR U1591 ( .A(p_input[344]), .B(n1656), .Z(n1659) );
  XNOR U1592 ( .A(n1656), .B(n1496), .Z(n1658) );
  IV U1593 ( .A(p_input[328]), .Z(n1496) );
  XOR U1594 ( .A(n1660), .B(n1661), .Z(n1656) );
  AND U1595 ( .A(n1662), .B(n1663), .Z(n1661) );
  XNOR U1596 ( .A(p_input[343]), .B(n1660), .Z(n1663) );
  XNOR U1597 ( .A(n1660), .B(n1505), .Z(n1662) );
  IV U1598 ( .A(p_input[327]), .Z(n1505) );
  XOR U1599 ( .A(n1664), .B(n1665), .Z(n1660) );
  AND U1600 ( .A(n1666), .B(n1667), .Z(n1665) );
  XNOR U1601 ( .A(p_input[342]), .B(n1664), .Z(n1667) );
  XNOR U1602 ( .A(n1664), .B(n1514), .Z(n1666) );
  IV U1603 ( .A(p_input[326]), .Z(n1514) );
  XOR U1604 ( .A(n1668), .B(n1669), .Z(n1664) );
  AND U1605 ( .A(n1670), .B(n1671), .Z(n1669) );
  XNOR U1606 ( .A(p_input[341]), .B(n1668), .Z(n1671) );
  XNOR U1607 ( .A(n1668), .B(n1523), .Z(n1670) );
  IV U1608 ( .A(p_input[325]), .Z(n1523) );
  XOR U1609 ( .A(n1672), .B(n1673), .Z(n1668) );
  AND U1610 ( .A(n1674), .B(n1675), .Z(n1673) );
  XNOR U1611 ( .A(p_input[340]), .B(n1672), .Z(n1675) );
  XNOR U1612 ( .A(n1672), .B(n1532), .Z(n1674) );
  IV U1613 ( .A(p_input[324]), .Z(n1532) );
  XOR U1614 ( .A(n1676), .B(n1677), .Z(n1672) );
  AND U1615 ( .A(n1678), .B(n1679), .Z(n1677) );
  XNOR U1616 ( .A(p_input[339]), .B(n1676), .Z(n1679) );
  XNOR U1617 ( .A(n1676), .B(n1541), .Z(n1678) );
  IV U1618 ( .A(p_input[323]), .Z(n1541) );
  XOR U1619 ( .A(n1680), .B(n1681), .Z(n1676) );
  AND U1620 ( .A(n1682), .B(n1683), .Z(n1681) );
  XNOR U1621 ( .A(p_input[338]), .B(n1680), .Z(n1683) );
  XNOR U1622 ( .A(n1680), .B(n1550), .Z(n1682) );
  IV U1623 ( .A(p_input[322]), .Z(n1550) );
  XNOR U1624 ( .A(n1684), .B(n1685), .Z(n1680) );
  AND U1625 ( .A(n1686), .B(n1687), .Z(n1685) );
  XOR U1626 ( .A(p_input[337]), .B(n1684), .Z(n1687) );
  XNOR U1627 ( .A(p_input[321]), .B(n1684), .Z(n1686) );
  AND U1628 ( .A(p_input[336]), .B(n1688), .Z(n1684) );
  IV U1629 ( .A(p_input[320]), .Z(n1688) );
  XOR U1630 ( .A(n1689), .B(n1690), .Z(n1247) );
  AND U1631 ( .A(n122), .B(n1691), .Z(n1690) );
  XNOR U1632 ( .A(n1692), .B(n1689), .Z(n1691) );
  XOR U1633 ( .A(n1693), .B(n1694), .Z(n122) );
  AND U1634 ( .A(n1695), .B(n1696), .Z(n1694) );
  XNOR U1635 ( .A(n1258), .B(n1693), .Z(n1696) );
  AND U1636 ( .A(p_input[319]), .B(p_input[303]), .Z(n1258) );
  XOR U1637 ( .A(n1693), .B(n1257), .Z(n1695) );
  AND U1638 ( .A(p_input[271]), .B(p_input[287]), .Z(n1257) );
  XOR U1639 ( .A(n1697), .B(n1698), .Z(n1693) );
  AND U1640 ( .A(n1699), .B(n1700), .Z(n1698) );
  XOR U1641 ( .A(n1697), .B(n1270), .Z(n1700) );
  XNOR U1642 ( .A(p_input[302]), .B(n1701), .Z(n1270) );
  AND U1643 ( .A(n109), .B(n1702), .Z(n1701) );
  XOR U1644 ( .A(p_input[318]), .B(p_input[302]), .Z(n1702) );
  XNOR U1645 ( .A(n1267), .B(n1697), .Z(n1699) );
  XOR U1646 ( .A(n1703), .B(n1704), .Z(n1267) );
  AND U1647 ( .A(n106), .B(n1705), .Z(n1704) );
  XOR U1648 ( .A(p_input[286]), .B(p_input[270]), .Z(n1705) );
  XOR U1649 ( .A(n1706), .B(n1707), .Z(n1697) );
  AND U1650 ( .A(n1708), .B(n1709), .Z(n1707) );
  XOR U1651 ( .A(n1706), .B(n1282), .Z(n1709) );
  XNOR U1652 ( .A(p_input[301]), .B(n1710), .Z(n1282) );
  AND U1653 ( .A(n109), .B(n1711), .Z(n1710) );
  XOR U1654 ( .A(p_input[317]), .B(p_input[301]), .Z(n1711) );
  XNOR U1655 ( .A(n1279), .B(n1706), .Z(n1708) );
  XOR U1656 ( .A(n1712), .B(n1713), .Z(n1279) );
  AND U1657 ( .A(n106), .B(n1714), .Z(n1713) );
  XOR U1658 ( .A(p_input[285]), .B(p_input[269]), .Z(n1714) );
  XOR U1659 ( .A(n1715), .B(n1716), .Z(n1706) );
  AND U1660 ( .A(n1717), .B(n1718), .Z(n1716) );
  XOR U1661 ( .A(n1715), .B(n1294), .Z(n1718) );
  XNOR U1662 ( .A(p_input[300]), .B(n1719), .Z(n1294) );
  AND U1663 ( .A(n109), .B(n1720), .Z(n1719) );
  XOR U1664 ( .A(p_input[316]), .B(p_input[300]), .Z(n1720) );
  XNOR U1665 ( .A(n1291), .B(n1715), .Z(n1717) );
  XOR U1666 ( .A(n1721), .B(n1722), .Z(n1291) );
  AND U1667 ( .A(n106), .B(n1723), .Z(n1722) );
  XOR U1668 ( .A(p_input[284]), .B(p_input[268]), .Z(n1723) );
  XOR U1669 ( .A(n1724), .B(n1725), .Z(n1715) );
  AND U1670 ( .A(n1726), .B(n1727), .Z(n1725) );
  XOR U1671 ( .A(n1724), .B(n1306), .Z(n1727) );
  XNOR U1672 ( .A(p_input[299]), .B(n1728), .Z(n1306) );
  AND U1673 ( .A(n109), .B(n1729), .Z(n1728) );
  XOR U1674 ( .A(p_input[315]), .B(p_input[299]), .Z(n1729) );
  XNOR U1675 ( .A(n1303), .B(n1724), .Z(n1726) );
  XOR U1676 ( .A(n1730), .B(n1731), .Z(n1303) );
  AND U1677 ( .A(n106), .B(n1732), .Z(n1731) );
  XOR U1678 ( .A(p_input[283]), .B(p_input[267]), .Z(n1732) );
  XOR U1679 ( .A(n1733), .B(n1734), .Z(n1724) );
  AND U1680 ( .A(n1735), .B(n1736), .Z(n1734) );
  XOR U1681 ( .A(n1733), .B(n1318), .Z(n1736) );
  XNOR U1682 ( .A(p_input[298]), .B(n1737), .Z(n1318) );
  AND U1683 ( .A(n109), .B(n1738), .Z(n1737) );
  XOR U1684 ( .A(p_input[314]), .B(p_input[298]), .Z(n1738) );
  XNOR U1685 ( .A(n1315), .B(n1733), .Z(n1735) );
  XOR U1686 ( .A(n1739), .B(n1740), .Z(n1315) );
  AND U1687 ( .A(n106), .B(n1741), .Z(n1740) );
  XOR U1688 ( .A(p_input[282]), .B(p_input[266]), .Z(n1741) );
  XOR U1689 ( .A(n1742), .B(n1743), .Z(n1733) );
  AND U1690 ( .A(n1744), .B(n1745), .Z(n1743) );
  XOR U1691 ( .A(n1742), .B(n1330), .Z(n1745) );
  XNOR U1692 ( .A(p_input[297]), .B(n1746), .Z(n1330) );
  AND U1693 ( .A(n109), .B(n1747), .Z(n1746) );
  XOR U1694 ( .A(p_input[313]), .B(p_input[297]), .Z(n1747) );
  XNOR U1695 ( .A(n1327), .B(n1742), .Z(n1744) );
  XOR U1696 ( .A(n1748), .B(n1749), .Z(n1327) );
  AND U1697 ( .A(n106), .B(n1750), .Z(n1749) );
  XOR U1698 ( .A(p_input[281]), .B(p_input[265]), .Z(n1750) );
  XOR U1699 ( .A(n1751), .B(n1752), .Z(n1742) );
  AND U1700 ( .A(n1753), .B(n1754), .Z(n1752) );
  XOR U1701 ( .A(n1751), .B(n1342), .Z(n1754) );
  XNOR U1702 ( .A(p_input[296]), .B(n1755), .Z(n1342) );
  AND U1703 ( .A(n109), .B(n1756), .Z(n1755) );
  XOR U1704 ( .A(p_input[312]), .B(p_input[296]), .Z(n1756) );
  XNOR U1705 ( .A(n1339), .B(n1751), .Z(n1753) );
  XOR U1706 ( .A(n1757), .B(n1758), .Z(n1339) );
  AND U1707 ( .A(n106), .B(n1759), .Z(n1758) );
  XOR U1708 ( .A(p_input[280]), .B(p_input[264]), .Z(n1759) );
  XOR U1709 ( .A(n1760), .B(n1761), .Z(n1751) );
  AND U1710 ( .A(n1762), .B(n1763), .Z(n1761) );
  XOR U1711 ( .A(n1760), .B(n1354), .Z(n1763) );
  XNOR U1712 ( .A(p_input[295]), .B(n1764), .Z(n1354) );
  AND U1713 ( .A(n109), .B(n1765), .Z(n1764) );
  XOR U1714 ( .A(p_input[311]), .B(p_input[295]), .Z(n1765) );
  XNOR U1715 ( .A(n1351), .B(n1760), .Z(n1762) );
  XOR U1716 ( .A(n1766), .B(n1767), .Z(n1351) );
  AND U1717 ( .A(n106), .B(n1768), .Z(n1767) );
  XOR U1718 ( .A(p_input[279]), .B(p_input[263]), .Z(n1768) );
  XOR U1719 ( .A(n1769), .B(n1770), .Z(n1760) );
  AND U1720 ( .A(n1771), .B(n1772), .Z(n1770) );
  XOR U1721 ( .A(n1769), .B(n1366), .Z(n1772) );
  XNOR U1722 ( .A(p_input[294]), .B(n1773), .Z(n1366) );
  AND U1723 ( .A(n109), .B(n1774), .Z(n1773) );
  XOR U1724 ( .A(p_input[310]), .B(p_input[294]), .Z(n1774) );
  XNOR U1725 ( .A(n1363), .B(n1769), .Z(n1771) );
  XOR U1726 ( .A(n1775), .B(n1776), .Z(n1363) );
  AND U1727 ( .A(n106), .B(n1777), .Z(n1776) );
  XOR U1728 ( .A(p_input[278]), .B(p_input[262]), .Z(n1777) );
  XOR U1729 ( .A(n1778), .B(n1779), .Z(n1769) );
  AND U1730 ( .A(n1780), .B(n1781), .Z(n1779) );
  XOR U1731 ( .A(n1778), .B(n1378), .Z(n1781) );
  XNOR U1732 ( .A(p_input[293]), .B(n1782), .Z(n1378) );
  AND U1733 ( .A(n109), .B(n1783), .Z(n1782) );
  XOR U1734 ( .A(p_input[309]), .B(p_input[293]), .Z(n1783) );
  XNOR U1735 ( .A(n1375), .B(n1778), .Z(n1780) );
  XOR U1736 ( .A(n1784), .B(n1785), .Z(n1375) );
  AND U1737 ( .A(n106), .B(n1786), .Z(n1785) );
  XOR U1738 ( .A(p_input[277]), .B(p_input[261]), .Z(n1786) );
  XOR U1739 ( .A(n1787), .B(n1788), .Z(n1778) );
  AND U1740 ( .A(n1789), .B(n1790), .Z(n1788) );
  XOR U1741 ( .A(n1390), .B(n1787), .Z(n1790) );
  XNOR U1742 ( .A(p_input[292]), .B(n1791), .Z(n1390) );
  AND U1743 ( .A(n109), .B(n1792), .Z(n1791) );
  XOR U1744 ( .A(p_input[308]), .B(p_input[292]), .Z(n1792) );
  XNOR U1745 ( .A(n1787), .B(n1387), .Z(n1789) );
  XOR U1746 ( .A(n1793), .B(n1794), .Z(n1387) );
  AND U1747 ( .A(n106), .B(n1795), .Z(n1794) );
  XOR U1748 ( .A(p_input[276]), .B(p_input[260]), .Z(n1795) );
  XOR U1749 ( .A(n1796), .B(n1797), .Z(n1787) );
  AND U1750 ( .A(n1798), .B(n1799), .Z(n1797) );
  XOR U1751 ( .A(n1796), .B(n1402), .Z(n1799) );
  XNOR U1752 ( .A(p_input[291]), .B(n1800), .Z(n1402) );
  AND U1753 ( .A(n109), .B(n1801), .Z(n1800) );
  XOR U1754 ( .A(p_input[307]), .B(p_input[291]), .Z(n1801) );
  XNOR U1755 ( .A(n1399), .B(n1796), .Z(n1798) );
  XOR U1756 ( .A(n1802), .B(n1803), .Z(n1399) );
  AND U1757 ( .A(n106), .B(n1804), .Z(n1803) );
  XOR U1758 ( .A(p_input[275]), .B(p_input[259]), .Z(n1804) );
  XOR U1759 ( .A(n1805), .B(n1806), .Z(n1796) );
  AND U1760 ( .A(n1807), .B(n1808), .Z(n1806) );
  XOR U1761 ( .A(n1805), .B(n1414), .Z(n1808) );
  XNOR U1762 ( .A(p_input[290]), .B(n1809), .Z(n1414) );
  AND U1763 ( .A(n109), .B(n1810), .Z(n1809) );
  XOR U1764 ( .A(p_input[306]), .B(p_input[290]), .Z(n1810) );
  XNOR U1765 ( .A(n1411), .B(n1805), .Z(n1807) );
  XOR U1766 ( .A(n1811), .B(n1812), .Z(n1411) );
  AND U1767 ( .A(n106), .B(n1813), .Z(n1812) );
  XOR U1768 ( .A(p_input[274]), .B(p_input[258]), .Z(n1813) );
  XOR U1769 ( .A(n1814), .B(n1815), .Z(n1805) );
  AND U1770 ( .A(n1816), .B(n1817), .Z(n1815) );
  XNOR U1771 ( .A(n1818), .B(n1427), .Z(n1817) );
  XNOR U1772 ( .A(p_input[289]), .B(n1819), .Z(n1427) );
  AND U1773 ( .A(n109), .B(n1820), .Z(n1819) );
  XNOR U1774 ( .A(p_input[305]), .B(n1821), .Z(n1820) );
  IV U1775 ( .A(p_input[289]), .Z(n1821) );
  XNOR U1776 ( .A(n1424), .B(n1814), .Z(n1816) );
  XNOR U1777 ( .A(p_input[257]), .B(n1822), .Z(n1424) );
  AND U1778 ( .A(n106), .B(n1823), .Z(n1822) );
  XOR U1779 ( .A(p_input[273]), .B(p_input[257]), .Z(n1823) );
  IV U1780 ( .A(n1818), .Z(n1814) );
  AND U1781 ( .A(n1689), .B(n1692), .Z(n1818) );
  XOR U1782 ( .A(p_input[288]), .B(n1824), .Z(n1692) );
  AND U1783 ( .A(n109), .B(n1825), .Z(n1824) );
  XOR U1784 ( .A(p_input[304]), .B(p_input[288]), .Z(n1825) );
  XOR U1785 ( .A(n1826), .B(n1827), .Z(n109) );
  AND U1786 ( .A(n1828), .B(n1829), .Z(n1827) );
  XNOR U1787 ( .A(p_input[319]), .B(n1826), .Z(n1829) );
  XOR U1788 ( .A(n1826), .B(p_input[303]), .Z(n1828) );
  XOR U1789 ( .A(n1830), .B(n1831), .Z(n1826) );
  AND U1790 ( .A(n1832), .B(n1833), .Z(n1831) );
  XNOR U1791 ( .A(p_input[318]), .B(n1830), .Z(n1833) );
  XOR U1792 ( .A(n1830), .B(p_input[302]), .Z(n1832) );
  XOR U1793 ( .A(n1834), .B(n1835), .Z(n1830) );
  AND U1794 ( .A(n1836), .B(n1837), .Z(n1835) );
  XNOR U1795 ( .A(p_input[317]), .B(n1834), .Z(n1837) );
  XOR U1796 ( .A(n1834), .B(p_input[301]), .Z(n1836) );
  XOR U1797 ( .A(n1838), .B(n1839), .Z(n1834) );
  AND U1798 ( .A(n1840), .B(n1841), .Z(n1839) );
  XNOR U1799 ( .A(p_input[316]), .B(n1838), .Z(n1841) );
  XOR U1800 ( .A(n1838), .B(p_input[300]), .Z(n1840) );
  XOR U1801 ( .A(n1842), .B(n1843), .Z(n1838) );
  AND U1802 ( .A(n1844), .B(n1845), .Z(n1843) );
  XNOR U1803 ( .A(p_input[315]), .B(n1842), .Z(n1845) );
  XOR U1804 ( .A(n1842), .B(p_input[299]), .Z(n1844) );
  XOR U1805 ( .A(n1846), .B(n1847), .Z(n1842) );
  AND U1806 ( .A(n1848), .B(n1849), .Z(n1847) );
  XNOR U1807 ( .A(p_input[314]), .B(n1846), .Z(n1849) );
  XOR U1808 ( .A(n1846), .B(p_input[298]), .Z(n1848) );
  XOR U1809 ( .A(n1850), .B(n1851), .Z(n1846) );
  AND U1810 ( .A(n1852), .B(n1853), .Z(n1851) );
  XNOR U1811 ( .A(p_input[313]), .B(n1850), .Z(n1853) );
  XOR U1812 ( .A(n1850), .B(p_input[297]), .Z(n1852) );
  XOR U1813 ( .A(n1854), .B(n1855), .Z(n1850) );
  AND U1814 ( .A(n1856), .B(n1857), .Z(n1855) );
  XNOR U1815 ( .A(p_input[312]), .B(n1854), .Z(n1857) );
  XOR U1816 ( .A(n1854), .B(p_input[296]), .Z(n1856) );
  XOR U1817 ( .A(n1858), .B(n1859), .Z(n1854) );
  AND U1818 ( .A(n1860), .B(n1861), .Z(n1859) );
  XNOR U1819 ( .A(p_input[311]), .B(n1858), .Z(n1861) );
  XOR U1820 ( .A(n1858), .B(p_input[295]), .Z(n1860) );
  XOR U1821 ( .A(n1862), .B(n1863), .Z(n1858) );
  AND U1822 ( .A(n1864), .B(n1865), .Z(n1863) );
  XNOR U1823 ( .A(p_input[310]), .B(n1862), .Z(n1865) );
  XOR U1824 ( .A(n1862), .B(p_input[294]), .Z(n1864) );
  XOR U1825 ( .A(n1866), .B(n1867), .Z(n1862) );
  AND U1826 ( .A(n1868), .B(n1869), .Z(n1867) );
  XNOR U1827 ( .A(p_input[309]), .B(n1866), .Z(n1869) );
  XOR U1828 ( .A(n1866), .B(p_input[293]), .Z(n1868) );
  XOR U1829 ( .A(n1870), .B(n1871), .Z(n1866) );
  AND U1830 ( .A(n1872), .B(n1873), .Z(n1871) );
  XNOR U1831 ( .A(p_input[308]), .B(n1870), .Z(n1873) );
  XOR U1832 ( .A(n1870), .B(p_input[292]), .Z(n1872) );
  XOR U1833 ( .A(n1874), .B(n1875), .Z(n1870) );
  AND U1834 ( .A(n1876), .B(n1877), .Z(n1875) );
  XNOR U1835 ( .A(p_input[307]), .B(n1874), .Z(n1877) );
  XOR U1836 ( .A(n1874), .B(p_input[291]), .Z(n1876) );
  XOR U1837 ( .A(n1878), .B(n1879), .Z(n1874) );
  AND U1838 ( .A(n1880), .B(n1881), .Z(n1879) );
  XNOR U1839 ( .A(p_input[306]), .B(n1878), .Z(n1881) );
  XOR U1840 ( .A(n1878), .B(p_input[290]), .Z(n1880) );
  XNOR U1841 ( .A(n1882), .B(n1883), .Z(n1878) );
  AND U1842 ( .A(n1884), .B(n1885), .Z(n1883) );
  XOR U1843 ( .A(p_input[305]), .B(n1882), .Z(n1885) );
  XNOR U1844 ( .A(p_input[289]), .B(n1882), .Z(n1884) );
  AND U1845 ( .A(p_input[304]), .B(n1886), .Z(n1882) );
  IV U1846 ( .A(p_input[288]), .Z(n1886) );
  XNOR U1847 ( .A(p_input[256]), .B(n1887), .Z(n1689) );
  AND U1848 ( .A(n106), .B(n1888), .Z(n1887) );
  XOR U1849 ( .A(p_input[272]), .B(p_input[256]), .Z(n1888) );
  XOR U1850 ( .A(n1889), .B(n1890), .Z(n106) );
  AND U1851 ( .A(n1891), .B(n1892), .Z(n1890) );
  XNOR U1852 ( .A(p_input[287]), .B(n1889), .Z(n1892) );
  XOR U1853 ( .A(n1889), .B(p_input[271]), .Z(n1891) );
  XOR U1854 ( .A(n1893), .B(n1894), .Z(n1889) );
  AND U1855 ( .A(n1895), .B(n1896), .Z(n1894) );
  XNOR U1856 ( .A(p_input[286]), .B(n1893), .Z(n1896) );
  XNOR U1857 ( .A(n1893), .B(n1703), .Z(n1895) );
  IV U1858 ( .A(p_input[270]), .Z(n1703) );
  XOR U1859 ( .A(n1897), .B(n1898), .Z(n1893) );
  AND U1860 ( .A(n1899), .B(n1900), .Z(n1898) );
  XNOR U1861 ( .A(p_input[285]), .B(n1897), .Z(n1900) );
  XNOR U1862 ( .A(n1897), .B(n1712), .Z(n1899) );
  IV U1863 ( .A(p_input[269]), .Z(n1712) );
  XOR U1864 ( .A(n1901), .B(n1902), .Z(n1897) );
  AND U1865 ( .A(n1903), .B(n1904), .Z(n1902) );
  XNOR U1866 ( .A(p_input[284]), .B(n1901), .Z(n1904) );
  XNOR U1867 ( .A(n1901), .B(n1721), .Z(n1903) );
  IV U1868 ( .A(p_input[268]), .Z(n1721) );
  XOR U1869 ( .A(n1905), .B(n1906), .Z(n1901) );
  AND U1870 ( .A(n1907), .B(n1908), .Z(n1906) );
  XNOR U1871 ( .A(p_input[283]), .B(n1905), .Z(n1908) );
  XNOR U1872 ( .A(n1905), .B(n1730), .Z(n1907) );
  IV U1873 ( .A(p_input[267]), .Z(n1730) );
  XOR U1874 ( .A(n1909), .B(n1910), .Z(n1905) );
  AND U1875 ( .A(n1911), .B(n1912), .Z(n1910) );
  XNOR U1876 ( .A(p_input[282]), .B(n1909), .Z(n1912) );
  XNOR U1877 ( .A(n1909), .B(n1739), .Z(n1911) );
  IV U1878 ( .A(p_input[266]), .Z(n1739) );
  XOR U1879 ( .A(n1913), .B(n1914), .Z(n1909) );
  AND U1880 ( .A(n1915), .B(n1916), .Z(n1914) );
  XNOR U1881 ( .A(p_input[281]), .B(n1913), .Z(n1916) );
  XNOR U1882 ( .A(n1913), .B(n1748), .Z(n1915) );
  IV U1883 ( .A(p_input[265]), .Z(n1748) );
  XOR U1884 ( .A(n1917), .B(n1918), .Z(n1913) );
  AND U1885 ( .A(n1919), .B(n1920), .Z(n1918) );
  XNOR U1886 ( .A(p_input[280]), .B(n1917), .Z(n1920) );
  XNOR U1887 ( .A(n1917), .B(n1757), .Z(n1919) );
  IV U1888 ( .A(p_input[264]), .Z(n1757) );
  XOR U1889 ( .A(n1921), .B(n1922), .Z(n1917) );
  AND U1890 ( .A(n1923), .B(n1924), .Z(n1922) );
  XNOR U1891 ( .A(p_input[279]), .B(n1921), .Z(n1924) );
  XNOR U1892 ( .A(n1921), .B(n1766), .Z(n1923) );
  IV U1893 ( .A(p_input[263]), .Z(n1766) );
  XOR U1894 ( .A(n1925), .B(n1926), .Z(n1921) );
  AND U1895 ( .A(n1927), .B(n1928), .Z(n1926) );
  XNOR U1896 ( .A(p_input[278]), .B(n1925), .Z(n1928) );
  XNOR U1897 ( .A(n1925), .B(n1775), .Z(n1927) );
  IV U1898 ( .A(p_input[262]), .Z(n1775) );
  XOR U1899 ( .A(n1929), .B(n1930), .Z(n1925) );
  AND U1900 ( .A(n1931), .B(n1932), .Z(n1930) );
  XNOR U1901 ( .A(p_input[277]), .B(n1929), .Z(n1932) );
  XNOR U1902 ( .A(n1929), .B(n1784), .Z(n1931) );
  IV U1903 ( .A(p_input[261]), .Z(n1784) );
  XOR U1904 ( .A(n1933), .B(n1934), .Z(n1929) );
  AND U1905 ( .A(n1935), .B(n1936), .Z(n1934) );
  XNOR U1906 ( .A(p_input[276]), .B(n1933), .Z(n1936) );
  XNOR U1907 ( .A(n1933), .B(n1793), .Z(n1935) );
  IV U1908 ( .A(p_input[260]), .Z(n1793) );
  XOR U1909 ( .A(n1937), .B(n1938), .Z(n1933) );
  AND U1910 ( .A(n1939), .B(n1940), .Z(n1938) );
  XNOR U1911 ( .A(p_input[275]), .B(n1937), .Z(n1940) );
  XNOR U1912 ( .A(n1937), .B(n1802), .Z(n1939) );
  IV U1913 ( .A(p_input[259]), .Z(n1802) );
  XOR U1914 ( .A(n1941), .B(n1942), .Z(n1937) );
  AND U1915 ( .A(n1943), .B(n1944), .Z(n1942) );
  XNOR U1916 ( .A(p_input[274]), .B(n1941), .Z(n1944) );
  XNOR U1917 ( .A(n1941), .B(n1811), .Z(n1943) );
  IV U1918 ( .A(p_input[258]), .Z(n1811) );
  XNOR U1919 ( .A(n1945), .B(n1946), .Z(n1941) );
  AND U1920 ( .A(n1947), .B(n1948), .Z(n1946) );
  XOR U1921 ( .A(p_input[273]), .B(n1945), .Z(n1948) );
  XNOR U1922 ( .A(p_input[257]), .B(n1945), .Z(n1947) );
  AND U1923 ( .A(p_input[272]), .B(n1949), .Z(n1945) );
  IV U1924 ( .A(p_input[256]), .Z(n1949) );
  XOR U1925 ( .A(n1950), .B(n1951), .Z(n21) );
  AND U1926 ( .A(n174), .B(n1952), .Z(n1951) );
  XNOR U1927 ( .A(n1953), .B(n1950), .Z(n1952) );
  XOR U1928 ( .A(n1954), .B(n1955), .Z(n174) );
  AND U1929 ( .A(n1956), .B(n1957), .Z(n1955) );
  XNOR U1930 ( .A(n193), .B(n1954), .Z(n1957) );
  AND U1931 ( .A(n1958), .B(n1959), .Z(n193) );
  XNOR U1932 ( .A(n1954), .B(n190), .Z(n1956) );
  IV U1933 ( .A(n1960), .Z(n190) );
  AND U1934 ( .A(n1961), .B(n1962), .Z(n1960) );
  XOR U1935 ( .A(n1963), .B(n1964), .Z(n1954) );
  AND U1936 ( .A(n1965), .B(n1966), .Z(n1964) );
  XOR U1937 ( .A(n1963), .B(n205), .Z(n1966) );
  XOR U1938 ( .A(n1967), .B(n1968), .Z(n205) );
  AND U1939 ( .A(n165), .B(n1969), .Z(n1968) );
  XOR U1940 ( .A(n1970), .B(n1967), .Z(n1969) );
  XNOR U1941 ( .A(n202), .B(n1963), .Z(n1965) );
  XOR U1942 ( .A(n1971), .B(n1972), .Z(n202) );
  AND U1943 ( .A(n162), .B(n1973), .Z(n1972) );
  XOR U1944 ( .A(n1974), .B(n1971), .Z(n1973) );
  XOR U1945 ( .A(n1975), .B(n1976), .Z(n1963) );
  AND U1946 ( .A(n1977), .B(n1978), .Z(n1976) );
  XOR U1947 ( .A(n1975), .B(n217), .Z(n1978) );
  XOR U1948 ( .A(n1979), .B(n1980), .Z(n217) );
  AND U1949 ( .A(n165), .B(n1981), .Z(n1980) );
  XOR U1950 ( .A(n1982), .B(n1979), .Z(n1981) );
  XNOR U1951 ( .A(n214), .B(n1975), .Z(n1977) );
  XOR U1952 ( .A(n1983), .B(n1984), .Z(n214) );
  AND U1953 ( .A(n162), .B(n1985), .Z(n1984) );
  XOR U1954 ( .A(n1986), .B(n1983), .Z(n1985) );
  XOR U1955 ( .A(n1987), .B(n1988), .Z(n1975) );
  AND U1956 ( .A(n1989), .B(n1990), .Z(n1988) );
  XOR U1957 ( .A(n1987), .B(n229), .Z(n1990) );
  XOR U1958 ( .A(n1991), .B(n1992), .Z(n229) );
  AND U1959 ( .A(n165), .B(n1993), .Z(n1992) );
  XOR U1960 ( .A(n1994), .B(n1991), .Z(n1993) );
  XNOR U1961 ( .A(n226), .B(n1987), .Z(n1989) );
  XOR U1962 ( .A(n1995), .B(n1996), .Z(n226) );
  AND U1963 ( .A(n162), .B(n1997), .Z(n1996) );
  XOR U1964 ( .A(n1998), .B(n1995), .Z(n1997) );
  XOR U1965 ( .A(n1999), .B(n2000), .Z(n1987) );
  AND U1966 ( .A(n2001), .B(n2002), .Z(n2000) );
  XOR U1967 ( .A(n1999), .B(n241), .Z(n2002) );
  XOR U1968 ( .A(n2003), .B(n2004), .Z(n241) );
  AND U1969 ( .A(n165), .B(n2005), .Z(n2004) );
  XOR U1970 ( .A(n2006), .B(n2003), .Z(n2005) );
  XNOR U1971 ( .A(n238), .B(n1999), .Z(n2001) );
  XOR U1972 ( .A(n2007), .B(n2008), .Z(n238) );
  AND U1973 ( .A(n162), .B(n2009), .Z(n2008) );
  XOR U1974 ( .A(n2010), .B(n2007), .Z(n2009) );
  XOR U1975 ( .A(n2011), .B(n2012), .Z(n1999) );
  AND U1976 ( .A(n2013), .B(n2014), .Z(n2012) );
  XOR U1977 ( .A(n2011), .B(n253), .Z(n2014) );
  XOR U1978 ( .A(n2015), .B(n2016), .Z(n253) );
  AND U1979 ( .A(n165), .B(n2017), .Z(n2016) );
  XOR U1980 ( .A(n2018), .B(n2015), .Z(n2017) );
  XNOR U1981 ( .A(n250), .B(n2011), .Z(n2013) );
  XOR U1982 ( .A(n2019), .B(n2020), .Z(n250) );
  AND U1983 ( .A(n162), .B(n2021), .Z(n2020) );
  XOR U1984 ( .A(n2022), .B(n2019), .Z(n2021) );
  XOR U1985 ( .A(n2023), .B(n2024), .Z(n2011) );
  AND U1986 ( .A(n2025), .B(n2026), .Z(n2024) );
  XOR U1987 ( .A(n2023), .B(n265), .Z(n2026) );
  XOR U1988 ( .A(n2027), .B(n2028), .Z(n265) );
  AND U1989 ( .A(n165), .B(n2029), .Z(n2028) );
  XOR U1990 ( .A(n2030), .B(n2027), .Z(n2029) );
  XNOR U1991 ( .A(n262), .B(n2023), .Z(n2025) );
  XOR U1992 ( .A(n2031), .B(n2032), .Z(n262) );
  AND U1993 ( .A(n162), .B(n2033), .Z(n2032) );
  XOR U1994 ( .A(n2034), .B(n2031), .Z(n2033) );
  XOR U1995 ( .A(n2035), .B(n2036), .Z(n2023) );
  AND U1996 ( .A(n2037), .B(n2038), .Z(n2036) );
  XOR U1997 ( .A(n2035), .B(n277), .Z(n2038) );
  XOR U1998 ( .A(n2039), .B(n2040), .Z(n277) );
  AND U1999 ( .A(n165), .B(n2041), .Z(n2040) );
  XOR U2000 ( .A(n2042), .B(n2039), .Z(n2041) );
  XNOR U2001 ( .A(n274), .B(n2035), .Z(n2037) );
  XOR U2002 ( .A(n2043), .B(n2044), .Z(n274) );
  AND U2003 ( .A(n162), .B(n2045), .Z(n2044) );
  XOR U2004 ( .A(n2046), .B(n2043), .Z(n2045) );
  XOR U2005 ( .A(n2047), .B(n2048), .Z(n2035) );
  AND U2006 ( .A(n2049), .B(n2050), .Z(n2048) );
  XOR U2007 ( .A(n2047), .B(n289), .Z(n2050) );
  XOR U2008 ( .A(n2051), .B(n2052), .Z(n289) );
  AND U2009 ( .A(n165), .B(n2053), .Z(n2052) );
  XOR U2010 ( .A(n2054), .B(n2051), .Z(n2053) );
  XNOR U2011 ( .A(n286), .B(n2047), .Z(n2049) );
  XOR U2012 ( .A(n2055), .B(n2056), .Z(n286) );
  AND U2013 ( .A(n162), .B(n2057), .Z(n2056) );
  XOR U2014 ( .A(n2058), .B(n2055), .Z(n2057) );
  XOR U2015 ( .A(n2059), .B(n2060), .Z(n2047) );
  AND U2016 ( .A(n2061), .B(n2062), .Z(n2060) );
  XOR U2017 ( .A(n2059), .B(n301), .Z(n2062) );
  XOR U2018 ( .A(n2063), .B(n2064), .Z(n301) );
  AND U2019 ( .A(n165), .B(n2065), .Z(n2064) );
  XOR U2020 ( .A(n2066), .B(n2063), .Z(n2065) );
  XNOR U2021 ( .A(n298), .B(n2059), .Z(n2061) );
  XOR U2022 ( .A(n2067), .B(n2068), .Z(n298) );
  AND U2023 ( .A(n162), .B(n2069), .Z(n2068) );
  XOR U2024 ( .A(n2070), .B(n2067), .Z(n2069) );
  XOR U2025 ( .A(n2071), .B(n2072), .Z(n2059) );
  AND U2026 ( .A(n2073), .B(n2074), .Z(n2072) );
  XOR U2027 ( .A(n2071), .B(n313), .Z(n2074) );
  XOR U2028 ( .A(n2075), .B(n2076), .Z(n313) );
  AND U2029 ( .A(n165), .B(n2077), .Z(n2076) );
  XOR U2030 ( .A(n2078), .B(n2075), .Z(n2077) );
  XNOR U2031 ( .A(n310), .B(n2071), .Z(n2073) );
  XOR U2032 ( .A(n2079), .B(n2080), .Z(n310) );
  AND U2033 ( .A(n162), .B(n2081), .Z(n2080) );
  XOR U2034 ( .A(n2082), .B(n2079), .Z(n2081) );
  XOR U2035 ( .A(n2083), .B(n2084), .Z(n2071) );
  AND U2036 ( .A(n2085), .B(n2086), .Z(n2084) );
  XOR U2037 ( .A(n325), .B(n2083), .Z(n2086) );
  XOR U2038 ( .A(n2087), .B(n2088), .Z(n325) );
  AND U2039 ( .A(n165), .B(n2089), .Z(n2088) );
  XOR U2040 ( .A(n2087), .B(n2090), .Z(n2089) );
  XNOR U2041 ( .A(n2083), .B(n322), .Z(n2085) );
  XOR U2042 ( .A(n2091), .B(n2092), .Z(n322) );
  AND U2043 ( .A(n162), .B(n2093), .Z(n2092) );
  XOR U2044 ( .A(n2091), .B(n2094), .Z(n2093) );
  XOR U2045 ( .A(n2095), .B(n2096), .Z(n2083) );
  AND U2046 ( .A(n2097), .B(n2098), .Z(n2096) );
  XOR U2047 ( .A(n2095), .B(n337), .Z(n2098) );
  XOR U2048 ( .A(n2099), .B(n2100), .Z(n337) );
  AND U2049 ( .A(n165), .B(n2101), .Z(n2100) );
  XOR U2050 ( .A(n2102), .B(n2099), .Z(n2101) );
  XNOR U2051 ( .A(n334), .B(n2095), .Z(n2097) );
  XOR U2052 ( .A(n2103), .B(n2104), .Z(n334) );
  AND U2053 ( .A(n162), .B(n2105), .Z(n2104) );
  XOR U2054 ( .A(n2106), .B(n2103), .Z(n2105) );
  XOR U2055 ( .A(n2107), .B(n2108), .Z(n2095) );
  AND U2056 ( .A(n2109), .B(n2110), .Z(n2108) );
  XOR U2057 ( .A(n2107), .B(n349), .Z(n2110) );
  XOR U2058 ( .A(n2111), .B(n2112), .Z(n349) );
  AND U2059 ( .A(n165), .B(n2113), .Z(n2112) );
  XOR U2060 ( .A(n2114), .B(n2111), .Z(n2113) );
  XNOR U2061 ( .A(n346), .B(n2107), .Z(n2109) );
  XOR U2062 ( .A(n2115), .B(n2116), .Z(n346) );
  AND U2063 ( .A(n162), .B(n2117), .Z(n2116) );
  XOR U2064 ( .A(n2118), .B(n2115), .Z(n2117) );
  XOR U2065 ( .A(n2119), .B(n2120), .Z(n2107) );
  AND U2066 ( .A(n2121), .B(n2122), .Z(n2120) );
  XNOR U2067 ( .A(n2123), .B(n361), .Z(n2122) );
  XOR U2068 ( .A(n2124), .B(n2125), .Z(n361) );
  AND U2069 ( .A(n165), .B(n2126), .Z(n2125) );
  XOR U2070 ( .A(n2127), .B(n2124), .Z(n2126) );
  XNOR U2071 ( .A(n358), .B(n2119), .Z(n2121) );
  XOR U2072 ( .A(n2128), .B(n2129), .Z(n358) );
  AND U2073 ( .A(n162), .B(n2130), .Z(n2129) );
  XOR U2074 ( .A(n2131), .B(n2128), .Z(n2130) );
  IV U2075 ( .A(n2123), .Z(n2119) );
  AND U2076 ( .A(n1950), .B(n1953), .Z(n2123) );
  XNOR U2077 ( .A(n2132), .B(n2133), .Z(n1953) );
  AND U2078 ( .A(n165), .B(n2134), .Z(n2133) );
  XNOR U2079 ( .A(n2135), .B(n2132), .Z(n2134) );
  XOR U2080 ( .A(n2136), .B(n2137), .Z(n165) );
  AND U2081 ( .A(n2138), .B(n2139), .Z(n2137) );
  XNOR U2082 ( .A(n1958), .B(n2136), .Z(n2139) );
  AND U2083 ( .A(n2140), .B(n2141), .Z(n1958) );
  XOR U2084 ( .A(n2136), .B(n1959), .Z(n2138) );
  AND U2085 ( .A(n2142), .B(n2143), .Z(n1959) );
  XOR U2086 ( .A(n2144), .B(n2145), .Z(n2136) );
  AND U2087 ( .A(n2146), .B(n2147), .Z(n2145) );
  XOR U2088 ( .A(n2144), .B(n1970), .Z(n2147) );
  XOR U2089 ( .A(n2148), .B(n2149), .Z(n1970) );
  AND U2090 ( .A(n133), .B(n2150), .Z(n2149) );
  XOR U2091 ( .A(n2151), .B(n2148), .Z(n2150) );
  XNOR U2092 ( .A(n1967), .B(n2144), .Z(n2146) );
  XOR U2093 ( .A(n2152), .B(n2153), .Z(n1967) );
  AND U2094 ( .A(n131), .B(n2154), .Z(n2153) );
  XOR U2095 ( .A(n2155), .B(n2152), .Z(n2154) );
  XOR U2096 ( .A(n2156), .B(n2157), .Z(n2144) );
  AND U2097 ( .A(n2158), .B(n2159), .Z(n2157) );
  XOR U2098 ( .A(n2156), .B(n1982), .Z(n2159) );
  XOR U2099 ( .A(n2160), .B(n2161), .Z(n1982) );
  AND U2100 ( .A(n133), .B(n2162), .Z(n2161) );
  XOR U2101 ( .A(n2163), .B(n2160), .Z(n2162) );
  XNOR U2102 ( .A(n1979), .B(n2156), .Z(n2158) );
  XOR U2103 ( .A(n2164), .B(n2165), .Z(n1979) );
  AND U2104 ( .A(n131), .B(n2166), .Z(n2165) );
  XOR U2105 ( .A(n2167), .B(n2164), .Z(n2166) );
  XOR U2106 ( .A(n2168), .B(n2169), .Z(n2156) );
  AND U2107 ( .A(n2170), .B(n2171), .Z(n2169) );
  XOR U2108 ( .A(n2168), .B(n1994), .Z(n2171) );
  XOR U2109 ( .A(n2172), .B(n2173), .Z(n1994) );
  AND U2110 ( .A(n133), .B(n2174), .Z(n2173) );
  XOR U2111 ( .A(n2175), .B(n2172), .Z(n2174) );
  XNOR U2112 ( .A(n1991), .B(n2168), .Z(n2170) );
  XOR U2113 ( .A(n2176), .B(n2177), .Z(n1991) );
  AND U2114 ( .A(n131), .B(n2178), .Z(n2177) );
  XOR U2115 ( .A(n2179), .B(n2176), .Z(n2178) );
  XOR U2116 ( .A(n2180), .B(n2181), .Z(n2168) );
  AND U2117 ( .A(n2182), .B(n2183), .Z(n2181) );
  XOR U2118 ( .A(n2180), .B(n2006), .Z(n2183) );
  XOR U2119 ( .A(n2184), .B(n2185), .Z(n2006) );
  AND U2120 ( .A(n133), .B(n2186), .Z(n2185) );
  XOR U2121 ( .A(n2187), .B(n2184), .Z(n2186) );
  XNOR U2122 ( .A(n2003), .B(n2180), .Z(n2182) );
  XOR U2123 ( .A(n2188), .B(n2189), .Z(n2003) );
  AND U2124 ( .A(n131), .B(n2190), .Z(n2189) );
  XOR U2125 ( .A(n2191), .B(n2188), .Z(n2190) );
  XOR U2126 ( .A(n2192), .B(n2193), .Z(n2180) );
  AND U2127 ( .A(n2194), .B(n2195), .Z(n2193) );
  XOR U2128 ( .A(n2192), .B(n2018), .Z(n2195) );
  XOR U2129 ( .A(n2196), .B(n2197), .Z(n2018) );
  AND U2130 ( .A(n133), .B(n2198), .Z(n2197) );
  XOR U2131 ( .A(n2199), .B(n2196), .Z(n2198) );
  XNOR U2132 ( .A(n2015), .B(n2192), .Z(n2194) );
  XOR U2133 ( .A(n2200), .B(n2201), .Z(n2015) );
  AND U2134 ( .A(n131), .B(n2202), .Z(n2201) );
  XOR U2135 ( .A(n2203), .B(n2200), .Z(n2202) );
  XOR U2136 ( .A(n2204), .B(n2205), .Z(n2192) );
  AND U2137 ( .A(n2206), .B(n2207), .Z(n2205) );
  XOR U2138 ( .A(n2204), .B(n2030), .Z(n2207) );
  XOR U2139 ( .A(n2208), .B(n2209), .Z(n2030) );
  AND U2140 ( .A(n133), .B(n2210), .Z(n2209) );
  XOR U2141 ( .A(n2211), .B(n2208), .Z(n2210) );
  XNOR U2142 ( .A(n2027), .B(n2204), .Z(n2206) );
  XOR U2143 ( .A(n2212), .B(n2213), .Z(n2027) );
  AND U2144 ( .A(n131), .B(n2214), .Z(n2213) );
  XOR U2145 ( .A(n2215), .B(n2212), .Z(n2214) );
  XOR U2146 ( .A(n2216), .B(n2217), .Z(n2204) );
  AND U2147 ( .A(n2218), .B(n2219), .Z(n2217) );
  XOR U2148 ( .A(n2216), .B(n2042), .Z(n2219) );
  XOR U2149 ( .A(n2220), .B(n2221), .Z(n2042) );
  AND U2150 ( .A(n133), .B(n2222), .Z(n2221) );
  XOR U2151 ( .A(n2223), .B(n2220), .Z(n2222) );
  XNOR U2152 ( .A(n2039), .B(n2216), .Z(n2218) );
  XOR U2153 ( .A(n2224), .B(n2225), .Z(n2039) );
  AND U2154 ( .A(n131), .B(n2226), .Z(n2225) );
  XOR U2155 ( .A(n2227), .B(n2224), .Z(n2226) );
  XOR U2156 ( .A(n2228), .B(n2229), .Z(n2216) );
  AND U2157 ( .A(n2230), .B(n2231), .Z(n2229) );
  XOR U2158 ( .A(n2228), .B(n2054), .Z(n2231) );
  XOR U2159 ( .A(n2232), .B(n2233), .Z(n2054) );
  AND U2160 ( .A(n133), .B(n2234), .Z(n2233) );
  XOR U2161 ( .A(n2235), .B(n2232), .Z(n2234) );
  XNOR U2162 ( .A(n2051), .B(n2228), .Z(n2230) );
  XOR U2163 ( .A(n2236), .B(n2237), .Z(n2051) );
  AND U2164 ( .A(n131), .B(n2238), .Z(n2237) );
  XOR U2165 ( .A(n2239), .B(n2236), .Z(n2238) );
  XOR U2166 ( .A(n2240), .B(n2241), .Z(n2228) );
  AND U2167 ( .A(n2242), .B(n2243), .Z(n2241) );
  XOR U2168 ( .A(n2240), .B(n2066), .Z(n2243) );
  XOR U2169 ( .A(n2244), .B(n2245), .Z(n2066) );
  AND U2170 ( .A(n133), .B(n2246), .Z(n2245) );
  XOR U2171 ( .A(n2247), .B(n2244), .Z(n2246) );
  XNOR U2172 ( .A(n2063), .B(n2240), .Z(n2242) );
  XOR U2173 ( .A(n2248), .B(n2249), .Z(n2063) );
  AND U2174 ( .A(n131), .B(n2250), .Z(n2249) );
  XOR U2175 ( .A(n2251), .B(n2248), .Z(n2250) );
  XOR U2176 ( .A(n2252), .B(n2253), .Z(n2240) );
  AND U2177 ( .A(n2254), .B(n2255), .Z(n2253) );
  XOR U2178 ( .A(n2252), .B(n2078), .Z(n2255) );
  XOR U2179 ( .A(n2256), .B(n2257), .Z(n2078) );
  AND U2180 ( .A(n133), .B(n2258), .Z(n2257) );
  XOR U2181 ( .A(n2259), .B(n2256), .Z(n2258) );
  XNOR U2182 ( .A(n2075), .B(n2252), .Z(n2254) );
  XOR U2183 ( .A(n2260), .B(n2261), .Z(n2075) );
  AND U2184 ( .A(n131), .B(n2262), .Z(n2261) );
  XOR U2185 ( .A(n2263), .B(n2260), .Z(n2262) );
  XOR U2186 ( .A(n2264), .B(n2265), .Z(n2252) );
  AND U2187 ( .A(n2266), .B(n2267), .Z(n2265) );
  XOR U2188 ( .A(n2090), .B(n2264), .Z(n2267) );
  XOR U2189 ( .A(n2268), .B(n2269), .Z(n2090) );
  AND U2190 ( .A(n133), .B(n2270), .Z(n2269) );
  XOR U2191 ( .A(n2268), .B(n2271), .Z(n2270) );
  XNOR U2192 ( .A(n2264), .B(n2087), .Z(n2266) );
  XOR U2193 ( .A(n2272), .B(n2273), .Z(n2087) );
  AND U2194 ( .A(n131), .B(n2274), .Z(n2273) );
  XOR U2195 ( .A(n2272), .B(n2275), .Z(n2274) );
  XOR U2196 ( .A(n2276), .B(n2277), .Z(n2264) );
  AND U2197 ( .A(n2278), .B(n2279), .Z(n2277) );
  XOR U2198 ( .A(n2276), .B(n2102), .Z(n2279) );
  XOR U2199 ( .A(n2280), .B(n2281), .Z(n2102) );
  AND U2200 ( .A(n133), .B(n2282), .Z(n2281) );
  XOR U2201 ( .A(n2283), .B(n2280), .Z(n2282) );
  XNOR U2202 ( .A(n2099), .B(n2276), .Z(n2278) );
  XOR U2203 ( .A(n2284), .B(n2285), .Z(n2099) );
  AND U2204 ( .A(n131), .B(n2286), .Z(n2285) );
  XOR U2205 ( .A(n2287), .B(n2284), .Z(n2286) );
  XOR U2206 ( .A(n2288), .B(n2289), .Z(n2276) );
  AND U2207 ( .A(n2290), .B(n2291), .Z(n2289) );
  XOR U2208 ( .A(n2288), .B(n2114), .Z(n2291) );
  XOR U2209 ( .A(n2292), .B(n2293), .Z(n2114) );
  AND U2210 ( .A(n133), .B(n2294), .Z(n2293) );
  XOR U2211 ( .A(n2295), .B(n2292), .Z(n2294) );
  XNOR U2212 ( .A(n2111), .B(n2288), .Z(n2290) );
  XOR U2213 ( .A(n2296), .B(n2297), .Z(n2111) );
  AND U2214 ( .A(n131), .B(n2298), .Z(n2297) );
  XOR U2215 ( .A(n2299), .B(n2296), .Z(n2298) );
  XOR U2216 ( .A(n2300), .B(n2301), .Z(n2288) );
  AND U2217 ( .A(n2302), .B(n2303), .Z(n2301) );
  XNOR U2218 ( .A(n2304), .B(n2127), .Z(n2303) );
  XOR U2219 ( .A(n2305), .B(n2306), .Z(n2127) );
  AND U2220 ( .A(n133), .B(n2307), .Z(n2306) );
  XOR U2221 ( .A(n2308), .B(n2305), .Z(n2307) );
  XNOR U2222 ( .A(n2124), .B(n2300), .Z(n2302) );
  XOR U2223 ( .A(n2309), .B(n2310), .Z(n2124) );
  AND U2224 ( .A(n131), .B(n2311), .Z(n2310) );
  XOR U2225 ( .A(n2312), .B(n2309), .Z(n2311) );
  IV U2226 ( .A(n2304), .Z(n2300) );
  AND U2227 ( .A(n2132), .B(n2135), .Z(n2304) );
  XNOR U2228 ( .A(n2313), .B(n2314), .Z(n2135) );
  AND U2229 ( .A(n133), .B(n2315), .Z(n2314) );
  XNOR U2230 ( .A(n2316), .B(n2313), .Z(n2315) );
  XOR U2231 ( .A(n2317), .B(n2318), .Z(n133) );
  AND U2232 ( .A(n2319), .B(n2320), .Z(n2318) );
  XNOR U2233 ( .A(n2140), .B(n2317), .Z(n2320) );
  AND U2234 ( .A(p_input[255]), .B(p_input[239]), .Z(n2140) );
  XOR U2235 ( .A(n2317), .B(n2141), .Z(n2319) );
  AND U2236 ( .A(p_input[223]), .B(p_input[207]), .Z(n2141) );
  XOR U2237 ( .A(n2321), .B(n2322), .Z(n2317) );
  AND U2238 ( .A(n2323), .B(n2324), .Z(n2322) );
  XOR U2239 ( .A(n2321), .B(n2151), .Z(n2324) );
  XNOR U2240 ( .A(p_input[238]), .B(n2325), .Z(n2151) );
  AND U2241 ( .A(n149), .B(n2326), .Z(n2325) );
  XOR U2242 ( .A(p_input[254]), .B(p_input[238]), .Z(n2326) );
  XNOR U2243 ( .A(n2148), .B(n2321), .Z(n2323) );
  XOR U2244 ( .A(n2327), .B(n2328), .Z(n2148) );
  AND U2245 ( .A(n147), .B(n2329), .Z(n2328) );
  XOR U2246 ( .A(p_input[222]), .B(p_input[206]), .Z(n2329) );
  XOR U2247 ( .A(n2330), .B(n2331), .Z(n2321) );
  AND U2248 ( .A(n2332), .B(n2333), .Z(n2331) );
  XOR U2249 ( .A(n2330), .B(n2163), .Z(n2333) );
  XNOR U2250 ( .A(p_input[237]), .B(n2334), .Z(n2163) );
  AND U2251 ( .A(n149), .B(n2335), .Z(n2334) );
  XOR U2252 ( .A(p_input[253]), .B(p_input[237]), .Z(n2335) );
  XNOR U2253 ( .A(n2160), .B(n2330), .Z(n2332) );
  XOR U2254 ( .A(n2336), .B(n2337), .Z(n2160) );
  AND U2255 ( .A(n147), .B(n2338), .Z(n2337) );
  XOR U2256 ( .A(p_input[221]), .B(p_input[205]), .Z(n2338) );
  XOR U2257 ( .A(n2339), .B(n2340), .Z(n2330) );
  AND U2258 ( .A(n2341), .B(n2342), .Z(n2340) );
  XOR U2259 ( .A(n2339), .B(n2175), .Z(n2342) );
  XNOR U2260 ( .A(p_input[236]), .B(n2343), .Z(n2175) );
  AND U2261 ( .A(n149), .B(n2344), .Z(n2343) );
  XOR U2262 ( .A(p_input[252]), .B(p_input[236]), .Z(n2344) );
  XNOR U2263 ( .A(n2172), .B(n2339), .Z(n2341) );
  XOR U2264 ( .A(n2345), .B(n2346), .Z(n2172) );
  AND U2265 ( .A(n147), .B(n2347), .Z(n2346) );
  XOR U2266 ( .A(p_input[220]), .B(p_input[204]), .Z(n2347) );
  XOR U2267 ( .A(n2348), .B(n2349), .Z(n2339) );
  AND U2268 ( .A(n2350), .B(n2351), .Z(n2349) );
  XOR U2269 ( .A(n2348), .B(n2187), .Z(n2351) );
  XNOR U2270 ( .A(p_input[235]), .B(n2352), .Z(n2187) );
  AND U2271 ( .A(n149), .B(n2353), .Z(n2352) );
  XOR U2272 ( .A(p_input[251]), .B(p_input[235]), .Z(n2353) );
  XNOR U2273 ( .A(n2184), .B(n2348), .Z(n2350) );
  XOR U2274 ( .A(n2354), .B(n2355), .Z(n2184) );
  AND U2275 ( .A(n147), .B(n2356), .Z(n2355) );
  XOR U2276 ( .A(p_input[219]), .B(p_input[203]), .Z(n2356) );
  XOR U2277 ( .A(n2357), .B(n2358), .Z(n2348) );
  AND U2278 ( .A(n2359), .B(n2360), .Z(n2358) );
  XOR U2279 ( .A(n2357), .B(n2199), .Z(n2360) );
  XNOR U2280 ( .A(p_input[234]), .B(n2361), .Z(n2199) );
  AND U2281 ( .A(n149), .B(n2362), .Z(n2361) );
  XOR U2282 ( .A(p_input[250]), .B(p_input[234]), .Z(n2362) );
  XNOR U2283 ( .A(n2196), .B(n2357), .Z(n2359) );
  XOR U2284 ( .A(n2363), .B(n2364), .Z(n2196) );
  AND U2285 ( .A(n147), .B(n2365), .Z(n2364) );
  XOR U2286 ( .A(p_input[218]), .B(p_input[202]), .Z(n2365) );
  XOR U2287 ( .A(n2366), .B(n2367), .Z(n2357) );
  AND U2288 ( .A(n2368), .B(n2369), .Z(n2367) );
  XOR U2289 ( .A(n2366), .B(n2211), .Z(n2369) );
  XNOR U2290 ( .A(p_input[233]), .B(n2370), .Z(n2211) );
  AND U2291 ( .A(n149), .B(n2371), .Z(n2370) );
  XOR U2292 ( .A(p_input[249]), .B(p_input[233]), .Z(n2371) );
  XNOR U2293 ( .A(n2208), .B(n2366), .Z(n2368) );
  XOR U2294 ( .A(n2372), .B(n2373), .Z(n2208) );
  AND U2295 ( .A(n147), .B(n2374), .Z(n2373) );
  XOR U2296 ( .A(p_input[217]), .B(p_input[201]), .Z(n2374) );
  XOR U2297 ( .A(n2375), .B(n2376), .Z(n2366) );
  AND U2298 ( .A(n2377), .B(n2378), .Z(n2376) );
  XOR U2299 ( .A(n2375), .B(n2223), .Z(n2378) );
  XNOR U2300 ( .A(p_input[232]), .B(n2379), .Z(n2223) );
  AND U2301 ( .A(n149), .B(n2380), .Z(n2379) );
  XOR U2302 ( .A(p_input[248]), .B(p_input[232]), .Z(n2380) );
  XNOR U2303 ( .A(n2220), .B(n2375), .Z(n2377) );
  XOR U2304 ( .A(n2381), .B(n2382), .Z(n2220) );
  AND U2305 ( .A(n147), .B(n2383), .Z(n2382) );
  XOR U2306 ( .A(p_input[216]), .B(p_input[200]), .Z(n2383) );
  XOR U2307 ( .A(n2384), .B(n2385), .Z(n2375) );
  AND U2308 ( .A(n2386), .B(n2387), .Z(n2385) );
  XOR U2309 ( .A(n2384), .B(n2235), .Z(n2387) );
  XNOR U2310 ( .A(p_input[231]), .B(n2388), .Z(n2235) );
  AND U2311 ( .A(n149), .B(n2389), .Z(n2388) );
  XOR U2312 ( .A(p_input[247]), .B(p_input[231]), .Z(n2389) );
  XNOR U2313 ( .A(n2232), .B(n2384), .Z(n2386) );
  XOR U2314 ( .A(n2390), .B(n2391), .Z(n2232) );
  AND U2315 ( .A(n147), .B(n2392), .Z(n2391) );
  XOR U2316 ( .A(p_input[215]), .B(p_input[199]), .Z(n2392) );
  XOR U2317 ( .A(n2393), .B(n2394), .Z(n2384) );
  AND U2318 ( .A(n2395), .B(n2396), .Z(n2394) );
  XOR U2319 ( .A(n2393), .B(n2247), .Z(n2396) );
  XNOR U2320 ( .A(p_input[230]), .B(n2397), .Z(n2247) );
  AND U2321 ( .A(n149), .B(n2398), .Z(n2397) );
  XOR U2322 ( .A(p_input[246]), .B(p_input[230]), .Z(n2398) );
  XNOR U2323 ( .A(n2244), .B(n2393), .Z(n2395) );
  XOR U2324 ( .A(n2399), .B(n2400), .Z(n2244) );
  AND U2325 ( .A(n147), .B(n2401), .Z(n2400) );
  XOR U2326 ( .A(p_input[214]), .B(p_input[198]), .Z(n2401) );
  XOR U2327 ( .A(n2402), .B(n2403), .Z(n2393) );
  AND U2328 ( .A(n2404), .B(n2405), .Z(n2403) );
  XOR U2329 ( .A(n2402), .B(n2259), .Z(n2405) );
  XNOR U2330 ( .A(p_input[229]), .B(n2406), .Z(n2259) );
  AND U2331 ( .A(n149), .B(n2407), .Z(n2406) );
  XOR U2332 ( .A(p_input[245]), .B(p_input[229]), .Z(n2407) );
  XNOR U2333 ( .A(n2256), .B(n2402), .Z(n2404) );
  XOR U2334 ( .A(n2408), .B(n2409), .Z(n2256) );
  AND U2335 ( .A(n147), .B(n2410), .Z(n2409) );
  XOR U2336 ( .A(p_input[213]), .B(p_input[197]), .Z(n2410) );
  XOR U2337 ( .A(n2411), .B(n2412), .Z(n2402) );
  AND U2338 ( .A(n2413), .B(n2414), .Z(n2412) );
  XOR U2339 ( .A(n2271), .B(n2411), .Z(n2414) );
  XNOR U2340 ( .A(p_input[228]), .B(n2415), .Z(n2271) );
  AND U2341 ( .A(n149), .B(n2416), .Z(n2415) );
  XOR U2342 ( .A(p_input[244]), .B(p_input[228]), .Z(n2416) );
  XNOR U2343 ( .A(n2411), .B(n2268), .Z(n2413) );
  XOR U2344 ( .A(n2417), .B(n2418), .Z(n2268) );
  AND U2345 ( .A(n147), .B(n2419), .Z(n2418) );
  XOR U2346 ( .A(p_input[212]), .B(p_input[196]), .Z(n2419) );
  XOR U2347 ( .A(n2420), .B(n2421), .Z(n2411) );
  AND U2348 ( .A(n2422), .B(n2423), .Z(n2421) );
  XOR U2349 ( .A(n2420), .B(n2283), .Z(n2423) );
  XNOR U2350 ( .A(p_input[227]), .B(n2424), .Z(n2283) );
  AND U2351 ( .A(n149), .B(n2425), .Z(n2424) );
  XOR U2352 ( .A(p_input[243]), .B(p_input[227]), .Z(n2425) );
  XNOR U2353 ( .A(n2280), .B(n2420), .Z(n2422) );
  XOR U2354 ( .A(n2426), .B(n2427), .Z(n2280) );
  AND U2355 ( .A(n147), .B(n2428), .Z(n2427) );
  XOR U2356 ( .A(p_input[211]), .B(p_input[195]), .Z(n2428) );
  XOR U2357 ( .A(n2429), .B(n2430), .Z(n2420) );
  AND U2358 ( .A(n2431), .B(n2432), .Z(n2430) );
  XOR U2359 ( .A(n2429), .B(n2295), .Z(n2432) );
  XNOR U2360 ( .A(p_input[226]), .B(n2433), .Z(n2295) );
  AND U2361 ( .A(n149), .B(n2434), .Z(n2433) );
  XOR U2362 ( .A(p_input[242]), .B(p_input[226]), .Z(n2434) );
  XNOR U2363 ( .A(n2292), .B(n2429), .Z(n2431) );
  XOR U2364 ( .A(n2435), .B(n2436), .Z(n2292) );
  AND U2365 ( .A(n147), .B(n2437), .Z(n2436) );
  XOR U2366 ( .A(p_input[210]), .B(p_input[194]), .Z(n2437) );
  XOR U2367 ( .A(n2438), .B(n2439), .Z(n2429) );
  AND U2368 ( .A(n2440), .B(n2441), .Z(n2439) );
  XNOR U2369 ( .A(n2442), .B(n2308), .Z(n2441) );
  XNOR U2370 ( .A(p_input[225]), .B(n2443), .Z(n2308) );
  AND U2371 ( .A(n149), .B(n2444), .Z(n2443) );
  XNOR U2372 ( .A(p_input[241]), .B(n2445), .Z(n2444) );
  IV U2373 ( .A(p_input[225]), .Z(n2445) );
  XNOR U2374 ( .A(n2305), .B(n2438), .Z(n2440) );
  XNOR U2375 ( .A(p_input[193]), .B(n2446), .Z(n2305) );
  AND U2376 ( .A(n147), .B(n2447), .Z(n2446) );
  XOR U2377 ( .A(p_input[209]), .B(p_input[193]), .Z(n2447) );
  IV U2378 ( .A(n2442), .Z(n2438) );
  AND U2379 ( .A(n2313), .B(n2316), .Z(n2442) );
  XOR U2380 ( .A(p_input[224]), .B(n2448), .Z(n2316) );
  AND U2381 ( .A(n149), .B(n2449), .Z(n2448) );
  XOR U2382 ( .A(p_input[240]), .B(p_input[224]), .Z(n2449) );
  XOR U2383 ( .A(n2450), .B(n2451), .Z(n149) );
  AND U2384 ( .A(n2452), .B(n2453), .Z(n2451) );
  XNOR U2385 ( .A(p_input[255]), .B(n2450), .Z(n2453) );
  XOR U2386 ( .A(n2450), .B(p_input[239]), .Z(n2452) );
  XOR U2387 ( .A(n2454), .B(n2455), .Z(n2450) );
  AND U2388 ( .A(n2456), .B(n2457), .Z(n2455) );
  XNOR U2389 ( .A(p_input[254]), .B(n2454), .Z(n2457) );
  XOR U2390 ( .A(n2454), .B(p_input[238]), .Z(n2456) );
  XOR U2391 ( .A(n2458), .B(n2459), .Z(n2454) );
  AND U2392 ( .A(n2460), .B(n2461), .Z(n2459) );
  XNOR U2393 ( .A(p_input[253]), .B(n2458), .Z(n2461) );
  XOR U2394 ( .A(n2458), .B(p_input[237]), .Z(n2460) );
  XOR U2395 ( .A(n2462), .B(n2463), .Z(n2458) );
  AND U2396 ( .A(n2464), .B(n2465), .Z(n2463) );
  XNOR U2397 ( .A(p_input[252]), .B(n2462), .Z(n2465) );
  XOR U2398 ( .A(n2462), .B(p_input[236]), .Z(n2464) );
  XOR U2399 ( .A(n2466), .B(n2467), .Z(n2462) );
  AND U2400 ( .A(n2468), .B(n2469), .Z(n2467) );
  XNOR U2401 ( .A(p_input[251]), .B(n2466), .Z(n2469) );
  XOR U2402 ( .A(n2466), .B(p_input[235]), .Z(n2468) );
  XOR U2403 ( .A(n2470), .B(n2471), .Z(n2466) );
  AND U2404 ( .A(n2472), .B(n2473), .Z(n2471) );
  XNOR U2405 ( .A(p_input[250]), .B(n2470), .Z(n2473) );
  XOR U2406 ( .A(n2470), .B(p_input[234]), .Z(n2472) );
  XOR U2407 ( .A(n2474), .B(n2475), .Z(n2470) );
  AND U2408 ( .A(n2476), .B(n2477), .Z(n2475) );
  XNOR U2409 ( .A(p_input[249]), .B(n2474), .Z(n2477) );
  XOR U2410 ( .A(n2474), .B(p_input[233]), .Z(n2476) );
  XOR U2411 ( .A(n2478), .B(n2479), .Z(n2474) );
  AND U2412 ( .A(n2480), .B(n2481), .Z(n2479) );
  XNOR U2413 ( .A(p_input[248]), .B(n2478), .Z(n2481) );
  XOR U2414 ( .A(n2478), .B(p_input[232]), .Z(n2480) );
  XOR U2415 ( .A(n2482), .B(n2483), .Z(n2478) );
  AND U2416 ( .A(n2484), .B(n2485), .Z(n2483) );
  XNOR U2417 ( .A(p_input[247]), .B(n2482), .Z(n2485) );
  XOR U2418 ( .A(n2482), .B(p_input[231]), .Z(n2484) );
  XOR U2419 ( .A(n2486), .B(n2487), .Z(n2482) );
  AND U2420 ( .A(n2488), .B(n2489), .Z(n2487) );
  XNOR U2421 ( .A(p_input[246]), .B(n2486), .Z(n2489) );
  XOR U2422 ( .A(n2486), .B(p_input[230]), .Z(n2488) );
  XOR U2423 ( .A(n2490), .B(n2491), .Z(n2486) );
  AND U2424 ( .A(n2492), .B(n2493), .Z(n2491) );
  XNOR U2425 ( .A(p_input[245]), .B(n2490), .Z(n2493) );
  XOR U2426 ( .A(n2490), .B(p_input[229]), .Z(n2492) );
  XOR U2427 ( .A(n2494), .B(n2495), .Z(n2490) );
  AND U2428 ( .A(n2496), .B(n2497), .Z(n2495) );
  XNOR U2429 ( .A(p_input[244]), .B(n2494), .Z(n2497) );
  XOR U2430 ( .A(n2494), .B(p_input[228]), .Z(n2496) );
  XOR U2431 ( .A(n2498), .B(n2499), .Z(n2494) );
  AND U2432 ( .A(n2500), .B(n2501), .Z(n2499) );
  XNOR U2433 ( .A(p_input[243]), .B(n2498), .Z(n2501) );
  XOR U2434 ( .A(n2498), .B(p_input[227]), .Z(n2500) );
  XOR U2435 ( .A(n2502), .B(n2503), .Z(n2498) );
  AND U2436 ( .A(n2504), .B(n2505), .Z(n2503) );
  XNOR U2437 ( .A(p_input[242]), .B(n2502), .Z(n2505) );
  XOR U2438 ( .A(n2502), .B(p_input[226]), .Z(n2504) );
  XNOR U2439 ( .A(n2506), .B(n2507), .Z(n2502) );
  AND U2440 ( .A(n2508), .B(n2509), .Z(n2507) );
  XOR U2441 ( .A(p_input[241]), .B(n2506), .Z(n2509) );
  XNOR U2442 ( .A(p_input[225]), .B(n2506), .Z(n2508) );
  AND U2443 ( .A(p_input[240]), .B(n2510), .Z(n2506) );
  IV U2444 ( .A(p_input[224]), .Z(n2510) );
  XNOR U2445 ( .A(p_input[192]), .B(n2511), .Z(n2313) );
  AND U2446 ( .A(n147), .B(n2512), .Z(n2511) );
  XOR U2447 ( .A(p_input[208]), .B(p_input[192]), .Z(n2512) );
  XOR U2448 ( .A(n2513), .B(n2514), .Z(n147) );
  AND U2449 ( .A(n2515), .B(n2516), .Z(n2514) );
  XNOR U2450 ( .A(p_input[223]), .B(n2513), .Z(n2516) );
  XOR U2451 ( .A(n2513), .B(p_input[207]), .Z(n2515) );
  XOR U2452 ( .A(n2517), .B(n2518), .Z(n2513) );
  AND U2453 ( .A(n2519), .B(n2520), .Z(n2518) );
  XNOR U2454 ( .A(p_input[222]), .B(n2517), .Z(n2520) );
  XNOR U2455 ( .A(n2517), .B(n2327), .Z(n2519) );
  IV U2456 ( .A(p_input[206]), .Z(n2327) );
  XOR U2457 ( .A(n2521), .B(n2522), .Z(n2517) );
  AND U2458 ( .A(n2523), .B(n2524), .Z(n2522) );
  XNOR U2459 ( .A(p_input[221]), .B(n2521), .Z(n2524) );
  XNOR U2460 ( .A(n2521), .B(n2336), .Z(n2523) );
  IV U2461 ( .A(p_input[205]), .Z(n2336) );
  XOR U2462 ( .A(n2525), .B(n2526), .Z(n2521) );
  AND U2463 ( .A(n2527), .B(n2528), .Z(n2526) );
  XNOR U2464 ( .A(p_input[220]), .B(n2525), .Z(n2528) );
  XNOR U2465 ( .A(n2525), .B(n2345), .Z(n2527) );
  IV U2466 ( .A(p_input[204]), .Z(n2345) );
  XOR U2467 ( .A(n2529), .B(n2530), .Z(n2525) );
  AND U2468 ( .A(n2531), .B(n2532), .Z(n2530) );
  XNOR U2469 ( .A(p_input[219]), .B(n2529), .Z(n2532) );
  XNOR U2470 ( .A(n2529), .B(n2354), .Z(n2531) );
  IV U2471 ( .A(p_input[203]), .Z(n2354) );
  XOR U2472 ( .A(n2533), .B(n2534), .Z(n2529) );
  AND U2473 ( .A(n2535), .B(n2536), .Z(n2534) );
  XNOR U2474 ( .A(p_input[218]), .B(n2533), .Z(n2536) );
  XNOR U2475 ( .A(n2533), .B(n2363), .Z(n2535) );
  IV U2476 ( .A(p_input[202]), .Z(n2363) );
  XOR U2477 ( .A(n2537), .B(n2538), .Z(n2533) );
  AND U2478 ( .A(n2539), .B(n2540), .Z(n2538) );
  XNOR U2479 ( .A(p_input[217]), .B(n2537), .Z(n2540) );
  XNOR U2480 ( .A(n2537), .B(n2372), .Z(n2539) );
  IV U2481 ( .A(p_input[201]), .Z(n2372) );
  XOR U2482 ( .A(n2541), .B(n2542), .Z(n2537) );
  AND U2483 ( .A(n2543), .B(n2544), .Z(n2542) );
  XNOR U2484 ( .A(p_input[216]), .B(n2541), .Z(n2544) );
  XNOR U2485 ( .A(n2541), .B(n2381), .Z(n2543) );
  IV U2486 ( .A(p_input[200]), .Z(n2381) );
  XOR U2487 ( .A(n2545), .B(n2546), .Z(n2541) );
  AND U2488 ( .A(n2547), .B(n2548), .Z(n2546) );
  XNOR U2489 ( .A(p_input[215]), .B(n2545), .Z(n2548) );
  XNOR U2490 ( .A(n2545), .B(n2390), .Z(n2547) );
  IV U2491 ( .A(p_input[199]), .Z(n2390) );
  XOR U2492 ( .A(n2549), .B(n2550), .Z(n2545) );
  AND U2493 ( .A(n2551), .B(n2552), .Z(n2550) );
  XNOR U2494 ( .A(p_input[214]), .B(n2549), .Z(n2552) );
  XNOR U2495 ( .A(n2549), .B(n2399), .Z(n2551) );
  IV U2496 ( .A(p_input[198]), .Z(n2399) );
  XOR U2497 ( .A(n2553), .B(n2554), .Z(n2549) );
  AND U2498 ( .A(n2555), .B(n2556), .Z(n2554) );
  XNOR U2499 ( .A(p_input[213]), .B(n2553), .Z(n2556) );
  XNOR U2500 ( .A(n2553), .B(n2408), .Z(n2555) );
  IV U2501 ( .A(p_input[197]), .Z(n2408) );
  XOR U2502 ( .A(n2557), .B(n2558), .Z(n2553) );
  AND U2503 ( .A(n2559), .B(n2560), .Z(n2558) );
  XNOR U2504 ( .A(p_input[212]), .B(n2557), .Z(n2560) );
  XNOR U2505 ( .A(n2557), .B(n2417), .Z(n2559) );
  IV U2506 ( .A(p_input[196]), .Z(n2417) );
  XOR U2507 ( .A(n2561), .B(n2562), .Z(n2557) );
  AND U2508 ( .A(n2563), .B(n2564), .Z(n2562) );
  XNOR U2509 ( .A(p_input[211]), .B(n2561), .Z(n2564) );
  XNOR U2510 ( .A(n2561), .B(n2426), .Z(n2563) );
  IV U2511 ( .A(p_input[195]), .Z(n2426) );
  XOR U2512 ( .A(n2565), .B(n2566), .Z(n2561) );
  AND U2513 ( .A(n2567), .B(n2568), .Z(n2566) );
  XNOR U2514 ( .A(p_input[210]), .B(n2565), .Z(n2568) );
  XNOR U2515 ( .A(n2565), .B(n2435), .Z(n2567) );
  IV U2516 ( .A(p_input[194]), .Z(n2435) );
  XNOR U2517 ( .A(n2569), .B(n2570), .Z(n2565) );
  AND U2518 ( .A(n2571), .B(n2572), .Z(n2570) );
  XOR U2519 ( .A(p_input[209]), .B(n2569), .Z(n2572) );
  XNOR U2520 ( .A(p_input[193]), .B(n2569), .Z(n2571) );
  AND U2521 ( .A(p_input[208]), .B(n2573), .Z(n2569) );
  IV U2522 ( .A(p_input[192]), .Z(n2573) );
  XOR U2523 ( .A(n2574), .B(n2575), .Z(n2132) );
  AND U2524 ( .A(n131), .B(n2576), .Z(n2575) );
  XNOR U2525 ( .A(n2577), .B(n2574), .Z(n2576) );
  XOR U2526 ( .A(n2578), .B(n2579), .Z(n131) );
  AND U2527 ( .A(n2580), .B(n2581), .Z(n2579) );
  XNOR U2528 ( .A(n2142), .B(n2578), .Z(n2581) );
  AND U2529 ( .A(p_input[191]), .B(p_input[175]), .Z(n2142) );
  XOR U2530 ( .A(n2578), .B(n2143), .Z(n2580) );
  AND U2531 ( .A(p_input[159]), .B(p_input[143]), .Z(n2143) );
  XOR U2532 ( .A(n2582), .B(n2583), .Z(n2578) );
  AND U2533 ( .A(n2584), .B(n2585), .Z(n2583) );
  XOR U2534 ( .A(n2582), .B(n2155), .Z(n2585) );
  XNOR U2535 ( .A(p_input[174]), .B(n2586), .Z(n2155) );
  AND U2536 ( .A(n153), .B(n2587), .Z(n2586) );
  XOR U2537 ( .A(p_input[190]), .B(p_input[174]), .Z(n2587) );
  XNOR U2538 ( .A(n2152), .B(n2582), .Z(n2584) );
  XOR U2539 ( .A(n2588), .B(n2589), .Z(n2152) );
  AND U2540 ( .A(n150), .B(n2590), .Z(n2589) );
  XOR U2541 ( .A(p_input[158]), .B(p_input[142]), .Z(n2590) );
  XOR U2542 ( .A(n2591), .B(n2592), .Z(n2582) );
  AND U2543 ( .A(n2593), .B(n2594), .Z(n2592) );
  XOR U2544 ( .A(n2591), .B(n2167), .Z(n2594) );
  XNOR U2545 ( .A(p_input[173]), .B(n2595), .Z(n2167) );
  AND U2546 ( .A(n153), .B(n2596), .Z(n2595) );
  XOR U2547 ( .A(p_input[189]), .B(p_input[173]), .Z(n2596) );
  XNOR U2548 ( .A(n2164), .B(n2591), .Z(n2593) );
  XOR U2549 ( .A(n2597), .B(n2598), .Z(n2164) );
  AND U2550 ( .A(n150), .B(n2599), .Z(n2598) );
  XOR U2551 ( .A(p_input[157]), .B(p_input[141]), .Z(n2599) );
  XOR U2552 ( .A(n2600), .B(n2601), .Z(n2591) );
  AND U2553 ( .A(n2602), .B(n2603), .Z(n2601) );
  XOR U2554 ( .A(n2600), .B(n2179), .Z(n2603) );
  XNOR U2555 ( .A(p_input[172]), .B(n2604), .Z(n2179) );
  AND U2556 ( .A(n153), .B(n2605), .Z(n2604) );
  XOR U2557 ( .A(p_input[188]), .B(p_input[172]), .Z(n2605) );
  XNOR U2558 ( .A(n2176), .B(n2600), .Z(n2602) );
  XOR U2559 ( .A(n2606), .B(n2607), .Z(n2176) );
  AND U2560 ( .A(n150), .B(n2608), .Z(n2607) );
  XOR U2561 ( .A(p_input[156]), .B(p_input[140]), .Z(n2608) );
  XOR U2562 ( .A(n2609), .B(n2610), .Z(n2600) );
  AND U2563 ( .A(n2611), .B(n2612), .Z(n2610) );
  XOR U2564 ( .A(n2609), .B(n2191), .Z(n2612) );
  XNOR U2565 ( .A(p_input[171]), .B(n2613), .Z(n2191) );
  AND U2566 ( .A(n153), .B(n2614), .Z(n2613) );
  XOR U2567 ( .A(p_input[187]), .B(p_input[171]), .Z(n2614) );
  XNOR U2568 ( .A(n2188), .B(n2609), .Z(n2611) );
  XOR U2569 ( .A(n2615), .B(n2616), .Z(n2188) );
  AND U2570 ( .A(n150), .B(n2617), .Z(n2616) );
  XOR U2571 ( .A(p_input[155]), .B(p_input[139]), .Z(n2617) );
  XOR U2572 ( .A(n2618), .B(n2619), .Z(n2609) );
  AND U2573 ( .A(n2620), .B(n2621), .Z(n2619) );
  XOR U2574 ( .A(n2618), .B(n2203), .Z(n2621) );
  XNOR U2575 ( .A(p_input[170]), .B(n2622), .Z(n2203) );
  AND U2576 ( .A(n153), .B(n2623), .Z(n2622) );
  XOR U2577 ( .A(p_input[186]), .B(p_input[170]), .Z(n2623) );
  XNOR U2578 ( .A(n2200), .B(n2618), .Z(n2620) );
  XOR U2579 ( .A(n2624), .B(n2625), .Z(n2200) );
  AND U2580 ( .A(n150), .B(n2626), .Z(n2625) );
  XOR U2581 ( .A(p_input[154]), .B(p_input[138]), .Z(n2626) );
  XOR U2582 ( .A(n2627), .B(n2628), .Z(n2618) );
  AND U2583 ( .A(n2629), .B(n2630), .Z(n2628) );
  XOR U2584 ( .A(n2627), .B(n2215), .Z(n2630) );
  XNOR U2585 ( .A(p_input[169]), .B(n2631), .Z(n2215) );
  AND U2586 ( .A(n153), .B(n2632), .Z(n2631) );
  XOR U2587 ( .A(p_input[185]), .B(p_input[169]), .Z(n2632) );
  XNOR U2588 ( .A(n2212), .B(n2627), .Z(n2629) );
  XOR U2589 ( .A(n2633), .B(n2634), .Z(n2212) );
  AND U2590 ( .A(n150), .B(n2635), .Z(n2634) );
  XOR U2591 ( .A(p_input[153]), .B(p_input[137]), .Z(n2635) );
  XOR U2592 ( .A(n2636), .B(n2637), .Z(n2627) );
  AND U2593 ( .A(n2638), .B(n2639), .Z(n2637) );
  XOR U2594 ( .A(n2636), .B(n2227), .Z(n2639) );
  XNOR U2595 ( .A(p_input[168]), .B(n2640), .Z(n2227) );
  AND U2596 ( .A(n153), .B(n2641), .Z(n2640) );
  XOR U2597 ( .A(p_input[184]), .B(p_input[168]), .Z(n2641) );
  XNOR U2598 ( .A(n2224), .B(n2636), .Z(n2638) );
  XOR U2599 ( .A(n2642), .B(n2643), .Z(n2224) );
  AND U2600 ( .A(n150), .B(n2644), .Z(n2643) );
  XOR U2601 ( .A(p_input[152]), .B(p_input[136]), .Z(n2644) );
  XOR U2602 ( .A(n2645), .B(n2646), .Z(n2636) );
  AND U2603 ( .A(n2647), .B(n2648), .Z(n2646) );
  XOR U2604 ( .A(n2645), .B(n2239), .Z(n2648) );
  XNOR U2605 ( .A(p_input[167]), .B(n2649), .Z(n2239) );
  AND U2606 ( .A(n153), .B(n2650), .Z(n2649) );
  XOR U2607 ( .A(p_input[183]), .B(p_input[167]), .Z(n2650) );
  XNOR U2608 ( .A(n2236), .B(n2645), .Z(n2647) );
  XOR U2609 ( .A(n2651), .B(n2652), .Z(n2236) );
  AND U2610 ( .A(n150), .B(n2653), .Z(n2652) );
  XOR U2611 ( .A(p_input[151]), .B(p_input[135]), .Z(n2653) );
  XOR U2612 ( .A(n2654), .B(n2655), .Z(n2645) );
  AND U2613 ( .A(n2656), .B(n2657), .Z(n2655) );
  XOR U2614 ( .A(n2654), .B(n2251), .Z(n2657) );
  XNOR U2615 ( .A(p_input[166]), .B(n2658), .Z(n2251) );
  AND U2616 ( .A(n153), .B(n2659), .Z(n2658) );
  XOR U2617 ( .A(p_input[182]), .B(p_input[166]), .Z(n2659) );
  XNOR U2618 ( .A(n2248), .B(n2654), .Z(n2656) );
  XOR U2619 ( .A(n2660), .B(n2661), .Z(n2248) );
  AND U2620 ( .A(n150), .B(n2662), .Z(n2661) );
  XOR U2621 ( .A(p_input[150]), .B(p_input[134]), .Z(n2662) );
  XOR U2622 ( .A(n2663), .B(n2664), .Z(n2654) );
  AND U2623 ( .A(n2665), .B(n2666), .Z(n2664) );
  XOR U2624 ( .A(n2663), .B(n2263), .Z(n2666) );
  XNOR U2625 ( .A(p_input[165]), .B(n2667), .Z(n2263) );
  AND U2626 ( .A(n153), .B(n2668), .Z(n2667) );
  XOR U2627 ( .A(p_input[181]), .B(p_input[165]), .Z(n2668) );
  XNOR U2628 ( .A(n2260), .B(n2663), .Z(n2665) );
  XOR U2629 ( .A(n2669), .B(n2670), .Z(n2260) );
  AND U2630 ( .A(n150), .B(n2671), .Z(n2670) );
  XOR U2631 ( .A(p_input[149]), .B(p_input[133]), .Z(n2671) );
  XOR U2632 ( .A(n2672), .B(n2673), .Z(n2663) );
  AND U2633 ( .A(n2674), .B(n2675), .Z(n2673) );
  XOR U2634 ( .A(n2275), .B(n2672), .Z(n2675) );
  XNOR U2635 ( .A(p_input[164]), .B(n2676), .Z(n2275) );
  AND U2636 ( .A(n153), .B(n2677), .Z(n2676) );
  XOR U2637 ( .A(p_input[180]), .B(p_input[164]), .Z(n2677) );
  XNOR U2638 ( .A(n2672), .B(n2272), .Z(n2674) );
  XOR U2639 ( .A(n2678), .B(n2679), .Z(n2272) );
  AND U2640 ( .A(n150), .B(n2680), .Z(n2679) );
  XOR U2641 ( .A(p_input[148]), .B(p_input[132]), .Z(n2680) );
  XOR U2642 ( .A(n2681), .B(n2682), .Z(n2672) );
  AND U2643 ( .A(n2683), .B(n2684), .Z(n2682) );
  XOR U2644 ( .A(n2681), .B(n2287), .Z(n2684) );
  XNOR U2645 ( .A(p_input[163]), .B(n2685), .Z(n2287) );
  AND U2646 ( .A(n153), .B(n2686), .Z(n2685) );
  XOR U2647 ( .A(p_input[179]), .B(p_input[163]), .Z(n2686) );
  XNOR U2648 ( .A(n2284), .B(n2681), .Z(n2683) );
  XOR U2649 ( .A(n2687), .B(n2688), .Z(n2284) );
  AND U2650 ( .A(n150), .B(n2689), .Z(n2688) );
  XOR U2651 ( .A(p_input[147]), .B(p_input[131]), .Z(n2689) );
  XOR U2652 ( .A(n2690), .B(n2691), .Z(n2681) );
  AND U2653 ( .A(n2692), .B(n2693), .Z(n2691) );
  XOR U2654 ( .A(n2690), .B(n2299), .Z(n2693) );
  XNOR U2655 ( .A(p_input[162]), .B(n2694), .Z(n2299) );
  AND U2656 ( .A(n153), .B(n2695), .Z(n2694) );
  XOR U2657 ( .A(p_input[178]), .B(p_input[162]), .Z(n2695) );
  XNOR U2658 ( .A(n2296), .B(n2690), .Z(n2692) );
  XOR U2659 ( .A(n2696), .B(n2697), .Z(n2296) );
  AND U2660 ( .A(n150), .B(n2698), .Z(n2697) );
  XOR U2661 ( .A(p_input[146]), .B(p_input[130]), .Z(n2698) );
  XOR U2662 ( .A(n2699), .B(n2700), .Z(n2690) );
  AND U2663 ( .A(n2701), .B(n2702), .Z(n2700) );
  XNOR U2664 ( .A(n2703), .B(n2312), .Z(n2702) );
  XNOR U2665 ( .A(p_input[161]), .B(n2704), .Z(n2312) );
  AND U2666 ( .A(n153), .B(n2705), .Z(n2704) );
  XNOR U2667 ( .A(p_input[177]), .B(n2706), .Z(n2705) );
  IV U2668 ( .A(p_input[161]), .Z(n2706) );
  XNOR U2669 ( .A(n2309), .B(n2699), .Z(n2701) );
  XNOR U2670 ( .A(p_input[129]), .B(n2707), .Z(n2309) );
  AND U2671 ( .A(n150), .B(n2708), .Z(n2707) );
  XOR U2672 ( .A(p_input[145]), .B(p_input[129]), .Z(n2708) );
  IV U2673 ( .A(n2703), .Z(n2699) );
  AND U2674 ( .A(n2574), .B(n2577), .Z(n2703) );
  XOR U2675 ( .A(p_input[160]), .B(n2709), .Z(n2577) );
  AND U2676 ( .A(n153), .B(n2710), .Z(n2709) );
  XOR U2677 ( .A(p_input[176]), .B(p_input[160]), .Z(n2710) );
  XOR U2678 ( .A(n2711), .B(n2712), .Z(n153) );
  AND U2679 ( .A(n2713), .B(n2714), .Z(n2712) );
  XNOR U2680 ( .A(p_input[191]), .B(n2711), .Z(n2714) );
  XOR U2681 ( .A(n2711), .B(p_input[175]), .Z(n2713) );
  XOR U2682 ( .A(n2715), .B(n2716), .Z(n2711) );
  AND U2683 ( .A(n2717), .B(n2718), .Z(n2716) );
  XNOR U2684 ( .A(p_input[190]), .B(n2715), .Z(n2718) );
  XOR U2685 ( .A(n2715), .B(p_input[174]), .Z(n2717) );
  XOR U2686 ( .A(n2719), .B(n2720), .Z(n2715) );
  AND U2687 ( .A(n2721), .B(n2722), .Z(n2720) );
  XNOR U2688 ( .A(p_input[189]), .B(n2719), .Z(n2722) );
  XOR U2689 ( .A(n2719), .B(p_input[173]), .Z(n2721) );
  XOR U2690 ( .A(n2723), .B(n2724), .Z(n2719) );
  AND U2691 ( .A(n2725), .B(n2726), .Z(n2724) );
  XNOR U2692 ( .A(p_input[188]), .B(n2723), .Z(n2726) );
  XOR U2693 ( .A(n2723), .B(p_input[172]), .Z(n2725) );
  XOR U2694 ( .A(n2727), .B(n2728), .Z(n2723) );
  AND U2695 ( .A(n2729), .B(n2730), .Z(n2728) );
  XNOR U2696 ( .A(p_input[187]), .B(n2727), .Z(n2730) );
  XOR U2697 ( .A(n2727), .B(p_input[171]), .Z(n2729) );
  XOR U2698 ( .A(n2731), .B(n2732), .Z(n2727) );
  AND U2699 ( .A(n2733), .B(n2734), .Z(n2732) );
  XNOR U2700 ( .A(p_input[186]), .B(n2731), .Z(n2734) );
  XOR U2701 ( .A(n2731), .B(p_input[170]), .Z(n2733) );
  XOR U2702 ( .A(n2735), .B(n2736), .Z(n2731) );
  AND U2703 ( .A(n2737), .B(n2738), .Z(n2736) );
  XNOR U2704 ( .A(p_input[185]), .B(n2735), .Z(n2738) );
  XOR U2705 ( .A(n2735), .B(p_input[169]), .Z(n2737) );
  XOR U2706 ( .A(n2739), .B(n2740), .Z(n2735) );
  AND U2707 ( .A(n2741), .B(n2742), .Z(n2740) );
  XNOR U2708 ( .A(p_input[184]), .B(n2739), .Z(n2742) );
  XOR U2709 ( .A(n2739), .B(p_input[168]), .Z(n2741) );
  XOR U2710 ( .A(n2743), .B(n2744), .Z(n2739) );
  AND U2711 ( .A(n2745), .B(n2746), .Z(n2744) );
  XNOR U2712 ( .A(p_input[183]), .B(n2743), .Z(n2746) );
  XOR U2713 ( .A(n2743), .B(p_input[167]), .Z(n2745) );
  XOR U2714 ( .A(n2747), .B(n2748), .Z(n2743) );
  AND U2715 ( .A(n2749), .B(n2750), .Z(n2748) );
  XNOR U2716 ( .A(p_input[182]), .B(n2747), .Z(n2750) );
  XOR U2717 ( .A(n2747), .B(p_input[166]), .Z(n2749) );
  XOR U2718 ( .A(n2751), .B(n2752), .Z(n2747) );
  AND U2719 ( .A(n2753), .B(n2754), .Z(n2752) );
  XNOR U2720 ( .A(p_input[181]), .B(n2751), .Z(n2754) );
  XOR U2721 ( .A(n2751), .B(p_input[165]), .Z(n2753) );
  XOR U2722 ( .A(n2755), .B(n2756), .Z(n2751) );
  AND U2723 ( .A(n2757), .B(n2758), .Z(n2756) );
  XNOR U2724 ( .A(p_input[180]), .B(n2755), .Z(n2758) );
  XOR U2725 ( .A(n2755), .B(p_input[164]), .Z(n2757) );
  XOR U2726 ( .A(n2759), .B(n2760), .Z(n2755) );
  AND U2727 ( .A(n2761), .B(n2762), .Z(n2760) );
  XNOR U2728 ( .A(p_input[179]), .B(n2759), .Z(n2762) );
  XOR U2729 ( .A(n2759), .B(p_input[163]), .Z(n2761) );
  XOR U2730 ( .A(n2763), .B(n2764), .Z(n2759) );
  AND U2731 ( .A(n2765), .B(n2766), .Z(n2764) );
  XNOR U2732 ( .A(p_input[178]), .B(n2763), .Z(n2766) );
  XOR U2733 ( .A(n2763), .B(p_input[162]), .Z(n2765) );
  XNOR U2734 ( .A(n2767), .B(n2768), .Z(n2763) );
  AND U2735 ( .A(n2769), .B(n2770), .Z(n2768) );
  XOR U2736 ( .A(p_input[177]), .B(n2767), .Z(n2770) );
  XNOR U2737 ( .A(p_input[161]), .B(n2767), .Z(n2769) );
  AND U2738 ( .A(p_input[176]), .B(n2771), .Z(n2767) );
  IV U2739 ( .A(p_input[160]), .Z(n2771) );
  XNOR U2740 ( .A(p_input[128]), .B(n2772), .Z(n2574) );
  AND U2741 ( .A(n150), .B(n2773), .Z(n2772) );
  XOR U2742 ( .A(p_input[144]), .B(p_input[128]), .Z(n2773) );
  XOR U2743 ( .A(n2774), .B(n2775), .Z(n150) );
  AND U2744 ( .A(n2776), .B(n2777), .Z(n2775) );
  XNOR U2745 ( .A(p_input[159]), .B(n2774), .Z(n2777) );
  XOR U2746 ( .A(n2774), .B(p_input[143]), .Z(n2776) );
  XOR U2747 ( .A(n2778), .B(n2779), .Z(n2774) );
  AND U2748 ( .A(n2780), .B(n2781), .Z(n2779) );
  XNOR U2749 ( .A(p_input[158]), .B(n2778), .Z(n2781) );
  XNOR U2750 ( .A(n2778), .B(n2588), .Z(n2780) );
  IV U2751 ( .A(p_input[142]), .Z(n2588) );
  XOR U2752 ( .A(n2782), .B(n2783), .Z(n2778) );
  AND U2753 ( .A(n2784), .B(n2785), .Z(n2783) );
  XNOR U2754 ( .A(p_input[157]), .B(n2782), .Z(n2785) );
  XNOR U2755 ( .A(n2782), .B(n2597), .Z(n2784) );
  IV U2756 ( .A(p_input[141]), .Z(n2597) );
  XOR U2757 ( .A(n2786), .B(n2787), .Z(n2782) );
  AND U2758 ( .A(n2788), .B(n2789), .Z(n2787) );
  XNOR U2759 ( .A(p_input[156]), .B(n2786), .Z(n2789) );
  XNOR U2760 ( .A(n2786), .B(n2606), .Z(n2788) );
  IV U2761 ( .A(p_input[140]), .Z(n2606) );
  XOR U2762 ( .A(n2790), .B(n2791), .Z(n2786) );
  AND U2763 ( .A(n2792), .B(n2793), .Z(n2791) );
  XNOR U2764 ( .A(p_input[155]), .B(n2790), .Z(n2793) );
  XNOR U2765 ( .A(n2790), .B(n2615), .Z(n2792) );
  IV U2766 ( .A(p_input[139]), .Z(n2615) );
  XOR U2767 ( .A(n2794), .B(n2795), .Z(n2790) );
  AND U2768 ( .A(n2796), .B(n2797), .Z(n2795) );
  XNOR U2769 ( .A(p_input[154]), .B(n2794), .Z(n2797) );
  XNOR U2770 ( .A(n2794), .B(n2624), .Z(n2796) );
  IV U2771 ( .A(p_input[138]), .Z(n2624) );
  XOR U2772 ( .A(n2798), .B(n2799), .Z(n2794) );
  AND U2773 ( .A(n2800), .B(n2801), .Z(n2799) );
  XNOR U2774 ( .A(p_input[153]), .B(n2798), .Z(n2801) );
  XNOR U2775 ( .A(n2798), .B(n2633), .Z(n2800) );
  IV U2776 ( .A(p_input[137]), .Z(n2633) );
  XOR U2777 ( .A(n2802), .B(n2803), .Z(n2798) );
  AND U2778 ( .A(n2804), .B(n2805), .Z(n2803) );
  XNOR U2779 ( .A(p_input[152]), .B(n2802), .Z(n2805) );
  XNOR U2780 ( .A(n2802), .B(n2642), .Z(n2804) );
  IV U2781 ( .A(p_input[136]), .Z(n2642) );
  XOR U2782 ( .A(n2806), .B(n2807), .Z(n2802) );
  AND U2783 ( .A(n2808), .B(n2809), .Z(n2807) );
  XNOR U2784 ( .A(p_input[151]), .B(n2806), .Z(n2809) );
  XNOR U2785 ( .A(n2806), .B(n2651), .Z(n2808) );
  IV U2786 ( .A(p_input[135]), .Z(n2651) );
  XOR U2787 ( .A(n2810), .B(n2811), .Z(n2806) );
  AND U2788 ( .A(n2812), .B(n2813), .Z(n2811) );
  XNOR U2789 ( .A(p_input[150]), .B(n2810), .Z(n2813) );
  XNOR U2790 ( .A(n2810), .B(n2660), .Z(n2812) );
  IV U2791 ( .A(p_input[134]), .Z(n2660) );
  XOR U2792 ( .A(n2814), .B(n2815), .Z(n2810) );
  AND U2793 ( .A(n2816), .B(n2817), .Z(n2815) );
  XNOR U2794 ( .A(p_input[149]), .B(n2814), .Z(n2817) );
  XNOR U2795 ( .A(n2814), .B(n2669), .Z(n2816) );
  IV U2796 ( .A(p_input[133]), .Z(n2669) );
  XOR U2797 ( .A(n2818), .B(n2819), .Z(n2814) );
  AND U2798 ( .A(n2820), .B(n2821), .Z(n2819) );
  XNOR U2799 ( .A(p_input[148]), .B(n2818), .Z(n2821) );
  XNOR U2800 ( .A(n2818), .B(n2678), .Z(n2820) );
  IV U2801 ( .A(p_input[132]), .Z(n2678) );
  XOR U2802 ( .A(n2822), .B(n2823), .Z(n2818) );
  AND U2803 ( .A(n2824), .B(n2825), .Z(n2823) );
  XNOR U2804 ( .A(p_input[147]), .B(n2822), .Z(n2825) );
  XNOR U2805 ( .A(n2822), .B(n2687), .Z(n2824) );
  IV U2806 ( .A(p_input[131]), .Z(n2687) );
  XOR U2807 ( .A(n2826), .B(n2827), .Z(n2822) );
  AND U2808 ( .A(n2828), .B(n2829), .Z(n2827) );
  XNOR U2809 ( .A(p_input[146]), .B(n2826), .Z(n2829) );
  XNOR U2810 ( .A(n2826), .B(n2696), .Z(n2828) );
  IV U2811 ( .A(p_input[130]), .Z(n2696) );
  XNOR U2812 ( .A(n2830), .B(n2831), .Z(n2826) );
  AND U2813 ( .A(n2832), .B(n2833), .Z(n2831) );
  XOR U2814 ( .A(p_input[145]), .B(n2830), .Z(n2833) );
  XNOR U2815 ( .A(p_input[129]), .B(n2830), .Z(n2832) );
  AND U2816 ( .A(p_input[144]), .B(n2834), .Z(n2830) );
  IV U2817 ( .A(p_input[128]), .Z(n2834) );
  XOR U2818 ( .A(n2835), .B(n2836), .Z(n1950) );
  AND U2819 ( .A(n162), .B(n2837), .Z(n2836) );
  XNOR U2820 ( .A(n2838), .B(n2835), .Z(n2837) );
  XOR U2821 ( .A(n2839), .B(n2840), .Z(n162) );
  AND U2822 ( .A(n2841), .B(n2842), .Z(n2840) );
  XNOR U2823 ( .A(n1962), .B(n2839), .Z(n2842) );
  AND U2824 ( .A(n2843), .B(n2844), .Z(n1962) );
  XOR U2825 ( .A(n2839), .B(n1961), .Z(n2841) );
  AND U2826 ( .A(n2845), .B(n2846), .Z(n1961) );
  XOR U2827 ( .A(n2847), .B(n2848), .Z(n2839) );
  AND U2828 ( .A(n2849), .B(n2850), .Z(n2848) );
  XOR U2829 ( .A(n2847), .B(n1974), .Z(n2850) );
  XOR U2830 ( .A(n2851), .B(n2852), .Z(n1974) );
  AND U2831 ( .A(n137), .B(n2853), .Z(n2852) );
  XOR U2832 ( .A(n2854), .B(n2851), .Z(n2853) );
  XNOR U2833 ( .A(n1971), .B(n2847), .Z(n2849) );
  XOR U2834 ( .A(n2855), .B(n2856), .Z(n1971) );
  AND U2835 ( .A(n134), .B(n2857), .Z(n2856) );
  XOR U2836 ( .A(n2858), .B(n2855), .Z(n2857) );
  XOR U2837 ( .A(n2859), .B(n2860), .Z(n2847) );
  AND U2838 ( .A(n2861), .B(n2862), .Z(n2860) );
  XOR U2839 ( .A(n2859), .B(n1986), .Z(n2862) );
  XOR U2840 ( .A(n2863), .B(n2864), .Z(n1986) );
  AND U2841 ( .A(n137), .B(n2865), .Z(n2864) );
  XOR U2842 ( .A(n2866), .B(n2863), .Z(n2865) );
  XNOR U2843 ( .A(n1983), .B(n2859), .Z(n2861) );
  XOR U2844 ( .A(n2867), .B(n2868), .Z(n1983) );
  AND U2845 ( .A(n134), .B(n2869), .Z(n2868) );
  XOR U2846 ( .A(n2870), .B(n2867), .Z(n2869) );
  XOR U2847 ( .A(n2871), .B(n2872), .Z(n2859) );
  AND U2848 ( .A(n2873), .B(n2874), .Z(n2872) );
  XOR U2849 ( .A(n2871), .B(n1998), .Z(n2874) );
  XOR U2850 ( .A(n2875), .B(n2876), .Z(n1998) );
  AND U2851 ( .A(n137), .B(n2877), .Z(n2876) );
  XOR U2852 ( .A(n2878), .B(n2875), .Z(n2877) );
  XNOR U2853 ( .A(n1995), .B(n2871), .Z(n2873) );
  XOR U2854 ( .A(n2879), .B(n2880), .Z(n1995) );
  AND U2855 ( .A(n134), .B(n2881), .Z(n2880) );
  XOR U2856 ( .A(n2882), .B(n2879), .Z(n2881) );
  XOR U2857 ( .A(n2883), .B(n2884), .Z(n2871) );
  AND U2858 ( .A(n2885), .B(n2886), .Z(n2884) );
  XOR U2859 ( .A(n2883), .B(n2010), .Z(n2886) );
  XOR U2860 ( .A(n2887), .B(n2888), .Z(n2010) );
  AND U2861 ( .A(n137), .B(n2889), .Z(n2888) );
  XOR U2862 ( .A(n2890), .B(n2887), .Z(n2889) );
  XNOR U2863 ( .A(n2007), .B(n2883), .Z(n2885) );
  XOR U2864 ( .A(n2891), .B(n2892), .Z(n2007) );
  AND U2865 ( .A(n134), .B(n2893), .Z(n2892) );
  XOR U2866 ( .A(n2894), .B(n2891), .Z(n2893) );
  XOR U2867 ( .A(n2895), .B(n2896), .Z(n2883) );
  AND U2868 ( .A(n2897), .B(n2898), .Z(n2896) );
  XOR U2869 ( .A(n2895), .B(n2022), .Z(n2898) );
  XOR U2870 ( .A(n2899), .B(n2900), .Z(n2022) );
  AND U2871 ( .A(n137), .B(n2901), .Z(n2900) );
  XOR U2872 ( .A(n2902), .B(n2899), .Z(n2901) );
  XNOR U2873 ( .A(n2019), .B(n2895), .Z(n2897) );
  XOR U2874 ( .A(n2903), .B(n2904), .Z(n2019) );
  AND U2875 ( .A(n134), .B(n2905), .Z(n2904) );
  XOR U2876 ( .A(n2906), .B(n2903), .Z(n2905) );
  XOR U2877 ( .A(n2907), .B(n2908), .Z(n2895) );
  AND U2878 ( .A(n2909), .B(n2910), .Z(n2908) );
  XOR U2879 ( .A(n2907), .B(n2034), .Z(n2910) );
  XOR U2880 ( .A(n2911), .B(n2912), .Z(n2034) );
  AND U2881 ( .A(n137), .B(n2913), .Z(n2912) );
  XOR U2882 ( .A(n2914), .B(n2911), .Z(n2913) );
  XNOR U2883 ( .A(n2031), .B(n2907), .Z(n2909) );
  XOR U2884 ( .A(n2915), .B(n2916), .Z(n2031) );
  AND U2885 ( .A(n134), .B(n2917), .Z(n2916) );
  XOR U2886 ( .A(n2918), .B(n2915), .Z(n2917) );
  XOR U2887 ( .A(n2919), .B(n2920), .Z(n2907) );
  AND U2888 ( .A(n2921), .B(n2922), .Z(n2920) );
  XOR U2889 ( .A(n2919), .B(n2046), .Z(n2922) );
  XOR U2890 ( .A(n2923), .B(n2924), .Z(n2046) );
  AND U2891 ( .A(n137), .B(n2925), .Z(n2924) );
  XOR U2892 ( .A(n2926), .B(n2923), .Z(n2925) );
  XNOR U2893 ( .A(n2043), .B(n2919), .Z(n2921) );
  XOR U2894 ( .A(n2927), .B(n2928), .Z(n2043) );
  AND U2895 ( .A(n134), .B(n2929), .Z(n2928) );
  XOR U2896 ( .A(n2930), .B(n2927), .Z(n2929) );
  XOR U2897 ( .A(n2931), .B(n2932), .Z(n2919) );
  AND U2898 ( .A(n2933), .B(n2934), .Z(n2932) );
  XOR U2899 ( .A(n2931), .B(n2058), .Z(n2934) );
  XOR U2900 ( .A(n2935), .B(n2936), .Z(n2058) );
  AND U2901 ( .A(n137), .B(n2937), .Z(n2936) );
  XOR U2902 ( .A(n2938), .B(n2935), .Z(n2937) );
  XNOR U2903 ( .A(n2055), .B(n2931), .Z(n2933) );
  XOR U2904 ( .A(n2939), .B(n2940), .Z(n2055) );
  AND U2905 ( .A(n134), .B(n2941), .Z(n2940) );
  XOR U2906 ( .A(n2942), .B(n2939), .Z(n2941) );
  XOR U2907 ( .A(n2943), .B(n2944), .Z(n2931) );
  AND U2908 ( .A(n2945), .B(n2946), .Z(n2944) );
  XOR U2909 ( .A(n2943), .B(n2070), .Z(n2946) );
  XOR U2910 ( .A(n2947), .B(n2948), .Z(n2070) );
  AND U2911 ( .A(n137), .B(n2949), .Z(n2948) );
  XOR U2912 ( .A(n2950), .B(n2947), .Z(n2949) );
  XNOR U2913 ( .A(n2067), .B(n2943), .Z(n2945) );
  XOR U2914 ( .A(n2951), .B(n2952), .Z(n2067) );
  AND U2915 ( .A(n134), .B(n2953), .Z(n2952) );
  XOR U2916 ( .A(n2954), .B(n2951), .Z(n2953) );
  XOR U2917 ( .A(n2955), .B(n2956), .Z(n2943) );
  AND U2918 ( .A(n2957), .B(n2958), .Z(n2956) );
  XOR U2919 ( .A(n2955), .B(n2082), .Z(n2958) );
  XOR U2920 ( .A(n2959), .B(n2960), .Z(n2082) );
  AND U2921 ( .A(n137), .B(n2961), .Z(n2960) );
  XOR U2922 ( .A(n2962), .B(n2959), .Z(n2961) );
  XNOR U2923 ( .A(n2079), .B(n2955), .Z(n2957) );
  XOR U2924 ( .A(n2963), .B(n2964), .Z(n2079) );
  AND U2925 ( .A(n134), .B(n2965), .Z(n2964) );
  XOR U2926 ( .A(n2966), .B(n2963), .Z(n2965) );
  XOR U2927 ( .A(n2967), .B(n2968), .Z(n2955) );
  AND U2928 ( .A(n2969), .B(n2970), .Z(n2968) );
  XOR U2929 ( .A(n2094), .B(n2967), .Z(n2970) );
  XOR U2930 ( .A(n2971), .B(n2972), .Z(n2094) );
  AND U2931 ( .A(n137), .B(n2973), .Z(n2972) );
  XOR U2932 ( .A(n2971), .B(n2974), .Z(n2973) );
  XNOR U2933 ( .A(n2967), .B(n2091), .Z(n2969) );
  XOR U2934 ( .A(n2975), .B(n2976), .Z(n2091) );
  AND U2935 ( .A(n134), .B(n2977), .Z(n2976) );
  XOR U2936 ( .A(n2975), .B(n2978), .Z(n2977) );
  XOR U2937 ( .A(n2979), .B(n2980), .Z(n2967) );
  AND U2938 ( .A(n2981), .B(n2982), .Z(n2980) );
  XOR U2939 ( .A(n2979), .B(n2106), .Z(n2982) );
  XOR U2940 ( .A(n2983), .B(n2984), .Z(n2106) );
  AND U2941 ( .A(n137), .B(n2985), .Z(n2984) );
  XOR U2942 ( .A(n2986), .B(n2983), .Z(n2985) );
  XNOR U2943 ( .A(n2103), .B(n2979), .Z(n2981) );
  XOR U2944 ( .A(n2987), .B(n2988), .Z(n2103) );
  AND U2945 ( .A(n134), .B(n2989), .Z(n2988) );
  XOR U2946 ( .A(n2990), .B(n2987), .Z(n2989) );
  XOR U2947 ( .A(n2991), .B(n2992), .Z(n2979) );
  AND U2948 ( .A(n2993), .B(n2994), .Z(n2992) );
  XOR U2949 ( .A(n2991), .B(n2118), .Z(n2994) );
  XOR U2950 ( .A(n2995), .B(n2996), .Z(n2118) );
  AND U2951 ( .A(n137), .B(n2997), .Z(n2996) );
  XOR U2952 ( .A(n2998), .B(n2995), .Z(n2997) );
  XNOR U2953 ( .A(n2115), .B(n2991), .Z(n2993) );
  XOR U2954 ( .A(n2999), .B(n3000), .Z(n2115) );
  AND U2955 ( .A(n134), .B(n3001), .Z(n3000) );
  XOR U2956 ( .A(n3002), .B(n2999), .Z(n3001) );
  XOR U2957 ( .A(n3003), .B(n3004), .Z(n2991) );
  AND U2958 ( .A(n3005), .B(n3006), .Z(n3004) );
  XNOR U2959 ( .A(n3007), .B(n2131), .Z(n3006) );
  XOR U2960 ( .A(n3008), .B(n3009), .Z(n2131) );
  AND U2961 ( .A(n137), .B(n3010), .Z(n3009) );
  XOR U2962 ( .A(n3011), .B(n3008), .Z(n3010) );
  XNOR U2963 ( .A(n2128), .B(n3003), .Z(n3005) );
  XOR U2964 ( .A(n3012), .B(n3013), .Z(n2128) );
  AND U2965 ( .A(n134), .B(n3014), .Z(n3013) );
  XOR U2966 ( .A(n3015), .B(n3012), .Z(n3014) );
  IV U2967 ( .A(n3007), .Z(n3003) );
  AND U2968 ( .A(n2835), .B(n2838), .Z(n3007) );
  XNOR U2969 ( .A(n3016), .B(n3017), .Z(n2838) );
  AND U2970 ( .A(n137), .B(n3018), .Z(n3017) );
  XNOR U2971 ( .A(n3019), .B(n3016), .Z(n3018) );
  XOR U2972 ( .A(n3020), .B(n3021), .Z(n137) );
  AND U2973 ( .A(n3022), .B(n3023), .Z(n3021) );
  XNOR U2974 ( .A(n2843), .B(n3020), .Z(n3023) );
  AND U2975 ( .A(p_input[127]), .B(p_input[111]), .Z(n2843) );
  XOR U2976 ( .A(n3020), .B(n2844), .Z(n3022) );
  AND U2977 ( .A(p_input[95]), .B(p_input[79]), .Z(n2844) );
  XOR U2978 ( .A(n3024), .B(n3025), .Z(n3020) );
  AND U2979 ( .A(n3026), .B(n3027), .Z(n3025) );
  XOR U2980 ( .A(n3024), .B(n2854), .Z(n3027) );
  XNOR U2981 ( .A(p_input[110]), .B(n3028), .Z(n2854) );
  AND U2982 ( .A(n173), .B(n3029), .Z(n3028) );
  XOR U2983 ( .A(p_input[126]), .B(p_input[110]), .Z(n3029) );
  XNOR U2984 ( .A(n2851), .B(n3024), .Z(n3026) );
  XOR U2985 ( .A(n3030), .B(n3031), .Z(n2851) );
  AND U2986 ( .A(n171), .B(n3032), .Z(n3031) );
  XOR U2987 ( .A(p_input[94]), .B(p_input[78]), .Z(n3032) );
  XOR U2988 ( .A(n3033), .B(n3034), .Z(n3024) );
  AND U2989 ( .A(n3035), .B(n3036), .Z(n3034) );
  XOR U2990 ( .A(n3033), .B(n2866), .Z(n3036) );
  XNOR U2991 ( .A(p_input[109]), .B(n3037), .Z(n2866) );
  AND U2992 ( .A(n173), .B(n3038), .Z(n3037) );
  XOR U2993 ( .A(p_input[125]), .B(p_input[109]), .Z(n3038) );
  XNOR U2994 ( .A(n2863), .B(n3033), .Z(n3035) );
  XOR U2995 ( .A(n3039), .B(n3040), .Z(n2863) );
  AND U2996 ( .A(n171), .B(n3041), .Z(n3040) );
  XOR U2997 ( .A(p_input[93]), .B(p_input[77]), .Z(n3041) );
  XOR U2998 ( .A(n3042), .B(n3043), .Z(n3033) );
  AND U2999 ( .A(n3044), .B(n3045), .Z(n3043) );
  XOR U3000 ( .A(n3042), .B(n2878), .Z(n3045) );
  XNOR U3001 ( .A(p_input[108]), .B(n3046), .Z(n2878) );
  AND U3002 ( .A(n173), .B(n3047), .Z(n3046) );
  XOR U3003 ( .A(p_input[124]), .B(p_input[108]), .Z(n3047) );
  XNOR U3004 ( .A(n2875), .B(n3042), .Z(n3044) );
  XOR U3005 ( .A(n3048), .B(n3049), .Z(n2875) );
  AND U3006 ( .A(n171), .B(n3050), .Z(n3049) );
  XOR U3007 ( .A(p_input[92]), .B(p_input[76]), .Z(n3050) );
  XOR U3008 ( .A(n3051), .B(n3052), .Z(n3042) );
  AND U3009 ( .A(n3053), .B(n3054), .Z(n3052) );
  XOR U3010 ( .A(n3051), .B(n2890), .Z(n3054) );
  XNOR U3011 ( .A(p_input[107]), .B(n3055), .Z(n2890) );
  AND U3012 ( .A(n173), .B(n3056), .Z(n3055) );
  XOR U3013 ( .A(p_input[123]), .B(p_input[107]), .Z(n3056) );
  XNOR U3014 ( .A(n2887), .B(n3051), .Z(n3053) );
  XOR U3015 ( .A(n3057), .B(n3058), .Z(n2887) );
  AND U3016 ( .A(n171), .B(n3059), .Z(n3058) );
  XOR U3017 ( .A(p_input[91]), .B(p_input[75]), .Z(n3059) );
  XOR U3018 ( .A(n3060), .B(n3061), .Z(n3051) );
  AND U3019 ( .A(n3062), .B(n3063), .Z(n3061) );
  XOR U3020 ( .A(n3060), .B(n2902), .Z(n3063) );
  XNOR U3021 ( .A(p_input[106]), .B(n3064), .Z(n2902) );
  AND U3022 ( .A(n173), .B(n3065), .Z(n3064) );
  XOR U3023 ( .A(p_input[122]), .B(p_input[106]), .Z(n3065) );
  XNOR U3024 ( .A(n2899), .B(n3060), .Z(n3062) );
  XOR U3025 ( .A(n3066), .B(n3067), .Z(n2899) );
  AND U3026 ( .A(n171), .B(n3068), .Z(n3067) );
  XOR U3027 ( .A(p_input[90]), .B(p_input[74]), .Z(n3068) );
  XOR U3028 ( .A(n3069), .B(n3070), .Z(n3060) );
  AND U3029 ( .A(n3071), .B(n3072), .Z(n3070) );
  XOR U3030 ( .A(n3069), .B(n2914), .Z(n3072) );
  XNOR U3031 ( .A(p_input[105]), .B(n3073), .Z(n2914) );
  AND U3032 ( .A(n173), .B(n3074), .Z(n3073) );
  XOR U3033 ( .A(p_input[121]), .B(p_input[105]), .Z(n3074) );
  XNOR U3034 ( .A(n2911), .B(n3069), .Z(n3071) );
  XOR U3035 ( .A(n3075), .B(n3076), .Z(n2911) );
  AND U3036 ( .A(n171), .B(n3077), .Z(n3076) );
  XOR U3037 ( .A(p_input[89]), .B(p_input[73]), .Z(n3077) );
  XOR U3038 ( .A(n3078), .B(n3079), .Z(n3069) );
  AND U3039 ( .A(n3080), .B(n3081), .Z(n3079) );
  XOR U3040 ( .A(n3078), .B(n2926), .Z(n3081) );
  XNOR U3041 ( .A(p_input[104]), .B(n3082), .Z(n2926) );
  AND U3042 ( .A(n173), .B(n3083), .Z(n3082) );
  XOR U3043 ( .A(p_input[120]), .B(p_input[104]), .Z(n3083) );
  XNOR U3044 ( .A(n2923), .B(n3078), .Z(n3080) );
  XOR U3045 ( .A(n3084), .B(n3085), .Z(n2923) );
  AND U3046 ( .A(n171), .B(n3086), .Z(n3085) );
  XOR U3047 ( .A(p_input[88]), .B(p_input[72]), .Z(n3086) );
  XOR U3048 ( .A(n3087), .B(n3088), .Z(n3078) );
  AND U3049 ( .A(n3089), .B(n3090), .Z(n3088) );
  XOR U3050 ( .A(n3087), .B(n2938), .Z(n3090) );
  XNOR U3051 ( .A(p_input[103]), .B(n3091), .Z(n2938) );
  AND U3052 ( .A(n173), .B(n3092), .Z(n3091) );
  XOR U3053 ( .A(p_input[119]), .B(p_input[103]), .Z(n3092) );
  XNOR U3054 ( .A(n2935), .B(n3087), .Z(n3089) );
  XOR U3055 ( .A(n3093), .B(n3094), .Z(n2935) );
  AND U3056 ( .A(n171), .B(n3095), .Z(n3094) );
  XOR U3057 ( .A(p_input[87]), .B(p_input[71]), .Z(n3095) );
  XOR U3058 ( .A(n3096), .B(n3097), .Z(n3087) );
  AND U3059 ( .A(n3098), .B(n3099), .Z(n3097) );
  XOR U3060 ( .A(n3096), .B(n2950), .Z(n3099) );
  XNOR U3061 ( .A(p_input[102]), .B(n3100), .Z(n2950) );
  AND U3062 ( .A(n173), .B(n3101), .Z(n3100) );
  XOR U3063 ( .A(p_input[118]), .B(p_input[102]), .Z(n3101) );
  XNOR U3064 ( .A(n2947), .B(n3096), .Z(n3098) );
  XOR U3065 ( .A(n3102), .B(n3103), .Z(n2947) );
  AND U3066 ( .A(n171), .B(n3104), .Z(n3103) );
  XOR U3067 ( .A(p_input[86]), .B(p_input[70]), .Z(n3104) );
  XOR U3068 ( .A(n3105), .B(n3106), .Z(n3096) );
  AND U3069 ( .A(n3107), .B(n3108), .Z(n3106) );
  XOR U3070 ( .A(n3105), .B(n2962), .Z(n3108) );
  XNOR U3071 ( .A(p_input[101]), .B(n3109), .Z(n2962) );
  AND U3072 ( .A(n173), .B(n3110), .Z(n3109) );
  XOR U3073 ( .A(p_input[117]), .B(p_input[101]), .Z(n3110) );
  XNOR U3074 ( .A(n2959), .B(n3105), .Z(n3107) );
  XOR U3075 ( .A(n3111), .B(n3112), .Z(n2959) );
  AND U3076 ( .A(n171), .B(n3113), .Z(n3112) );
  XOR U3077 ( .A(p_input[85]), .B(p_input[69]), .Z(n3113) );
  XOR U3078 ( .A(n3114), .B(n3115), .Z(n3105) );
  AND U3079 ( .A(n3116), .B(n3117), .Z(n3115) );
  XOR U3080 ( .A(n2974), .B(n3114), .Z(n3117) );
  XNOR U3081 ( .A(p_input[100]), .B(n3118), .Z(n2974) );
  AND U3082 ( .A(n173), .B(n3119), .Z(n3118) );
  XOR U3083 ( .A(p_input[116]), .B(p_input[100]), .Z(n3119) );
  XNOR U3084 ( .A(n3114), .B(n2971), .Z(n3116) );
  XOR U3085 ( .A(n3120), .B(n3121), .Z(n2971) );
  AND U3086 ( .A(n171), .B(n3122), .Z(n3121) );
  XOR U3087 ( .A(p_input[84]), .B(p_input[68]), .Z(n3122) );
  XOR U3088 ( .A(n3123), .B(n3124), .Z(n3114) );
  AND U3089 ( .A(n3125), .B(n3126), .Z(n3124) );
  XOR U3090 ( .A(n3123), .B(n2986), .Z(n3126) );
  XNOR U3091 ( .A(p_input[99]), .B(n3127), .Z(n2986) );
  AND U3092 ( .A(n173), .B(n3128), .Z(n3127) );
  XOR U3093 ( .A(p_input[99]), .B(p_input[115]), .Z(n3128) );
  XNOR U3094 ( .A(n2983), .B(n3123), .Z(n3125) );
  XOR U3095 ( .A(n3129), .B(n3130), .Z(n2983) );
  AND U3096 ( .A(n171), .B(n3131), .Z(n3130) );
  XOR U3097 ( .A(p_input[83]), .B(p_input[67]), .Z(n3131) );
  XOR U3098 ( .A(n3132), .B(n3133), .Z(n3123) );
  AND U3099 ( .A(n3134), .B(n3135), .Z(n3133) );
  XOR U3100 ( .A(n3132), .B(n2998), .Z(n3135) );
  XNOR U3101 ( .A(p_input[98]), .B(n3136), .Z(n2998) );
  AND U3102 ( .A(n173), .B(n3137), .Z(n3136) );
  XOR U3103 ( .A(p_input[98]), .B(p_input[114]), .Z(n3137) );
  XNOR U3104 ( .A(n2995), .B(n3132), .Z(n3134) );
  XOR U3105 ( .A(n3138), .B(n3139), .Z(n2995) );
  AND U3106 ( .A(n171), .B(n3140), .Z(n3139) );
  XOR U3107 ( .A(p_input[82]), .B(p_input[66]), .Z(n3140) );
  XOR U3108 ( .A(n3141), .B(n3142), .Z(n3132) );
  AND U3109 ( .A(n3143), .B(n3144), .Z(n3142) );
  XNOR U3110 ( .A(n3145), .B(n3011), .Z(n3144) );
  XNOR U3111 ( .A(p_input[97]), .B(n3146), .Z(n3011) );
  AND U3112 ( .A(n173), .B(n3147), .Z(n3146) );
  XNOR U3113 ( .A(n3148), .B(p_input[113]), .Z(n3147) );
  IV U3114 ( .A(p_input[97]), .Z(n3148) );
  XNOR U3115 ( .A(n3008), .B(n3141), .Z(n3143) );
  XNOR U3116 ( .A(p_input[65]), .B(n3149), .Z(n3008) );
  AND U3117 ( .A(n171), .B(n3150), .Z(n3149) );
  XOR U3118 ( .A(p_input[81]), .B(p_input[65]), .Z(n3150) );
  IV U3119 ( .A(n3145), .Z(n3141) );
  AND U3120 ( .A(n3016), .B(n3019), .Z(n3145) );
  XOR U3121 ( .A(p_input[96]), .B(n3151), .Z(n3019) );
  AND U3122 ( .A(n173), .B(n3152), .Z(n3151) );
  XOR U3123 ( .A(p_input[96]), .B(p_input[112]), .Z(n3152) );
  XOR U3124 ( .A(n3153), .B(n3154), .Z(n173) );
  AND U3125 ( .A(n3155), .B(n3156), .Z(n3154) );
  XNOR U3126 ( .A(p_input[127]), .B(n3153), .Z(n3156) );
  XOR U3127 ( .A(n3153), .B(p_input[111]), .Z(n3155) );
  XOR U3128 ( .A(n3157), .B(n3158), .Z(n3153) );
  AND U3129 ( .A(n3159), .B(n3160), .Z(n3158) );
  XNOR U3130 ( .A(p_input[126]), .B(n3157), .Z(n3160) );
  XOR U3131 ( .A(n3157), .B(p_input[110]), .Z(n3159) );
  XOR U3132 ( .A(n3161), .B(n3162), .Z(n3157) );
  AND U3133 ( .A(n3163), .B(n3164), .Z(n3162) );
  XNOR U3134 ( .A(p_input[125]), .B(n3161), .Z(n3164) );
  XOR U3135 ( .A(n3161), .B(p_input[109]), .Z(n3163) );
  XOR U3136 ( .A(n3165), .B(n3166), .Z(n3161) );
  AND U3137 ( .A(n3167), .B(n3168), .Z(n3166) );
  XNOR U3138 ( .A(p_input[124]), .B(n3165), .Z(n3168) );
  XOR U3139 ( .A(n3165), .B(p_input[108]), .Z(n3167) );
  XOR U3140 ( .A(n3169), .B(n3170), .Z(n3165) );
  AND U3141 ( .A(n3171), .B(n3172), .Z(n3170) );
  XNOR U3142 ( .A(p_input[123]), .B(n3169), .Z(n3172) );
  XOR U3143 ( .A(n3169), .B(p_input[107]), .Z(n3171) );
  XOR U3144 ( .A(n3173), .B(n3174), .Z(n3169) );
  AND U3145 ( .A(n3175), .B(n3176), .Z(n3174) );
  XNOR U3146 ( .A(p_input[122]), .B(n3173), .Z(n3176) );
  XOR U3147 ( .A(n3173), .B(p_input[106]), .Z(n3175) );
  XOR U3148 ( .A(n3177), .B(n3178), .Z(n3173) );
  AND U3149 ( .A(n3179), .B(n3180), .Z(n3178) );
  XNOR U3150 ( .A(p_input[121]), .B(n3177), .Z(n3180) );
  XOR U3151 ( .A(n3177), .B(p_input[105]), .Z(n3179) );
  XOR U3152 ( .A(n3181), .B(n3182), .Z(n3177) );
  AND U3153 ( .A(n3183), .B(n3184), .Z(n3182) );
  XNOR U3154 ( .A(p_input[120]), .B(n3181), .Z(n3184) );
  XOR U3155 ( .A(n3181), .B(p_input[104]), .Z(n3183) );
  XOR U3156 ( .A(n3185), .B(n3186), .Z(n3181) );
  AND U3157 ( .A(n3187), .B(n3188), .Z(n3186) );
  XNOR U3158 ( .A(p_input[119]), .B(n3185), .Z(n3188) );
  XOR U3159 ( .A(n3185), .B(p_input[103]), .Z(n3187) );
  XOR U3160 ( .A(n3189), .B(n3190), .Z(n3185) );
  AND U3161 ( .A(n3191), .B(n3192), .Z(n3190) );
  XNOR U3162 ( .A(p_input[118]), .B(n3189), .Z(n3192) );
  XOR U3163 ( .A(n3189), .B(p_input[102]), .Z(n3191) );
  XOR U3164 ( .A(n3193), .B(n3194), .Z(n3189) );
  AND U3165 ( .A(n3195), .B(n3196), .Z(n3194) );
  XNOR U3166 ( .A(p_input[117]), .B(n3193), .Z(n3196) );
  XOR U3167 ( .A(n3193), .B(p_input[101]), .Z(n3195) );
  XOR U3168 ( .A(n3197), .B(n3198), .Z(n3193) );
  AND U3169 ( .A(n3199), .B(n3200), .Z(n3198) );
  XNOR U3170 ( .A(p_input[116]), .B(n3197), .Z(n3200) );
  XOR U3171 ( .A(n3197), .B(p_input[100]), .Z(n3199) );
  XOR U3172 ( .A(n3201), .B(n3202), .Z(n3197) );
  AND U3173 ( .A(n3203), .B(n3204), .Z(n3202) );
  XNOR U3174 ( .A(p_input[115]), .B(n3201), .Z(n3204) );
  XOR U3175 ( .A(n3201), .B(p_input[99]), .Z(n3203) );
  XOR U3176 ( .A(n3205), .B(n3206), .Z(n3201) );
  AND U3177 ( .A(n3207), .B(n3208), .Z(n3206) );
  XNOR U3178 ( .A(p_input[114]), .B(n3205), .Z(n3208) );
  XOR U3179 ( .A(n3205), .B(p_input[98]), .Z(n3207) );
  XNOR U3180 ( .A(n3209), .B(n3210), .Z(n3205) );
  AND U3181 ( .A(n3211), .B(n3212), .Z(n3210) );
  XOR U3182 ( .A(p_input[113]), .B(n3209), .Z(n3212) );
  XNOR U3183 ( .A(p_input[97]), .B(n3209), .Z(n3211) );
  AND U3184 ( .A(p_input[112]), .B(n3213), .Z(n3209) );
  IV U3185 ( .A(p_input[96]), .Z(n3213) );
  XNOR U3186 ( .A(p_input[64]), .B(n3214), .Z(n3016) );
  AND U3187 ( .A(n171), .B(n3215), .Z(n3214) );
  XOR U3188 ( .A(p_input[80]), .B(p_input[64]), .Z(n3215) );
  XOR U3189 ( .A(n3216), .B(n3217), .Z(n171) );
  AND U3190 ( .A(n3218), .B(n3219), .Z(n3217) );
  XNOR U3191 ( .A(p_input[95]), .B(n3216), .Z(n3219) );
  XOR U3192 ( .A(n3216), .B(p_input[79]), .Z(n3218) );
  XOR U3193 ( .A(n3220), .B(n3221), .Z(n3216) );
  AND U3194 ( .A(n3222), .B(n3223), .Z(n3221) );
  XNOR U3195 ( .A(p_input[94]), .B(n3220), .Z(n3223) );
  XNOR U3196 ( .A(n3220), .B(n3030), .Z(n3222) );
  IV U3197 ( .A(p_input[78]), .Z(n3030) );
  XOR U3198 ( .A(n3224), .B(n3225), .Z(n3220) );
  AND U3199 ( .A(n3226), .B(n3227), .Z(n3225) );
  XNOR U3200 ( .A(p_input[93]), .B(n3224), .Z(n3227) );
  XNOR U3201 ( .A(n3224), .B(n3039), .Z(n3226) );
  IV U3202 ( .A(p_input[77]), .Z(n3039) );
  XOR U3203 ( .A(n3228), .B(n3229), .Z(n3224) );
  AND U3204 ( .A(n3230), .B(n3231), .Z(n3229) );
  XNOR U3205 ( .A(p_input[92]), .B(n3228), .Z(n3231) );
  XNOR U3206 ( .A(n3228), .B(n3048), .Z(n3230) );
  IV U3207 ( .A(p_input[76]), .Z(n3048) );
  XOR U3208 ( .A(n3232), .B(n3233), .Z(n3228) );
  AND U3209 ( .A(n3234), .B(n3235), .Z(n3233) );
  XNOR U3210 ( .A(p_input[91]), .B(n3232), .Z(n3235) );
  XNOR U3211 ( .A(n3232), .B(n3057), .Z(n3234) );
  IV U3212 ( .A(p_input[75]), .Z(n3057) );
  XOR U3213 ( .A(n3236), .B(n3237), .Z(n3232) );
  AND U3214 ( .A(n3238), .B(n3239), .Z(n3237) );
  XNOR U3215 ( .A(p_input[90]), .B(n3236), .Z(n3239) );
  XNOR U3216 ( .A(n3236), .B(n3066), .Z(n3238) );
  IV U3217 ( .A(p_input[74]), .Z(n3066) );
  XOR U3218 ( .A(n3240), .B(n3241), .Z(n3236) );
  AND U3219 ( .A(n3242), .B(n3243), .Z(n3241) );
  XNOR U3220 ( .A(p_input[89]), .B(n3240), .Z(n3243) );
  XNOR U3221 ( .A(n3240), .B(n3075), .Z(n3242) );
  IV U3222 ( .A(p_input[73]), .Z(n3075) );
  XOR U3223 ( .A(n3244), .B(n3245), .Z(n3240) );
  AND U3224 ( .A(n3246), .B(n3247), .Z(n3245) );
  XNOR U3225 ( .A(p_input[88]), .B(n3244), .Z(n3247) );
  XNOR U3226 ( .A(n3244), .B(n3084), .Z(n3246) );
  IV U3227 ( .A(p_input[72]), .Z(n3084) );
  XOR U3228 ( .A(n3248), .B(n3249), .Z(n3244) );
  AND U3229 ( .A(n3250), .B(n3251), .Z(n3249) );
  XNOR U3230 ( .A(p_input[87]), .B(n3248), .Z(n3251) );
  XNOR U3231 ( .A(n3248), .B(n3093), .Z(n3250) );
  IV U3232 ( .A(p_input[71]), .Z(n3093) );
  XOR U3233 ( .A(n3252), .B(n3253), .Z(n3248) );
  AND U3234 ( .A(n3254), .B(n3255), .Z(n3253) );
  XNOR U3235 ( .A(p_input[86]), .B(n3252), .Z(n3255) );
  XNOR U3236 ( .A(n3252), .B(n3102), .Z(n3254) );
  IV U3237 ( .A(p_input[70]), .Z(n3102) );
  XOR U3238 ( .A(n3256), .B(n3257), .Z(n3252) );
  AND U3239 ( .A(n3258), .B(n3259), .Z(n3257) );
  XNOR U3240 ( .A(p_input[85]), .B(n3256), .Z(n3259) );
  XNOR U3241 ( .A(n3256), .B(n3111), .Z(n3258) );
  IV U3242 ( .A(p_input[69]), .Z(n3111) );
  XOR U3243 ( .A(n3260), .B(n3261), .Z(n3256) );
  AND U3244 ( .A(n3262), .B(n3263), .Z(n3261) );
  XNOR U3245 ( .A(p_input[84]), .B(n3260), .Z(n3263) );
  XNOR U3246 ( .A(n3260), .B(n3120), .Z(n3262) );
  IV U3247 ( .A(p_input[68]), .Z(n3120) );
  XOR U3248 ( .A(n3264), .B(n3265), .Z(n3260) );
  AND U3249 ( .A(n3266), .B(n3267), .Z(n3265) );
  XNOR U3250 ( .A(p_input[83]), .B(n3264), .Z(n3267) );
  XNOR U3251 ( .A(n3264), .B(n3129), .Z(n3266) );
  IV U3252 ( .A(p_input[67]), .Z(n3129) );
  XOR U3253 ( .A(n3268), .B(n3269), .Z(n3264) );
  AND U3254 ( .A(n3270), .B(n3271), .Z(n3269) );
  XNOR U3255 ( .A(p_input[82]), .B(n3268), .Z(n3271) );
  XNOR U3256 ( .A(n3268), .B(n3138), .Z(n3270) );
  IV U3257 ( .A(p_input[66]), .Z(n3138) );
  XNOR U3258 ( .A(n3272), .B(n3273), .Z(n3268) );
  AND U3259 ( .A(n3274), .B(n3275), .Z(n3273) );
  XOR U3260 ( .A(p_input[81]), .B(n3272), .Z(n3275) );
  XNOR U3261 ( .A(p_input[65]), .B(n3272), .Z(n3274) );
  AND U3262 ( .A(p_input[80]), .B(n3276), .Z(n3272) );
  IV U3263 ( .A(p_input[64]), .Z(n3276) );
  XOR U3264 ( .A(n3277), .B(n3278), .Z(n2835) );
  AND U3265 ( .A(n134), .B(n3279), .Z(n3278) );
  XNOR U3266 ( .A(n3280), .B(n3277), .Z(n3279) );
  XOR U3267 ( .A(n3281), .B(n3282), .Z(n134) );
  AND U3268 ( .A(n3283), .B(n3284), .Z(n3282) );
  XNOR U3269 ( .A(n2846), .B(n3281), .Z(n3284) );
  AND U3270 ( .A(p_input[63]), .B(p_input[47]), .Z(n2846) );
  XOR U3271 ( .A(n3281), .B(n2845), .Z(n3283) );
  AND U3272 ( .A(p_input[15]), .B(p_input[31]), .Z(n2845) );
  XOR U3273 ( .A(n3285), .B(n3286), .Z(n3281) );
  AND U3274 ( .A(n3287), .B(n3288), .Z(n3286) );
  XOR U3275 ( .A(n3285), .B(n2858), .Z(n3288) );
  XNOR U3276 ( .A(p_input[46]), .B(n3289), .Z(n2858) );
  AND U3277 ( .A(n181), .B(n3290), .Z(n3289) );
  XOR U3278 ( .A(p_input[62]), .B(p_input[46]), .Z(n3290) );
  XNOR U3279 ( .A(n2855), .B(n3285), .Z(n3287) );
  XOR U3280 ( .A(n3291), .B(n3292), .Z(n2855) );
  AND U3281 ( .A(n178), .B(n3293), .Z(n3292) );
  XOR U3282 ( .A(p_input[30]), .B(p_input[14]), .Z(n3293) );
  XOR U3283 ( .A(n3294), .B(n3295), .Z(n3285) );
  AND U3284 ( .A(n3296), .B(n3297), .Z(n3295) );
  XOR U3285 ( .A(n3294), .B(n2870), .Z(n3297) );
  XNOR U3286 ( .A(p_input[45]), .B(n3298), .Z(n2870) );
  AND U3287 ( .A(n181), .B(n3299), .Z(n3298) );
  XOR U3288 ( .A(p_input[61]), .B(p_input[45]), .Z(n3299) );
  XNOR U3289 ( .A(n2867), .B(n3294), .Z(n3296) );
  XOR U3290 ( .A(n3300), .B(n3301), .Z(n2867) );
  AND U3291 ( .A(n178), .B(n3302), .Z(n3301) );
  XOR U3292 ( .A(p_input[29]), .B(p_input[13]), .Z(n3302) );
  XOR U3293 ( .A(n3303), .B(n3304), .Z(n3294) );
  AND U3294 ( .A(n3305), .B(n3306), .Z(n3304) );
  XOR U3295 ( .A(n3303), .B(n2882), .Z(n3306) );
  XNOR U3296 ( .A(p_input[44]), .B(n3307), .Z(n2882) );
  AND U3297 ( .A(n181), .B(n3308), .Z(n3307) );
  XOR U3298 ( .A(p_input[60]), .B(p_input[44]), .Z(n3308) );
  XNOR U3299 ( .A(n2879), .B(n3303), .Z(n3305) );
  XOR U3300 ( .A(n3309), .B(n3310), .Z(n2879) );
  AND U3301 ( .A(n178), .B(n3311), .Z(n3310) );
  XOR U3302 ( .A(p_input[28]), .B(p_input[12]), .Z(n3311) );
  XOR U3303 ( .A(n3312), .B(n3313), .Z(n3303) );
  AND U3304 ( .A(n3314), .B(n3315), .Z(n3313) );
  XOR U3305 ( .A(n3312), .B(n2894), .Z(n3315) );
  XNOR U3306 ( .A(p_input[43]), .B(n3316), .Z(n2894) );
  AND U3307 ( .A(n181), .B(n3317), .Z(n3316) );
  XOR U3308 ( .A(p_input[59]), .B(p_input[43]), .Z(n3317) );
  XNOR U3309 ( .A(n2891), .B(n3312), .Z(n3314) );
  XOR U3310 ( .A(n3318), .B(n3319), .Z(n2891) );
  AND U3311 ( .A(n178), .B(n3320), .Z(n3319) );
  XOR U3312 ( .A(p_input[27]), .B(p_input[11]), .Z(n3320) );
  XOR U3313 ( .A(n3321), .B(n3322), .Z(n3312) );
  AND U3314 ( .A(n3323), .B(n3324), .Z(n3322) );
  XOR U3315 ( .A(n3321), .B(n2906), .Z(n3324) );
  XNOR U3316 ( .A(p_input[42]), .B(n3325), .Z(n2906) );
  AND U3317 ( .A(n181), .B(n3326), .Z(n3325) );
  XOR U3318 ( .A(p_input[58]), .B(p_input[42]), .Z(n3326) );
  XNOR U3319 ( .A(n2903), .B(n3321), .Z(n3323) );
  XOR U3320 ( .A(n3327), .B(n3328), .Z(n2903) );
  AND U3321 ( .A(n178), .B(n3329), .Z(n3328) );
  XOR U3322 ( .A(p_input[26]), .B(p_input[10]), .Z(n3329) );
  XOR U3323 ( .A(n3330), .B(n3331), .Z(n3321) );
  AND U3324 ( .A(n3332), .B(n3333), .Z(n3331) );
  XOR U3325 ( .A(n3330), .B(n2918), .Z(n3333) );
  XNOR U3326 ( .A(p_input[41]), .B(n3334), .Z(n2918) );
  AND U3327 ( .A(n181), .B(n3335), .Z(n3334) );
  XOR U3328 ( .A(p_input[57]), .B(p_input[41]), .Z(n3335) );
  XNOR U3329 ( .A(n2915), .B(n3330), .Z(n3332) );
  XOR U3330 ( .A(n3336), .B(n3337), .Z(n2915) );
  AND U3331 ( .A(n178), .B(n3338), .Z(n3337) );
  XOR U3332 ( .A(p_input[9]), .B(p_input[25]), .Z(n3338) );
  XOR U3333 ( .A(n3339), .B(n3340), .Z(n3330) );
  AND U3334 ( .A(n3341), .B(n3342), .Z(n3340) );
  XOR U3335 ( .A(n3339), .B(n2930), .Z(n3342) );
  XNOR U3336 ( .A(p_input[40]), .B(n3343), .Z(n2930) );
  AND U3337 ( .A(n181), .B(n3344), .Z(n3343) );
  XOR U3338 ( .A(p_input[56]), .B(p_input[40]), .Z(n3344) );
  XNOR U3339 ( .A(n2927), .B(n3339), .Z(n3341) );
  XOR U3340 ( .A(n3345), .B(n3346), .Z(n2927) );
  AND U3341 ( .A(n178), .B(n3347), .Z(n3346) );
  XOR U3342 ( .A(p_input[8]), .B(p_input[24]), .Z(n3347) );
  XOR U3343 ( .A(n3348), .B(n3349), .Z(n3339) );
  AND U3344 ( .A(n3350), .B(n3351), .Z(n3349) );
  XOR U3345 ( .A(n3348), .B(n2942), .Z(n3351) );
  XNOR U3346 ( .A(p_input[39]), .B(n3352), .Z(n2942) );
  AND U3347 ( .A(n181), .B(n3353), .Z(n3352) );
  XOR U3348 ( .A(p_input[55]), .B(p_input[39]), .Z(n3353) );
  XNOR U3349 ( .A(n2939), .B(n3348), .Z(n3350) );
  XOR U3350 ( .A(n3354), .B(n3355), .Z(n2939) );
  AND U3351 ( .A(n178), .B(n3356), .Z(n3355) );
  XOR U3352 ( .A(p_input[7]), .B(p_input[23]), .Z(n3356) );
  XOR U3353 ( .A(n3357), .B(n3358), .Z(n3348) );
  AND U3354 ( .A(n3359), .B(n3360), .Z(n3358) );
  XOR U3355 ( .A(n3357), .B(n2954), .Z(n3360) );
  XNOR U3356 ( .A(p_input[38]), .B(n3361), .Z(n2954) );
  AND U3357 ( .A(n181), .B(n3362), .Z(n3361) );
  XOR U3358 ( .A(p_input[54]), .B(p_input[38]), .Z(n3362) );
  XNOR U3359 ( .A(n2951), .B(n3357), .Z(n3359) );
  XOR U3360 ( .A(n3363), .B(n3364), .Z(n2951) );
  AND U3361 ( .A(n178), .B(n3365), .Z(n3364) );
  XOR U3362 ( .A(p_input[6]), .B(p_input[22]), .Z(n3365) );
  XOR U3363 ( .A(n3366), .B(n3367), .Z(n3357) );
  AND U3364 ( .A(n3368), .B(n3369), .Z(n3367) );
  XOR U3365 ( .A(n3366), .B(n2966), .Z(n3369) );
  XNOR U3366 ( .A(p_input[37]), .B(n3370), .Z(n2966) );
  AND U3367 ( .A(n181), .B(n3371), .Z(n3370) );
  XOR U3368 ( .A(p_input[53]), .B(p_input[37]), .Z(n3371) );
  XNOR U3369 ( .A(n2963), .B(n3366), .Z(n3368) );
  XOR U3370 ( .A(n3372), .B(n3373), .Z(n2963) );
  AND U3371 ( .A(n178), .B(n3374), .Z(n3373) );
  XOR U3372 ( .A(p_input[5]), .B(p_input[21]), .Z(n3374) );
  XOR U3373 ( .A(n3375), .B(n3376), .Z(n3366) );
  AND U3374 ( .A(n3377), .B(n3378), .Z(n3376) );
  XOR U3375 ( .A(n2978), .B(n3375), .Z(n3378) );
  XNOR U3376 ( .A(p_input[36]), .B(n3379), .Z(n2978) );
  AND U3377 ( .A(n181), .B(n3380), .Z(n3379) );
  XOR U3378 ( .A(p_input[52]), .B(p_input[36]), .Z(n3380) );
  XNOR U3379 ( .A(n3375), .B(n2975), .Z(n3377) );
  XOR U3380 ( .A(n3381), .B(n3382), .Z(n2975) );
  AND U3381 ( .A(n178), .B(n3383), .Z(n3382) );
  XOR U3382 ( .A(p_input[4]), .B(p_input[20]), .Z(n3383) );
  XOR U3383 ( .A(n3384), .B(n3385), .Z(n3375) );
  AND U3384 ( .A(n3386), .B(n3387), .Z(n3385) );
  XOR U3385 ( .A(n3384), .B(n2990), .Z(n3387) );
  XNOR U3386 ( .A(p_input[35]), .B(n3388), .Z(n2990) );
  AND U3387 ( .A(n181), .B(n3389), .Z(n3388) );
  XOR U3388 ( .A(p_input[51]), .B(p_input[35]), .Z(n3389) );
  XNOR U3389 ( .A(n2987), .B(n3384), .Z(n3386) );
  XOR U3390 ( .A(n3390), .B(n3391), .Z(n2987) );
  AND U3391 ( .A(n178), .B(n3392), .Z(n3391) );
  XOR U3392 ( .A(p_input[3]), .B(p_input[19]), .Z(n3392) );
  XOR U3393 ( .A(n3393), .B(n3394), .Z(n3384) );
  AND U3394 ( .A(n3395), .B(n3396), .Z(n3394) );
  XOR U3395 ( .A(n3393), .B(n3002), .Z(n3396) );
  XNOR U3396 ( .A(p_input[34]), .B(n3397), .Z(n3002) );
  AND U3397 ( .A(n181), .B(n3398), .Z(n3397) );
  XOR U3398 ( .A(p_input[50]), .B(p_input[34]), .Z(n3398) );
  XNOR U3399 ( .A(n2999), .B(n3393), .Z(n3395) );
  XOR U3400 ( .A(n3399), .B(n3400), .Z(n2999) );
  AND U3401 ( .A(n178), .B(n3401), .Z(n3400) );
  XOR U3402 ( .A(p_input[2]), .B(p_input[18]), .Z(n3401) );
  XOR U3403 ( .A(n3402), .B(n3403), .Z(n3393) );
  AND U3404 ( .A(n3404), .B(n3405), .Z(n3403) );
  XNOR U3405 ( .A(n3406), .B(n3015), .Z(n3405) );
  XNOR U3406 ( .A(p_input[33]), .B(n3407), .Z(n3015) );
  AND U3407 ( .A(n181), .B(n3408), .Z(n3407) );
  XNOR U3408 ( .A(p_input[49]), .B(n3409), .Z(n3408) );
  IV U3409 ( .A(p_input[33]), .Z(n3409) );
  XNOR U3410 ( .A(n3012), .B(n3402), .Z(n3404) );
  XNOR U3411 ( .A(p_input[1]), .B(n3410), .Z(n3012) );
  AND U3412 ( .A(n178), .B(n3411), .Z(n3410) );
  XOR U3413 ( .A(p_input[1]), .B(p_input[17]), .Z(n3411) );
  IV U3414 ( .A(n3406), .Z(n3402) );
  AND U3415 ( .A(n3277), .B(n3280), .Z(n3406) );
  XOR U3416 ( .A(p_input[32]), .B(n3412), .Z(n3280) );
  AND U3417 ( .A(n181), .B(n3413), .Z(n3412) );
  XOR U3418 ( .A(p_input[48]), .B(p_input[32]), .Z(n3413) );
  XOR U3419 ( .A(n3414), .B(n3415), .Z(n181) );
  AND U3420 ( .A(n3416), .B(n3417), .Z(n3415) );
  XNOR U3421 ( .A(p_input[63]), .B(n3414), .Z(n3417) );
  XOR U3422 ( .A(n3414), .B(p_input[47]), .Z(n3416) );
  XOR U3423 ( .A(n3418), .B(n3419), .Z(n3414) );
  AND U3424 ( .A(n3420), .B(n3421), .Z(n3419) );
  XNOR U3425 ( .A(p_input[62]), .B(n3418), .Z(n3421) );
  XOR U3426 ( .A(n3418), .B(p_input[46]), .Z(n3420) );
  XOR U3427 ( .A(n3422), .B(n3423), .Z(n3418) );
  AND U3428 ( .A(n3424), .B(n3425), .Z(n3423) );
  XNOR U3429 ( .A(p_input[61]), .B(n3422), .Z(n3425) );
  XOR U3430 ( .A(n3422), .B(p_input[45]), .Z(n3424) );
  XOR U3431 ( .A(n3426), .B(n3427), .Z(n3422) );
  AND U3432 ( .A(n3428), .B(n3429), .Z(n3427) );
  XNOR U3433 ( .A(p_input[60]), .B(n3426), .Z(n3429) );
  XOR U3434 ( .A(n3426), .B(p_input[44]), .Z(n3428) );
  XOR U3435 ( .A(n3430), .B(n3431), .Z(n3426) );
  AND U3436 ( .A(n3432), .B(n3433), .Z(n3431) );
  XNOR U3437 ( .A(p_input[59]), .B(n3430), .Z(n3433) );
  XOR U3438 ( .A(n3430), .B(p_input[43]), .Z(n3432) );
  XOR U3439 ( .A(n3434), .B(n3435), .Z(n3430) );
  AND U3440 ( .A(n3436), .B(n3437), .Z(n3435) );
  XNOR U3441 ( .A(p_input[58]), .B(n3434), .Z(n3437) );
  XOR U3442 ( .A(n3434), .B(p_input[42]), .Z(n3436) );
  XOR U3443 ( .A(n3438), .B(n3439), .Z(n3434) );
  AND U3444 ( .A(n3440), .B(n3441), .Z(n3439) );
  XNOR U3445 ( .A(p_input[57]), .B(n3438), .Z(n3441) );
  XOR U3446 ( .A(n3438), .B(p_input[41]), .Z(n3440) );
  XOR U3447 ( .A(n3442), .B(n3443), .Z(n3438) );
  AND U3448 ( .A(n3444), .B(n3445), .Z(n3443) );
  XNOR U3449 ( .A(p_input[56]), .B(n3442), .Z(n3445) );
  XOR U3450 ( .A(n3442), .B(p_input[40]), .Z(n3444) );
  XOR U3451 ( .A(n3446), .B(n3447), .Z(n3442) );
  AND U3452 ( .A(n3448), .B(n3449), .Z(n3447) );
  XNOR U3453 ( .A(p_input[55]), .B(n3446), .Z(n3449) );
  XOR U3454 ( .A(n3446), .B(p_input[39]), .Z(n3448) );
  XOR U3455 ( .A(n3450), .B(n3451), .Z(n3446) );
  AND U3456 ( .A(n3452), .B(n3453), .Z(n3451) );
  XNOR U3457 ( .A(p_input[54]), .B(n3450), .Z(n3453) );
  XOR U3458 ( .A(n3450), .B(p_input[38]), .Z(n3452) );
  XOR U3459 ( .A(n3454), .B(n3455), .Z(n3450) );
  AND U3460 ( .A(n3456), .B(n3457), .Z(n3455) );
  XNOR U3461 ( .A(p_input[53]), .B(n3454), .Z(n3457) );
  XOR U3462 ( .A(n3454), .B(p_input[37]), .Z(n3456) );
  XOR U3463 ( .A(n3458), .B(n3459), .Z(n3454) );
  AND U3464 ( .A(n3460), .B(n3461), .Z(n3459) );
  XNOR U3465 ( .A(p_input[52]), .B(n3458), .Z(n3461) );
  XOR U3466 ( .A(n3458), .B(p_input[36]), .Z(n3460) );
  XOR U3467 ( .A(n3462), .B(n3463), .Z(n3458) );
  AND U3468 ( .A(n3464), .B(n3465), .Z(n3463) );
  XNOR U3469 ( .A(p_input[51]), .B(n3462), .Z(n3465) );
  XOR U3470 ( .A(n3462), .B(p_input[35]), .Z(n3464) );
  XOR U3471 ( .A(n3466), .B(n3467), .Z(n3462) );
  AND U3472 ( .A(n3468), .B(n3469), .Z(n3467) );
  XNOR U3473 ( .A(p_input[50]), .B(n3466), .Z(n3469) );
  XOR U3474 ( .A(n3466), .B(p_input[34]), .Z(n3468) );
  XNOR U3475 ( .A(n3470), .B(n3471), .Z(n3466) );
  AND U3476 ( .A(n3472), .B(n3473), .Z(n3471) );
  XOR U3477 ( .A(p_input[49]), .B(n3470), .Z(n3473) );
  XNOR U3478 ( .A(p_input[33]), .B(n3470), .Z(n3472) );
  AND U3479 ( .A(p_input[48]), .B(n3474), .Z(n3470) );
  IV U3480 ( .A(p_input[32]), .Z(n3474) );
  XNOR U3481 ( .A(p_input[0]), .B(n3475), .Z(n3277) );
  AND U3482 ( .A(n178), .B(n3476), .Z(n3475) );
  XOR U3483 ( .A(p_input[16]), .B(p_input[0]), .Z(n3476) );
  XOR U3484 ( .A(n3477), .B(n3478), .Z(n178) );
  AND U3485 ( .A(n3479), .B(n3480), .Z(n3478) );
  XNOR U3486 ( .A(p_input[31]), .B(n3477), .Z(n3480) );
  XOR U3487 ( .A(n3477), .B(p_input[15]), .Z(n3479) );
  XOR U3488 ( .A(n3481), .B(n3482), .Z(n3477) );
  AND U3489 ( .A(n3483), .B(n3484), .Z(n3482) );
  XNOR U3490 ( .A(p_input[30]), .B(n3481), .Z(n3484) );
  XNOR U3491 ( .A(n3481), .B(n3291), .Z(n3483) );
  IV U3492 ( .A(p_input[14]), .Z(n3291) );
  XOR U3493 ( .A(n3485), .B(n3486), .Z(n3481) );
  AND U3494 ( .A(n3487), .B(n3488), .Z(n3486) );
  XNOR U3495 ( .A(p_input[29]), .B(n3485), .Z(n3488) );
  XNOR U3496 ( .A(n3485), .B(n3300), .Z(n3487) );
  IV U3497 ( .A(p_input[13]), .Z(n3300) );
  XOR U3498 ( .A(n3489), .B(n3490), .Z(n3485) );
  AND U3499 ( .A(n3491), .B(n3492), .Z(n3490) );
  XNOR U3500 ( .A(p_input[28]), .B(n3489), .Z(n3492) );
  XNOR U3501 ( .A(n3489), .B(n3309), .Z(n3491) );
  IV U3502 ( .A(p_input[12]), .Z(n3309) );
  XOR U3503 ( .A(n3493), .B(n3494), .Z(n3489) );
  AND U3504 ( .A(n3495), .B(n3496), .Z(n3494) );
  XNOR U3505 ( .A(p_input[27]), .B(n3493), .Z(n3496) );
  XNOR U3506 ( .A(n3493), .B(n3318), .Z(n3495) );
  IV U3507 ( .A(p_input[11]), .Z(n3318) );
  XOR U3508 ( .A(n3497), .B(n3498), .Z(n3493) );
  AND U3509 ( .A(n3499), .B(n3500), .Z(n3498) );
  XNOR U3510 ( .A(p_input[26]), .B(n3497), .Z(n3500) );
  XNOR U3511 ( .A(n3497), .B(n3327), .Z(n3499) );
  IV U3512 ( .A(p_input[10]), .Z(n3327) );
  XOR U3513 ( .A(n3501), .B(n3502), .Z(n3497) );
  AND U3514 ( .A(n3503), .B(n3504), .Z(n3502) );
  XNOR U3515 ( .A(p_input[25]), .B(n3501), .Z(n3504) );
  XNOR U3516 ( .A(n3501), .B(n3336), .Z(n3503) );
  IV U3517 ( .A(p_input[9]), .Z(n3336) );
  XOR U3518 ( .A(n3505), .B(n3506), .Z(n3501) );
  AND U3519 ( .A(n3507), .B(n3508), .Z(n3506) );
  XNOR U3520 ( .A(p_input[24]), .B(n3505), .Z(n3508) );
  XNOR U3521 ( .A(n3505), .B(n3345), .Z(n3507) );
  IV U3522 ( .A(p_input[8]), .Z(n3345) );
  XOR U3523 ( .A(n3509), .B(n3510), .Z(n3505) );
  AND U3524 ( .A(n3511), .B(n3512), .Z(n3510) );
  XNOR U3525 ( .A(p_input[23]), .B(n3509), .Z(n3512) );
  XNOR U3526 ( .A(n3509), .B(n3354), .Z(n3511) );
  IV U3527 ( .A(p_input[7]), .Z(n3354) );
  XOR U3528 ( .A(n3513), .B(n3514), .Z(n3509) );
  AND U3529 ( .A(n3515), .B(n3516), .Z(n3514) );
  XNOR U3530 ( .A(p_input[22]), .B(n3513), .Z(n3516) );
  XNOR U3531 ( .A(n3513), .B(n3363), .Z(n3515) );
  IV U3532 ( .A(p_input[6]), .Z(n3363) );
  XOR U3533 ( .A(n3517), .B(n3518), .Z(n3513) );
  AND U3534 ( .A(n3519), .B(n3520), .Z(n3518) );
  XNOR U3535 ( .A(p_input[21]), .B(n3517), .Z(n3520) );
  XNOR U3536 ( .A(n3517), .B(n3372), .Z(n3519) );
  IV U3537 ( .A(p_input[5]), .Z(n3372) );
  XOR U3538 ( .A(n3521), .B(n3522), .Z(n3517) );
  AND U3539 ( .A(n3523), .B(n3524), .Z(n3522) );
  XNOR U3540 ( .A(p_input[20]), .B(n3521), .Z(n3524) );
  XNOR U3541 ( .A(n3521), .B(n3381), .Z(n3523) );
  IV U3542 ( .A(p_input[4]), .Z(n3381) );
  XOR U3543 ( .A(n3525), .B(n3526), .Z(n3521) );
  AND U3544 ( .A(n3527), .B(n3528), .Z(n3526) );
  XNOR U3545 ( .A(p_input[19]), .B(n3525), .Z(n3528) );
  XNOR U3546 ( .A(n3525), .B(n3390), .Z(n3527) );
  IV U3547 ( .A(p_input[3]), .Z(n3390) );
  XOR U3548 ( .A(n3529), .B(n3530), .Z(n3525) );
  AND U3549 ( .A(n3531), .B(n3532), .Z(n3530) );
  XNOR U3550 ( .A(p_input[18]), .B(n3529), .Z(n3532) );
  XNOR U3551 ( .A(n3529), .B(n3399), .Z(n3531) );
  IV U3552 ( .A(p_input[2]), .Z(n3399) );
  XNOR U3553 ( .A(n3533), .B(n3534), .Z(n3529) );
  AND U3554 ( .A(n3535), .B(n3536), .Z(n3534) );
  XOR U3555 ( .A(p_input[17]), .B(n3533), .Z(n3536) );
  XNOR U3556 ( .A(p_input[1]), .B(n3533), .Z(n3535) );
  AND U3557 ( .A(p_input[16]), .B(n3537), .Z(n3533) );
  IV U3558 ( .A(p_input[0]), .Z(n3537) );
endmodule

